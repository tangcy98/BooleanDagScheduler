module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 ;
  assign n192 = x126 | x127 ;
  assign n271 = x126 & x127 ;
  assign n272 = x124 | x125 ;
  assign n31331 = ~x126 ;
  assign n273 = n31331 & n272 ;
  assign n191 = n271 | n273 ;
  assign n276 = x124 & n191 ;
  assign n277 = x122 | x123 ;
  assign n278 = x124 | n277 ;
  assign n31332 = ~n276 ;
  assign n279 = n31332 & n278 ;
  assign n31333 = ~x124 ;
  assign n275 = n31333 & n191 ;
  assign n31334 = ~n275 ;
  assign n280 = x125 & n31334 ;
  assign n31335 = ~n272 ;
  assign n281 = n31335 & n191 ;
  assign n282 = n280 | n281 ;
  assign n283 = n279 | n282 ;
  assign n31336 = ~n192 ;
  assign n284 = n31336 & n283 ;
  assign n31337 = ~x127 ;
  assign n274 = x126 & n31337 ;
  assign n286 = x126 | n272 ;
  assign n31338 = ~n274 ;
  assign n287 = n31338 & n286 ;
  assign n31339 = ~n287 ;
  assign n288 = x124 & n31339 ;
  assign n289 = n31333 & n277 ;
  assign n290 = n288 | n289 ;
  assign n291 = n282 & n290 ;
  assign n285 = x126 & n31335 ;
  assign n31340 = ~n273 ;
  assign n292 = x127 & n31340 ;
  assign n31341 = ~n285 ;
  assign n293 = n31341 & n292 ;
  assign n294 = n291 | n293 ;
  assign n190 = n284 | n294 ;
  assign n296 = x122 & n190 ;
  assign n298 = x120 | x121 ;
  assign n299 = x122 | n298 ;
  assign n31342 = ~n296 ;
  assign n300 = n31342 & n299 ;
  assign n31343 = ~n300 ;
  assign n301 = n191 & n31343 ;
  assign n31344 = ~n271 ;
  assign n302 = n31344 & n299 ;
  assign n303 = n31340 & n302 ;
  assign n304 = n31342 & n303 ;
  assign n305 = n282 | n290 ;
  assign n306 = n31336 & n305 ;
  assign n307 = n294 | n306 ;
  assign n31345 = ~n277 ;
  assign n308 = n31345 & n307 ;
  assign n31346 = ~x122 ;
  assign n309 = n31346 & n190 ;
  assign n31347 = ~n309 ;
  assign n310 = x123 & n31347 ;
  assign n311 = n308 | n310 ;
  assign n312 = n304 | n311 ;
  assign n31348 = ~n301 ;
  assign n313 = n31348 & n312 ;
  assign n31349 = ~n283 ;
  assign n322 = n31349 & n190 ;
  assign n323 = n291 | n322 ;
  assign n314 = n31345 & n190 ;
  assign n31350 = ~n293 ;
  assign n315 = n287 & n31350 ;
  assign n31351 = ~n291 ;
  assign n316 = n31351 & n315 ;
  assign n31352 = ~n284 ;
  assign n317 = n31352 & n316 ;
  assign n318 = n314 | n317 ;
  assign n319 = x124 & n318 ;
  assign n320 = x124 | n317 ;
  assign n321 = n314 | n320 ;
  assign n31353 = ~n319 ;
  assign n324 = n31353 & n321 ;
  assign n325 = n323 | n324 ;
  assign n326 = n313 | n325 ;
  assign n327 = n31336 & n326 ;
  assign n31354 = ~n282 ;
  assign n336 = n31354 & n190 ;
  assign n31355 = ~n336 ;
  assign n337 = n290 & n31355 ;
  assign n338 = n192 & n283 ;
  assign n31356 = ~n337 ;
  assign n339 = n31356 & n338 ;
  assign n340 = n282 & n31350 ;
  assign n341 = n31351 & n340 ;
  assign n342 = n31352 & n341 ;
  assign n343 = n339 | n342 ;
  assign n31357 = ~n190 ;
  assign n297 = x122 & n31357 ;
  assign n328 = n31346 & n298 ;
  assign n329 = n297 | n328 ;
  assign n31358 = ~n329 ;
  assign n333 = n287 & n31358 ;
  assign n330 = n31346 & n307 ;
  assign n31359 = ~n330 ;
  assign n331 = x123 & n31359 ;
  assign n332 = n314 | n331 ;
  assign n334 = n304 | n332 ;
  assign n31360 = ~n333 ;
  assign n335 = n31360 & n334 ;
  assign n344 = n324 & n335 ;
  assign n345 = n343 | n344 ;
  assign n189 = n327 | n345 ;
  assign n386 = n301 | n304 ;
  assign n31361 = ~n386 ;
  assign n387 = n332 & n31361 ;
  assign n389 = n189 & n387 ;
  assign n388 = n189 & n31361 ;
  assign n390 = n332 | n388 ;
  assign n31362 = ~n389 ;
  assign n391 = n31362 & n390 ;
  assign n392 = n313 & n324 ;
  assign n393 = n313 | n324 ;
  assign n31363 = ~n393 ;
  assign n394 = n189 & n31363 ;
  assign n395 = n392 | n394 ;
  assign n396 = n391 | n395 ;
  assign n348 = x120 & n189 ;
  assign n350 = x118 | x119 ;
  assign n351 = x120 | n350 ;
  assign n31364 = ~n348 ;
  assign n352 = n31364 & n351 ;
  assign n31365 = ~n352 ;
  assign n353 = n190 & n31365 ;
  assign n31366 = ~n298 ;
  assign n349 = n31366 & n189 ;
  assign n354 = n308 | n317 ;
  assign n355 = x124 & n354 ;
  assign n31367 = ~n355 ;
  assign n356 = n321 & n31367 ;
  assign n31368 = ~n305 ;
  assign n357 = n190 & n31368 ;
  assign n358 = n291 | n357 ;
  assign n359 = n356 | n358 ;
  assign n360 = n335 | n359 ;
  assign n361 = n31336 & n360 ;
  assign n362 = n345 | n361 ;
  assign n31369 = ~x120 ;
  assign n363 = n31369 & n362 ;
  assign n31370 = ~n363 ;
  assign n364 = x121 & n31370 ;
  assign n365 = n349 | n364 ;
  assign n367 = n31350 & n351 ;
  assign n368 = n31351 & n367 ;
  assign n369 = n31352 & n368 ;
  assign n370 = n31364 & n369 ;
  assign n371 = n365 | n370 ;
  assign n31371 = ~n353 ;
  assign n372 = n31371 & n371 ;
  assign n31372 = ~n372 ;
  assign n373 = n191 & n31372 ;
  assign n374 = n191 | n353 ;
  assign n31373 = ~n374 ;
  assign n375 = n371 & n31373 ;
  assign n31374 = ~n342 ;
  assign n376 = n190 & n31374 ;
  assign n31375 = ~n339 ;
  assign n377 = n31375 & n376 ;
  assign n31376 = ~n344 ;
  assign n378 = n31376 & n377 ;
  assign n31377 = ~n361 ;
  assign n379 = n31377 & n378 ;
  assign n380 = n349 | n379 ;
  assign n381 = x122 & n380 ;
  assign n382 = x122 | n379 ;
  assign n383 = n349 | n382 ;
  assign n31378 = ~n381 ;
  assign n384 = n31378 & n383 ;
  assign n385 = n375 | n384 ;
  assign n31379 = ~n373 ;
  assign n397 = n31379 & n385 ;
  assign n398 = n396 | n397 ;
  assign n399 = n31336 & n398 ;
  assign n347 = n313 & n189 ;
  assign n402 = n324 | n347 ;
  assign n31380 = ~n392 ;
  assign n403 = n192 & n31380 ;
  assign n404 = n402 & n403 ;
  assign n405 = n321 & n31374 ;
  assign n406 = n31353 & n405 ;
  assign n407 = n31375 & n406 ;
  assign n408 = n31380 & n407 ;
  assign n31381 = ~n327 ;
  assign n409 = n31381 & n408 ;
  assign n410 = n404 | n409 ;
  assign n400 = n287 & n31372 ;
  assign n31382 = ~n400 ;
  assign n401 = n391 & n31382 ;
  assign n411 = n385 & n401 ;
  assign n412 = n410 | n411 ;
  assign n413 = n399 | n412 ;
  assign n31383 = ~n189 ;
  assign n366 = x120 & n31383 ;
  assign n433 = n31369 & n350 ;
  assign n434 = n366 | n433 ;
  assign n31384 = ~n434 ;
  assign n435 = n190 & n31384 ;
  assign n436 = n287 | n435 ;
  assign n31385 = ~n436 ;
  assign n437 = n371 & n31385 ;
  assign n31386 = ~n437 ;
  assign n486 = n384 & n31386 ;
  assign n487 = n31379 & n486 ;
  assign n488 = n413 & n487 ;
  assign n438 = n384 | n437 ;
  assign n441 = n343 | n392 ;
  assign n442 = n327 | n441 ;
  assign n443 = n31369 & n442 ;
  assign n31387 = ~n443 ;
  assign n444 = x121 & n31387 ;
  assign n445 = n349 | n444 ;
  assign n446 = n370 | n445 ;
  assign n31388 = ~n435 ;
  assign n447 = n31388 & n446 ;
  assign n31389 = ~n447 ;
  assign n448 = n191 & n31389 ;
  assign n31390 = ~n448 ;
  assign n449 = n391 & n31390 ;
  assign n450 = n438 & n449 ;
  assign n451 = n410 | n450 ;
  assign n439 = n31382 & n438 ;
  assign n440 = n396 | n439 ;
  assign n452 = n31336 & n440 ;
  assign n188 = n451 | n452 ;
  assign n489 = n373 | n437 ;
  assign n31391 = ~n489 ;
  assign n490 = n188 & n31391 ;
  assign n491 = n384 | n490 ;
  assign n31392 = ~n488 ;
  assign n492 = n31392 & n491 ;
  assign n493 = n391 | n397 ;
  assign n31393 = ~n493 ;
  assign n494 = n413 & n31393 ;
  assign n495 = n411 | n494 ;
  assign n496 = n492 | n495 ;
  assign n31394 = ~n413 ;
  assign n414 = x118 & n31394 ;
  assign n415 = x116 | x117 ;
  assign n31395 = ~x118 ;
  assign n417 = n31395 & n415 ;
  assign n418 = n414 | n417 ;
  assign n31396 = ~n418 ;
  assign n429 = n189 & n31396 ;
  assign n419 = x118 & n413 ;
  assign n416 = x118 | n415 ;
  assign n420 = n31374 & n416 ;
  assign n421 = n31375 & n420 ;
  assign n422 = n31380 & n421 ;
  assign n423 = n31381 & n422 ;
  assign n31397 = ~n419 ;
  assign n424 = n31397 & n423 ;
  assign n425 = n31395 & n413 ;
  assign n31398 = ~n425 ;
  assign n426 = x119 & n31398 ;
  assign n31399 = ~n350 ;
  assign n427 = n31399 & n413 ;
  assign n428 = n426 | n427 ;
  assign n430 = n424 | n428 ;
  assign n31400 = ~n429 ;
  assign n431 = n31400 & n430 ;
  assign n31401 = ~n431 ;
  assign n432 = n190 & n31401 ;
  assign n454 = x118 & n188 ;
  assign n31402 = ~n454 ;
  assign n455 = n416 & n31402 ;
  assign n31403 = ~n455 ;
  assign n456 = n189 & n31403 ;
  assign n457 = n190 | n456 ;
  assign n31404 = ~n457 ;
  assign n458 = n430 & n31404 ;
  assign n31405 = ~n409 ;
  assign n460 = n189 & n31405 ;
  assign n31406 = ~n404 ;
  assign n461 = n31406 & n460 ;
  assign n31407 = ~n411 ;
  assign n462 = n31407 & n461 ;
  assign n31408 = ~n399 ;
  assign n463 = n31408 & n462 ;
  assign n464 = n427 | n463 ;
  assign n466 = x120 & n464 ;
  assign n465 = x120 | n463 ;
  assign n467 = n427 | n465 ;
  assign n31409 = ~n466 ;
  assign n468 = n31409 & n467 ;
  assign n469 = n458 | n468 ;
  assign n31410 = ~n432 ;
  assign n470 = n31410 & n469 ;
  assign n31411 = ~n470 ;
  assign n517 = n191 & n31411 ;
  assign n31412 = ~n370 ;
  assign n476 = n365 & n31412 ;
  assign n477 = n31388 & n476 ;
  assign n478 = n413 & n477 ;
  assign n479 = n370 | n435 ;
  assign n31413 = ~n479 ;
  assign n480 = n188 & n31413 ;
  assign n481 = n445 | n480 ;
  assign n31414 = ~n478 ;
  assign n483 = n31414 & n481 ;
  assign n472 = n190 | n429 ;
  assign n31415 = ~n472 ;
  assign n473 = n430 & n31415 ;
  assign n474 = n468 | n473 ;
  assign n518 = n191 | n432 ;
  assign n31416 = ~n518 ;
  assign n519 = n474 & n31416 ;
  assign n521 = n483 | n519 ;
  assign n31417 = ~n517 ;
  assign n522 = n31417 & n521 ;
  assign n523 = n496 | n522 ;
  assign n524 = n31336 & n523 ;
  assign n459 = n192 & n31407 ;
  assign n502 = n397 & n413 ;
  assign n503 = n391 | n502 ;
  assign n504 = n459 & n503 ;
  assign n505 = n389 | n409 ;
  assign n31418 = ~n505 ;
  assign n506 = n390 & n31418 ;
  assign n507 = n31406 & n506 ;
  assign n508 = n31407 & n507 ;
  assign n509 = n31408 & n508 ;
  assign n511 = n504 | n509 ;
  assign n471 = n287 & n31411 ;
  assign n31419 = ~n471 ;
  assign n525 = n31419 & n492 ;
  assign n526 = n521 & n525 ;
  assign n527 = n511 | n526 ;
  assign n528 = n524 | n527 ;
  assign n31420 = ~n528 ;
  assign n529 = x116 & n31420 ;
  assign n530 = x114 | x115 ;
  assign n31421 = ~x116 ;
  assign n532 = n31421 & n530 ;
  assign n533 = n529 | n532 ;
  assign n31422 = ~n533 ;
  assign n544 = n413 & n31422 ;
  assign n534 = x116 & n528 ;
  assign n531 = x116 | n530 ;
  assign n535 = n31405 & n531 ;
  assign n536 = n31406 & n535 ;
  assign n537 = n31407 & n536 ;
  assign n538 = n31408 & n537 ;
  assign n31423 = ~n534 ;
  assign n539 = n31423 & n538 ;
  assign n540 = n31421 & n528 ;
  assign n31424 = ~n540 ;
  assign n541 = x117 & n31424 ;
  assign n31425 = ~n415 ;
  assign n542 = n31425 & n528 ;
  assign n543 = n541 | n542 ;
  assign n545 = n539 | n543 ;
  assign n31426 = ~n544 ;
  assign n546 = n31426 & n545 ;
  assign n31427 = ~n546 ;
  assign n547 = n189 & n31427 ;
  assign n475 = n287 | n432 ;
  assign n31428 = ~n475 ;
  assign n482 = n474 & n31428 ;
  assign n484 = n482 | n483 ;
  assign n498 = n31410 & n474 ;
  assign n31429 = ~n498 ;
  assign n499 = n191 & n31429 ;
  assign n31430 = ~n499 ;
  assign n500 = n492 & n31430 ;
  assign n501 = n484 & n500 ;
  assign n512 = n501 | n511 ;
  assign n485 = n31419 & n484 ;
  assign n497 = n485 | n496 ;
  assign n513 = n31336 & n497 ;
  assign n187 = n512 | n513 ;
  assign n515 = x116 & n187 ;
  assign n31431 = ~n515 ;
  assign n548 = n31431 & n531 ;
  assign n31432 = ~n548 ;
  assign n549 = n188 & n31432 ;
  assign n550 = n189 | n549 ;
  assign n31433 = ~n550 ;
  assign n551 = n545 & n31433 ;
  assign n552 = n484 & n525 ;
  assign n31434 = ~n509 ;
  assign n553 = n413 & n31434 ;
  assign n31435 = ~n504 ;
  assign n554 = n31435 & n553 ;
  assign n31436 = ~n552 ;
  assign n555 = n31436 & n554 ;
  assign n31437 = ~n513 ;
  assign n556 = n31437 & n555 ;
  assign n557 = n542 | n556 ;
  assign n559 = x118 & n557 ;
  assign n558 = x118 | n556 ;
  assign n560 = n542 | n558 ;
  assign n31438 = ~n559 ;
  assign n561 = n31438 & n560 ;
  assign n562 = n551 | n561 ;
  assign n31439 = ~n547 ;
  assign n563 = n31439 & n562 ;
  assign n31440 = ~n563 ;
  assign n564 = n190 & n31440 ;
  assign n568 = n424 | n429 ;
  assign n31441 = ~n568 ;
  assign n570 = n428 & n31441 ;
  assign n571 = n528 & n570 ;
  assign n569 = n187 & n31441 ;
  assign n572 = n428 | n569 ;
  assign n31442 = ~n571 ;
  assign n573 = n31442 & n572 ;
  assign n565 = n189 | n544 ;
  assign n31443 = ~n565 ;
  assign n566 = n545 & n31443 ;
  assign n567 = n561 | n566 ;
  assign n574 = n190 | n547 ;
  assign n31444 = ~n574 ;
  assign n575 = n567 & n31444 ;
  assign n576 = n573 | n575 ;
  assign n31445 = ~n564 ;
  assign n577 = n31445 & n576 ;
  assign n31446 = ~n577 ;
  assign n578 = n191 & n31446 ;
  assign n31447 = ~n473 ;
  assign n579 = n468 & n31447 ;
  assign n580 = n31410 & n579 ;
  assign n581 = n187 & n580 ;
  assign n582 = n432 | n473 ;
  assign n31448 = ~n582 ;
  assign n583 = n187 & n31448 ;
  assign n584 = n468 | n583 ;
  assign n31449 = ~n581 ;
  assign n585 = n31449 & n584 ;
  assign n586 = n287 | n564 ;
  assign n31450 = ~n586 ;
  assign n587 = n576 & n31450 ;
  assign n588 = n585 | n587 ;
  assign n31451 = ~n578 ;
  assign n589 = n31451 & n588 ;
  assign n520 = n31419 & n483 ;
  assign n31452 = ~n482 ;
  assign n590 = n31452 & n520 ;
  assign n591 = n528 & n590 ;
  assign n592 = n471 | n482 ;
  assign n31453 = ~n592 ;
  assign n593 = n187 & n31453 ;
  assign n594 = n483 | n593 ;
  assign n31454 = ~n591 ;
  assign n595 = n31454 & n594 ;
  assign n597 = n485 | n492 ;
  assign n31455 = ~n597 ;
  assign n598 = n528 & n31455 ;
  assign n599 = n552 | n598 ;
  assign n600 = n595 | n599 ;
  assign n601 = n589 | n600 ;
  assign n602 = n31336 & n601 ;
  assign n31456 = ~n492 ;
  assign n516 = n31456 & n187 ;
  assign n31457 = ~n516 ;
  assign n606 = n485 & n31457 ;
  assign n607 = n192 & n597 ;
  assign n31458 = ~n606 ;
  assign n608 = n31458 & n607 ;
  assign n510 = n488 | n509 ;
  assign n31459 = ~n510 ;
  assign n609 = n491 & n31459 ;
  assign n610 = n31435 & n609 ;
  assign n611 = n31436 & n610 ;
  assign n612 = n31437 & n611 ;
  assign n613 = n608 | n612 ;
  assign n604 = n287 & n31446 ;
  assign n31460 = ~n604 ;
  assign n605 = n595 & n31460 ;
  assign n614 = n588 & n605 ;
  assign n615 = n613 | n614 ;
  assign n186 = n602 | n615 ;
  assign n619 = x114 & n186 ;
  assign n620 = x112 | x113 ;
  assign n621 = x114 | n620 ;
  assign n31461 = ~n619 ;
  assign n622 = n31461 & n621 ;
  assign n31462 = ~n622 ;
  assign n623 = n187 & n31462 ;
  assign n624 = n31434 & n621 ;
  assign n625 = n31435 & n624 ;
  assign n626 = n31436 & n625 ;
  assign n627 = n31437 & n626 ;
  assign n628 = n31461 & n627 ;
  assign n31463 = ~n530 ;
  assign n618 = n31463 & n186 ;
  assign n31464 = ~x114 ;
  assign n629 = n31464 & n186 ;
  assign n31465 = ~n629 ;
  assign n630 = x115 & n31465 ;
  assign n631 = n618 | n630 ;
  assign n632 = n628 | n631 ;
  assign n31466 = ~n623 ;
  assign n633 = n31466 & n632 ;
  assign n31467 = ~n633 ;
  assign n634 = n413 & n31467 ;
  assign n31468 = ~n186 ;
  assign n617 = x114 & n31468 ;
  assign n635 = n31464 & n620 ;
  assign n636 = n617 | n635 ;
  assign n31469 = ~n636 ;
  assign n637 = n528 & n31469 ;
  assign n638 = n413 | n637 ;
  assign n31470 = ~n638 ;
  assign n647 = n632 & n31470 ;
  assign n31471 = ~n612 ;
  assign n639 = n528 & n31471 ;
  assign n31472 = ~n608 ;
  assign n640 = n31472 & n639 ;
  assign n31473 = ~n614 ;
  assign n641 = n31473 & n640 ;
  assign n31474 = ~n602 ;
  assign n642 = n31474 & n641 ;
  assign n643 = n618 | n642 ;
  assign n644 = x116 & n643 ;
  assign n645 = x116 | n642 ;
  assign n646 = n618 | n645 ;
  assign n31475 = ~n644 ;
  assign n648 = n31475 & n646 ;
  assign n649 = n647 | n648 ;
  assign n31476 = ~n634 ;
  assign n650 = n31476 & n649 ;
  assign n31477 = ~n650 ;
  assign n651 = n189 & n31477 ;
  assign n652 = n539 | n544 ;
  assign n31478 = ~n652 ;
  assign n653 = n543 & n31478 ;
  assign n655 = n186 & n653 ;
  assign n654 = n186 & n31478 ;
  assign n656 = n543 | n654 ;
  assign n31479 = ~n655 ;
  assign n657 = n31479 & n656 ;
  assign n658 = n189 | n634 ;
  assign n31480 = ~n658 ;
  assign n659 = n649 & n31480 ;
  assign n660 = n657 | n659 ;
  assign n31481 = ~n651 ;
  assign n661 = n31481 & n660 ;
  assign n31482 = ~n661 ;
  assign n662 = n190 & n31482 ;
  assign n31483 = ~n566 ;
  assign n663 = n561 & n31483 ;
  assign n664 = n31439 & n663 ;
  assign n667 = n186 & n664 ;
  assign n665 = n547 | n566 ;
  assign n31484 = ~n665 ;
  assign n666 = n186 & n31484 ;
  assign n668 = n561 | n666 ;
  assign n31485 = ~n667 ;
  assign n669 = n31485 & n668 ;
  assign n670 = n190 | n651 ;
  assign n31486 = ~n670 ;
  assign n671 = n660 & n31486 ;
  assign n672 = n669 | n671 ;
  assign n31487 = ~n662 ;
  assign n673 = n31487 & n672 ;
  assign n31488 = ~n673 ;
  assign n674 = n287 & n31488 ;
  assign n603 = n31445 & n573 ;
  assign n31489 = ~n575 ;
  assign n675 = n31489 & n603 ;
  assign n676 = n186 & n675 ;
  assign n677 = n564 | n575 ;
  assign n31490 = ~n677 ;
  assign n678 = n186 & n31490 ;
  assign n679 = n573 | n678 ;
  assign n31491 = ~n676 ;
  assign n680 = n31491 & n679 ;
  assign n681 = n188 & n31467 ;
  assign n682 = n188 | n623 ;
  assign n31492 = ~n682 ;
  assign n683 = n632 & n31492 ;
  assign n684 = n648 | n683 ;
  assign n31493 = ~n681 ;
  assign n685 = n31493 & n684 ;
  assign n31494 = ~n685 ;
  assign n686 = n189 & n31494 ;
  assign n687 = n31480 & n684 ;
  assign n688 = n657 | n687 ;
  assign n31495 = ~n686 ;
  assign n689 = n31495 & n688 ;
  assign n31496 = ~n689 ;
  assign n690 = n190 & n31496 ;
  assign n691 = n287 | n690 ;
  assign n31497 = ~n691 ;
  assign n692 = n672 & n31497 ;
  assign n693 = n680 | n692 ;
  assign n31498 = ~n674 ;
  assign n694 = n31498 & n693 ;
  assign n31499 = ~n587 ;
  assign n695 = n585 & n31499 ;
  assign n696 = n31460 & n695 ;
  assign n697 = n186 & n696 ;
  assign n698 = n587 | n604 ;
  assign n31500 = ~n698 ;
  assign n699 = n186 & n31500 ;
  assign n700 = n585 | n699 ;
  assign n31501 = ~n697 ;
  assign n701 = n31501 & n700 ;
  assign n596 = n589 | n595 ;
  assign n31502 = ~n596 ;
  assign n703 = n31502 & n186 ;
  assign n704 = n614 | n703 ;
  assign n705 = n701 | n704 ;
  assign n706 = n694 | n705 ;
  assign n707 = n31336 & n706 ;
  assign n710 = n192 & n596 ;
  assign n31503 = ~n595 ;
  assign n709 = n31503 & n186 ;
  assign n31504 = ~n709 ;
  assign n711 = n589 & n31504 ;
  assign n31505 = ~n711 ;
  assign n712 = n710 & n31505 ;
  assign n713 = n591 | n612 ;
  assign n31506 = ~n713 ;
  assign n714 = n594 & n31506 ;
  assign n715 = n31472 & n714 ;
  assign n716 = n31473 & n715 ;
  assign n717 = n31474 & n716 ;
  assign n718 = n712 | n717 ;
  assign n708 = n31498 & n701 ;
  assign n719 = n693 & n708 ;
  assign n720 = n718 | n719 ;
  assign n185 = n707 | n720 ;
  assign n702 = n694 | n701 ;
  assign n827 = n192 & n702 ;
  assign n31507 = ~n701 ;
  assign n826 = n31507 & n185 ;
  assign n31508 = ~n826 ;
  assign n828 = n694 & n31508 ;
  assign n31509 = ~n828 ;
  assign n829 = n827 & n31509 ;
  assign n830 = n697 | n717 ;
  assign n31510 = ~n830 ;
  assign n831 = n700 & n31510 ;
  assign n31511 = ~n712 ;
  assign n832 = n31511 & n831 ;
  assign n31512 = ~n719 ;
  assign n833 = n31512 & n832 ;
  assign n31513 = ~n707 ;
  assign n834 = n31513 & n833 ;
  assign n835 = n829 | n834 ;
  assign n722 = x112 & n185 ;
  assign n724 = x110 | x111 ;
  assign n725 = x112 | n724 ;
  assign n31514 = ~n722 ;
  assign n726 = n31514 & n725 ;
  assign n31515 = ~n726 ;
  assign n727 = n186 & n31515 ;
  assign n31516 = ~n620 ;
  assign n723 = n31516 & n185 ;
  assign n31517 = ~x112 ;
  assign n728 = n31517 & n185 ;
  assign n31518 = ~n728 ;
  assign n729 = x113 & n31518 ;
  assign n730 = n723 | n729 ;
  assign n732 = n31471 & n725 ;
  assign n733 = n31472 & n732 ;
  assign n734 = n31473 & n733 ;
  assign n735 = n31474 & n734 ;
  assign n736 = n31514 & n735 ;
  assign n737 = n730 | n736 ;
  assign n31519 = ~n727 ;
  assign n738 = n31519 & n737 ;
  assign n31520 = ~n738 ;
  assign n739 = n528 & n31520 ;
  assign n31521 = ~n717 ;
  assign n744 = n186 & n31521 ;
  assign n745 = n31511 & n744 ;
  assign n746 = n31512 & n745 ;
  assign n747 = n31513 & n746 ;
  assign n748 = n723 | n747 ;
  assign n750 = x114 & n748 ;
  assign n749 = x114 | n747 ;
  assign n751 = n723 | n749 ;
  assign n31522 = ~n750 ;
  assign n752 = n31522 & n751 ;
  assign n31523 = ~n185 ;
  assign n731 = x112 & n31523 ;
  assign n740 = n31517 & n724 ;
  assign n741 = n731 | n740 ;
  assign n31524 = ~n741 ;
  assign n742 = n186 & n31524 ;
  assign n743 = n528 | n742 ;
  assign n31525 = ~n743 ;
  assign n753 = n737 & n31525 ;
  assign n754 = n752 | n753 ;
  assign n31526 = ~n739 ;
  assign n755 = n31526 & n754 ;
  assign n31527 = ~n755 ;
  assign n756 = n413 & n31527 ;
  assign n757 = n628 | n637 ;
  assign n31528 = ~n757 ;
  assign n758 = n631 & n31528 ;
  assign n759 = n185 & n758 ;
  assign n760 = n185 & n31528 ;
  assign n761 = n631 | n760 ;
  assign n31529 = ~n759 ;
  assign n762 = n31529 & n761 ;
  assign n763 = n413 | n739 ;
  assign n31530 = ~n763 ;
  assign n764 = n754 & n31530 ;
  assign n765 = n762 | n764 ;
  assign n31531 = ~n756 ;
  assign n766 = n31531 & n765 ;
  assign n31532 = ~n766 ;
  assign n767 = n189 & n31532 ;
  assign n31533 = ~n647 ;
  assign n768 = n31533 & n648 ;
  assign n770 = n31476 & n768 ;
  assign n772 = n185 & n770 ;
  assign n769 = n634 | n647 ;
  assign n31534 = ~n769 ;
  assign n771 = n185 & n31534 ;
  assign n773 = n648 | n771 ;
  assign n31535 = ~n772 ;
  assign n774 = n31535 & n773 ;
  assign n775 = n189 | n756 ;
  assign n31536 = ~n775 ;
  assign n776 = n765 & n31536 ;
  assign n777 = n774 | n776 ;
  assign n31537 = ~n767 ;
  assign n778 = n31537 & n777 ;
  assign n31538 = ~n778 ;
  assign n779 = n190 & n31538 ;
  assign n780 = n31481 & n657 ;
  assign n31539 = ~n659 ;
  assign n781 = n31539 & n780 ;
  assign n782 = n185 & n781 ;
  assign n783 = n651 | n659 ;
  assign n31540 = ~n783 ;
  assign n784 = n185 & n31540 ;
  assign n785 = n657 | n784 ;
  assign n31541 = ~n782 ;
  assign n786 = n31541 & n785 ;
  assign n787 = n187 & n31520 ;
  assign n788 = n187 | n727 ;
  assign n31542 = ~n788 ;
  assign n789 = n737 & n31542 ;
  assign n790 = n752 | n789 ;
  assign n31543 = ~n787 ;
  assign n791 = n31543 & n790 ;
  assign n31544 = ~n791 ;
  assign n792 = n188 & n31544 ;
  assign n793 = n31530 & n790 ;
  assign n794 = n762 | n793 ;
  assign n31545 = ~n792 ;
  assign n795 = n31545 & n794 ;
  assign n31546 = ~n795 ;
  assign n796 = n189 & n31546 ;
  assign n797 = n190 | n796 ;
  assign n31547 = ~n797 ;
  assign n798 = n777 & n31547 ;
  assign n799 = n786 | n798 ;
  assign n31548 = ~n779 ;
  assign n800 = n31548 & n799 ;
  assign n31549 = ~n800 ;
  assign n801 = n191 & n31549 ;
  assign n812 = n31498 & n680 ;
  assign n31550 = ~n692 ;
  assign n813 = n31550 & n812 ;
  assign n814 = n185 & n813 ;
  assign n815 = n674 | n692 ;
  assign n31551 = ~n815 ;
  assign n816 = n185 & n31551 ;
  assign n817 = n680 | n816 ;
  assign n31552 = ~n814 ;
  assign n818 = n31552 & n817 ;
  assign n31553 = ~n801 ;
  assign n825 = n31553 & n818 ;
  assign n31554 = ~n671 ;
  assign n802 = n669 & n31554 ;
  assign n803 = n31487 & n802 ;
  assign n804 = n185 & n803 ;
  assign n805 = n671 | n690 ;
  assign n31555 = ~n805 ;
  assign n806 = n185 & n31555 ;
  assign n807 = n669 | n806 ;
  assign n31556 = ~n804 ;
  assign n808 = n31556 & n807 ;
  assign n858 = n191 | n779 ;
  assign n31557 = ~n858 ;
  assign n859 = n799 & n31557 ;
  assign n860 = n808 | n859 ;
  assign n863 = n825 & n860 ;
  assign n864 = n835 | n863 ;
  assign n31558 = ~n702 ;
  assign n819 = n31558 & n185 ;
  assign n820 = n719 | n819 ;
  assign n821 = n818 | n820 ;
  assign n861 = n31553 & n860 ;
  assign n862 = n821 | n861 ;
  assign n865 = n31336 & n862 ;
  assign n184 = n864 | n865 ;
  assign n809 = n287 | n779 ;
  assign n31559 = ~n809 ;
  assign n810 = n799 & n31559 ;
  assign n811 = n808 | n810 ;
  assign n822 = n31553 & n811 ;
  assign n823 = n821 | n822 ;
  assign n824 = n31336 & n823 ;
  assign n836 = n811 & n825 ;
  assign n837 = n835 | n836 ;
  assign n838 = n824 | n837 ;
  assign n31560 = ~n859 ;
  assign n958 = n808 & n31560 ;
  assign n959 = n31553 & n958 ;
  assign n960 = n838 & n959 ;
  assign n961 = n801 | n859 ;
  assign n31561 = ~n961 ;
  assign n962 = n184 & n31561 ;
  assign n963 = n808 | n962 ;
  assign n31562 = ~n960 ;
  assign n964 = n31562 & n963 ;
  assign n965 = n818 | n822 ;
  assign n31563 = ~n965 ;
  assign n966 = n184 & n31563 ;
  assign n967 = n836 | n966 ;
  assign n968 = n964 | n967 ;
  assign n31564 = ~n838 ;
  assign n839 = x110 & n31564 ;
  assign n840 = x108 | x109 ;
  assign n31565 = ~x110 ;
  assign n842 = n31565 & n840 ;
  assign n843 = n839 | n842 ;
  assign n31566 = ~n843 ;
  assign n844 = n185 & n31566 ;
  assign n845 = x110 & n838 ;
  assign n841 = x110 | n840 ;
  assign n846 = n31521 & n841 ;
  assign n847 = n31511 & n846 ;
  assign n848 = n31512 & n847 ;
  assign n849 = n31513 & n848 ;
  assign n31567 = ~n845 ;
  assign n850 = n31567 & n849 ;
  assign n851 = n31565 & n838 ;
  assign n31568 = ~n851 ;
  assign n852 = x111 & n31568 ;
  assign n31569 = ~n724 ;
  assign n853 = n31569 & n838 ;
  assign n854 = n852 | n853 ;
  assign n855 = n850 | n854 ;
  assign n31570 = ~n844 ;
  assign n856 = n31570 & n855 ;
  assign n31571 = ~n856 ;
  assign n857 = n186 & n31571 ;
  assign n867 = x110 & n184 ;
  assign n31572 = ~n867 ;
  assign n868 = n841 & n31572 ;
  assign n31573 = ~n868 ;
  assign n869 = n185 & n31573 ;
  assign n870 = n186 | n869 ;
  assign n31574 = ~n870 ;
  assign n871 = n855 & n31574 ;
  assign n31575 = ~n834 ;
  assign n872 = n185 & n31575 ;
  assign n31576 = ~n829 ;
  assign n873 = n31576 & n872 ;
  assign n31577 = ~n836 ;
  assign n874 = n31577 & n873 ;
  assign n31578 = ~n824 ;
  assign n875 = n31578 & n874 ;
  assign n876 = n853 | n875 ;
  assign n878 = x112 & n876 ;
  assign n877 = x112 | n875 ;
  assign n879 = n853 | n877 ;
  assign n31579 = ~n878 ;
  assign n880 = n31579 & n879 ;
  assign n881 = n871 | n880 ;
  assign n31580 = ~n857 ;
  assign n882 = n31580 & n881 ;
  assign n31581 = ~n882 ;
  assign n883 = n528 & n31581 ;
  assign n31582 = ~n736 ;
  assign n890 = n730 & n31582 ;
  assign n31583 = ~n742 ;
  assign n891 = n31583 & n890 ;
  assign n892 = n838 & n891 ;
  assign n893 = n736 | n742 ;
  assign n31584 = ~n893 ;
  assign n894 = n184 & n31584 ;
  assign n895 = n730 | n894 ;
  assign n31585 = ~n892 ;
  assign n896 = n31585 & n895 ;
  assign n884 = n186 | n844 ;
  assign n31586 = ~n884 ;
  assign n885 = n855 & n31586 ;
  assign n886 = n880 | n885 ;
  assign n31587 = ~n869 ;
  assign n887 = n855 & n31587 ;
  assign n31588 = ~n887 ;
  assign n888 = n186 & n31588 ;
  assign n889 = n528 | n888 ;
  assign n31589 = ~n889 ;
  assign n897 = n886 & n31589 ;
  assign n898 = n896 | n897 ;
  assign n31590 = ~n883 ;
  assign n899 = n31590 & n898 ;
  assign n31591 = ~n899 ;
  assign n900 = n413 & n31591 ;
  assign n31592 = ~n753 ;
  assign n901 = n752 & n31592 ;
  assign n902 = n31526 & n901 ;
  assign n903 = n838 & n902 ;
  assign n904 = n739 | n753 ;
  assign n31593 = ~n904 ;
  assign n905 = n184 & n31593 ;
  assign n906 = n752 | n905 ;
  assign n31594 = ~n903 ;
  assign n907 = n31594 & n906 ;
  assign n908 = n413 | n883 ;
  assign n31595 = ~n908 ;
  assign n909 = n898 & n31595 ;
  assign n910 = n907 | n909 ;
  assign n31596 = ~n900 ;
  assign n911 = n31596 & n910 ;
  assign n31597 = ~n911 ;
  assign n912 = n189 & n31597 ;
  assign n913 = n31531 & n762 ;
  assign n31598 = ~n764 ;
  assign n914 = n31598 & n913 ;
  assign n915 = n838 & n914 ;
  assign n916 = n756 | n764 ;
  assign n31599 = ~n916 ;
  assign n917 = n838 & n31599 ;
  assign n918 = n762 | n917 ;
  assign n31600 = ~n915 ;
  assign n919 = n31600 & n918 ;
  assign n920 = n189 | n900 ;
  assign n31601 = ~n920 ;
  assign n921 = n910 & n31601 ;
  assign n922 = n919 | n921 ;
  assign n31602 = ~n912 ;
  assign n923 = n31602 & n922 ;
  assign n31603 = ~n923 ;
  assign n924 = n190 & n31603 ;
  assign n31604 = ~n776 ;
  assign n925 = n774 & n31604 ;
  assign n926 = n31537 & n925 ;
  assign n927 = n184 & n926 ;
  assign n928 = n767 | n776 ;
  assign n31605 = ~n928 ;
  assign n929 = n184 & n31605 ;
  assign n930 = n774 | n929 ;
  assign n31606 = ~n927 ;
  assign n931 = n31606 & n930 ;
  assign n932 = n187 & n31581 ;
  assign n933 = n187 | n857 ;
  assign n31607 = ~n933 ;
  assign n934 = n886 & n31607 ;
  assign n935 = n896 | n934 ;
  assign n31608 = ~n932 ;
  assign n936 = n31608 & n935 ;
  assign n31609 = ~n936 ;
  assign n937 = n188 & n31609 ;
  assign n938 = n31595 & n935 ;
  assign n939 = n907 | n938 ;
  assign n31610 = ~n937 ;
  assign n940 = n31610 & n939 ;
  assign n31611 = ~n940 ;
  assign n941 = n189 & n31611 ;
  assign n942 = n190 | n941 ;
  assign n31612 = ~n942 ;
  assign n943 = n922 & n31612 ;
  assign n944 = n931 | n943 ;
  assign n31613 = ~n924 ;
  assign n945 = n31613 & n944 ;
  assign n31614 = ~n945 ;
  assign n946 = n191 & n31614 ;
  assign n947 = n31548 & n786 ;
  assign n31615 = ~n798 ;
  assign n948 = n31615 & n947 ;
  assign n949 = n838 & n948 ;
  assign n950 = n779 | n798 ;
  assign n31616 = ~n950 ;
  assign n951 = n184 & n31616 ;
  assign n952 = n786 | n951 ;
  assign n31617 = ~n949 ;
  assign n953 = n31617 & n952 ;
  assign n988 = n287 | n924 ;
  assign n31618 = ~n988 ;
  assign n989 = n944 & n31618 ;
  assign n990 = n953 | n989 ;
  assign n31619 = ~n946 ;
  assign n991 = n31619 & n990 ;
  assign n992 = n968 | n991 ;
  assign n993 = n31336 & n992 ;
  assign n31620 = ~n818 ;
  assign n972 = n31620 & n838 ;
  assign n31621 = ~n972 ;
  assign n973 = n822 & n31621 ;
  assign n974 = n192 & n965 ;
  assign n31622 = ~n973 ;
  assign n975 = n31622 & n974 ;
  assign n976 = n814 | n834 ;
  assign n31623 = ~n976 ;
  assign n977 = n817 & n31623 ;
  assign n978 = n31576 & n977 ;
  assign n979 = n31577 & n978 ;
  assign n980 = n31578 & n979 ;
  assign n981 = n975 | n980 ;
  assign n970 = n31619 & n964 ;
  assign n994 = n970 & n990 ;
  assign n995 = n981 | n994 ;
  assign n996 = n993 | n995 ;
  assign n31624 = ~n996 ;
  assign n997 = x108 & n31624 ;
  assign n998 = x106 | x107 ;
  assign n31625 = ~x108 ;
  assign n1000 = n31625 & n998 ;
  assign n1001 = n997 | n1000 ;
  assign n31626 = ~n1001 ;
  assign n1010 = n838 & n31626 ;
  assign n954 = n191 | n924 ;
  assign n31627 = ~n954 ;
  assign n955 = n944 & n31627 ;
  assign n956 = n953 | n955 ;
  assign n971 = n956 & n970 ;
  assign n982 = n971 | n981 ;
  assign n957 = n31619 & n956 ;
  assign n969 = n957 | n968 ;
  assign n983 = n31336 & n969 ;
  assign n183 = n982 | n983 ;
  assign n986 = x108 & n183 ;
  assign n999 = x108 | n998 ;
  assign n1002 = n31575 & n999 ;
  assign n1003 = n31576 & n1002 ;
  assign n1004 = n31577 & n1003 ;
  assign n1005 = n31578 & n1004 ;
  assign n31628 = ~n986 ;
  assign n1006 = n31628 & n1005 ;
  assign n987 = n31625 & n183 ;
  assign n31629 = ~n987 ;
  assign n1007 = x109 & n31629 ;
  assign n31630 = ~n840 ;
  assign n1008 = n31630 & n183 ;
  assign n1009 = n1007 | n1008 ;
  assign n1011 = n1006 | n1009 ;
  assign n31631 = ~n1010 ;
  assign n1012 = n31631 & n1011 ;
  assign n31632 = ~n1012 ;
  assign n1013 = n185 & n31632 ;
  assign n1014 = n31628 & n999 ;
  assign n31633 = ~n1014 ;
  assign n1015 = n184 & n31633 ;
  assign n1016 = n185 | n1015 ;
  assign n31634 = ~n1016 ;
  assign n1017 = n1011 & n31634 ;
  assign n31635 = ~n980 ;
  assign n1018 = n838 & n31635 ;
  assign n31636 = ~n975 ;
  assign n1019 = n31636 & n1018 ;
  assign n31637 = ~n971 ;
  assign n1020 = n31637 & n1019 ;
  assign n31638 = ~n983 ;
  assign n1021 = n31638 & n1020 ;
  assign n1022 = n1008 | n1021 ;
  assign n1024 = x110 & n1022 ;
  assign n1023 = x110 | n1021 ;
  assign n1025 = n1008 | n1023 ;
  assign n31639 = ~n1024 ;
  assign n1026 = n31639 & n1025 ;
  assign n1027 = n1017 | n1026 ;
  assign n31640 = ~n1013 ;
  assign n1028 = n31640 & n1027 ;
  assign n31641 = ~n1028 ;
  assign n1029 = n186 & n31641 ;
  assign n1033 = n844 | n850 ;
  assign n31642 = ~n1033 ;
  assign n1035 = n854 & n31642 ;
  assign n1036 = n183 & n1035 ;
  assign n1034 = n183 & n31642 ;
  assign n1037 = n854 | n1034 ;
  assign n31643 = ~n1036 ;
  assign n1038 = n31643 & n1037 ;
  assign n1030 = n185 | n1010 ;
  assign n31644 = ~n1030 ;
  assign n1031 = n1011 & n31644 ;
  assign n1032 = n1026 | n1031 ;
  assign n1040 = n186 | n1013 ;
  assign n31645 = ~n1040 ;
  assign n1041 = n1032 & n31645 ;
  assign n1042 = n1038 | n1041 ;
  assign n31646 = ~n1029 ;
  assign n1043 = n31646 & n1042 ;
  assign n31647 = ~n1043 ;
  assign n1044 = n528 & n31647 ;
  assign n31648 = ~n885 ;
  assign n1045 = n880 & n31648 ;
  assign n31649 = ~n888 ;
  assign n1046 = n31649 & n1045 ;
  assign n1047 = n183 & n1046 ;
  assign n1048 = n885 | n888 ;
  assign n31650 = ~n1048 ;
  assign n1049 = n183 & n31650 ;
  assign n1050 = n880 | n1049 ;
  assign n31651 = ~n1047 ;
  assign n1051 = n31651 & n1050 ;
  assign n1052 = n528 | n1029 ;
  assign n31652 = ~n1052 ;
  assign n1053 = n1042 & n31652 ;
  assign n1054 = n1051 | n1053 ;
  assign n31653 = ~n1044 ;
  assign n1055 = n31653 & n1054 ;
  assign n31654 = ~n1055 ;
  assign n1056 = n188 & n31654 ;
  assign n1058 = n896 & n31608 ;
  assign n31655 = ~n897 ;
  assign n1059 = n31655 & n1058 ;
  assign n1060 = n183 & n1059 ;
  assign n1061 = n883 | n897 ;
  assign n31656 = ~n1061 ;
  assign n1062 = n183 & n31656 ;
  assign n1063 = n896 | n1062 ;
  assign n31657 = ~n1060 ;
  assign n1064 = n31657 & n1063 ;
  assign n1057 = n413 | n1044 ;
  assign n31658 = ~n1057 ;
  assign n1065 = n1054 & n31658 ;
  assign n1066 = n1064 | n1065 ;
  assign n31659 = ~n1056 ;
  assign n1067 = n31659 & n1066 ;
  assign n31660 = ~n1067 ;
  assign n1068 = n189 & n31660 ;
  assign n31661 = ~n909 ;
  assign n1069 = n907 & n31661 ;
  assign n1070 = n31596 & n1069 ;
  assign n1071 = n183 & n1070 ;
  assign n1072 = n900 | n909 ;
  assign n31662 = ~n1072 ;
  assign n1073 = n183 & n31662 ;
  assign n1074 = n907 | n1073 ;
  assign n31663 = ~n1071 ;
  assign n1075 = n31663 & n1074 ;
  assign n1076 = n187 & n31647 ;
  assign n31664 = ~n1076 ;
  assign n1077 = n1054 & n31664 ;
  assign n31665 = ~n1077 ;
  assign n1078 = n413 & n31665 ;
  assign n1079 = n189 | n1078 ;
  assign n31666 = ~n1079 ;
  assign n1080 = n1066 & n31666 ;
  assign n1081 = n1075 | n1080 ;
  assign n31667 = ~n1068 ;
  assign n1082 = n31667 & n1081 ;
  assign n31668 = ~n1082 ;
  assign n1083 = n190 & n31668 ;
  assign n31669 = ~n941 ;
  assign n1086 = n919 & n31669 ;
  assign n31670 = ~n921 ;
  assign n1087 = n31670 & n1086 ;
  assign n1088 = n183 & n1087 ;
  assign n1084 = n912 | n921 ;
  assign n31671 = ~n1084 ;
  assign n1085 = n183 & n31671 ;
  assign n1089 = n919 | n1085 ;
  assign n31672 = ~n1088 ;
  assign n1090 = n31672 & n1089 ;
  assign n1091 = n190 | n1068 ;
  assign n31673 = ~n1091 ;
  assign n1092 = n1081 & n31673 ;
  assign n1093 = n1090 | n1092 ;
  assign n31674 = ~n1083 ;
  assign n1094 = n31674 & n1093 ;
  assign n31675 = ~n1094 ;
  assign n1095 = n287 & n31675 ;
  assign n31676 = ~n943 ;
  assign n1096 = n931 & n31676 ;
  assign n1097 = n31613 & n1096 ;
  assign n1098 = n183 & n1097 ;
  assign n1099 = n924 | n943 ;
  assign n31677 = ~n1099 ;
  assign n1100 = n996 & n31677 ;
  assign n1101 = n931 | n1100 ;
  assign n31678 = ~n1098 ;
  assign n1102 = n31678 & n1101 ;
  assign n31679 = ~n1078 ;
  assign n1103 = n1066 & n31679 ;
  assign n31680 = ~n1103 ;
  assign n1104 = n189 & n31680 ;
  assign n31681 = ~n1104 ;
  assign n1105 = n1081 & n31681 ;
  assign n31682 = ~n1105 ;
  assign n1106 = n190 & n31682 ;
  assign n1107 = n287 | n1106 ;
  assign n31683 = ~n1107 ;
  assign n1108 = n1093 & n31683 ;
  assign n1109 = n1102 | n1108 ;
  assign n31684 = ~n1095 ;
  assign n1110 = n31684 & n1109 ;
  assign n1111 = n31619 & n953 ;
  assign n31685 = ~n955 ;
  assign n1112 = n31685 & n1111 ;
  assign n1113 = n183 & n1112 ;
  assign n1114 = n946 | n955 ;
  assign n31686 = ~n1114 ;
  assign n1115 = n183 & n31686 ;
  assign n1116 = n953 | n1115 ;
  assign n31687 = ~n1113 ;
  assign n1117 = n31687 & n1116 ;
  assign n1119 = n957 | n964 ;
  assign n31688 = ~n1119 ;
  assign n1120 = n183 & n31688 ;
  assign n1121 = n971 | n1120 ;
  assign n1122 = n1117 | n1121 ;
  assign n1123 = n1110 | n1122 ;
  assign n1124 = n31336 & n1123 ;
  assign n31689 = ~n964 ;
  assign n985 = n31689 & n183 ;
  assign n31690 = ~n985 ;
  assign n1126 = n957 & n31690 ;
  assign n1127 = n192 & n1119 ;
  assign n31691 = ~n1126 ;
  assign n1128 = n31691 & n1127 ;
  assign n1129 = n960 | n980 ;
  assign n31692 = ~n1129 ;
  assign n1130 = n963 & n31692 ;
  assign n1131 = n31636 & n1130 ;
  assign n1132 = n31637 & n1131 ;
  assign n1133 = n31638 & n1132 ;
  assign n1134 = n1128 | n1133 ;
  assign n1125 = n31684 & n1117 ;
  assign n1135 = n1109 & n1125 ;
  assign n1136 = n1134 | n1135 ;
  assign n182 = n1124 | n1136 ;
  assign n1140 = x106 & n182 ;
  assign n1141 = x104 | x105 ;
  assign n1142 = x106 | n1141 ;
  assign n31693 = ~n1140 ;
  assign n1143 = n31693 & n1142 ;
  assign n31694 = ~n1143 ;
  assign n1144 = n183 & n31694 ;
  assign n1145 = n31635 & n1142 ;
  assign n1146 = n31636 & n1145 ;
  assign n1147 = n31637 & n1146 ;
  assign n1148 = n31638 & n1147 ;
  assign n1149 = n31693 & n1148 ;
  assign n31695 = ~n998 ;
  assign n1139 = n31695 & n182 ;
  assign n31696 = ~x106 ;
  assign n1150 = n31696 & n182 ;
  assign n31697 = ~n1150 ;
  assign n1151 = x107 & n31697 ;
  assign n1152 = n1139 | n1151 ;
  assign n1153 = n1149 | n1152 ;
  assign n31698 = ~n1144 ;
  assign n1154 = n31698 & n1153 ;
  assign n31699 = ~n1154 ;
  assign n1155 = n838 & n31699 ;
  assign n31700 = ~n1133 ;
  assign n1160 = n996 & n31700 ;
  assign n31701 = ~n1128 ;
  assign n1161 = n31701 & n1160 ;
  assign n31702 = ~n1135 ;
  assign n1162 = n31702 & n1161 ;
  assign n31703 = ~n1124 ;
  assign n1163 = n31703 & n1162 ;
  assign n1164 = n1139 | n1163 ;
  assign n1166 = x108 & n1164 ;
  assign n1165 = x108 | n1163 ;
  assign n1167 = n1139 | n1165 ;
  assign n31704 = ~n1166 ;
  assign n1168 = n31704 & n1167 ;
  assign n31705 = ~n182 ;
  assign n1138 = x106 & n31705 ;
  assign n1156 = n31696 & n1141 ;
  assign n1157 = n1138 | n1156 ;
  assign n31706 = ~n1157 ;
  assign n1158 = n996 & n31706 ;
  assign n1159 = n838 | n1158 ;
  assign n31707 = ~n1159 ;
  assign n1169 = n1153 & n31707 ;
  assign n1170 = n1168 | n1169 ;
  assign n31708 = ~n1155 ;
  assign n1171 = n31708 & n1170 ;
  assign n31709 = ~n1171 ;
  assign n1172 = n185 & n31709 ;
  assign n1173 = n1006 | n1010 ;
  assign n31710 = ~n1173 ;
  assign n1174 = n1009 & n31710 ;
  assign n1176 = n182 & n1174 ;
  assign n1175 = n182 & n31710 ;
  assign n1177 = n1009 | n1175 ;
  assign n31711 = ~n1176 ;
  assign n1178 = n31711 & n1177 ;
  assign n1179 = n185 | n1155 ;
  assign n31712 = ~n1179 ;
  assign n1180 = n1170 & n31712 ;
  assign n1181 = n1178 | n1180 ;
  assign n31713 = ~n1172 ;
  assign n1182 = n31713 & n1181 ;
  assign n31714 = ~n1182 ;
  assign n1183 = n186 & n31714 ;
  assign n31715 = ~n1031 ;
  assign n1184 = n1026 & n31715 ;
  assign n1185 = n31640 & n1184 ;
  assign n1186 = n182 & n1185 ;
  assign n1187 = n1013 | n1031 ;
  assign n31716 = ~n1187 ;
  assign n1188 = n182 & n31716 ;
  assign n1189 = n1026 | n1188 ;
  assign n31717 = ~n1186 ;
  assign n1190 = n31717 & n1189 ;
  assign n1191 = n186 | n1172 ;
  assign n31718 = ~n1191 ;
  assign n1192 = n1181 & n31718 ;
  assign n1193 = n1190 | n1192 ;
  assign n31719 = ~n1183 ;
  assign n1194 = n31719 & n1193 ;
  assign n31720 = ~n1194 ;
  assign n1195 = n528 & n31720 ;
  assign n1039 = n31646 & n1038 ;
  assign n31721 = ~n1041 ;
  assign n1196 = n1039 & n31721 ;
  assign n1199 = n182 & n1196 ;
  assign n1197 = n1029 | n1041 ;
  assign n31722 = ~n1197 ;
  assign n1198 = n182 & n31722 ;
  assign n1200 = n1038 | n1198 ;
  assign n31723 = ~n1199 ;
  assign n1201 = n31723 & n1200 ;
  assign n1202 = n184 & n31699 ;
  assign n1203 = n184 | n1144 ;
  assign n31724 = ~n1203 ;
  assign n1204 = n1153 & n31724 ;
  assign n1205 = n1168 | n1204 ;
  assign n31725 = ~n1202 ;
  assign n1206 = n31725 & n1205 ;
  assign n31726 = ~n1206 ;
  assign n1207 = n185 & n31726 ;
  assign n1208 = n31712 & n1205 ;
  assign n1209 = n1178 | n1208 ;
  assign n31727 = ~n1207 ;
  assign n1210 = n31727 & n1209 ;
  assign n31728 = ~n1210 ;
  assign n1211 = n186 & n31728 ;
  assign n1212 = n528 | n1211 ;
  assign n31729 = ~n1212 ;
  assign n1213 = n1193 & n31729 ;
  assign n1214 = n1201 | n1213 ;
  assign n31730 = ~n1195 ;
  assign n1215 = n31730 & n1214 ;
  assign n31731 = ~n1215 ;
  assign n1216 = n188 & n31731 ;
  assign n31732 = ~n1053 ;
  assign n1217 = n1051 & n31732 ;
  assign n1218 = n31653 & n1217 ;
  assign n1219 = n182 & n1218 ;
  assign n1220 = n1044 | n1053 ;
  assign n31733 = ~n1220 ;
  assign n1221 = n182 & n31733 ;
  assign n1222 = n1051 | n1221 ;
  assign n31734 = ~n1219 ;
  assign n1223 = n31734 & n1222 ;
  assign n1224 = n413 | n1195 ;
  assign n31735 = ~n1224 ;
  assign n1225 = n1214 & n31735 ;
  assign n1226 = n1223 | n1225 ;
  assign n31736 = ~n1216 ;
  assign n1227 = n31736 & n1226 ;
  assign n31737 = ~n1227 ;
  assign n1228 = n189 & n31737 ;
  assign n1229 = n31718 & n1209 ;
  assign n1230 = n1190 | n1229 ;
  assign n31738 = ~n1211 ;
  assign n1231 = n31738 & n1230 ;
  assign n31739 = ~n1231 ;
  assign n1232 = n187 & n31739 ;
  assign n1233 = n31729 & n1230 ;
  assign n1234 = n1201 | n1233 ;
  assign n31740 = ~n1232 ;
  assign n1235 = n31740 & n1234 ;
  assign n31741 = ~n1235 ;
  assign n1236 = n413 & n31741 ;
  assign n1237 = n189 | n1236 ;
  assign n31742 = ~n1237 ;
  assign n1238 = n1226 & n31742 ;
  assign n1239 = n1064 & n31679 ;
  assign n31743 = ~n1065 ;
  assign n1240 = n31743 & n1239 ;
  assign n1241 = n182 & n1240 ;
  assign n1242 = n1056 | n1065 ;
  assign n31744 = ~n1242 ;
  assign n1243 = n182 & n31744 ;
  assign n1244 = n1064 | n1243 ;
  assign n31745 = ~n1241 ;
  assign n1245 = n31745 & n1244 ;
  assign n1246 = n1238 | n1245 ;
  assign n31746 = ~n1228 ;
  assign n1247 = n31746 & n1246 ;
  assign n31747 = ~n1247 ;
  assign n1248 = n190 & n31747 ;
  assign n31748 = ~n1080 ;
  assign n1249 = n1075 & n31748 ;
  assign n1250 = n31667 & n1249 ;
  assign n1251 = n182 & n1250 ;
  assign n1252 = n1068 | n1080 ;
  assign n31749 = ~n1252 ;
  assign n1253 = n182 & n31749 ;
  assign n1254 = n1075 | n1253 ;
  assign n31750 = ~n1251 ;
  assign n1255 = n31750 & n1254 ;
  assign n1256 = n190 | n1228 ;
  assign n31751 = ~n1256 ;
  assign n1257 = n1246 & n31751 ;
  assign n1258 = n1255 | n1257 ;
  assign n31752 = ~n1248 ;
  assign n1259 = n31752 & n1258 ;
  assign n31753 = ~n1259 ;
  assign n1260 = n287 & n31753 ;
  assign n31754 = ~n1106 ;
  assign n1263 = n1090 & n31754 ;
  assign n31755 = ~n1092 ;
  assign n1264 = n31755 & n1263 ;
  assign n1265 = n182 & n1264 ;
  assign n1261 = n1083 | n1092 ;
  assign n31756 = ~n1261 ;
  assign n1262 = n182 & n31756 ;
  assign n1266 = n1090 | n1262 ;
  assign n31757 = ~n1265 ;
  assign n1267 = n31757 & n1266 ;
  assign n1268 = n31735 & n1234 ;
  assign n1269 = n1223 | n1268 ;
  assign n31758 = ~n1236 ;
  assign n1270 = n31758 & n1269 ;
  assign n31759 = ~n1270 ;
  assign n1271 = n189 & n31759 ;
  assign n1272 = n31742 & n1269 ;
  assign n1273 = n1245 | n1272 ;
  assign n31760 = ~n1271 ;
  assign n1274 = n31760 & n1273 ;
  assign n31761 = ~n1274 ;
  assign n1275 = n190 & n31761 ;
  assign n1276 = n287 | n1275 ;
  assign n31762 = ~n1276 ;
  assign n1277 = n1258 & n31762 ;
  assign n1278 = n1267 | n1277 ;
  assign n31763 = ~n1260 ;
  assign n1279 = n31763 & n1278 ;
  assign n31764 = ~n1108 ;
  assign n1280 = n1102 & n31764 ;
  assign n1281 = n31684 & n1280 ;
  assign n1282 = n182 & n1281 ;
  assign n1283 = n1095 | n1108 ;
  assign n31765 = ~n1283 ;
  assign n1284 = n182 & n31765 ;
  assign n1285 = n1102 | n1284 ;
  assign n31766 = ~n1282 ;
  assign n1286 = n31766 & n1285 ;
  assign n1118 = n1110 | n1117 ;
  assign n31767 = ~n1118 ;
  assign n1288 = n31767 & n182 ;
  assign n1289 = n1135 | n1288 ;
  assign n1290 = n1286 | n1289 ;
  assign n1291 = n1279 | n1290 ;
  assign n1292 = n31336 & n1291 ;
  assign n1295 = n192 & n1118 ;
  assign n31768 = ~n1117 ;
  assign n1294 = n31768 & n182 ;
  assign n31769 = ~n1294 ;
  assign n1296 = n1110 & n31769 ;
  assign n31770 = ~n1296 ;
  assign n1297 = n1295 & n31770 ;
  assign n1298 = n1113 | n1133 ;
  assign n31771 = ~n1298 ;
  assign n1299 = n1116 & n31771 ;
  assign n1300 = n31701 & n1299 ;
  assign n1301 = n31702 & n1300 ;
  assign n1302 = n31703 & n1301 ;
  assign n1303 = n1297 | n1302 ;
  assign n1293 = n31763 & n1286 ;
  assign n1304 = n1278 & n1293 ;
  assign n1305 = n1303 | n1304 ;
  assign n181 = n1292 | n1305 ;
  assign n1287 = n1279 | n1286 ;
  assign n1476 = n192 & n1287 ;
  assign n31772 = ~n1286 ;
  assign n1475 = n31772 & n181 ;
  assign n31773 = ~n1475 ;
  assign n1477 = n1279 & n31773 ;
  assign n31774 = ~n1477 ;
  assign n1478 = n1476 & n31774 ;
  assign n1479 = n1282 | n1302 ;
  assign n31775 = ~n1479 ;
  assign n1480 = n1285 & n31775 ;
  assign n31776 = ~n1297 ;
  assign n1481 = n31776 & n1480 ;
  assign n31777 = ~n1304 ;
  assign n1482 = n31777 & n1481 ;
  assign n31778 = ~n1292 ;
  assign n1483 = n31778 & n1482 ;
  assign n1484 = n1478 | n1483 ;
  assign n1307 = x104 & n181 ;
  assign n1309 = x102 | x103 ;
  assign n1310 = x104 | n1309 ;
  assign n31779 = ~n1307 ;
  assign n1311 = n31779 & n1310 ;
  assign n31780 = ~n1311 ;
  assign n1312 = n182 & n31780 ;
  assign n1314 = n31700 & n1310 ;
  assign n1315 = n31701 & n1314 ;
  assign n1316 = n31702 & n1315 ;
  assign n1317 = n31703 & n1316 ;
  assign n1318 = n31779 & n1317 ;
  assign n31781 = ~n1141 ;
  assign n1308 = n31781 & n181 ;
  assign n31782 = ~x104 ;
  assign n1319 = n31782 & n181 ;
  assign n31783 = ~n1319 ;
  assign n1320 = x105 & n31783 ;
  assign n1321 = n1308 | n1320 ;
  assign n1322 = n1318 | n1321 ;
  assign n31784 = ~n1312 ;
  assign n1323 = n31784 & n1322 ;
  assign n31785 = ~n1323 ;
  assign n1324 = n996 & n31785 ;
  assign n31786 = ~n1302 ;
  assign n1329 = n182 & n31786 ;
  assign n1330 = n31776 & n1329 ;
  assign n1331 = n31777 & n1330 ;
  assign n1332 = n31778 & n1331 ;
  assign n1333 = n1308 | n1332 ;
  assign n1335 = x106 & n1333 ;
  assign n1334 = x106 | n1332 ;
  assign n1336 = n1308 | n1334 ;
  assign n31787 = ~n1335 ;
  assign n1337 = n31787 & n1336 ;
  assign n31788 = ~n181 ;
  assign n1313 = x104 & n31788 ;
  assign n1325 = n31782 & n1309 ;
  assign n1326 = n1313 | n1325 ;
  assign n31789 = ~n1326 ;
  assign n1327 = n182 & n31789 ;
  assign n1328 = n996 | n1327 ;
  assign n31790 = ~n1328 ;
  assign n1338 = n1322 & n31790 ;
  assign n1339 = n1337 | n1338 ;
  assign n31791 = ~n1324 ;
  assign n1340 = n31791 & n1339 ;
  assign n31792 = ~n1340 ;
  assign n1341 = n838 & n31792 ;
  assign n1342 = n1149 | n1158 ;
  assign n31793 = ~n1342 ;
  assign n1343 = n1152 & n31793 ;
  assign n1344 = n181 & n1343 ;
  assign n1345 = n181 & n31793 ;
  assign n1346 = n1152 | n1345 ;
  assign n31794 = ~n1344 ;
  assign n1347 = n31794 & n1346 ;
  assign n1348 = n838 | n1324 ;
  assign n31795 = ~n1348 ;
  assign n1349 = n1339 & n31795 ;
  assign n1350 = n1347 | n1349 ;
  assign n31796 = ~n1341 ;
  assign n1351 = n31796 & n1350 ;
  assign n31797 = ~n1351 ;
  assign n1352 = n185 & n31797 ;
  assign n31798 = ~n1169 ;
  assign n1353 = n1168 & n31798 ;
  assign n1355 = n31708 & n1353 ;
  assign n1356 = n181 & n1355 ;
  assign n1354 = n1155 | n1169 ;
  assign n31799 = ~n1354 ;
  assign n1357 = n181 & n31799 ;
  assign n1358 = n1168 | n1357 ;
  assign n31800 = ~n1356 ;
  assign n1359 = n31800 & n1358 ;
  assign n1360 = n185 | n1341 ;
  assign n31801 = ~n1360 ;
  assign n1361 = n1350 & n31801 ;
  assign n1362 = n1359 | n1361 ;
  assign n31802 = ~n1352 ;
  assign n1363 = n31802 & n1362 ;
  assign n31803 = ~n1363 ;
  assign n1364 = n186 & n31803 ;
  assign n1365 = n31713 & n1178 ;
  assign n31804 = ~n1180 ;
  assign n1366 = n31804 & n1365 ;
  assign n1367 = n181 & n1366 ;
  assign n1368 = n1172 | n1180 ;
  assign n31805 = ~n1368 ;
  assign n1369 = n181 & n31805 ;
  assign n1370 = n1178 | n1369 ;
  assign n31806 = ~n1367 ;
  assign n1371 = n31806 & n1370 ;
  assign n1372 = n183 & n31785 ;
  assign n1373 = n183 | n1312 ;
  assign n31807 = ~n1373 ;
  assign n1374 = n1322 & n31807 ;
  assign n1375 = n1337 | n1374 ;
  assign n31808 = ~n1372 ;
  assign n1376 = n31808 & n1375 ;
  assign n31809 = ~n1376 ;
  assign n1377 = n184 & n31809 ;
  assign n1378 = n31795 & n1375 ;
  assign n1379 = n1347 | n1378 ;
  assign n31810 = ~n1377 ;
  assign n1380 = n31810 & n1379 ;
  assign n31811 = ~n1380 ;
  assign n1381 = n185 & n31811 ;
  assign n1382 = n186 | n1381 ;
  assign n31812 = ~n1382 ;
  assign n1383 = n1362 & n31812 ;
  assign n1384 = n1371 | n1383 ;
  assign n31813 = ~n1364 ;
  assign n1385 = n31813 & n1384 ;
  assign n31814 = ~n1385 ;
  assign n1386 = n187 & n31814 ;
  assign n31815 = ~n1192 ;
  assign n1387 = n1190 & n31815 ;
  assign n1388 = n31719 & n1387 ;
  assign n1389 = n181 & n1388 ;
  assign n1390 = n1192 | n1211 ;
  assign n31816 = ~n1390 ;
  assign n1391 = n181 & n31816 ;
  assign n1392 = n1190 | n1391 ;
  assign n31817 = ~n1389 ;
  assign n1393 = n31817 & n1392 ;
  assign n1394 = n528 | n1364 ;
  assign n31818 = ~n1394 ;
  assign n1395 = n1384 & n31818 ;
  assign n1396 = n1393 | n1395 ;
  assign n31819 = ~n1386 ;
  assign n1397 = n31819 & n1396 ;
  assign n31820 = ~n1397 ;
  assign n1398 = n413 & n31820 ;
  assign n1399 = n31730 & n1201 ;
  assign n31821 = ~n1213 ;
  assign n1400 = n31821 & n1399 ;
  assign n1401 = n181 & n1400 ;
  assign n1402 = n1195 | n1213 ;
  assign n31822 = ~n1402 ;
  assign n1403 = n181 & n31822 ;
  assign n1404 = n1201 | n1403 ;
  assign n31823 = ~n1401 ;
  assign n1405 = n31823 & n1404 ;
  assign n1406 = n31801 & n1379 ;
  assign n1407 = n1359 | n1406 ;
  assign n31824 = ~n1381 ;
  assign n1408 = n31824 & n1407 ;
  assign n31825 = ~n1408 ;
  assign n1409 = n186 & n31825 ;
  assign n1410 = n31812 & n1407 ;
  assign n1411 = n1371 | n1410 ;
  assign n31826 = ~n1409 ;
  assign n1412 = n31826 & n1411 ;
  assign n31827 = ~n1412 ;
  assign n1413 = n528 & n31827 ;
  assign n1414 = n413 | n1413 ;
  assign n31828 = ~n1414 ;
  assign n1415 = n1396 & n31828 ;
  assign n1416 = n1405 | n1415 ;
  assign n31829 = ~n1398 ;
  assign n1417 = n31829 & n1416 ;
  assign n31830 = ~n1417 ;
  assign n1418 = n189 & n31830 ;
  assign n31831 = ~n1225 ;
  assign n1419 = n1223 & n31831 ;
  assign n1420 = n31736 & n1419 ;
  assign n1421 = n181 & n1420 ;
  assign n1422 = n1225 | n1236 ;
  assign n31832 = ~n1422 ;
  assign n1423 = n181 & n31832 ;
  assign n1424 = n1223 | n1423 ;
  assign n31833 = ~n1421 ;
  assign n1425 = n31833 & n1424 ;
  assign n1426 = n189 | n1398 ;
  assign n31834 = ~n1426 ;
  assign n1427 = n1416 & n31834 ;
  assign n1428 = n1425 | n1427 ;
  assign n31835 = ~n1418 ;
  assign n1429 = n31835 & n1428 ;
  assign n31836 = ~n1429 ;
  assign n1430 = n190 & n31836 ;
  assign n1431 = n31818 & n1411 ;
  assign n1432 = n1393 | n1431 ;
  assign n31837 = ~n1413 ;
  assign n1433 = n31837 & n1432 ;
  assign n31838 = ~n1433 ;
  assign n1434 = n188 & n31838 ;
  assign n1435 = n31828 & n1432 ;
  assign n1436 = n1405 | n1435 ;
  assign n31839 = ~n1434 ;
  assign n1437 = n31839 & n1436 ;
  assign n31840 = ~n1437 ;
  assign n1438 = n189 & n31840 ;
  assign n1439 = n190 | n1438 ;
  assign n31841 = ~n1439 ;
  assign n1440 = n1428 & n31841 ;
  assign n1441 = n31746 & n1245 ;
  assign n31842 = ~n1238 ;
  assign n1442 = n31842 & n1441 ;
  assign n1443 = n181 & n1442 ;
  assign n1444 = n1228 | n1238 ;
  assign n31843 = ~n1444 ;
  assign n1445 = n181 & n31843 ;
  assign n1446 = n1245 | n1445 ;
  assign n31844 = ~n1443 ;
  assign n1447 = n31844 & n1446 ;
  assign n1448 = n1440 | n1447 ;
  assign n31845 = ~n1430 ;
  assign n1449 = n31845 & n1448 ;
  assign n31846 = ~n1449 ;
  assign n1450 = n191 & n31846 ;
  assign n1461 = n31763 & n1267 ;
  assign n31847 = ~n1277 ;
  assign n1462 = n31847 & n1461 ;
  assign n1463 = n181 & n1462 ;
  assign n1464 = n1260 | n1277 ;
  assign n31848 = ~n1464 ;
  assign n1465 = n181 & n31848 ;
  assign n1466 = n1267 | n1465 ;
  assign n31849 = ~n1463 ;
  assign n1467 = n31849 & n1466 ;
  assign n31850 = ~n1450 ;
  assign n1474 = n31850 & n1467 ;
  assign n31851 = ~n1257 ;
  assign n1451 = n1255 & n31851 ;
  assign n1452 = n31752 & n1451 ;
  assign n1453 = n181 & n1452 ;
  assign n1454 = n1257 | n1275 ;
  assign n31852 = ~n1454 ;
  assign n1455 = n181 & n31852 ;
  assign n1456 = n1255 | n1455 ;
  assign n31853 = ~n1453 ;
  assign n1457 = n31853 & n1456 ;
  assign n1507 = n191 | n1430 ;
  assign n31854 = ~n1507 ;
  assign n1508 = n1448 & n31854 ;
  assign n1509 = n1457 | n1508 ;
  assign n1512 = n1474 & n1509 ;
  assign n1513 = n1484 | n1512 ;
  assign n31855 = ~n1287 ;
  assign n1468 = n31855 & n181 ;
  assign n1469 = n1304 | n1468 ;
  assign n1470 = n1467 | n1469 ;
  assign n1510 = n31850 & n1509 ;
  assign n1511 = n1470 | n1510 ;
  assign n1514 = n31336 & n1511 ;
  assign n180 = n1513 | n1514 ;
  assign n1458 = n287 | n1430 ;
  assign n31856 = ~n1458 ;
  assign n1459 = n1448 & n31856 ;
  assign n1460 = n1457 | n1459 ;
  assign n1471 = n31850 & n1460 ;
  assign n1472 = n1470 | n1471 ;
  assign n1473 = n31336 & n1472 ;
  assign n1485 = n1460 & n1474 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = n1473 | n1486 ;
  assign n31857 = ~n1508 ;
  assign n1671 = n1457 & n31857 ;
  assign n1672 = n31850 & n1671 ;
  assign n1673 = n1487 & n1672 ;
  assign n1674 = n1450 | n1508 ;
  assign n31858 = ~n1674 ;
  assign n1675 = n180 & n31858 ;
  assign n1676 = n1457 | n1675 ;
  assign n31859 = ~n1673 ;
  assign n1677 = n31859 & n1676 ;
  assign n1678 = n1467 | n1471 ;
  assign n31860 = ~n1678 ;
  assign n1679 = n180 & n31860 ;
  assign n1680 = n1485 | n1679 ;
  assign n1681 = n1677 | n1680 ;
  assign n31861 = ~n1487 ;
  assign n1488 = x102 & n31861 ;
  assign n1489 = x100 | x101 ;
  assign n31862 = ~x102 ;
  assign n1491 = n31862 & n1489 ;
  assign n1492 = n1488 | n1491 ;
  assign n31863 = ~n1492 ;
  assign n1493 = n181 & n31863 ;
  assign n1494 = x102 & n1487 ;
  assign n1490 = x102 | n1489 ;
  assign n1495 = n31786 & n1490 ;
  assign n1496 = n31776 & n1495 ;
  assign n1497 = n31777 & n1496 ;
  assign n1498 = n31778 & n1497 ;
  assign n31864 = ~n1494 ;
  assign n1499 = n31864 & n1498 ;
  assign n1500 = n31862 & n1487 ;
  assign n31865 = ~n1500 ;
  assign n1501 = x103 & n31865 ;
  assign n31866 = ~n1309 ;
  assign n1502 = n31866 & n1487 ;
  assign n1503 = n1501 | n1502 ;
  assign n1504 = n1499 | n1503 ;
  assign n31867 = ~n1493 ;
  assign n1505 = n31867 & n1504 ;
  assign n31868 = ~n1505 ;
  assign n1506 = n182 & n31868 ;
  assign n1516 = x102 & n180 ;
  assign n31869 = ~n1516 ;
  assign n1517 = n1490 & n31869 ;
  assign n31870 = ~n1517 ;
  assign n1518 = n181 & n31870 ;
  assign n1519 = n182 | n1518 ;
  assign n31871 = ~n1519 ;
  assign n1520 = n1504 & n31871 ;
  assign n31872 = ~n1483 ;
  assign n1521 = n181 & n31872 ;
  assign n31873 = ~n1478 ;
  assign n1522 = n31873 & n1521 ;
  assign n31874 = ~n1485 ;
  assign n1523 = n31874 & n1522 ;
  assign n31875 = ~n1473 ;
  assign n1524 = n31875 & n1523 ;
  assign n1525 = n1502 | n1524 ;
  assign n1527 = x104 & n1525 ;
  assign n1526 = x104 | n1524 ;
  assign n1528 = n1502 | n1526 ;
  assign n31876 = ~n1527 ;
  assign n1529 = n31876 & n1528 ;
  assign n1530 = n1520 | n1529 ;
  assign n31877 = ~n1506 ;
  assign n1531 = n31877 & n1530 ;
  assign n31878 = ~n1531 ;
  assign n1532 = n996 & n31878 ;
  assign n1536 = n1312 | n1318 ;
  assign n31879 = ~n1536 ;
  assign n1538 = n1321 & n31879 ;
  assign n1539 = n1487 & n1538 ;
  assign n1537 = n180 & n31879 ;
  assign n1540 = n1321 | n1537 ;
  assign n31880 = ~n1539 ;
  assign n1541 = n31880 & n1540 ;
  assign n1533 = n182 | n1493 ;
  assign n31881 = ~n1533 ;
  assign n1534 = n1504 & n31881 ;
  assign n1535 = n1529 | n1534 ;
  assign n31882 = ~n1518 ;
  assign n1543 = n1504 & n31882 ;
  assign n31883 = ~n1543 ;
  assign n1544 = n182 & n31883 ;
  assign n1545 = n996 | n1544 ;
  assign n31884 = ~n1545 ;
  assign n1546 = n1535 & n31884 ;
  assign n1547 = n1541 | n1546 ;
  assign n31885 = ~n1532 ;
  assign n1548 = n31885 & n1547 ;
  assign n31886 = ~n1548 ;
  assign n1549 = n838 & n31886 ;
  assign n31887 = ~n1338 ;
  assign n1550 = n1337 & n31887 ;
  assign n1551 = n31791 & n1550 ;
  assign n1552 = n1487 & n1551 ;
  assign n1553 = n1324 | n1338 ;
  assign n31888 = ~n1553 ;
  assign n1554 = n180 & n31888 ;
  assign n1555 = n1337 | n1554 ;
  assign n31889 = ~n1552 ;
  assign n1556 = n31889 & n1555 ;
  assign n1557 = n838 | n1532 ;
  assign n31890 = ~n1557 ;
  assign n1558 = n1547 & n31890 ;
  assign n1559 = n1556 | n1558 ;
  assign n31891 = ~n1549 ;
  assign n1560 = n31891 & n1559 ;
  assign n31892 = ~n1560 ;
  assign n1561 = n185 & n31892 ;
  assign n1562 = n31796 & n1347 ;
  assign n31893 = ~n1349 ;
  assign n1563 = n31893 & n1562 ;
  assign n1566 = n1487 & n1563 ;
  assign n1564 = n1341 | n1349 ;
  assign n31894 = ~n1564 ;
  assign n1565 = n1487 & n31894 ;
  assign n1567 = n1347 | n1565 ;
  assign n31895 = ~n1566 ;
  assign n1568 = n31895 & n1567 ;
  assign n1569 = n185 | n1549 ;
  assign n31896 = ~n1569 ;
  assign n1570 = n1559 & n31896 ;
  assign n1571 = n1568 | n1570 ;
  assign n31897 = ~n1561 ;
  assign n1572 = n31897 & n1571 ;
  assign n31898 = ~n1572 ;
  assign n1573 = n186 & n31898 ;
  assign n31899 = ~n1361 ;
  assign n1574 = n1359 & n31899 ;
  assign n1575 = n31802 & n1574 ;
  assign n1576 = n1487 & n1575 ;
  assign n1577 = n1352 | n1361 ;
  assign n31900 = ~n1577 ;
  assign n1578 = n180 & n31900 ;
  assign n1579 = n1359 | n1578 ;
  assign n31901 = ~n1576 ;
  assign n1580 = n31901 & n1579 ;
  assign n1581 = n183 & n31878 ;
  assign n1582 = n183 | n1506 ;
  assign n31902 = ~n1582 ;
  assign n1583 = n1535 & n31902 ;
  assign n1584 = n1541 | n1583 ;
  assign n31903 = ~n1581 ;
  assign n1585 = n31903 & n1584 ;
  assign n31904 = ~n1585 ;
  assign n1586 = n184 & n31904 ;
  assign n1587 = n31890 & n1584 ;
  assign n1588 = n1556 | n1587 ;
  assign n31905 = ~n1586 ;
  assign n1589 = n31905 & n1588 ;
  assign n31906 = ~n1589 ;
  assign n1590 = n185 & n31906 ;
  assign n1591 = n186 | n1590 ;
  assign n31907 = ~n1591 ;
  assign n1592 = n1571 & n31907 ;
  assign n1593 = n1580 | n1592 ;
  assign n31908 = ~n1573 ;
  assign n1594 = n31908 & n1593 ;
  assign n31909 = ~n1594 ;
  assign n1595 = n187 & n31909 ;
  assign n1596 = n31813 & n1371 ;
  assign n31910 = ~n1383 ;
  assign n1597 = n31910 & n1596 ;
  assign n1598 = n1487 & n1597 ;
  assign n1599 = n1364 | n1383 ;
  assign n31911 = ~n1599 ;
  assign n1600 = n180 & n31911 ;
  assign n1601 = n1371 | n1600 ;
  assign n31912 = ~n1598 ;
  assign n1602 = n31912 & n1601 ;
  assign n1603 = n528 | n1573 ;
  assign n31913 = ~n1603 ;
  assign n1604 = n1593 & n31913 ;
  assign n1605 = n1602 | n1604 ;
  assign n31914 = ~n1595 ;
  assign n1606 = n31914 & n1605 ;
  assign n31915 = ~n1606 ;
  assign n1607 = n413 & n31915 ;
  assign n31916 = ~n1395 ;
  assign n1608 = n1393 & n31916 ;
  assign n1609 = n31819 & n1608 ;
  assign n1610 = n1487 & n1609 ;
  assign n1611 = n1386 | n1395 ;
  assign n31917 = ~n1611 ;
  assign n1612 = n180 & n31917 ;
  assign n1613 = n1393 | n1612 ;
  assign n31918 = ~n1610 ;
  assign n1614 = n31918 & n1613 ;
  assign n1615 = n31896 & n1588 ;
  assign n1616 = n1568 | n1615 ;
  assign n31919 = ~n1590 ;
  assign n1617 = n31919 & n1616 ;
  assign n31920 = ~n1617 ;
  assign n1618 = n186 & n31920 ;
  assign n1619 = n31907 & n1616 ;
  assign n1620 = n1580 | n1619 ;
  assign n31921 = ~n1618 ;
  assign n1621 = n31921 & n1620 ;
  assign n31922 = ~n1621 ;
  assign n1622 = n528 & n31922 ;
  assign n1623 = n413 | n1622 ;
  assign n31923 = ~n1623 ;
  assign n1624 = n1605 & n31923 ;
  assign n1625 = n1614 | n1624 ;
  assign n31924 = ~n1607 ;
  assign n1626 = n31924 & n1625 ;
  assign n31925 = ~n1626 ;
  assign n1627 = n189 & n31925 ;
  assign n1628 = n31829 & n1405 ;
  assign n31926 = ~n1415 ;
  assign n1629 = n31926 & n1628 ;
  assign n1630 = n1487 & n1629 ;
  assign n1631 = n1398 | n1415 ;
  assign n31927 = ~n1631 ;
  assign n1632 = n180 & n31927 ;
  assign n1633 = n1405 | n1632 ;
  assign n31928 = ~n1630 ;
  assign n1634 = n31928 & n1633 ;
  assign n1635 = n189 | n1607 ;
  assign n31929 = ~n1635 ;
  assign n1636 = n1625 & n31929 ;
  assign n1637 = n1634 | n1636 ;
  assign n31930 = ~n1627 ;
  assign n1638 = n31930 & n1637 ;
  assign n31931 = ~n1638 ;
  assign n1639 = n190 & n31931 ;
  assign n31932 = ~n1427 ;
  assign n1640 = n1425 & n31932 ;
  assign n1641 = n31835 & n1640 ;
  assign n1642 = n180 & n1641 ;
  assign n1643 = n1418 | n1427 ;
  assign n31933 = ~n1643 ;
  assign n1644 = n180 & n31933 ;
  assign n1645 = n1425 | n1644 ;
  assign n31934 = ~n1642 ;
  assign n1646 = n31934 & n1645 ;
  assign n1647 = n31913 & n1620 ;
  assign n1648 = n1602 | n1647 ;
  assign n31935 = ~n1622 ;
  assign n1649 = n31935 & n1648 ;
  assign n31936 = ~n1649 ;
  assign n1650 = n188 & n31936 ;
  assign n1651 = n31923 & n1648 ;
  assign n1652 = n1614 | n1651 ;
  assign n31937 = ~n1650 ;
  assign n1653 = n31937 & n1652 ;
  assign n31938 = ~n1653 ;
  assign n1654 = n189 & n31938 ;
  assign n1655 = n190 | n1654 ;
  assign n31939 = ~n1655 ;
  assign n1656 = n1637 & n31939 ;
  assign n1657 = n1646 | n1656 ;
  assign n31940 = ~n1639 ;
  assign n1658 = n31940 & n1657 ;
  assign n31941 = ~n1658 ;
  assign n1659 = n191 & n31941 ;
  assign n1661 = n31845 & n1447 ;
  assign n31942 = ~n1440 ;
  assign n1662 = n31942 & n1661 ;
  assign n1663 = n1487 & n1662 ;
  assign n1664 = n1430 | n1440 ;
  assign n31943 = ~n1664 ;
  assign n1665 = n180 & n31943 ;
  assign n1666 = n1447 | n1665 ;
  assign n31944 = ~n1663 ;
  assign n1667 = n31944 & n1666 ;
  assign n1699 = n287 | n1639 ;
  assign n31945 = ~n1699 ;
  assign n1700 = n1657 & n31945 ;
  assign n1701 = n1667 | n1700 ;
  assign n31946 = ~n1659 ;
  assign n1702 = n31946 & n1701 ;
  assign n1703 = n1681 | n1702 ;
  assign n1704 = n31336 & n1703 ;
  assign n31947 = ~n1467 ;
  assign n1685 = n31947 & n1487 ;
  assign n31948 = ~n1685 ;
  assign n1686 = n1471 & n31948 ;
  assign n1687 = n192 & n1678 ;
  assign n31949 = ~n1686 ;
  assign n1688 = n31949 & n1687 ;
  assign n1689 = n1463 | n1483 ;
  assign n31950 = ~n1689 ;
  assign n1690 = n1466 & n31950 ;
  assign n1691 = n31873 & n1690 ;
  assign n1692 = n31874 & n1691 ;
  assign n1693 = n31875 & n1692 ;
  assign n1694 = n1688 | n1693 ;
  assign n1683 = n31946 & n1677 ;
  assign n1705 = n1683 & n1701 ;
  assign n1706 = n1694 | n1705 ;
  assign n1707 = n1704 | n1706 ;
  assign n31951 = ~n1707 ;
  assign n1708 = x100 & n31951 ;
  assign n1709 = x98 | x99 ;
  assign n31952 = ~x100 ;
  assign n1711 = n31952 & n1709 ;
  assign n1712 = n1708 | n1711 ;
  assign n31953 = ~n1712 ;
  assign n1723 = n1487 & n31953 ;
  assign n1713 = x100 & n1707 ;
  assign n1710 = x100 | n1709 ;
  assign n1714 = n31872 & n1710 ;
  assign n1715 = n31873 & n1714 ;
  assign n1716 = n31874 & n1715 ;
  assign n1717 = n31875 & n1716 ;
  assign n31954 = ~n1713 ;
  assign n1718 = n31954 & n1717 ;
  assign n1719 = n31952 & n1707 ;
  assign n31955 = ~n1719 ;
  assign n1720 = x101 & n31955 ;
  assign n31956 = ~n1489 ;
  assign n1721 = n31956 & n1707 ;
  assign n1722 = n1720 | n1721 ;
  assign n1724 = n1718 | n1722 ;
  assign n31957 = ~n1723 ;
  assign n1725 = n31957 & n1724 ;
  assign n31958 = ~n1725 ;
  assign n1726 = n181 & n31958 ;
  assign n1660 = n191 | n1639 ;
  assign n31959 = ~n1660 ;
  assign n1668 = n1657 & n31959 ;
  assign n1669 = n1667 | n1668 ;
  assign n1684 = n1669 & n1683 ;
  assign n1695 = n1684 | n1694 ;
  assign n1670 = n31946 & n1669 ;
  assign n1682 = n1670 | n1681 ;
  assign n1696 = n31336 & n1682 ;
  assign n179 = n1695 | n1696 ;
  assign n1698 = x100 & n179 ;
  assign n31960 = ~n1698 ;
  assign n1727 = n31960 & n1710 ;
  assign n31961 = ~n1727 ;
  assign n1728 = n180 & n31961 ;
  assign n1729 = n181 | n1728 ;
  assign n31962 = ~n1729 ;
  assign n1730 = n1724 & n31962 ;
  assign n31963 = ~n1693 ;
  assign n1731 = n1487 & n31963 ;
  assign n31964 = ~n1688 ;
  assign n1732 = n31964 & n1731 ;
  assign n31965 = ~n1705 ;
  assign n1733 = n31965 & n1732 ;
  assign n31966 = ~n1704 ;
  assign n1734 = n31966 & n1733 ;
  assign n1735 = n1721 | n1734 ;
  assign n1737 = x102 & n1735 ;
  assign n1736 = x102 | n1734 ;
  assign n1738 = n1721 | n1736 ;
  assign n31967 = ~n1737 ;
  assign n1739 = n31967 & n1738 ;
  assign n1740 = n1730 | n1739 ;
  assign n31968 = ~n1726 ;
  assign n1741 = n31968 & n1740 ;
  assign n31969 = ~n1741 ;
  assign n1742 = n182 & n31969 ;
  assign n1746 = n1493 | n1499 ;
  assign n31970 = ~n1746 ;
  assign n1748 = n1503 & n31970 ;
  assign n1749 = n1707 & n1748 ;
  assign n1747 = n179 & n31970 ;
  assign n1750 = n1503 | n1747 ;
  assign n31971 = ~n1749 ;
  assign n1751 = n31971 & n1750 ;
  assign n1743 = n181 | n1723 ;
  assign n31972 = ~n1743 ;
  assign n1744 = n1724 & n31972 ;
  assign n1745 = n1739 | n1744 ;
  assign n1753 = n182 | n1726 ;
  assign n31973 = ~n1753 ;
  assign n1754 = n1745 & n31973 ;
  assign n1755 = n1751 | n1754 ;
  assign n31974 = ~n1742 ;
  assign n1756 = n31974 & n1755 ;
  assign n31975 = ~n1756 ;
  assign n1757 = n996 & n31975 ;
  assign n31976 = ~n1534 ;
  assign n1758 = n1529 & n31976 ;
  assign n31977 = ~n1544 ;
  assign n1759 = n31977 & n1758 ;
  assign n1760 = n1707 & n1759 ;
  assign n1761 = n1534 | n1544 ;
  assign n31978 = ~n1761 ;
  assign n1762 = n179 & n31978 ;
  assign n1763 = n1529 | n1762 ;
  assign n31979 = ~n1760 ;
  assign n1764 = n31979 & n1763 ;
  assign n1765 = n996 | n1742 ;
  assign n31980 = ~n1765 ;
  assign n1766 = n1755 & n31980 ;
  assign n1767 = n1764 | n1766 ;
  assign n31981 = ~n1757 ;
  assign n1768 = n31981 & n1767 ;
  assign n31982 = ~n1768 ;
  assign n1769 = n184 & n31982 ;
  assign n1542 = n31885 & n1541 ;
  assign n31983 = ~n1546 ;
  assign n1770 = n1542 & n31983 ;
  assign n1771 = n1707 & n1770 ;
  assign n1772 = n1532 | n1546 ;
  assign n31984 = ~n1772 ;
  assign n1773 = n179 & n31984 ;
  assign n1774 = n1541 | n1773 ;
  assign n31985 = ~n1771 ;
  assign n1775 = n31985 & n1774 ;
  assign n1776 = n838 | n1757 ;
  assign n31986 = ~n1776 ;
  assign n1777 = n1767 & n31986 ;
  assign n1778 = n1775 | n1777 ;
  assign n31987 = ~n1769 ;
  assign n1779 = n31987 & n1778 ;
  assign n31988 = ~n1779 ;
  assign n1780 = n185 & n31988 ;
  assign n31989 = ~n1558 ;
  assign n1781 = n1556 & n31989 ;
  assign n1782 = n31891 & n1781 ;
  assign n1783 = n1707 & n1782 ;
  assign n1784 = n1549 | n1558 ;
  assign n31990 = ~n1784 ;
  assign n1785 = n179 & n31990 ;
  assign n1786 = n1556 | n1785 ;
  assign n31991 = ~n1783 ;
  assign n1787 = n31991 & n1786 ;
  assign n1788 = n183 & n31975 ;
  assign n31992 = ~n1788 ;
  assign n1789 = n1767 & n31992 ;
  assign n31993 = ~n1789 ;
  assign n1790 = n838 & n31993 ;
  assign n1791 = n185 | n1790 ;
  assign n31994 = ~n1791 ;
  assign n1792 = n1778 & n31994 ;
  assign n1793 = n1787 | n1792 ;
  assign n31995 = ~n1780 ;
  assign n1794 = n31995 & n1793 ;
  assign n31996 = ~n1794 ;
  assign n1795 = n186 & n31996 ;
  assign n1798 = n1568 & n31919 ;
  assign n31997 = ~n1570 ;
  assign n1799 = n31997 & n1798 ;
  assign n1800 = n1707 & n1799 ;
  assign n1796 = n1561 | n1570 ;
  assign n31998 = ~n1796 ;
  assign n1797 = n179 & n31998 ;
  assign n1801 = n1568 | n1797 ;
  assign n31999 = ~n1800 ;
  assign n1802 = n31999 & n1801 ;
  assign n1803 = n186 | n1780 ;
  assign n32000 = ~n1803 ;
  assign n1804 = n1793 & n32000 ;
  assign n1805 = n1802 | n1804 ;
  assign n32001 = ~n1795 ;
  assign n1806 = n32001 & n1805 ;
  assign n32002 = ~n1806 ;
  assign n1807 = n528 & n32002 ;
  assign n32003 = ~n1592 ;
  assign n1808 = n1580 & n32003 ;
  assign n1809 = n31908 & n1808 ;
  assign n1810 = n1707 & n1809 ;
  assign n1811 = n1573 | n1592 ;
  assign n32004 = ~n1811 ;
  assign n1812 = n179 & n32004 ;
  assign n1813 = n1580 | n1812 ;
  assign n32005 = ~n1810 ;
  assign n1814 = n32005 & n1813 ;
  assign n32006 = ~n1790 ;
  assign n1815 = n1778 & n32006 ;
  assign n32007 = ~n1815 ;
  assign n1816 = n185 & n32007 ;
  assign n32008 = ~n1816 ;
  assign n1817 = n1793 & n32008 ;
  assign n32009 = ~n1817 ;
  assign n1818 = n186 & n32009 ;
  assign n1819 = n528 | n1818 ;
  assign n32010 = ~n1819 ;
  assign n1820 = n1805 & n32010 ;
  assign n1821 = n1814 | n1820 ;
  assign n32011 = ~n1807 ;
  assign n1822 = n32011 & n1821 ;
  assign n32012 = ~n1822 ;
  assign n1823 = n188 & n32012 ;
  assign n1826 = n1602 & n31935 ;
  assign n32013 = ~n1604 ;
  assign n1827 = n32013 & n1826 ;
  assign n1828 = n1707 & n1827 ;
  assign n1824 = n1595 | n1604 ;
  assign n32014 = ~n1824 ;
  assign n1825 = n179 & n32014 ;
  assign n1829 = n1602 | n1825 ;
  assign n32015 = ~n1828 ;
  assign n1830 = n32015 & n1829 ;
  assign n1831 = n413 | n1807 ;
  assign n32016 = ~n1831 ;
  assign n1832 = n1821 & n32016 ;
  assign n1833 = n1830 | n1832 ;
  assign n32017 = ~n1823 ;
  assign n1834 = n32017 & n1833 ;
  assign n32018 = ~n1834 ;
  assign n1835 = n189 & n32018 ;
  assign n32019 = ~n1624 ;
  assign n1836 = n1614 & n32019 ;
  assign n1837 = n31924 & n1836 ;
  assign n1838 = n1707 & n1837 ;
  assign n1839 = n1607 | n1624 ;
  assign n32020 = ~n1839 ;
  assign n1840 = n179 & n32020 ;
  assign n1841 = n1614 | n1840 ;
  assign n32021 = ~n1838 ;
  assign n1842 = n32021 & n1841 ;
  assign n32022 = ~n1818 ;
  assign n1843 = n1805 & n32022 ;
  assign n32023 = ~n1843 ;
  assign n1844 = n187 & n32023 ;
  assign n32024 = ~n1844 ;
  assign n1845 = n1821 & n32024 ;
  assign n32025 = ~n1845 ;
  assign n1846 = n413 & n32025 ;
  assign n1847 = n189 | n1846 ;
  assign n32026 = ~n1847 ;
  assign n1848 = n1833 & n32026 ;
  assign n1849 = n1842 | n1848 ;
  assign n32027 = ~n1835 ;
  assign n1850 = n32027 & n1849 ;
  assign n32028 = ~n1850 ;
  assign n1851 = n190 & n32028 ;
  assign n32029 = ~n1654 ;
  assign n1852 = n1634 & n32029 ;
  assign n32030 = ~n1636 ;
  assign n1853 = n32030 & n1852 ;
  assign n1854 = n179 & n1853 ;
  assign n1855 = n1627 | n1636 ;
  assign n32031 = ~n1855 ;
  assign n1856 = n179 & n32031 ;
  assign n1857 = n1634 | n1856 ;
  assign n32032 = ~n1854 ;
  assign n1858 = n32032 & n1857 ;
  assign n1859 = n190 | n1835 ;
  assign n32033 = ~n1859 ;
  assign n1860 = n1849 & n32033 ;
  assign n1861 = n1858 | n1860 ;
  assign n32034 = ~n1851 ;
  assign n1862 = n32034 & n1861 ;
  assign n32035 = ~n1862 ;
  assign n1863 = n287 & n32035 ;
  assign n32036 = ~n1656 ;
  assign n1864 = n1646 & n32036 ;
  assign n1865 = n31940 & n1864 ;
  assign n1866 = n179 & n1865 ;
  assign n1867 = n1639 | n1656 ;
  assign n32037 = ~n1867 ;
  assign n1868 = n179 & n32037 ;
  assign n1869 = n1646 | n1868 ;
  assign n32038 = ~n1866 ;
  assign n1870 = n32038 & n1869 ;
  assign n32039 = ~n1846 ;
  assign n1871 = n1833 & n32039 ;
  assign n32040 = ~n1871 ;
  assign n1872 = n189 & n32040 ;
  assign n32041 = ~n1872 ;
  assign n1873 = n1849 & n32041 ;
  assign n32042 = ~n1873 ;
  assign n1874 = n190 & n32042 ;
  assign n1875 = n287 | n1874 ;
  assign n32043 = ~n1875 ;
  assign n1876 = n1861 & n32043 ;
  assign n1877 = n1870 | n1876 ;
  assign n32044 = ~n1863 ;
  assign n1878 = n32044 & n1877 ;
  assign n1879 = n31946 & n1667 ;
  assign n32045 = ~n1668 ;
  assign n1880 = n32045 & n1879 ;
  assign n1881 = n1707 & n1880 ;
  assign n1882 = n1659 | n1668 ;
  assign n32046 = ~n1882 ;
  assign n1883 = n179 & n32046 ;
  assign n1884 = n1667 | n1883 ;
  assign n32047 = ~n1881 ;
  assign n1885 = n32047 & n1884 ;
  assign n1887 = n1677 | n1702 ;
  assign n32048 = ~n1887 ;
  assign n1888 = n1707 & n32048 ;
  assign n1889 = n1705 | n1888 ;
  assign n1890 = n1885 | n1889 ;
  assign n1891 = n1878 | n1890 ;
  assign n1892 = n31336 & n1891 ;
  assign n1895 = n192 & n1887 ;
  assign n32049 = ~n1677 ;
  assign n1894 = n32049 & n1707 ;
  assign n32050 = ~n1894 ;
  assign n1896 = n1702 & n32050 ;
  assign n32051 = ~n1896 ;
  assign n1897 = n1895 & n32051 ;
  assign n1898 = n1673 | n1693 ;
  assign n32052 = ~n1898 ;
  assign n1899 = n1676 & n32052 ;
  assign n1900 = n31964 & n1899 ;
  assign n1901 = n31965 & n1900 ;
  assign n1902 = n31966 & n1901 ;
  assign n1903 = n1897 | n1902 ;
  assign n1893 = n32044 & n1885 ;
  assign n1904 = n1877 & n1893 ;
  assign n1905 = n1903 | n1904 ;
  assign n178 = n1892 | n1905 ;
  assign n1909 = x98 & n178 ;
  assign n1910 = x96 | x97 ;
  assign n1911 = x98 | n1910 ;
  assign n32053 = ~n1909 ;
  assign n1912 = n32053 & n1911 ;
  assign n32054 = ~n1912 ;
  assign n1913 = n179 & n32054 ;
  assign n1914 = n31963 & n1911 ;
  assign n1915 = n31964 & n1914 ;
  assign n1916 = n31965 & n1915 ;
  assign n1917 = n31966 & n1916 ;
  assign n1918 = n32053 & n1917 ;
  assign n32055 = ~n1709 ;
  assign n1908 = n32055 & n178 ;
  assign n32056 = ~x98 ;
  assign n1919 = n32056 & n178 ;
  assign n32057 = ~n1919 ;
  assign n1920 = x99 & n32057 ;
  assign n1921 = n1908 | n1920 ;
  assign n1922 = n1918 | n1921 ;
  assign n32058 = ~n1913 ;
  assign n1923 = n32058 & n1922 ;
  assign n32059 = ~n1923 ;
  assign n1924 = n1487 & n32059 ;
  assign n32060 = ~n1902 ;
  assign n1929 = n1707 & n32060 ;
  assign n32061 = ~n1897 ;
  assign n1930 = n32061 & n1929 ;
  assign n32062 = ~n1904 ;
  assign n1931 = n32062 & n1930 ;
  assign n32063 = ~n1892 ;
  assign n1932 = n32063 & n1931 ;
  assign n1933 = n1908 | n1932 ;
  assign n1935 = x100 & n1933 ;
  assign n1934 = x100 | n1932 ;
  assign n1936 = n1908 | n1934 ;
  assign n32064 = ~n1935 ;
  assign n1937 = n32064 & n1936 ;
  assign n32065 = ~n178 ;
  assign n1907 = x98 & n32065 ;
  assign n1925 = n32056 & n1910 ;
  assign n1926 = n1907 | n1925 ;
  assign n32066 = ~n1926 ;
  assign n1927 = n1707 & n32066 ;
  assign n1928 = n1487 | n1927 ;
  assign n32067 = ~n1928 ;
  assign n1938 = n1922 & n32067 ;
  assign n1939 = n1937 | n1938 ;
  assign n32068 = ~n1924 ;
  assign n1940 = n32068 & n1939 ;
  assign n32069 = ~n1940 ;
  assign n1941 = n181 & n32069 ;
  assign n1942 = n1718 | n1723 ;
  assign n32070 = ~n1942 ;
  assign n1943 = n1722 & n32070 ;
  assign n1944 = n178 & n1943 ;
  assign n1945 = n178 & n32070 ;
  assign n1946 = n1722 | n1945 ;
  assign n32071 = ~n1944 ;
  assign n1947 = n32071 & n1946 ;
  assign n1948 = n181 | n1924 ;
  assign n32072 = ~n1948 ;
  assign n1949 = n1939 & n32072 ;
  assign n1950 = n1947 | n1949 ;
  assign n32073 = ~n1941 ;
  assign n1951 = n32073 & n1950 ;
  assign n32074 = ~n1951 ;
  assign n1952 = n182 & n32074 ;
  assign n32075 = ~n1744 ;
  assign n1953 = n1739 & n32075 ;
  assign n1954 = n31968 & n1953 ;
  assign n1955 = n178 & n1954 ;
  assign n1956 = n1726 | n1744 ;
  assign n32076 = ~n1956 ;
  assign n1957 = n178 & n32076 ;
  assign n1958 = n1739 | n1957 ;
  assign n32077 = ~n1955 ;
  assign n1959 = n32077 & n1958 ;
  assign n1960 = n182 | n1941 ;
  assign n32078 = ~n1960 ;
  assign n1961 = n1950 & n32078 ;
  assign n1962 = n1959 | n1961 ;
  assign n32079 = ~n1952 ;
  assign n1963 = n32079 & n1962 ;
  assign n32080 = ~n1963 ;
  assign n1964 = n996 & n32080 ;
  assign n1752 = n31974 & n1751 ;
  assign n32081 = ~n1754 ;
  assign n1965 = n1752 & n32081 ;
  assign n1968 = n178 & n1965 ;
  assign n1966 = n1742 | n1754 ;
  assign n32082 = ~n1966 ;
  assign n1967 = n178 & n32082 ;
  assign n1969 = n1751 | n1967 ;
  assign n32083 = ~n1968 ;
  assign n1970 = n32083 & n1969 ;
  assign n1971 = n180 & n32059 ;
  assign n1972 = n180 | n1913 ;
  assign n32084 = ~n1972 ;
  assign n1973 = n1922 & n32084 ;
  assign n1974 = n1937 | n1973 ;
  assign n32085 = ~n1971 ;
  assign n1975 = n32085 & n1974 ;
  assign n32086 = ~n1975 ;
  assign n1976 = n181 & n32086 ;
  assign n1977 = n32072 & n1974 ;
  assign n1978 = n1947 | n1977 ;
  assign n32087 = ~n1976 ;
  assign n1979 = n32087 & n1978 ;
  assign n32088 = ~n1979 ;
  assign n1980 = n182 & n32088 ;
  assign n1981 = n183 | n1980 ;
  assign n32089 = ~n1981 ;
  assign n1982 = n1962 & n32089 ;
  assign n1983 = n1970 | n1982 ;
  assign n32090 = ~n1964 ;
  assign n1984 = n32090 & n1983 ;
  assign n32091 = ~n1984 ;
  assign n1985 = n184 & n32091 ;
  assign n32092 = ~n1766 ;
  assign n1986 = n1764 & n32092 ;
  assign n1987 = n31981 & n1986 ;
  assign n1988 = n178 & n1987 ;
  assign n1989 = n1757 | n1766 ;
  assign n32093 = ~n1989 ;
  assign n1990 = n178 & n32093 ;
  assign n1991 = n1764 | n1990 ;
  assign n32094 = ~n1988 ;
  assign n1992 = n32094 & n1991 ;
  assign n1993 = n838 | n1964 ;
  assign n32095 = ~n1993 ;
  assign n1994 = n1983 & n32095 ;
  assign n1995 = n1992 | n1994 ;
  assign n32096 = ~n1985 ;
  assign n1996 = n32096 & n1995 ;
  assign n32097 = ~n1996 ;
  assign n1997 = n185 & n32097 ;
  assign n1998 = n1775 & n32006 ;
  assign n32098 = ~n1777 ;
  assign n1999 = n32098 & n1998 ;
  assign n2000 = n178 & n1999 ;
  assign n2001 = n1769 | n1777 ;
  assign n32099 = ~n2001 ;
  assign n2002 = n178 & n32099 ;
  assign n2003 = n1775 | n2002 ;
  assign n32100 = ~n2000 ;
  assign n2004 = n32100 & n2003 ;
  assign n2005 = n32078 & n1978 ;
  assign n2006 = n1959 | n2005 ;
  assign n32101 = ~n1980 ;
  assign n2007 = n32101 & n2006 ;
  assign n32102 = ~n2007 ;
  assign n2008 = n183 & n32102 ;
  assign n2009 = n32089 & n2006 ;
  assign n2010 = n1970 | n2009 ;
  assign n32103 = ~n2008 ;
  assign n2011 = n32103 & n2010 ;
  assign n32104 = ~n2011 ;
  assign n2012 = n838 & n32104 ;
  assign n2013 = n185 | n2012 ;
  assign n32105 = ~n2013 ;
  assign n2014 = n1995 & n32105 ;
  assign n2015 = n2004 | n2014 ;
  assign n32106 = ~n1997 ;
  assign n2016 = n32106 & n2015 ;
  assign n32107 = ~n2016 ;
  assign n2017 = n186 & n32107 ;
  assign n32108 = ~n1792 ;
  assign n2018 = n1787 & n32108 ;
  assign n2019 = n31995 & n2018 ;
  assign n2020 = n178 & n2019 ;
  assign n2021 = n1780 | n1792 ;
  assign n32109 = ~n2021 ;
  assign n2022 = n178 & n32109 ;
  assign n2023 = n1787 | n2022 ;
  assign n32110 = ~n2020 ;
  assign n2024 = n32110 & n2023 ;
  assign n2025 = n186 | n1997 ;
  assign n32111 = ~n2025 ;
  assign n2026 = n2015 & n32111 ;
  assign n2027 = n2024 | n2026 ;
  assign n32112 = ~n2017 ;
  assign n2028 = n32112 & n2027 ;
  assign n32113 = ~n2028 ;
  assign n2029 = n528 & n32113 ;
  assign n2030 = n1802 & n32022 ;
  assign n32114 = ~n1804 ;
  assign n2031 = n32114 & n2030 ;
  assign n2032 = n178 & n2031 ;
  assign n2033 = n1795 | n1804 ;
  assign n32115 = ~n2033 ;
  assign n2034 = n178 & n32115 ;
  assign n2035 = n1802 | n2034 ;
  assign n32116 = ~n2032 ;
  assign n2036 = n32116 & n2035 ;
  assign n2037 = n32095 & n2010 ;
  assign n2038 = n1992 | n2037 ;
  assign n32117 = ~n2012 ;
  assign n2039 = n32117 & n2038 ;
  assign n32118 = ~n2039 ;
  assign n2040 = n185 & n32118 ;
  assign n2041 = n32105 & n2038 ;
  assign n2042 = n2004 | n2041 ;
  assign n32119 = ~n2040 ;
  assign n2043 = n32119 & n2042 ;
  assign n32120 = ~n2043 ;
  assign n2044 = n186 & n32120 ;
  assign n2045 = n528 | n2044 ;
  assign n32121 = ~n2045 ;
  assign n2046 = n2027 & n32121 ;
  assign n2048 = n2036 | n2046 ;
  assign n32122 = ~n2029 ;
  assign n2049 = n32122 & n2048 ;
  assign n32123 = ~n2049 ;
  assign n2050 = n188 & n32123 ;
  assign n32124 = ~n1820 ;
  assign n2051 = n1814 & n32124 ;
  assign n2052 = n32011 & n2051 ;
  assign n2053 = n178 & n2052 ;
  assign n2054 = n1807 | n1820 ;
  assign n32125 = ~n2054 ;
  assign n2055 = n178 & n32125 ;
  assign n2056 = n1814 | n2055 ;
  assign n32126 = ~n2053 ;
  assign n2057 = n32126 & n2056 ;
  assign n2058 = n413 | n2029 ;
  assign n32127 = ~n2058 ;
  assign n2059 = n2048 & n32127 ;
  assign n2062 = n2057 | n2059 ;
  assign n32128 = ~n2050 ;
  assign n2063 = n32128 & n2062 ;
  assign n32129 = ~n2063 ;
  assign n2064 = n189 & n32129 ;
  assign n2067 = n1830 & n32039 ;
  assign n32130 = ~n1832 ;
  assign n2068 = n32130 & n2067 ;
  assign n2069 = n178 & n2068 ;
  assign n2065 = n1823 | n1832 ;
  assign n32131 = ~n2065 ;
  assign n2066 = n178 & n32131 ;
  assign n2070 = n1830 | n2066 ;
  assign n32132 = ~n2069 ;
  assign n2071 = n32132 & n2070 ;
  assign n2073 = n32111 & n2042 ;
  assign n2074 = n2024 | n2073 ;
  assign n32133 = ~n2044 ;
  assign n2075 = n32133 & n2074 ;
  assign n32134 = ~n2075 ;
  assign n2076 = n187 & n32134 ;
  assign n2077 = n32121 & n2074 ;
  assign n2078 = n2036 | n2077 ;
  assign n32135 = ~n2076 ;
  assign n2079 = n32135 & n2078 ;
  assign n32136 = ~n2079 ;
  assign n2080 = n413 & n32136 ;
  assign n2082 = n189 | n2080 ;
  assign n32137 = ~n2082 ;
  assign n2083 = n2062 & n32137 ;
  assign n2086 = n2071 | n2083 ;
  assign n32138 = ~n2064 ;
  assign n2087 = n32138 & n2086 ;
  assign n32139 = ~n2087 ;
  assign n2088 = n190 & n32139 ;
  assign n32140 = ~n1848 ;
  assign n2089 = n1842 & n32140 ;
  assign n2090 = n32027 & n2089 ;
  assign n2091 = n178 & n2090 ;
  assign n2092 = n1835 | n1848 ;
  assign n32141 = ~n2092 ;
  assign n2093 = n178 & n32141 ;
  assign n2094 = n1842 | n2093 ;
  assign n32142 = ~n2091 ;
  assign n2095 = n32142 & n2094 ;
  assign n2096 = n190 | n2064 ;
  assign n32143 = ~n2096 ;
  assign n2097 = n2086 & n32143 ;
  assign n2100 = n2095 | n2097 ;
  assign n32144 = ~n2088 ;
  assign n2101 = n32144 & n2100 ;
  assign n32145 = ~n2101 ;
  assign n2102 = n287 & n32145 ;
  assign n32146 = ~n1874 ;
  assign n2103 = n1858 & n32146 ;
  assign n32147 = ~n1860 ;
  assign n2104 = n32147 & n2103 ;
  assign n2105 = n178 & n2104 ;
  assign n2106 = n1851 | n1860 ;
  assign n32148 = ~n2106 ;
  assign n2107 = n178 & n32148 ;
  assign n2108 = n1858 | n2107 ;
  assign n32149 = ~n2105 ;
  assign n2109 = n32149 & n2108 ;
  assign n2111 = n32127 & n2078 ;
  assign n2112 = n2057 | n2111 ;
  assign n32150 = ~n2080 ;
  assign n2113 = n32150 & n2112 ;
  assign n32151 = ~n2113 ;
  assign n2114 = n189 & n32151 ;
  assign n2115 = n32137 & n2112 ;
  assign n2116 = n2071 | n2115 ;
  assign n32152 = ~n2114 ;
  assign n2117 = n32152 & n2116 ;
  assign n32153 = ~n2117 ;
  assign n2118 = n190 & n32153 ;
  assign n2120 = n287 | n2118 ;
  assign n32154 = ~n2120 ;
  assign n2121 = n2100 & n32154 ;
  assign n2124 = n2109 | n2121 ;
  assign n32155 = ~n2102 ;
  assign n2125 = n32155 & n2124 ;
  assign n32156 = ~n1876 ;
  assign n2126 = n1870 & n32156 ;
  assign n2127 = n32044 & n2126 ;
  assign n2128 = n178 & n2127 ;
  assign n2129 = n1863 | n1876 ;
  assign n32157 = ~n2129 ;
  assign n2130 = n178 & n32157 ;
  assign n2131 = n1870 | n2130 ;
  assign n32158 = ~n2128 ;
  assign n2132 = n32158 & n2131 ;
  assign n1886 = n1878 | n1885 ;
  assign n32159 = ~n1886 ;
  assign n2135 = n32159 & n178 ;
  assign n2136 = n1904 | n2135 ;
  assign n2137 = n2132 | n2136 ;
  assign n2138 = n2125 | n2137 ;
  assign n2139 = n31336 & n2138 ;
  assign n2140 = n32155 & n2132 ;
  assign n2141 = n2124 & n2140 ;
  assign n2143 = n192 & n1886 ;
  assign n32160 = ~n1885 ;
  assign n2142 = n32160 & n178 ;
  assign n32161 = ~n2142 ;
  assign n2144 = n1878 & n32161 ;
  assign n32162 = ~n2144 ;
  assign n2145 = n2143 & n32162 ;
  assign n2146 = n1881 | n1902 ;
  assign n32163 = ~n2146 ;
  assign n2147 = n1884 & n32163 ;
  assign n2148 = n32061 & n2147 ;
  assign n2149 = n32062 & n2148 ;
  assign n2150 = n32063 & n2149 ;
  assign n2161 = n2145 | n2150 ;
  assign n2162 = n2141 | n2161 ;
  assign n177 = n2139 | n2162 ;
  assign n2110 = n32155 & n2109 ;
  assign n32164 = ~n2121 ;
  assign n2122 = n2110 & n32164 ;
  assign n2164 = n2122 & n177 ;
  assign n2123 = n2102 | n2121 ;
  assign n32165 = ~n2123 ;
  assign n2166 = n32165 & n177 ;
  assign n2167 = n2109 | n2166 ;
  assign n32166 = ~n2164 ;
  assign n2168 = n32166 & n2167 ;
  assign n2133 = n2125 | n2132 ;
  assign n32167 = ~n2133 ;
  assign n2201 = n32167 & n177 ;
  assign n2202 = n2141 | n2201 ;
  assign n2203 = n2168 | n2202 ;
  assign n2185 = x96 & n177 ;
  assign n2187 = x94 | x95 ;
  assign n2188 = x96 | n2187 ;
  assign n32168 = ~n2185 ;
  assign n2189 = n32168 & n2188 ;
  assign n32169 = ~n2189 ;
  assign n2190 = n178 & n32169 ;
  assign n32170 = ~n1910 ;
  assign n2186 = n32170 & n177 ;
  assign n32171 = ~x96 ;
  assign n2191 = n32171 & n177 ;
  assign n32172 = ~n2191 ;
  assign n2192 = x97 & n32172 ;
  assign n2193 = n2186 | n2192 ;
  assign n2205 = n32060 & n2188 ;
  assign n2206 = n32061 & n2205 ;
  assign n2207 = n32062 & n2206 ;
  assign n2208 = n32063 & n2207 ;
  assign n2209 = n32168 & n2208 ;
  assign n2211 = n2193 | n2209 ;
  assign n32173 = ~n2190 ;
  assign n2212 = n32173 & n2211 ;
  assign n32174 = ~n2212 ;
  assign n2213 = n1707 & n32174 ;
  assign n32175 = ~n177 ;
  assign n2204 = x96 & n32175 ;
  assign n2214 = n32171 & n2187 ;
  assign n2215 = n2204 | n2214 ;
  assign n32176 = ~n2215 ;
  assign n2216 = n178 & n32176 ;
  assign n2219 = n1707 | n2216 ;
  assign n32177 = ~n2219 ;
  assign n2220 = n2211 & n32177 ;
  assign n32178 = ~n2150 ;
  assign n2222 = n178 & n32178 ;
  assign n32179 = ~n2145 ;
  assign n2223 = n32179 & n2222 ;
  assign n32180 = ~n2141 ;
  assign n2224 = n32180 & n2223 ;
  assign n32181 = ~n2139 ;
  assign n2225 = n32181 & n2224 ;
  assign n2226 = n2186 | n2225 ;
  assign n2228 = x98 & n2226 ;
  assign n2227 = x98 | n2225 ;
  assign n2229 = n2186 | n2227 ;
  assign n32182 = ~n2228 ;
  assign n2230 = n32182 & n2229 ;
  assign n2233 = n2220 | n2230 ;
  assign n32183 = ~n2213 ;
  assign n2234 = n32183 & n2233 ;
  assign n32184 = ~n2234 ;
  assign n2235 = n1487 & n32184 ;
  assign n2236 = n1918 | n1927 ;
  assign n32185 = ~n2236 ;
  assign n2237 = n1921 & n32185 ;
  assign n2238 = n177 & n2237 ;
  assign n2239 = n177 & n32185 ;
  assign n2240 = n1921 | n2239 ;
  assign n32186 = ~n2238 ;
  assign n2241 = n32186 & n2240 ;
  assign n2243 = n1487 | n2213 ;
  assign n32187 = ~n2243 ;
  assign n2244 = n2233 & n32187 ;
  assign n2247 = n2241 | n2244 ;
  assign n32188 = ~n2235 ;
  assign n2248 = n32188 & n2247 ;
  assign n32189 = ~n2248 ;
  assign n2249 = n181 & n32189 ;
  assign n32190 = ~n1938 ;
  assign n2250 = n1937 & n32190 ;
  assign n2252 = n32068 & n2250 ;
  assign n2253 = n177 & n2252 ;
  assign n2251 = n1924 | n1938 ;
  assign n32191 = ~n2251 ;
  assign n2254 = n177 & n32191 ;
  assign n2255 = n1937 | n2254 ;
  assign n32192 = ~n2253 ;
  assign n2256 = n32192 & n2255 ;
  assign n2257 = n181 | n2235 ;
  assign n32193 = ~n2257 ;
  assign n2258 = n2247 & n32193 ;
  assign n2262 = n2256 | n2258 ;
  assign n32194 = ~n2249 ;
  assign n2263 = n32194 & n2262 ;
  assign n32195 = ~n2263 ;
  assign n2264 = n182 & n32195 ;
  assign n2265 = n32073 & n1947 ;
  assign n32196 = ~n1949 ;
  assign n2266 = n32196 & n2265 ;
  assign n2269 = n177 & n2266 ;
  assign n2267 = n1941 | n1949 ;
  assign n32197 = ~n2267 ;
  assign n2268 = n177 & n32197 ;
  assign n2270 = n1947 | n2268 ;
  assign n32198 = ~n2269 ;
  assign n2271 = n32198 & n2270 ;
  assign n2273 = n179 & n32174 ;
  assign n2274 = n179 | n2190 ;
  assign n32199 = ~n2274 ;
  assign n2275 = n2211 & n32199 ;
  assign n2276 = n2230 | n2275 ;
  assign n32200 = ~n2273 ;
  assign n2277 = n32200 & n2276 ;
  assign n32201 = ~n2277 ;
  assign n2278 = n180 & n32201 ;
  assign n2279 = n32187 & n2276 ;
  assign n2280 = n2241 | n2279 ;
  assign n32202 = ~n2278 ;
  assign n2281 = n32202 & n2280 ;
  assign n32203 = ~n2281 ;
  assign n2282 = n181 & n32203 ;
  assign n2283 = n182 | n2282 ;
  assign n32204 = ~n2283 ;
  assign n2284 = n2262 & n32204 ;
  assign n2287 = n2271 | n2284 ;
  assign n32205 = ~n2264 ;
  assign n2288 = n32205 & n2287 ;
  assign n32206 = ~n2288 ;
  assign n2289 = n183 & n32206 ;
  assign n32207 = ~n1961 ;
  assign n2290 = n1959 & n32207 ;
  assign n2291 = n32079 & n2290 ;
  assign n2292 = n177 & n2291 ;
  assign n2293 = n1961 | n1980 ;
  assign n32208 = ~n2293 ;
  assign n2294 = n177 & n32208 ;
  assign n2295 = n1959 | n2294 ;
  assign n32209 = ~n2292 ;
  assign n2296 = n32209 & n2295 ;
  assign n2297 = n183 | n2264 ;
  assign n32210 = ~n2297 ;
  assign n2298 = n2287 & n32210 ;
  assign n2302 = n2296 | n2298 ;
  assign n32211 = ~n2289 ;
  assign n2303 = n32211 & n2302 ;
  assign n32212 = ~n2303 ;
  assign n2304 = n838 & n32212 ;
  assign n2306 = n32090 & n1970 ;
  assign n32213 = ~n1982 ;
  assign n2307 = n32213 & n2306 ;
  assign n2308 = n177 & n2307 ;
  assign n2309 = n1964 | n1982 ;
  assign n32214 = ~n2309 ;
  assign n2310 = n177 & n32214 ;
  assign n2311 = n1970 | n2310 ;
  assign n32215 = ~n2308 ;
  assign n2312 = n32215 & n2311 ;
  assign n2314 = n32193 & n2280 ;
  assign n2315 = n2256 | n2314 ;
  assign n32216 = ~n2282 ;
  assign n2316 = n32216 & n2315 ;
  assign n32217 = ~n2316 ;
  assign n2317 = n182 & n32217 ;
  assign n2318 = n32204 & n2315 ;
  assign n2319 = n2271 | n2318 ;
  assign n32218 = ~n2317 ;
  assign n2320 = n32218 & n2319 ;
  assign n32219 = ~n2320 ;
  assign n2321 = n996 & n32219 ;
  assign n2322 = n838 | n2321 ;
  assign n32220 = ~n2322 ;
  assign n2323 = n2302 & n32220 ;
  assign n2326 = n2312 | n2323 ;
  assign n32221 = ~n2304 ;
  assign n2328 = n32221 & n2326 ;
  assign n32222 = ~n2328 ;
  assign n2329 = n185 & n32222 ;
  assign n2305 = n185 | n2304 ;
  assign n32223 = ~n2305 ;
  assign n2327 = n32223 & n2326 ;
  assign n32224 = ~n1994 ;
  assign n2331 = n1992 & n32224 ;
  assign n2332 = n32096 & n2331 ;
  assign n2333 = n177 & n2332 ;
  assign n2334 = n1994 | n2012 ;
  assign n32225 = ~n2334 ;
  assign n2335 = n177 & n32225 ;
  assign n2336 = n1992 | n2335 ;
  assign n32226 = ~n2333 ;
  assign n2337 = n32226 & n2336 ;
  assign n2340 = n2327 | n2337 ;
  assign n32227 = ~n2329 ;
  assign n2341 = n32227 & n2340 ;
  assign n32228 = ~n2341 ;
  assign n2342 = n186 & n32228 ;
  assign n2344 = n32106 & n2004 ;
  assign n32229 = ~n2014 ;
  assign n2345 = n32229 & n2344 ;
  assign n2346 = n177 & n2345 ;
  assign n2347 = n1997 | n2014 ;
  assign n32230 = ~n2347 ;
  assign n2348 = n177 & n32230 ;
  assign n2349 = n2004 | n2348 ;
  assign n32231 = ~n2346 ;
  assign n2350 = n32231 & n2349 ;
  assign n2352 = n32210 & n2319 ;
  assign n2353 = n2296 | n2352 ;
  assign n32232 = ~n2321 ;
  assign n2354 = n32232 & n2353 ;
  assign n32233 = ~n2354 ;
  assign n2355 = n184 & n32233 ;
  assign n2356 = n32220 & n2353 ;
  assign n2357 = n2312 | n2356 ;
  assign n32234 = ~n2355 ;
  assign n2360 = n32234 & n2357 ;
  assign n32235 = ~n2360 ;
  assign n2361 = n185 & n32235 ;
  assign n2364 = n186 | n2361 ;
  assign n32236 = ~n2364 ;
  assign n2371 = n2340 & n32236 ;
  assign n2374 = n2350 | n2371 ;
  assign n32237 = ~n2342 ;
  assign n2375 = n32237 & n2374 ;
  assign n32238 = ~n2375 ;
  assign n2376 = n187 & n32238 ;
  assign n32239 = ~n2026 ;
  assign n2377 = n2024 & n32239 ;
  assign n2378 = n32112 & n2377 ;
  assign n2379 = n177 & n2378 ;
  assign n2380 = n2026 | n2044 ;
  assign n32240 = ~n2380 ;
  assign n2381 = n177 & n32240 ;
  assign n2382 = n2024 | n2381 ;
  assign n32241 = ~n2379 ;
  assign n2383 = n32241 & n2382 ;
  assign n2343 = n528 | n2342 ;
  assign n32242 = ~n2343 ;
  assign n2388 = n32242 & n2374 ;
  assign n2392 = n2383 | n2388 ;
  assign n32243 = ~n2376 ;
  assign n2394 = n32243 & n2392 ;
  assign n32244 = ~n2394 ;
  assign n2395 = n413 & n32244 ;
  assign n2358 = n32223 & n2357 ;
  assign n2359 = n2337 | n2358 ;
  assign n32245 = ~n2361 ;
  assign n2362 = n2359 & n32245 ;
  assign n32246 = ~n2362 ;
  assign n2363 = n186 & n32246 ;
  assign n2365 = n2359 & n32236 ;
  assign n2366 = n2350 | n2365 ;
  assign n32247 = ~n2363 ;
  assign n2367 = n32247 & n2366 ;
  assign n32248 = ~n2367 ;
  assign n2368 = n528 & n32248 ;
  assign n2369 = n413 | n2368 ;
  assign n32249 = ~n2369 ;
  assign n2393 = n32249 & n2392 ;
  assign n2047 = n2029 | n2046 ;
  assign n32250 = ~n2047 ;
  assign n2181 = n32250 & n177 ;
  assign n2182 = n2036 | n2181 ;
  assign n2398 = n32122 & n2036 ;
  assign n32251 = ~n2046 ;
  assign n2399 = n32251 & n2398 ;
  assign n2400 = n177 & n2399 ;
  assign n32252 = ~n2400 ;
  assign n2401 = n2182 & n32252 ;
  assign n2402 = n2393 | n2401 ;
  assign n32253 = ~n2395 ;
  assign n2403 = n32253 & n2402 ;
  assign n32254 = ~n2403 ;
  assign n2404 = n189 & n32254 ;
  assign n2081 = n2059 | n2080 ;
  assign n32255 = ~n2081 ;
  assign n2177 = n32255 & n177 ;
  assign n2178 = n2057 | n2177 ;
  assign n32256 = ~n2059 ;
  assign n2060 = n2057 & n32256 ;
  assign n2061 = n32128 & n2060 ;
  assign n2179 = n2061 & n177 ;
  assign n32257 = ~n2179 ;
  assign n2180 = n2178 & n32257 ;
  assign n2396 = n189 | n2395 ;
  assign n32258 = ~n2396 ;
  assign n2405 = n32258 & n2402 ;
  assign n2406 = n2180 | n2405 ;
  assign n32259 = ~n2404 ;
  assign n2407 = n32259 & n2406 ;
  assign n32260 = ~n2407 ;
  assign n2408 = n190 & n32260 ;
  assign n2085 = n2064 | n2083 ;
  assign n32261 = ~n2085 ;
  assign n2175 = n32261 & n177 ;
  assign n2176 = n2071 | n2175 ;
  assign n2072 = n32138 & n2071 ;
  assign n32262 = ~n2083 ;
  assign n2084 = n2072 & n32262 ;
  assign n2183 = n2084 & n177 ;
  assign n32263 = ~n2183 ;
  assign n2184 = n2176 & n32263 ;
  assign n2370 = n32242 & n2366 ;
  assign n2384 = n2370 | n2383 ;
  assign n32264 = ~n2368 ;
  assign n2385 = n32264 & n2384 ;
  assign n32265 = ~n2385 ;
  assign n2386 = n188 & n32265 ;
  assign n2387 = n32249 & n2384 ;
  assign n2413 = n2387 | n2401 ;
  assign n32266 = ~n2386 ;
  assign n2414 = n32266 & n2413 ;
  assign n32267 = ~n2414 ;
  assign n2415 = n189 & n32267 ;
  assign n2416 = n190 | n2415 ;
  assign n32268 = ~n2416 ;
  assign n2417 = n2406 & n32268 ;
  assign n2418 = n2184 | n2417 ;
  assign n32269 = ~n2408 ;
  assign n2423 = n32269 & n2418 ;
  assign n32270 = ~n2423 ;
  assign n2424 = n191 & n32270 ;
  assign n32271 = ~n2097 ;
  assign n2098 = n2095 & n32271 ;
  assign n2099 = n32144 & n2098 ;
  assign n2170 = n2099 & n177 ;
  assign n2119 = n2097 | n2118 ;
  assign n32272 = ~n2119 ;
  assign n2171 = n32272 & n177 ;
  assign n2172 = n2095 | n2171 ;
  assign n32273 = ~n2170 ;
  assign n2173 = n32273 & n2172 ;
  assign n2410 = n191 | n2408 ;
  assign n32274 = ~n2410 ;
  assign n2487 = n32274 & n2418 ;
  assign n2488 = n2173 | n2487 ;
  assign n32275 = ~n2424 ;
  assign n2489 = n32275 & n2488 ;
  assign n2490 = n2203 | n2489 ;
  assign n2491 = n31336 & n2490 ;
  assign n2151 = n2128 | n2150 ;
  assign n32276 = ~n2151 ;
  assign n2152 = n2131 & n32276 ;
  assign n2153 = n32179 & n2152 ;
  assign n2154 = n32180 & n2153 ;
  assign n2155 = n32181 & n2154 ;
  assign n2134 = n192 & n2133 ;
  assign n32277 = ~n2132 ;
  assign n2194 = n32277 & n177 ;
  assign n32278 = ~n2194 ;
  assign n2195 = n2125 & n32278 ;
  assign n32279 = ~n2195 ;
  assign n2196 = n2134 & n32279 ;
  assign n2197 = n2155 | n2196 ;
  assign n2428 = n2168 & n32275 ;
  assign n2492 = n2428 & n2488 ;
  assign n2493 = n2197 | n2492 ;
  assign n176 = n2491 | n2493 ;
  assign n2409 = n287 | n2408 ;
  assign n32280 = ~n2409 ;
  assign n2419 = n32280 & n2418 ;
  assign n2420 = n2173 | n2419 ;
  assign n2425 = n2420 & n32275 ;
  assign n2426 = n2203 | n2425 ;
  assign n2427 = n31336 & n2426 ;
  assign n2165 = n2155 | n2164 ;
  assign n32281 = ~n2165 ;
  assign n2169 = n32281 & n2167 ;
  assign n32282 = ~n2196 ;
  assign n2199 = n2169 & n32282 ;
  assign n2429 = n2420 & n2428 ;
  assign n32283 = ~n2429 ;
  assign n2474 = n2199 & n32283 ;
  assign n32284 = ~n2427 ;
  assign n2475 = n32284 & n2474 ;
  assign n2430 = n2197 | n2429 ;
  assign n2431 = n2427 | n2430 ;
  assign n32285 = ~n2168 ;
  assign n2435 = n32285 & n2431 ;
  assign n32286 = ~n2435 ;
  assign n2478 = n2425 & n32286 ;
  assign n2479 = n2168 | n2425 ;
  assign n2482 = n192 & n2479 ;
  assign n32287 = ~n2478 ;
  assign n2483 = n32287 & n2482 ;
  assign n2484 = n2475 | n2483 ;
  assign n2411 = n2184 & n32269 ;
  assign n32288 = ~n2417 ;
  assign n2421 = n2411 & n32288 ;
  assign n2459 = n2421 & n2431 ;
  assign n2422 = n2408 | n2417 ;
  assign n32289 = ~n2422 ;
  assign n2501 = n32289 & n176 ;
  assign n2502 = n2184 | n2501 ;
  assign n32290 = ~n2459 ;
  assign n2503 = n32290 & n2502 ;
  assign n2672 = n2405 | n2415 ;
  assign n32291 = ~n2672 ;
  assign n2673 = n176 & n32291 ;
  assign n2674 = n2180 | n2673 ;
  assign n32292 = ~n2405 ;
  assign n2412 = n2180 & n32292 ;
  assign n32293 = ~n2415 ;
  assign n2675 = n2412 & n32293 ;
  assign n2676 = n176 & n2675 ;
  assign n32294 = ~n2676 ;
  assign n2677 = n2674 & n32294 ;
  assign n295 = x92 | x93 ;
  assign n32295 = ~x94 ;
  assign n453 = n32295 & n295 ;
  assign n32296 = ~n2431 ;
  assign n2432 = x94 & n32296 ;
  assign n2433 = n453 | n2432 ;
  assign n32297 = ~n2433 ;
  assign n2434 = n177 & n32297 ;
  assign n32298 = ~n2187 ;
  assign n2446 = n32298 & n2431 ;
  assign n2447 = n32295 & n2431 ;
  assign n32299 = ~n2447 ;
  assign n2448 = x95 & n32299 ;
  assign n2449 = n2446 | n2448 ;
  assign n346 = x94 | n295 ;
  assign n2157 = n346 & n32178 ;
  assign n2158 = n32179 & n2157 ;
  assign n2159 = n32180 & n2158 ;
  assign n2160 = n32181 & n2159 ;
  assign n2450 = x94 & n2431 ;
  assign n32300 = ~n2450 ;
  assign n2451 = n2160 & n32300 ;
  assign n2452 = n2449 | n2451 ;
  assign n32301 = ~n2434 ;
  assign n2453 = n32301 & n2452 ;
  assign n32302 = ~n2453 ;
  assign n2454 = n178 & n32302 ;
  assign n32303 = ~n2155 ;
  assign n2174 = n32303 & n177 ;
  assign n2198 = n2174 & n32282 ;
  assign n2465 = n2198 & n32283 ;
  assign n2466 = n32284 & n2465 ;
  assign n2467 = n2446 | n2466 ;
  assign n2468 = x96 & n2467 ;
  assign n2469 = x96 | n2466 ;
  assign n2470 = n2446 | n2469 ;
  assign n32304 = ~n2468 ;
  assign n2471 = n32304 & n2470 ;
  assign n2517 = x94 & n176 ;
  assign n32305 = ~n2517 ;
  assign n2518 = n346 & n32305 ;
  assign n32306 = ~n2518 ;
  assign n2519 = n177 & n32306 ;
  assign n2520 = n178 | n2519 ;
  assign n32307 = ~n2520 ;
  assign n2521 = n2452 & n32307 ;
  assign n2522 = n2471 | n2521 ;
  assign n32308 = ~n2454 ;
  assign n2523 = n32308 & n2522 ;
  assign n32309 = ~n2523 ;
  assign n2526 = n179 & n32309 ;
  assign n32310 = ~n2209 ;
  assign n2210 = n2193 & n32310 ;
  assign n32311 = ~n2216 ;
  assign n2217 = n2210 & n32311 ;
  assign n2458 = n2217 & n2431 ;
  assign n2218 = n2209 | n2216 ;
  assign n32312 = ~n2218 ;
  assign n2510 = n32312 & n176 ;
  assign n2511 = n2193 | n2510 ;
  assign n32313 = ~n2458 ;
  assign n2512 = n32313 & n2511 ;
  assign n2455 = n179 | n2454 ;
  assign n32314 = ~n2455 ;
  assign n2528 = n32314 & n2522 ;
  assign n2529 = n2512 | n2528 ;
  assign n32315 = ~n2526 ;
  assign n2530 = n32315 & n2529 ;
  assign n32316 = ~n2530 ;
  assign n2531 = n180 & n32316 ;
  assign n32317 = ~n2220 ;
  assign n2231 = n32317 & n2230 ;
  assign n2232 = n32183 & n2231 ;
  assign n2463 = n2232 & n2431 ;
  assign n2221 = n2213 | n2220 ;
  assign n32318 = ~n2221 ;
  assign n2507 = n32318 & n176 ;
  assign n2508 = n2230 | n2507 ;
  assign n32319 = ~n2463 ;
  assign n2509 = n32319 & n2508 ;
  assign n2524 = n1707 & n32309 ;
  assign n2527 = n1487 | n2524 ;
  assign n32320 = ~n2527 ;
  assign n2532 = n32320 & n2529 ;
  assign n2533 = n2509 | n2532 ;
  assign n32321 = ~n2531 ;
  assign n2534 = n32321 & n2533 ;
  assign n32322 = ~n2534 ;
  assign n2535 = n181 & n32322 ;
  assign n2242 = n32188 & n2241 ;
  assign n32323 = ~n2244 ;
  assign n2245 = n2242 & n32323 ;
  assign n2445 = n2245 & n2431 ;
  assign n2246 = n2235 | n2244 ;
  assign n32324 = ~n2246 ;
  assign n2460 = n32324 & n2431 ;
  assign n2461 = n2241 | n2460 ;
  assign n32325 = ~n2445 ;
  assign n2462 = n32325 & n2461 ;
  assign n32326 = ~n2519 ;
  assign n2539 = n2452 & n32326 ;
  assign n32327 = ~n2539 ;
  assign n2540 = n178 & n32327 ;
  assign n2541 = n1707 | n2540 ;
  assign n32328 = ~n2541 ;
  assign n2542 = n2522 & n32328 ;
  assign n2543 = n2512 | n2542 ;
  assign n32329 = ~n2524 ;
  assign n2544 = n32329 & n2543 ;
  assign n32330 = ~n2544 ;
  assign n2545 = n1487 & n32330 ;
  assign n2546 = n181 | n2545 ;
  assign n32331 = ~n2546 ;
  assign n2547 = n2533 & n32331 ;
  assign n2548 = n2462 | n2547 ;
  assign n32332 = ~n2535 ;
  assign n2549 = n32332 & n2548 ;
  assign n32333 = ~n2549 ;
  assign n2550 = n182 & n32333 ;
  assign n32334 = ~n2258 ;
  assign n2259 = n2256 & n32334 ;
  assign n2260 = n32194 & n2259 ;
  assign n2443 = n2260 & n2431 ;
  assign n2261 = n2249 | n2258 ;
  assign n32335 = ~n2261 ;
  assign n2514 = n32335 & n176 ;
  assign n2515 = n2256 | n2514 ;
  assign n32336 = ~n2443 ;
  assign n2516 = n32336 & n2515 ;
  assign n2536 = n182 | n2535 ;
  assign n32337 = ~n2536 ;
  assign n2551 = n32337 & n2548 ;
  assign n2552 = n2516 | n2551 ;
  assign n32338 = ~n2550 ;
  assign n2553 = n32338 & n2552 ;
  assign n32339 = ~n2553 ;
  assign n2554 = n996 & n32339 ;
  assign n2272 = n32205 & n2271 ;
  assign n32340 = ~n2284 ;
  assign n2285 = n2272 & n32340 ;
  assign n2444 = n2285 & n2431 ;
  assign n2286 = n2264 | n2284 ;
  assign n32341 = ~n2286 ;
  assign n2498 = n32341 & n176 ;
  assign n2499 = n2271 | n2498 ;
  assign n32342 = ~n2444 ;
  assign n2500 = n32342 & n2499 ;
  assign n2557 = n32320 & n2543 ;
  assign n2558 = n2509 | n2557 ;
  assign n32343 = ~n2545 ;
  assign n2559 = n32343 & n2558 ;
  assign n32344 = ~n2559 ;
  assign n2560 = n181 & n32344 ;
  assign n2561 = n32331 & n2558 ;
  assign n2562 = n2462 | n2561 ;
  assign n32345 = ~n2560 ;
  assign n2563 = n32345 & n2562 ;
  assign n32346 = ~n2563 ;
  assign n2564 = n182 & n32346 ;
  assign n2565 = n183 | n2564 ;
  assign n32347 = ~n2565 ;
  assign n2566 = n2552 & n32347 ;
  assign n2567 = n2500 | n2566 ;
  assign n32348 = ~n2554 ;
  assign n2568 = n32348 & n2567 ;
  assign n32349 = ~n2568 ;
  assign n2569 = n184 & n32349 ;
  assign n2555 = n838 | n2554 ;
  assign n32350 = ~n2555 ;
  assign n2570 = n32350 & n2567 ;
  assign n32351 = ~n2298 ;
  assign n2299 = n2296 & n32351 ;
  assign n2300 = n32211 & n2299 ;
  assign n2464 = n2300 & n2431 ;
  assign n2301 = n2289 | n2298 ;
  assign n32352 = ~n2301 ;
  assign n2599 = n32352 & n176 ;
  assign n2600 = n2296 | n2599 ;
  assign n32353 = ~n2464 ;
  assign n2601 = n32353 & n2600 ;
  assign n2602 = n2570 | n2601 ;
  assign n32354 = ~n2569 ;
  assign n2603 = n32354 & n2602 ;
  assign n32355 = ~n2603 ;
  assign n2604 = n185 & n32355 ;
  assign n2313 = n32221 & n2312 ;
  assign n32356 = ~n2323 ;
  assign n2324 = n2313 & n32356 ;
  assign n2442 = n2324 & n2431 ;
  assign n2325 = n2304 | n2323 ;
  assign n32357 = ~n2325 ;
  assign n2596 = n32357 & n176 ;
  assign n2597 = n2312 | n2596 ;
  assign n32358 = ~n2442 ;
  assign n2598 = n32358 & n2597 ;
  assign n2571 = n32337 & n2562 ;
  assign n2572 = n2516 | n2571 ;
  assign n32359 = ~n2564 ;
  assign n2573 = n32359 & n2572 ;
  assign n32360 = ~n2573 ;
  assign n2574 = n183 & n32360 ;
  assign n2575 = n32347 & n2572 ;
  assign n2576 = n2500 | n2575 ;
  assign n32361 = ~n2574 ;
  assign n2577 = n32361 & n2576 ;
  assign n32362 = ~n2577 ;
  assign n2578 = n838 & n32362 ;
  assign n2579 = n185 | n2578 ;
  assign n32363 = ~n2579 ;
  assign n2607 = n32363 & n2602 ;
  assign n2608 = n2598 | n2607 ;
  assign n32364 = ~n2604 ;
  assign n2609 = n32364 & n2608 ;
  assign n32365 = ~n2609 ;
  assign n2610 = n186 & n32365 ;
  assign n32366 = ~n2327 ;
  assign n2338 = n32366 & n2337 ;
  assign n2339 = n32227 & n2338 ;
  assign n2441 = n2339 & n2431 ;
  assign n2330 = n2327 | n2329 ;
  assign n32367 = ~n2330 ;
  assign n2495 = n32367 & n176 ;
  assign n2496 = n2337 | n2495 ;
  assign n32368 = ~n2441 ;
  assign n2497 = n32368 & n2496 ;
  assign n2605 = n186 | n2604 ;
  assign n32369 = ~n2605 ;
  assign n2611 = n32369 & n2608 ;
  assign n2612 = n2497 | n2611 ;
  assign n32370 = ~n2610 ;
  assign n2613 = n32370 & n2612 ;
  assign n32371 = ~n2613 ;
  assign n2614 = n528 & n32371 ;
  assign n2351 = n32237 & n2350 ;
  assign n32372 = ~n2371 ;
  assign n2372 = n2351 & n32372 ;
  assign n2440 = n2372 & n2431 ;
  assign n2373 = n2342 | n2371 ;
  assign n32373 = ~n2373 ;
  assign n2504 = n32373 & n176 ;
  assign n2505 = n2350 | n2504 ;
  assign n32374 = ~n2440 ;
  assign n2506 = n32374 & n2505 ;
  assign n2580 = n32350 & n2576 ;
  assign n2619 = n2580 | n2601 ;
  assign n32375 = ~n2578 ;
  assign n2620 = n32375 & n2619 ;
  assign n32376 = ~n2620 ;
  assign n2621 = n185 & n32376 ;
  assign n2622 = n32363 & n2619 ;
  assign n2623 = n2598 | n2622 ;
  assign n32377 = ~n2621 ;
  assign n2624 = n32377 & n2623 ;
  assign n32378 = ~n2624 ;
  assign n2625 = n186 & n32378 ;
  assign n2626 = n528 | n2625 ;
  assign n32379 = ~n2626 ;
  assign n2627 = n2612 & n32379 ;
  assign n2628 = n2506 | n2627 ;
  assign n32380 = ~n2614 ;
  assign n2629 = n32380 & n2628 ;
  assign n32381 = ~n2629 ;
  assign n2630 = n188 & n32381 ;
  assign n32382 = ~n2388 ;
  assign n2389 = n2383 & n32382 ;
  assign n2390 = n32243 & n2389 ;
  assign n2436 = n2390 & n2431 ;
  assign n2391 = n2376 | n2388 ;
  assign n32383 = ~n2391 ;
  assign n2437 = n32383 & n2431 ;
  assign n2438 = n2383 | n2437 ;
  assign n32384 = ~n2436 ;
  assign n2439 = n32384 & n2438 ;
  assign n2615 = n413 | n2614 ;
  assign n32385 = ~n2615 ;
  assign n2631 = n32385 & n2628 ;
  assign n2632 = n2439 | n2631 ;
  assign n32386 = ~n2630 ;
  assign n2633 = n32386 & n2632 ;
  assign n32387 = ~n2633 ;
  assign n2634 = n189 & n32387 ;
  assign n2635 = n190 | n2634 ;
  assign n2636 = n32369 & n2623 ;
  assign n2637 = n2497 | n2636 ;
  assign n32388 = ~n2625 ;
  assign n2638 = n32388 & n2637 ;
  assign n32389 = ~n2638 ;
  assign n2639 = n187 & n32389 ;
  assign n2640 = n32379 & n2637 ;
  assign n2641 = n2506 | n2640 ;
  assign n32390 = ~n2639 ;
  assign n2642 = n32390 & n2641 ;
  assign n32391 = ~n2642 ;
  assign n2643 = n413 & n32391 ;
  assign n2644 = n189 | n2643 ;
  assign n2645 = n32385 & n2641 ;
  assign n2646 = n2439 | n2645 ;
  assign n32392 = ~n2644 ;
  assign n2649 = n32392 & n2646 ;
  assign n2678 = n32253 & n2401 ;
  assign n32393 = ~n2393 ;
  assign n2679 = n32393 & n2678 ;
  assign n2680 = n2431 & n2679 ;
  assign n2397 = n2393 | n2395 ;
  assign n32394 = ~n2397 ;
  assign n2513 = n32394 & n176 ;
  assign n2681 = n2401 | n2513 ;
  assign n32395 = ~n2680 ;
  assign n2682 = n32395 & n2681 ;
  assign n2683 = n2649 | n2682 ;
  assign n32396 = ~n2635 ;
  assign n2684 = n32396 & n2683 ;
  assign n2685 = n2677 | n2684 ;
  assign n32397 = ~n2643 ;
  assign n2647 = n32397 & n2646 ;
  assign n32398 = ~n2647 ;
  assign n2648 = n189 & n32398 ;
  assign n32399 = ~n2648 ;
  assign n2687 = n32399 & n2683 ;
  assign n32400 = ~n2687 ;
  assign n2688 = n190 & n32400 ;
  assign n2690 = n287 | n2688 ;
  assign n32401 = ~n2690 ;
  assign n2691 = n2685 & n32401 ;
  assign n2692 = n2503 | n2691 ;
  assign n32402 = ~n2487 ;
  assign n2661 = n2173 & n32402 ;
  assign n2662 = n32275 & n2661 ;
  assign n2663 = n2431 & n2662 ;
  assign n2665 = n2424 | n2487 ;
  assign n32403 = ~n2665 ;
  assign n2666 = n176 & n32403 ;
  assign n2667 = n2173 | n2666 ;
  assign n32404 = ~n2663 ;
  assign n2668 = n32404 & n2667 ;
  assign n32405 = ~n2688 ;
  assign n2695 = n2685 & n32405 ;
  assign n32406 = ~n2695 ;
  assign n2696 = n191 & n32406 ;
  assign n32407 = ~n2696 ;
  assign n2697 = n2668 & n32407 ;
  assign n2698 = n2692 & n2697 ;
  assign n2699 = n2484 | n2698 ;
  assign n32408 = ~n2479 ;
  assign n2480 = n2431 & n32408 ;
  assign n2481 = n2429 | n2480 ;
  assign n2669 = n2481 | n2668 ;
  assign n2704 = n2692 & n32407 ;
  assign n2751 = n2669 | n2704 ;
  assign n2752 = n31336 & n2751 ;
  assign n2753 = n2699 | n2752 ;
  assign n2705 = n2668 | n2704 ;
  assign n32409 = ~n2705 ;
  assign n2795 = n32409 & n2753 ;
  assign n2796 = n2698 | n2795 ;
  assign n2703 = n2503 & n32407 ;
  assign n2689 = n191 | n2688 ;
  assign n32410 = ~n2689 ;
  assign n2707 = n2685 & n32410 ;
  assign n32411 = ~n2707 ;
  assign n2940 = n2703 & n32411 ;
  assign n2941 = n2753 & n2940 ;
  assign n2708 = n2503 | n2707 ;
  assign n2709 = n32407 & n2708 ;
  assign n2710 = n2669 | n2709 ;
  assign n2711 = n31336 & n2710 ;
  assign n2712 = n2697 & n2708 ;
  assign n2713 = n2484 | n2712 ;
  assign n175 = n2711 | n2713 ;
  assign n2943 = n2696 | n2707 ;
  assign n32412 = ~n2943 ;
  assign n2944 = n175 & n32412 ;
  assign n2945 = n2503 | n2944 ;
  assign n32413 = ~n2941 ;
  assign n2946 = n32413 & n2945 ;
  assign n2947 = n2796 | n2946 ;
  assign n32414 = ~n295 ;
  assign n2774 = n32414 & n2753 ;
  assign n32415 = ~x92 ;
  assign n2775 = n32415 & n2753 ;
  assign n32416 = ~n2775 ;
  assign n2776 = x93 & n32416 ;
  assign n2777 = n2774 | n2776 ;
  assign n514 = x90 | x91 ;
  assign n616 = x92 | n514 ;
  assign n2156 = n616 & n32303 ;
  assign n2200 = n2156 & n32282 ;
  assign n2472 = n2200 & n32283 ;
  assign n2473 = n32284 & n2472 ;
  assign n2778 = x92 & n2753 ;
  assign n32417 = ~n2778 ;
  assign n2779 = n2473 & n32417 ;
  assign n2780 = n2777 | n2779 ;
  assign n721 = n32415 & n514 ;
  assign n32418 = ~n2753 ;
  assign n2784 = x92 & n32418 ;
  assign n2785 = n721 | n2784 ;
  assign n32419 = ~n2785 ;
  assign n2786 = n2431 & n32419 ;
  assign n32420 = ~n2786 ;
  assign n2787 = n2780 & n32420 ;
  assign n32421 = ~n2787 ;
  assign n2788 = n177 & n32421 ;
  assign n2743 = x92 & n175 ;
  assign n32422 = ~n2743 ;
  assign n2744 = n616 & n32422 ;
  assign n32423 = ~n2744 ;
  assign n2745 = n176 & n32423 ;
  assign n2746 = n177 | n2745 ;
  assign n32424 = ~n2746 ;
  assign n2781 = n32424 & n2780 ;
  assign n32425 = ~n2475 ;
  assign n2476 = n2431 & n32425 ;
  assign n32426 = ~n2483 ;
  assign n2485 = n2476 & n32426 ;
  assign n32427 = ~n2698 ;
  assign n2700 = n2485 & n32427 ;
  assign n32428 = ~n2752 ;
  assign n2799 = n2700 & n32428 ;
  assign n2800 = n2774 | n2799 ;
  assign n2801 = x94 & n2800 ;
  assign n2802 = x94 | n2799 ;
  assign n2803 = n2774 | n2802 ;
  assign n32429 = ~n2801 ;
  assign n2804 = n32429 & n2803 ;
  assign n2805 = n2781 | n2804 ;
  assign n32430 = ~n2788 ;
  assign n2806 = n32430 & n2805 ;
  assign n32431 = ~n2806 ;
  assign n2807 = n178 & n32431 ;
  assign n2456 = n2434 | n2451 ;
  assign n32432 = ~n2456 ;
  assign n2728 = n32432 & n175 ;
  assign n2729 = n2449 | n2728 ;
  assign n2457 = n2449 & n32432 ;
  assign n2772 = n2457 & n2753 ;
  assign n32433 = ~n2772 ;
  assign n2773 = n2729 & n32433 ;
  assign n2789 = n178 | n2788 ;
  assign n2790 = n177 | n2786 ;
  assign n32434 = ~n2790 ;
  assign n2791 = n2780 & n32434 ;
  assign n2812 = n2791 | n2804 ;
  assign n32435 = ~n2789 ;
  assign n2813 = n32435 & n2812 ;
  assign n2814 = n2773 | n2813 ;
  assign n32436 = ~n2807 ;
  assign n2815 = n32436 & n2814 ;
  assign n32437 = ~n2815 ;
  assign n2816 = n1707 & n32437 ;
  assign n2595 = n2521 | n2540 ;
  assign n32438 = ~n2595 ;
  assign n2726 = n32438 & n175 ;
  assign n2727 = n2471 | n2726 ;
  assign n32439 = ~n2521 ;
  assign n2538 = n2471 & n32439 ;
  assign n32440 = ~n2540 ;
  assign n2594 = n2538 & n32440 ;
  assign n2770 = n2594 & n2753 ;
  assign n32441 = ~n2770 ;
  assign n2771 = n2727 & n32441 ;
  assign n2809 = n1707 | n2807 ;
  assign n32442 = ~n2809 ;
  assign n2818 = n32442 & n2814 ;
  assign n2819 = n2771 | n2818 ;
  assign n32443 = ~n2816 ;
  assign n2820 = n32443 & n2819 ;
  assign n32444 = ~n2820 ;
  assign n2821 = n180 & n32444 ;
  assign n2593 = n2524 | n2542 ;
  assign n32445 = ~n2593 ;
  assign n2739 = n32445 & n175 ;
  assign n2740 = n2512 | n2739 ;
  assign n2525 = n2512 & n32329 ;
  assign n32446 = ~n2542 ;
  assign n2592 = n2525 & n32446 ;
  assign n2768 = n2592 & n2753 ;
  assign n32447 = ~n2768 ;
  assign n2769 = n2740 & n32447 ;
  assign n2817 = n1487 | n2816 ;
  assign n32448 = ~n2817 ;
  assign n2822 = n32448 & n2819 ;
  assign n2823 = n2769 | n2822 ;
  assign n32449 = ~n2821 ;
  assign n2824 = n32449 & n2823 ;
  assign n32450 = ~n2824 ;
  assign n2825 = n181 & n32450 ;
  assign n2591 = n2545 | n2557 ;
  assign n32451 = ~n2591 ;
  assign n2717 = n32451 & n175 ;
  assign n2718 = n2509 | n2717 ;
  assign n32452 = ~n2557 ;
  assign n2589 = n2509 & n32452 ;
  assign n2590 = n32343 & n2589 ;
  assign n2766 = n2590 & n2753 ;
  assign n32453 = ~n2766 ;
  assign n2767 = n2718 & n32453 ;
  assign n2831 = n179 & n32437 ;
  assign n32454 = ~n2831 ;
  assign n2832 = n2819 & n32454 ;
  assign n32455 = ~n2832 ;
  assign n2833 = n1487 & n32455 ;
  assign n2834 = n181 | n2833 ;
  assign n32456 = ~n2834 ;
  assign n2835 = n2823 & n32456 ;
  assign n2836 = n2767 | n2835 ;
  assign n32457 = ~n2825 ;
  assign n2837 = n32457 & n2836 ;
  assign n32458 = ~n2837 ;
  assign n2838 = n182 & n32458 ;
  assign n2588 = n2560 | n2561 ;
  assign n32459 = ~n2588 ;
  assign n2730 = n32459 & n175 ;
  assign n2731 = n2462 | n2730 ;
  assign n2537 = n2462 & n32332 ;
  assign n32460 = ~n2561 ;
  assign n2587 = n2537 & n32460 ;
  assign n2764 = n2587 & n2753 ;
  assign n32461 = ~n2764 ;
  assign n2765 = n2731 & n32461 ;
  assign n2826 = n182 | n2825 ;
  assign n32462 = ~n2826 ;
  assign n2839 = n32462 & n2836 ;
  assign n2840 = n2765 | n2839 ;
  assign n32463 = ~n2838 ;
  assign n2841 = n32463 & n2840 ;
  assign n32464 = ~n2841 ;
  assign n2842 = n996 & n32464 ;
  assign n2586 = n2564 | n2571 ;
  assign n32465 = ~n2586 ;
  assign n2741 = n32465 & n175 ;
  assign n2742 = n2516 | n2741 ;
  assign n32466 = ~n2571 ;
  assign n2584 = n2516 & n32466 ;
  assign n2585 = n32359 & n2584 ;
  assign n2797 = n2585 & n2753 ;
  assign n32467 = ~n2797 ;
  assign n2798 = n2742 & n32467 ;
  assign n32468 = ~n2833 ;
  assign n2850 = n2823 & n32468 ;
  assign n32469 = ~n2850 ;
  assign n2851 = n181 & n32469 ;
  assign n32470 = ~n2851 ;
  assign n2852 = n2836 & n32470 ;
  assign n32471 = ~n2852 ;
  assign n2853 = n182 & n32471 ;
  assign n2854 = n183 | n2853 ;
  assign n32472 = ~n2854 ;
  assign n2855 = n2840 & n32472 ;
  assign n2856 = n2798 | n2855 ;
  assign n32473 = ~n2842 ;
  assign n2857 = n32473 & n2856 ;
  assign n32474 = ~n2857 ;
  assign n2858 = n184 & n32474 ;
  assign n2583 = n2574 | n2575 ;
  assign n32475 = ~n2583 ;
  assign n2732 = n32475 & n175 ;
  assign n2733 = n2500 | n2732 ;
  assign n2556 = n2500 & n32348 ;
  assign n32476 = ~n2575 ;
  assign n2582 = n2556 & n32476 ;
  assign n2754 = n2582 & n2753 ;
  assign n32477 = ~n2754 ;
  assign n2755 = n2733 & n32477 ;
  assign n2843 = n838 | n2842 ;
  assign n32478 = ~n2843 ;
  assign n2859 = n32478 & n2856 ;
  assign n2860 = n2755 | n2859 ;
  assign n32479 = ~n2858 ;
  assign n2861 = n32479 & n2860 ;
  assign n32480 = ~n2861 ;
  assign n2862 = n185 & n32480 ;
  assign n2581 = n2578 | n2580 ;
  assign n32481 = ~n2581 ;
  assign n2715 = n32481 & n175 ;
  assign n2716 = n2601 | n2715 ;
  assign n32482 = ~n2580 ;
  assign n2617 = n32482 & n2601 ;
  assign n2618 = n32375 & n2617 ;
  assign n2762 = n2618 & n2753 ;
  assign n32483 = ~n2762 ;
  assign n2763 = n2716 & n32483 ;
  assign n32484 = ~n2853 ;
  assign n2870 = n2840 & n32484 ;
  assign n32485 = ~n2870 ;
  assign n2871 = n183 & n32485 ;
  assign n32486 = ~n2871 ;
  assign n2872 = n2856 & n32486 ;
  assign n32487 = ~n2872 ;
  assign n2873 = n838 & n32487 ;
  assign n2874 = n185 | n2873 ;
  assign n32488 = ~n2874 ;
  assign n2875 = n2860 & n32488 ;
  assign n2876 = n2763 | n2875 ;
  assign n32489 = ~n2862 ;
  assign n2877 = n32489 & n2876 ;
  assign n32490 = ~n2877 ;
  assign n2878 = n186 & n32490 ;
  assign n2660 = n2621 | n2622 ;
  assign n32491 = ~n2660 ;
  assign n2719 = n32491 & n175 ;
  assign n2720 = n2598 | n2719 ;
  assign n2606 = n2598 & n32364 ;
  assign n32492 = ~n2622 ;
  assign n2659 = n2606 & n32492 ;
  assign n2760 = n2659 & n2753 ;
  assign n32493 = ~n2760 ;
  assign n2761 = n2720 & n32493 ;
  assign n2863 = n186 | n2862 ;
  assign n32494 = ~n2863 ;
  assign n2879 = n32494 & n2876 ;
  assign n2880 = n2761 | n2879 ;
  assign n32495 = ~n2878 ;
  assign n2881 = n32495 & n2880 ;
  assign n32496 = ~n2881 ;
  assign n2882 = n528 & n32496 ;
  assign n2658 = n2625 | n2636 ;
  assign n32497 = ~n2658 ;
  assign n2721 = n32497 & n175 ;
  assign n2722 = n2497 | n2721 ;
  assign n32498 = ~n2636 ;
  assign n2656 = n2497 & n32498 ;
  assign n2657 = n32388 & n2656 ;
  assign n2758 = n2657 & n2753 ;
  assign n32499 = ~n2758 ;
  assign n2759 = n2722 & n32499 ;
  assign n32500 = ~n2873 ;
  assign n2890 = n2860 & n32500 ;
  assign n32501 = ~n2890 ;
  assign n2891 = n185 & n32501 ;
  assign n32502 = ~n2891 ;
  assign n2892 = n2876 & n32502 ;
  assign n32503 = ~n2892 ;
  assign n2893 = n186 & n32503 ;
  assign n2894 = n528 | n2893 ;
  assign n32504 = ~n2894 ;
  assign n2895 = n2880 & n32504 ;
  assign n2896 = n2759 | n2895 ;
  assign n32505 = ~n2882 ;
  assign n2897 = n32505 & n2896 ;
  assign n32506 = ~n2897 ;
  assign n2898 = n188 & n32506 ;
  assign n2655 = n2639 | n2640 ;
  assign n32507 = ~n2655 ;
  assign n2724 = n32507 & n175 ;
  assign n2725 = n2506 | n2724 ;
  assign n2616 = n2506 & n32380 ;
  assign n32508 = ~n2640 ;
  assign n2654 = n2616 & n32508 ;
  assign n2782 = n2654 & n2753 ;
  assign n32509 = ~n2782 ;
  assign n2783 = n2725 & n32509 ;
  assign n2883 = n413 | n2882 ;
  assign n32510 = ~n2883 ;
  assign n2899 = n32510 & n2896 ;
  assign n2901 = n2783 | n2899 ;
  assign n32511 = ~n2898 ;
  assign n2902 = n32511 & n2901 ;
  assign n32512 = ~n2902 ;
  assign n2903 = n189 & n32512 ;
  assign n2653 = n2643 | n2645 ;
  assign n32513 = ~n2653 ;
  assign n2734 = n32513 & n175 ;
  assign n2735 = n2439 | n2734 ;
  assign n32514 = ~n2645 ;
  assign n2651 = n2439 & n32514 ;
  assign n2652 = n32397 & n2651 ;
  assign n2756 = n2652 & n2753 ;
  assign n32515 = ~n2756 ;
  assign n2757 = n2735 & n32515 ;
  assign n32516 = ~n2893 ;
  assign n2910 = n2880 & n32516 ;
  assign n32517 = ~n2910 ;
  assign n2911 = n187 & n32517 ;
  assign n32518 = ~n2911 ;
  assign n2912 = n2896 & n32518 ;
  assign n32519 = ~n2912 ;
  assign n2913 = n413 & n32519 ;
  assign n2914 = n189 | n2913 ;
  assign n32520 = ~n2914 ;
  assign n2915 = n2901 & n32520 ;
  assign n2916 = n2757 | n2915 ;
  assign n32521 = ~n2903 ;
  assign n2917 = n32521 & n2916 ;
  assign n32522 = ~n2917 ;
  assign n2918 = n190 & n32522 ;
  assign n2904 = n190 | n2903 ;
  assign n32523 = ~n2904 ;
  assign n2919 = n32523 & n2916 ;
  assign n32524 = ~n2634 ;
  assign n2950 = n32524 & n2682 ;
  assign n32525 = ~n2649 ;
  assign n2951 = n32525 & n2950 ;
  assign n2952 = n175 & n2951 ;
  assign n2650 = n2648 | n2649 ;
  assign n32526 = ~n2650 ;
  assign n2747 = n32526 & n175 ;
  assign n2953 = n2682 | n2747 ;
  assign n32527 = ~n2952 ;
  assign n2954 = n32527 & n2953 ;
  assign n2955 = n2919 | n2954 ;
  assign n32528 = ~n2918 ;
  assign n2958 = n32528 & n2955 ;
  assign n32529 = ~n2958 ;
  assign n2959 = n287 & n32529 ;
  assign n32530 = ~n2684 ;
  assign n2686 = n2677 & n32530 ;
  assign n2693 = n2686 & n32405 ;
  assign n2723 = n2693 & n175 ;
  assign n2694 = n2684 | n2688 ;
  assign n32531 = ~n2694 ;
  assign n2736 = n32531 & n175 ;
  assign n2737 = n2677 | n2736 ;
  assign n32532 = ~n2723 ;
  assign n2738 = n32532 & n2737 ;
  assign n32533 = ~n2913 ;
  assign n2926 = n2901 & n32533 ;
  assign n32534 = ~n2926 ;
  assign n2927 = n189 & n32534 ;
  assign n32535 = ~n2927 ;
  assign n2928 = n2916 & n32535 ;
  assign n32536 = ~n2928 ;
  assign n2929 = n190 & n32536 ;
  assign n2930 = n287 | n2929 ;
  assign n32537 = ~n2930 ;
  assign n2956 = n32537 & n2955 ;
  assign n2963 = n2738 | n2956 ;
  assign n32538 = ~n2959 ;
  assign n2964 = n32538 & n2963 ;
  assign n2965 = n2947 | n2964 ;
  assign n2966 = n31336 & n2965 ;
  assign n2706 = n192 & n2705 ;
  assign n32539 = ~n2668 ;
  assign n2748 = n32539 & n175 ;
  assign n32540 = ~n2748 ;
  assign n2749 = n2704 & n32540 ;
  assign n32541 = ~n2749 ;
  assign n2750 = n2706 & n32541 ;
  assign n2664 = n2475 | n2663 ;
  assign n32542 = ~n2664 ;
  assign n2670 = n32542 & n2667 ;
  assign n2671 = n32426 & n2670 ;
  assign n2701 = n2671 & n32427 ;
  assign n2933 = n2701 & n32428 ;
  assign n2934 = n2750 | n2933 ;
  assign n2961 = n2946 & n32538 ;
  assign n2969 = n2961 & n2963 ;
  assign n2973 = n2934 | n2969 ;
  assign n174 = n2966 | n2973 ;
  assign n2962 = n2956 | n2959 ;
  assign n32543 = ~n2962 ;
  assign n2993 = n32543 & n174 ;
  assign n2994 = n2738 | n2993 ;
  assign n32544 = ~n2956 ;
  assign n2957 = n2738 & n32544 ;
  assign n2960 = n2957 & n32538 ;
  assign n2996 = n2960 & n174 ;
  assign n32545 = ~n2996 ;
  assign n2997 = n2994 & n32545 ;
  assign n2967 = n2946 | n2964 ;
  assign n32546 = ~n2967 ;
  assign n2990 = n32546 & n174 ;
  assign n3242 = n2969 | n2990 ;
  assign n3243 = n2997 | n3242 ;
  assign n32547 = ~n2933 ;
  assign n2935 = n2753 & n32547 ;
  assign n32548 = ~n2750 ;
  assign n2936 = n32548 & n2935 ;
  assign n32549 = ~n2969 ;
  assign n2970 = n2936 & n32549 ;
  assign n32550 = ~n2966 ;
  assign n2971 = n32550 & n2970 ;
  assign n32551 = ~n514 ;
  assign n2978 = n32551 & n174 ;
  assign n2979 = n2971 | n2978 ;
  assign n2980 = x92 & n2979 ;
  assign n2972 = x92 | n2971 ;
  assign n2995 = n2972 | n2978 ;
  assign n32552 = ~n2980 ;
  assign n3019 = n32552 & n2995 ;
  assign n866 = x88 | x89 ;
  assign n32553 = ~x90 ;
  assign n1137 = n32553 & n866 ;
  assign n32554 = ~n174 ;
  assign n2981 = x90 & n32554 ;
  assign n2982 = n1137 | n2981 ;
  assign n32555 = ~n2982 ;
  assign n2983 = n2753 & n32555 ;
  assign n2984 = n2431 | n2983 ;
  assign n984 = x90 | n866 ;
  assign n2477 = n984 & n32425 ;
  assign n2486 = n2477 & n32426 ;
  assign n2702 = n2486 & n32427 ;
  assign n2939 = n2702 & n32428 ;
  assign n2976 = x90 & n174 ;
  assign n32556 = ~n2976 ;
  assign n2977 = n2939 & n32556 ;
  assign n3055 = n32553 & n174 ;
  assign n32557 = ~n3055 ;
  assign n3056 = x91 & n32557 ;
  assign n3057 = n2978 | n3056 ;
  assign n3058 = n2977 | n3057 ;
  assign n32558 = ~n2984 ;
  assign n3059 = n32558 & n3058 ;
  assign n3060 = n3019 | n3059 ;
  assign n3048 = n984 & n32556 ;
  assign n32559 = ~n3048 ;
  assign n3049 = n175 & n32559 ;
  assign n32560 = ~n3049 ;
  assign n3063 = n32560 & n3058 ;
  assign n32561 = ~n3063 ;
  assign n3064 = n2431 & n32561 ;
  assign n32562 = ~n3064 ;
  assign n3065 = n3060 & n32562 ;
  assign n32563 = ~n3065 ;
  assign n3066 = n177 & n32563 ;
  assign n2793 = n2779 | n2786 ;
  assign n32564 = ~n2793 ;
  assign n2794 = n2777 & n32564 ;
  assign n2975 = n2794 & n174 ;
  assign n3011 = n32564 & n174 ;
  assign n3012 = n2777 | n3011 ;
  assign n32565 = ~n2975 ;
  assign n3013 = n32565 & n3012 ;
  assign n3070 = n177 | n3064 ;
  assign n32566 = ~n3070 ;
  assign n3071 = n3060 & n32566 ;
  assign n3072 = n3013 | n3071 ;
  assign n32567 = ~n3066 ;
  assign n3073 = n32567 & n3072 ;
  assign n32568 = ~n3073 ;
  assign n3074 = n178 & n32568 ;
  assign n32569 = ~n2791 ;
  assign n2810 = n32569 & n2804 ;
  assign n2811 = n32430 & n2810 ;
  assign n3003 = n2811 & n174 ;
  assign n2792 = n2788 | n2791 ;
  assign n32570 = ~n2792 ;
  assign n3022 = n32570 & n174 ;
  assign n3023 = n2804 | n3022 ;
  assign n32571 = ~n3003 ;
  assign n3024 = n32571 & n3023 ;
  assign n3067 = n178 | n3066 ;
  assign n32572 = ~n3067 ;
  assign n3075 = n32572 & n3072 ;
  assign n3076 = n3024 | n3075 ;
  assign n32573 = ~n3074 ;
  assign n3077 = n32573 & n3076 ;
  assign n32574 = ~n3077 ;
  assign n3078 = n1707 & n32574 ;
  assign n2808 = n2773 & n32436 ;
  assign n32575 = ~n2813 ;
  assign n2931 = n2808 & n32575 ;
  assign n2989 = n2931 & n174 ;
  assign n2932 = n2807 | n2813 ;
  assign n32576 = ~n2932 ;
  assign n3025 = n32576 & n174 ;
  assign n3026 = n2773 | n3025 ;
  assign n32577 = ~n2989 ;
  assign n3027 = n32577 & n3026 ;
  assign n3085 = n176 & n32561 ;
  assign n3050 = n176 | n3049 ;
  assign n32578 = ~n3050 ;
  assign n3087 = n32578 & n3058 ;
  assign n3088 = n3019 | n3087 ;
  assign n32579 = ~n3085 ;
  assign n3089 = n32579 & n3088 ;
  assign n32580 = ~n3089 ;
  assign n3090 = n177 & n32580 ;
  assign n3091 = n32566 & n3088 ;
  assign n3092 = n3013 | n3091 ;
  assign n32581 = ~n3090 ;
  assign n3093 = n32581 & n3092 ;
  assign n32582 = ~n3093 ;
  assign n3094 = n178 & n32582 ;
  assign n3095 = n1707 | n3094 ;
  assign n32583 = ~n3095 ;
  assign n3096 = n3076 & n32583 ;
  assign n3097 = n3027 | n3096 ;
  assign n32584 = ~n3078 ;
  assign n3098 = n32584 & n3097 ;
  assign n32585 = ~n3098 ;
  assign n3099 = n180 & n32585 ;
  assign n2830 = n2816 | n2818 ;
  assign n32586 = ~n2830 ;
  assign n2991 = n32586 & n174 ;
  assign n2992 = n2771 | n2991 ;
  assign n32587 = ~n2818 ;
  assign n2828 = n2771 & n32587 ;
  assign n2829 = n32443 & n2828 ;
  assign n3014 = n2829 & n174 ;
  assign n32588 = ~n3014 ;
  assign n3015 = n2992 & n32588 ;
  assign n3079 = n1487 | n3078 ;
  assign n32589 = ~n3079 ;
  assign n3100 = n32589 & n3097 ;
  assign n3101 = n3015 | n3100 ;
  assign n32590 = ~n3099 ;
  assign n3102 = n32590 & n3101 ;
  assign n32591 = ~n3102 ;
  assign n3103 = n181 & n32591 ;
  assign n2848 = n2769 & n32468 ;
  assign n32592 = ~n2822 ;
  assign n2849 = n32592 & n2848 ;
  assign n2999 = n2849 & n174 ;
  assign n2827 = n2821 | n2822 ;
  assign n32593 = ~n2827 ;
  assign n3000 = n32593 & n174 ;
  assign n3001 = n2769 | n3000 ;
  assign n32594 = ~n2999 ;
  assign n3002 = n32594 & n3001 ;
  assign n3111 = n32572 & n3092 ;
  assign n3112 = n3024 | n3111 ;
  assign n32595 = ~n3094 ;
  assign n3113 = n32595 & n3112 ;
  assign n32596 = ~n3113 ;
  assign n3114 = n179 & n32596 ;
  assign n3115 = n32583 & n3112 ;
  assign n3116 = n3027 | n3115 ;
  assign n32597 = ~n3114 ;
  assign n3117 = n32597 & n3116 ;
  assign n32598 = ~n3117 ;
  assign n3118 = n1487 & n32598 ;
  assign n3119 = n181 | n3118 ;
  assign n32599 = ~n3119 ;
  assign n3120 = n3101 & n32599 ;
  assign n3121 = n3002 | n3120 ;
  assign n32600 = ~n3103 ;
  assign n3122 = n32600 & n3121 ;
  assign n32601 = ~n3122 ;
  assign n3123 = n182 & n32601 ;
  assign n2845 = n2825 | n2835 ;
  assign n32602 = ~n2845 ;
  assign n3034 = n32602 & n174 ;
  assign n3035 = n2767 | n3034 ;
  assign n32603 = ~n2835 ;
  assign n2846 = n2767 & n32603 ;
  assign n2847 = n32457 & n2846 ;
  assign n3036 = n2847 & n174 ;
  assign n32604 = ~n3036 ;
  assign n3037 = n3035 & n32604 ;
  assign n3104 = n182 | n3103 ;
  assign n32605 = ~n3104 ;
  assign n3124 = n32605 & n3121 ;
  assign n3125 = n3037 | n3124 ;
  assign n32606 = ~n3123 ;
  assign n3126 = n32606 & n3125 ;
  assign n32607 = ~n3126 ;
  assign n3127 = n996 & n32607 ;
  assign n2844 = n2838 | n2839 ;
  assign n32608 = ~n2844 ;
  assign n3016 = n32608 & n174 ;
  assign n3017 = n2765 | n3016 ;
  assign n2868 = n2765 & n32484 ;
  assign n32609 = ~n2839 ;
  assign n2869 = n32609 & n2868 ;
  assign n3038 = n2869 & n174 ;
  assign n32610 = ~n3038 ;
  assign n3039 = n3017 & n32610 ;
  assign n3135 = n32589 & n3116 ;
  assign n3136 = n3015 | n3135 ;
  assign n32611 = ~n3118 ;
  assign n3137 = n32611 & n3136 ;
  assign n32612 = ~n3137 ;
  assign n3138 = n181 & n32612 ;
  assign n3139 = n32599 & n3136 ;
  assign n3140 = n3002 | n3139 ;
  assign n32613 = ~n3138 ;
  assign n3141 = n32613 & n3140 ;
  assign n32614 = ~n3141 ;
  assign n3142 = n182 & n32614 ;
  assign n3143 = n183 | n3142 ;
  assign n32615 = ~n3143 ;
  assign n3144 = n3125 & n32615 ;
  assign n3145 = n3039 | n3144 ;
  assign n32616 = ~n3127 ;
  assign n3146 = n32616 & n3145 ;
  assign n32617 = ~n3146 ;
  assign n3147 = n184 & n32617 ;
  assign n2867 = n2842 | n2855 ;
  assign n32618 = ~n2867 ;
  assign n3007 = n32618 & n174 ;
  assign n3008 = n2798 | n3007 ;
  assign n32619 = ~n2855 ;
  assign n2865 = n2798 & n32619 ;
  assign n2866 = n32473 & n2865 ;
  assign n3029 = n2866 & n174 ;
  assign n32620 = ~n3029 ;
  assign n3030 = n3008 & n32620 ;
  assign n3129 = n838 | n3127 ;
  assign n32621 = ~n3129 ;
  assign n3148 = n32621 & n3145 ;
  assign n3151 = n3030 | n3148 ;
  assign n32622 = ~n3147 ;
  assign n3152 = n32622 & n3151 ;
  assign n32623 = ~n3152 ;
  assign n3153 = n185 & n32623 ;
  assign n2888 = n2755 & n32500 ;
  assign n32624 = ~n2859 ;
  assign n2889 = n32624 & n2888 ;
  assign n3021 = n2889 & n174 ;
  assign n2864 = n2858 | n2859 ;
  assign n32625 = ~n2864 ;
  assign n3040 = n32625 & n174 ;
  assign n3041 = n2755 | n3040 ;
  assign n32626 = ~n3021 ;
  assign n3042 = n32626 & n3041 ;
  assign n3159 = n32605 & n3140 ;
  assign n3160 = n3037 | n3159 ;
  assign n32627 = ~n3142 ;
  assign n3161 = n32627 & n3160 ;
  assign n32628 = ~n3161 ;
  assign n3162 = n183 & n32628 ;
  assign n3163 = n32615 & n3160 ;
  assign n3164 = n3039 | n3163 ;
  assign n32629 = ~n3162 ;
  assign n3165 = n32629 & n3164 ;
  assign n32630 = ~n3165 ;
  assign n3166 = n838 & n32630 ;
  assign n3167 = n185 | n3166 ;
  assign n32631 = ~n3167 ;
  assign n3168 = n3151 & n32631 ;
  assign n3169 = n3042 | n3168 ;
  assign n32632 = ~n3153 ;
  assign n3170 = n32632 & n3169 ;
  assign n32633 = ~n3170 ;
  assign n3171 = n186 & n32633 ;
  assign n32634 = ~n2875 ;
  assign n2885 = n2763 & n32634 ;
  assign n2886 = n32489 & n2885 ;
  assign n3018 = n2886 & n174 ;
  assign n2887 = n2862 | n2875 ;
  assign n32635 = ~n2887 ;
  assign n3031 = n32635 & n174 ;
  assign n3032 = n2763 | n3031 ;
  assign n32636 = ~n3018 ;
  assign n3033 = n32636 & n3032 ;
  assign n3154 = n186 | n3153 ;
  assign n32637 = ~n3154 ;
  assign n3172 = n32637 & n3169 ;
  assign n3173 = n3033 | n3172 ;
  assign n32638 = ~n3171 ;
  assign n3174 = n32638 & n3173 ;
  assign n32639 = ~n3174 ;
  assign n3175 = n528 & n32639 ;
  assign n2908 = n2761 & n32516 ;
  assign n32640 = ~n2879 ;
  assign n2909 = n32640 & n2908 ;
  assign n3020 = n2909 & n174 ;
  assign n2884 = n2878 | n2879 ;
  assign n32641 = ~n2884 ;
  assign n3043 = n32641 & n174 ;
  assign n3044 = n2761 | n3043 ;
  assign n32642 = ~n3020 ;
  assign n3045 = n32642 & n3044 ;
  assign n3183 = n32621 & n3164 ;
  assign n3184 = n3030 | n3183 ;
  assign n32643 = ~n3166 ;
  assign n3185 = n32643 & n3184 ;
  assign n32644 = ~n3185 ;
  assign n3186 = n185 & n32644 ;
  assign n3187 = n32631 & n3184 ;
  assign n3188 = n3042 | n3187 ;
  assign n32645 = ~n3186 ;
  assign n3189 = n32645 & n3188 ;
  assign n32646 = ~n3189 ;
  assign n3190 = n186 & n32646 ;
  assign n3191 = n528 | n3190 ;
  assign n32647 = ~n3191 ;
  assign n3192 = n3173 & n32647 ;
  assign n3193 = n3045 | n3192 ;
  assign n32648 = ~n3175 ;
  assign n3194 = n32648 & n3193 ;
  assign n32649 = ~n3194 ;
  assign n3195 = n188 & n32649 ;
  assign n2907 = n2882 | n2895 ;
  assign n32650 = ~n2907 ;
  assign n3046 = n32650 & n174 ;
  assign n3047 = n2759 | n3046 ;
  assign n32651 = ~n2895 ;
  assign n2905 = n2759 & n32651 ;
  assign n2906 = n32505 & n2905 ;
  assign n3051 = n2906 & n174 ;
  assign n32652 = ~n3051 ;
  assign n3052 = n3047 & n32652 ;
  assign n3176 = n413 | n3175 ;
  assign n32653 = ~n3176 ;
  assign n3196 = n32653 & n3193 ;
  assign n3197 = n3052 | n3196 ;
  assign n32654 = ~n3195 ;
  assign n3198 = n32654 & n3197 ;
  assign n32655 = ~n3198 ;
  assign n3199 = n189 & n32655 ;
  assign n2900 = n2898 | n2899 ;
  assign n32656 = ~n2900 ;
  assign n3009 = n32656 & n174 ;
  assign n3010 = n2783 | n3009 ;
  assign n2924 = n2783 & n32533 ;
  assign n32657 = ~n2899 ;
  assign n2925 = n32657 & n2924 ;
  assign n3053 = n2925 & n174 ;
  assign n32658 = ~n3053 ;
  assign n3054 = n3010 & n32658 ;
  assign n3207 = n32637 & n3188 ;
  assign n3208 = n3033 | n3207 ;
  assign n32659 = ~n3190 ;
  assign n3209 = n32659 & n3208 ;
  assign n32660 = ~n3209 ;
  assign n3210 = n187 & n32660 ;
  assign n3211 = n32647 & n3208 ;
  assign n3212 = n3045 | n3211 ;
  assign n32661 = ~n3210 ;
  assign n3213 = n32661 & n3212 ;
  assign n32662 = ~n3213 ;
  assign n3214 = n413 & n32662 ;
  assign n3215 = n189 | n3214 ;
  assign n32663 = ~n3215 ;
  assign n3216 = n3197 & n32663 ;
  assign n3217 = n3054 | n3216 ;
  assign n32664 = ~n3199 ;
  assign n3218 = n32664 & n3217 ;
  assign n32665 = ~n3218 ;
  assign n3219 = n190 & n32665 ;
  assign n32666 = ~n2915 ;
  assign n2921 = n2757 & n32666 ;
  assign n2922 = n32521 & n2921 ;
  assign n2998 = n2922 & n174 ;
  assign n2923 = n2903 | n2915 ;
  assign n32667 = ~n2923 ;
  assign n3004 = n32667 & n174 ;
  assign n3005 = n2757 | n3004 ;
  assign n32668 = ~n2998 ;
  assign n3006 = n32668 & n3005 ;
  assign n3200 = n190 | n3199 ;
  assign n32669 = ~n3200 ;
  assign n3220 = n32669 & n3217 ;
  assign n3221 = n3006 | n3220 ;
  assign n32670 = ~n3219 ;
  assign n3222 = n32670 & n3221 ;
  assign n32671 = ~n3222 ;
  assign n3223 = n287 & n32671 ;
  assign n3230 = n32653 & n3212 ;
  assign n3231 = n3052 | n3230 ;
  assign n32672 = ~n3214 ;
  assign n3232 = n32672 & n3231 ;
  assign n32673 = ~n3232 ;
  assign n3233 = n189 & n32673 ;
  assign n3234 = n32663 & n3231 ;
  assign n3235 = n3054 | n3234 ;
  assign n32674 = ~n3233 ;
  assign n3236 = n32674 & n3235 ;
  assign n32675 = ~n3236 ;
  assign n3237 = n190 & n32675 ;
  assign n3238 = n287 | n3237 ;
  assign n32676 = ~n3238 ;
  assign n3239 = n3221 & n32676 ;
  assign n32677 = ~n2929 ;
  assign n3256 = n32677 & n2954 ;
  assign n32678 = ~n2919 ;
  assign n3257 = n32678 & n3256 ;
  assign n3258 = n174 & n3257 ;
  assign n2920 = n2918 | n2919 ;
  assign n32679 = ~n2920 ;
  assign n3028 = n32679 & n174 ;
  assign n3259 = n2954 | n3028 ;
  assign n32680 = ~n3258 ;
  assign n3260 = n32680 & n3259 ;
  assign n3263 = n3239 | n3260 ;
  assign n32681 = ~n3223 ;
  assign n3264 = n32681 & n3263 ;
  assign n3267 = n3243 | n3264 ;
  assign n3268 = n31336 & n3267 ;
  assign n2968 = n192 & n2967 ;
  assign n32682 = ~n2946 ;
  assign n2986 = n32682 & n174 ;
  assign n32683 = ~n2986 ;
  assign n2987 = n2964 & n32683 ;
  assign n32684 = ~n2987 ;
  assign n2988 = n2968 & n32684 ;
  assign n2942 = n2933 | n2941 ;
  assign n32685 = ~n2942 ;
  assign n2948 = n32685 & n2945 ;
  assign n2949 = n32548 & n2948 ;
  assign n3244 = n2949 & n32549 ;
  assign n3245 = n32550 & n3244 ;
  assign n3246 = n2988 | n3245 ;
  assign n3224 = n2997 & n32681 ;
  assign n3269 = n3224 & n3263 ;
  assign n3270 = n3246 | n3269 ;
  assign n173 = n3268 | n3270 ;
  assign n1306 = x86 | x87 ;
  assign n1515 = x88 | n1306 ;
  assign n3278 = x88 & n173 ;
  assign n32686 = ~n3278 ;
  assign n3279 = n1515 & n32686 ;
  assign n32687 = ~n3279 ;
  assign n3280 = n174 & n32687 ;
  assign n2937 = n1515 & n32547 ;
  assign n2938 = n32548 & n2937 ;
  assign n3254 = n2938 & n32549 ;
  assign n3255 = n32550 & n3254 ;
  assign n3291 = n3255 & n32686 ;
  assign n32688 = ~n866 ;
  assign n3299 = n32688 & n173 ;
  assign n32689 = ~x88 ;
  assign n3353 = n32689 & n173 ;
  assign n32690 = ~n3353 ;
  assign n3354 = x89 & n32690 ;
  assign n3355 = n3299 | n3354 ;
  assign n3356 = n3291 | n3355 ;
  assign n32691 = ~n3280 ;
  assign n3357 = n32691 & n3356 ;
  assign n32692 = ~n3357 ;
  assign n3358 = n2753 & n32692 ;
  assign n1697 = n32689 & n1306 ;
  assign n32693 = ~n173 ;
  assign n3349 = x88 & n32693 ;
  assign n3350 = n1697 | n3349 ;
  assign n32694 = ~n3350 ;
  assign n3351 = n174 & n32694 ;
  assign n3352 = n2753 | n3351 ;
  assign n32695 = ~n3352 ;
  assign n3362 = n32695 & n3356 ;
  assign n32696 = ~n3245 ;
  assign n3247 = n174 & n32696 ;
  assign n32697 = ~n2988 ;
  assign n3248 = n32697 & n3247 ;
  assign n32698 = ~n3269 ;
  assign n3365 = n3248 & n32698 ;
  assign n32699 = ~n3268 ;
  assign n3366 = n32699 & n3365 ;
  assign n3367 = n3299 | n3366 ;
  assign n3368 = x90 & n3367 ;
  assign n3369 = x90 | n3366 ;
  assign n3370 = n3299 | n3369 ;
  assign n32700 = ~n3368 ;
  assign n3371 = n32700 & n3370 ;
  assign n3372 = n3362 | n3371 ;
  assign n32701 = ~n3358 ;
  assign n3373 = n32701 & n3372 ;
  assign n32702 = ~n3373 ;
  assign n3374 = n2431 & n32702 ;
  assign n2985 = n2977 | n2983 ;
  assign n32703 = ~n2985 ;
  assign n3311 = n32703 & n173 ;
  assign n3312 = n3057 | n3311 ;
  assign n3062 = n32703 & n3057 ;
  assign n3318 = n3062 & n173 ;
  assign n32704 = ~n3318 ;
  assign n3319 = n3312 & n32704 ;
  assign n3359 = n2431 | n3358 ;
  assign n32705 = ~n3359 ;
  assign n3377 = n32705 & n3372 ;
  assign n3378 = n3319 | n3377 ;
  assign n32706 = ~n3374 ;
  assign n3379 = n32706 & n3378 ;
  assign n32707 = ~n3379 ;
  assign n3380 = n177 & n32707 ;
  assign n3086 = n3059 | n3085 ;
  assign n32708 = ~n3086 ;
  assign n3293 = n32708 & n173 ;
  assign n3294 = n3019 | n3293 ;
  assign n32709 = ~n3059 ;
  assign n3061 = n3019 & n32709 ;
  assign n3069 = n3061 & n32562 ;
  assign n3343 = n3069 & n173 ;
  assign n32710 = ~n3343 ;
  assign n3344 = n3294 & n32710 ;
  assign n3375 = n177 | n3374 ;
  assign n32711 = ~n3375 ;
  assign n3381 = n32711 & n3378 ;
  assign n3382 = n3344 | n3381 ;
  assign n32712 = ~n3380 ;
  assign n3383 = n32712 & n3382 ;
  assign n32713 = ~n3383 ;
  assign n3384 = n178 & n32713 ;
  assign n3084 = n3066 | n3071 ;
  assign n32714 = ~n3084 ;
  assign n3297 = n32714 & n173 ;
  assign n3298 = n3013 | n3297 ;
  assign n3068 = n3013 & n32567 ;
  assign n32715 = ~n3071 ;
  assign n3083 = n3068 & n32715 ;
  assign n3341 = n3083 & n173 ;
  assign n32716 = ~n3341 ;
  assign n3342 = n3298 & n32716 ;
  assign n3360 = n175 & n32692 ;
  assign n3281 = n175 | n3280 ;
  assign n32717 = ~n3281 ;
  assign n3364 = n32717 & n3356 ;
  assign n3394 = n3364 | n3371 ;
  assign n32718 = ~n3360 ;
  assign n3395 = n32718 & n3394 ;
  assign n32719 = ~n3395 ;
  assign n3396 = n176 & n32719 ;
  assign n3397 = n32705 & n3394 ;
  assign n3398 = n3319 | n3397 ;
  assign n32720 = ~n3396 ;
  assign n3399 = n32720 & n3398 ;
  assign n32721 = ~n3399 ;
  assign n3400 = n177 & n32721 ;
  assign n3401 = n178 | n3400 ;
  assign n32722 = ~n3401 ;
  assign n3402 = n3382 & n32722 ;
  assign n3403 = n3342 | n3402 ;
  assign n32723 = ~n3384 ;
  assign n3404 = n32723 & n3403 ;
  assign n32724 = ~n3404 ;
  assign n3405 = n179 & n32724 ;
  assign n3110 = n3075 | n3094 ;
  assign n32725 = ~n3110 ;
  assign n3289 = n32725 & n173 ;
  assign n3290 = n3024 | n3289 ;
  assign n32726 = ~n3075 ;
  assign n3081 = n3024 & n32726 ;
  assign n3082 = n32573 & n3081 ;
  assign n3300 = n3082 & n173 ;
  assign n32727 = ~n3300 ;
  assign n3301 = n3290 & n32727 ;
  assign n3385 = n1707 | n3384 ;
  assign n32728 = ~n3385 ;
  assign n3406 = n32728 & n3403 ;
  assign n3407 = n3301 | n3406 ;
  assign n32729 = ~n3405 ;
  assign n3408 = n32729 & n3407 ;
  assign n32730 = ~n3408 ;
  assign n3409 = n1487 & n32730 ;
  assign n3109 = n3078 | n3096 ;
  assign n32731 = ~n3109 ;
  assign n3304 = n32731 & n173 ;
  assign n3305 = n3027 | n3304 ;
  assign n3080 = n3027 & n32584 ;
  assign n32732 = ~n3096 ;
  assign n3108 = n3080 & n32732 ;
  assign n3309 = n3108 & n173 ;
  assign n32733 = ~n3309 ;
  assign n3310 = n3305 & n32733 ;
  assign n3417 = n32711 & n3398 ;
  assign n3418 = n3344 | n3417 ;
  assign n32734 = ~n3400 ;
  assign n3419 = n32734 & n3418 ;
  assign n32735 = ~n3419 ;
  assign n3420 = n178 & n32735 ;
  assign n3421 = n32722 & n3418 ;
  assign n3422 = n3342 | n3421 ;
  assign n32736 = ~n3420 ;
  assign n3423 = n32736 & n3422 ;
  assign n32737 = ~n3423 ;
  assign n3424 = n1707 & n32737 ;
  assign n3425 = n1487 | n3424 ;
  assign n32738 = ~n3425 ;
  assign n3426 = n3407 & n32738 ;
  assign n3427 = n3310 | n3426 ;
  assign n32739 = ~n3409 ;
  assign n3428 = n32739 & n3427 ;
  assign n32740 = ~n3428 ;
  assign n3429 = n181 & n32740 ;
  assign n3134 = n3100 | n3118 ;
  assign n32741 = ~n3134 ;
  assign n3273 = n32741 & n173 ;
  assign n3274 = n3015 | n3273 ;
  assign n32742 = ~n3100 ;
  assign n3106 = n3015 & n32742 ;
  assign n3107 = n32590 & n3106 ;
  assign n3315 = n3107 & n173 ;
  assign n32743 = ~n3315 ;
  assign n3316 = n3274 & n32743 ;
  assign n3411 = n181 | n3409 ;
  assign n32744 = ~n3411 ;
  assign n3430 = n32744 & n3427 ;
  assign n3431 = n3316 | n3430 ;
  assign n32745 = ~n3429 ;
  assign n3432 = n32745 & n3431 ;
  assign n32746 = ~n3432 ;
  assign n3433 = n182 & n32746 ;
  assign n3133 = n3103 | n3120 ;
  assign n32747 = ~n3133 ;
  assign n3320 = n32747 & n173 ;
  assign n3321 = n3002 | n3320 ;
  assign n3105 = n3002 & n32600 ;
  assign n32748 = ~n3120 ;
  assign n3132 = n3105 & n32748 ;
  assign n3332 = n3132 & n173 ;
  assign n32749 = ~n3332 ;
  assign n3333 = n3321 & n32749 ;
  assign n3441 = n32728 & n3422 ;
  assign n3442 = n3301 | n3441 ;
  assign n32750 = ~n3424 ;
  assign n3443 = n32750 & n3442 ;
  assign n32751 = ~n3443 ;
  assign n3444 = n180 & n32751 ;
  assign n3445 = n32738 & n3442 ;
  assign n3446 = n3310 | n3445 ;
  assign n32752 = ~n3444 ;
  assign n3447 = n32752 & n3446 ;
  assign n32753 = ~n3447 ;
  assign n3448 = n181 & n32753 ;
  assign n3449 = n182 | n3448 ;
  assign n32754 = ~n3449 ;
  assign n3450 = n3431 & n32754 ;
  assign n3451 = n3333 | n3450 ;
  assign n32755 = ~n3433 ;
  assign n3452 = n32755 & n3451 ;
  assign n32756 = ~n3452 ;
  assign n3453 = n183 & n32756 ;
  assign n3158 = n3124 | n3142 ;
  assign n32757 = ~n3158 ;
  assign n3302 = n32757 & n173 ;
  assign n3303 = n3037 | n3302 ;
  assign n32758 = ~n3124 ;
  assign n3130 = n3037 & n32758 ;
  assign n3131 = n32606 & n3130 ;
  assign n3325 = n3131 & n173 ;
  assign n32759 = ~n3325 ;
  assign n3326 = n3303 & n32759 ;
  assign n3434 = n183 | n3433 ;
  assign n32760 = ~n3434 ;
  assign n3454 = n32760 & n3451 ;
  assign n3455 = n3326 | n3454 ;
  assign n32761 = ~n3453 ;
  assign n3456 = n32761 & n3455 ;
  assign n32762 = ~n3456 ;
  assign n3457 = n838 & n32762 ;
  assign n3128 = n3039 & n32616 ;
  assign n32763 = ~n3144 ;
  assign n3156 = n3128 & n32763 ;
  assign n3317 = n3156 & n173 ;
  assign n3157 = n3127 | n3144 ;
  assign n32764 = ~n3157 ;
  assign n3329 = n32764 & n173 ;
  assign n3330 = n3039 | n3329 ;
  assign n32765 = ~n3317 ;
  assign n3331 = n32765 & n3330 ;
  assign n3465 = n32744 & n3446 ;
  assign n3466 = n3316 | n3465 ;
  assign n32766 = ~n3448 ;
  assign n3467 = n32766 & n3466 ;
  assign n32767 = ~n3467 ;
  assign n3468 = n182 & n32767 ;
  assign n3469 = n32754 & n3466 ;
  assign n3470 = n3333 | n3469 ;
  assign n32768 = ~n3468 ;
  assign n3471 = n32768 & n3470 ;
  assign n32769 = ~n3471 ;
  assign n3472 = n996 & n32769 ;
  assign n3473 = n838 | n3472 ;
  assign n32770 = ~n3473 ;
  assign n3474 = n3455 & n32770 ;
  assign n3475 = n3331 | n3474 ;
  assign n32771 = ~n3457 ;
  assign n3476 = n32771 & n3475 ;
  assign n32772 = ~n3476 ;
  assign n3477 = n185 & n32772 ;
  assign n32773 = ~n3148 ;
  assign n3149 = n3030 & n32773 ;
  assign n3150 = n32622 & n3149 ;
  assign n3272 = n3150 & n173 ;
  assign n3182 = n3148 | n3166 ;
  assign n32774 = ~n3182 ;
  assign n3275 = n32774 & n173 ;
  assign n3276 = n3030 | n3275 ;
  assign n32775 = ~n3272 ;
  assign n3277 = n32775 & n3276 ;
  assign n3458 = n185 | n3457 ;
  assign n32776 = ~n3458 ;
  assign n3478 = n32776 & n3475 ;
  assign n3479 = n3277 | n3478 ;
  assign n32777 = ~n3477 ;
  assign n3480 = n32777 & n3479 ;
  assign n32778 = ~n3480 ;
  assign n3481 = n186 & n32778 ;
  assign n3155 = n3042 & n32632 ;
  assign n32779 = ~n3168 ;
  assign n3180 = n3155 & n32779 ;
  assign n3288 = n3180 & n173 ;
  assign n3181 = n3153 | n3168 ;
  assign n32780 = ~n3181 ;
  assign n3306 = n32780 & n173 ;
  assign n3307 = n3042 | n3306 ;
  assign n32781 = ~n3288 ;
  assign n3308 = n32781 & n3307 ;
  assign n3489 = n32760 & n3470 ;
  assign n3490 = n3326 | n3489 ;
  assign n32782 = ~n3472 ;
  assign n3491 = n32782 & n3490 ;
  assign n32783 = ~n3491 ;
  assign n3492 = n184 & n32783 ;
  assign n3493 = n32770 & n3490 ;
  assign n3494 = n3331 | n3493 ;
  assign n32784 = ~n3492 ;
  assign n3495 = n32784 & n3494 ;
  assign n32785 = ~n3495 ;
  assign n3496 = n185 & n32785 ;
  assign n3497 = n186 | n3496 ;
  assign n32786 = ~n3497 ;
  assign n3498 = n3479 & n32786 ;
  assign n3499 = n3308 | n3498 ;
  assign n32787 = ~n3481 ;
  assign n3500 = n32787 & n3499 ;
  assign n32788 = ~n3500 ;
  assign n3501 = n187 & n32788 ;
  assign n3206 = n3172 | n3190 ;
  assign n32789 = ~n3206 ;
  assign n3313 = n32789 & n173 ;
  assign n3314 = n3033 | n3313 ;
  assign n32790 = ~n3172 ;
  assign n3178 = n3033 & n32790 ;
  assign n3179 = n32638 & n3178 ;
  assign n3336 = n3179 & n173 ;
  assign n32791 = ~n3336 ;
  assign n3337 = n3314 & n32791 ;
  assign n3483 = n528 | n3481 ;
  assign n32792 = ~n3483 ;
  assign n3502 = n32792 & n3499 ;
  assign n3503 = n3337 | n3502 ;
  assign n32793 = ~n3501 ;
  assign n3504 = n32793 & n3503 ;
  assign n32794 = ~n3504 ;
  assign n3505 = n413 & n32794 ;
  assign n3205 = n3175 | n3192 ;
  assign n32795 = ~n3205 ;
  assign n3327 = n32795 & n173 ;
  assign n3328 = n3045 | n3327 ;
  assign n3177 = n3045 & n32648 ;
  assign n32796 = ~n3192 ;
  assign n3204 = n3177 & n32796 ;
  assign n3334 = n3204 & n173 ;
  assign n32797 = ~n3334 ;
  assign n3335 = n3328 & n32797 ;
  assign n3513 = n32776 & n3494 ;
  assign n3514 = n3277 | n3513 ;
  assign n32798 = ~n3496 ;
  assign n3515 = n32798 & n3514 ;
  assign n32799 = ~n3515 ;
  assign n3516 = n186 & n32799 ;
  assign n3517 = n32786 & n3514 ;
  assign n3518 = n3308 | n3517 ;
  assign n32800 = ~n3516 ;
  assign n3519 = n32800 & n3518 ;
  assign n32801 = ~n3519 ;
  assign n3520 = n528 & n32801 ;
  assign n3521 = n413 | n3520 ;
  assign n32802 = ~n3521 ;
  assign n3522 = n3503 & n32802 ;
  assign n3523 = n3335 | n3522 ;
  assign n32803 = ~n3505 ;
  assign n3524 = n32803 & n3523 ;
  assign n32804 = ~n3524 ;
  assign n3525 = n189 & n32804 ;
  assign n32805 = ~n3196 ;
  assign n3202 = n3052 & n32805 ;
  assign n3203 = n32654 & n3202 ;
  assign n3287 = n3203 & n173 ;
  assign n3229 = n3196 | n3214 ;
  assign n32806 = ~n3229 ;
  assign n3338 = n32806 & n173 ;
  assign n3339 = n3052 | n3338 ;
  assign n32807 = ~n3287 ;
  assign n3340 = n32807 & n3339 ;
  assign n3506 = n189 | n3505 ;
  assign n32808 = ~n3506 ;
  assign n3526 = n32808 & n3523 ;
  assign n3527 = n3340 | n3526 ;
  assign n32809 = ~n3525 ;
  assign n3528 = n32809 & n3527 ;
  assign n32810 = ~n3528 ;
  assign n3529 = n190 & n32810 ;
  assign n3228 = n3199 | n3216 ;
  assign n32811 = ~n3228 ;
  assign n3285 = n32811 & n173 ;
  assign n3286 = n3054 | n3285 ;
  assign n3201 = n3054 & n32664 ;
  assign n32812 = ~n3216 ;
  assign n3227 = n3201 & n32812 ;
  assign n3295 = n3227 & n173 ;
  assign n32813 = ~n3295 ;
  assign n3296 = n3286 & n32813 ;
  assign n3535 = n32792 & n3518 ;
  assign n3536 = n3337 | n3535 ;
  assign n32814 = ~n3520 ;
  assign n3537 = n32814 & n3536 ;
  assign n32815 = ~n3537 ;
  assign n3538 = n188 & n32815 ;
  assign n3539 = n32802 & n3536 ;
  assign n3540 = n3335 | n3539 ;
  assign n32816 = ~n3538 ;
  assign n3541 = n32816 & n3540 ;
  assign n32817 = ~n3541 ;
  assign n3542 = n189 & n32817 ;
  assign n3543 = n190 | n3542 ;
  assign n32818 = ~n3543 ;
  assign n3544 = n3527 & n32818 ;
  assign n3545 = n3296 | n3544 ;
  assign n32819 = ~n3529 ;
  assign n3550 = n32819 & n3545 ;
  assign n32820 = ~n3550 ;
  assign n3551 = n191 & n32820 ;
  assign n32821 = ~n3220 ;
  assign n3225 = n3006 & n32821 ;
  assign n3226 = n32670 & n3225 ;
  assign n3284 = n3226 & n173 ;
  assign n3241 = n3220 | n3237 ;
  assign n32822 = ~n3241 ;
  assign n3322 = n32822 & n173 ;
  assign n3323 = n3006 | n3322 ;
  assign n32823 = ~n3284 ;
  assign n3324 = n32823 & n3323 ;
  assign n3532 = n191 | n3529 ;
  assign n32824 = ~n3532 ;
  assign n3553 = n32824 & n3545 ;
  assign n3554 = n3324 | n3553 ;
  assign n32825 = ~n3551 ;
  assign n3555 = n32825 & n3554 ;
  assign n3265 = n2997 | n3264 ;
  assign n32826 = ~n3265 ;
  assign n3345 = n32826 & n173 ;
  assign n3563 = n3269 | n3345 ;
  assign n3261 = n32681 & n3260 ;
  assign n32827 = ~n3239 ;
  assign n3262 = n32827 & n3261 ;
  assign n3283 = n3262 & n173 ;
  assign n3240 = n3223 | n3239 ;
  assign n32828 = ~n3240 ;
  assign n3282 = n32828 & n173 ;
  assign n3574 = n3260 | n3282 ;
  assign n32829 = ~n3283 ;
  assign n3575 = n32829 & n3574 ;
  assign n3576 = n3563 | n3575 ;
  assign n3577 = n3555 | n3576 ;
  assign n3578 = n31336 & n3577 ;
  assign n3266 = n192 & n3265 ;
  assign n32830 = ~n2997 ;
  assign n3346 = n32830 & n173 ;
  assign n32831 = ~n3346 ;
  assign n3347 = n3264 & n32831 ;
  assign n32832 = ~n3347 ;
  assign n3348 = n3266 & n32832 ;
  assign n3249 = n2996 | n3245 ;
  assign n32833 = ~n3249 ;
  assign n3250 = n2994 & n32833 ;
  assign n3251 = n32697 & n3250 ;
  assign n3564 = n3251 & n32698 ;
  assign n3565 = n32699 & n3564 ;
  assign n3566 = n3348 | n3565 ;
  assign n3581 = n32825 & n3575 ;
  assign n3582 = n3554 & n3581 ;
  assign n3583 = n3566 | n3582 ;
  assign n172 = n3578 | n3583 ;
  assign n3530 = n287 | n3529 ;
  assign n32834 = ~n3530 ;
  assign n3546 = n32834 & n3545 ;
  assign n3547 = n3324 | n3546 ;
  assign n3552 = n3547 & n32825 ;
  assign n3579 = n3552 | n3576 ;
  assign n3580 = n31336 & n3579 ;
  assign n3629 = n3547 & n3581 ;
  assign n3630 = n3566 | n3629 ;
  assign n3631 = n3580 | n3630 ;
  assign n32835 = ~n1306 ;
  assign n3638 = n32835 & n3631 ;
  assign n32836 = ~x86 ;
  assign n3639 = n32836 & n3631 ;
  assign n32837 = ~n3639 ;
  assign n3640 = x87 & n32837 ;
  assign n3641 = n3638 | n3640 ;
  assign n1906 = x84 | x85 ;
  assign n2163 = x86 | n1906 ;
  assign n3252 = n2163 & n32696 ;
  assign n3253 = n32697 & n3252 ;
  assign n3572 = n3253 & n32698 ;
  assign n3573 = n32699 & n3572 ;
  assign n3646 = x86 & n3631 ;
  assign n32838 = ~n3646 ;
  assign n3647 = n3573 & n32838 ;
  assign n3648 = n3641 | n3647 ;
  assign n2494 = n32836 & n1906 ;
  assign n32839 = ~n3631 ;
  assign n3652 = x86 & n32839 ;
  assign n3653 = n2494 | n3652 ;
  assign n32840 = ~n3653 ;
  assign n3654 = n173 & n32840 ;
  assign n32841 = ~n3654 ;
  assign n3655 = n3648 & n32841 ;
  assign n32842 = ~n3655 ;
  assign n3656 = n174 & n32842 ;
  assign n3607 = x86 & n172 ;
  assign n32843 = ~n3607 ;
  assign n3608 = n2163 & n32843 ;
  assign n32844 = ~n3608 ;
  assign n3609 = n173 & n32844 ;
  assign n3610 = n174 | n3609 ;
  assign n32845 = ~n3610 ;
  assign n3649 = n32845 & n3648 ;
  assign n32846 = ~n3565 ;
  assign n3567 = n173 & n32846 ;
  assign n32847 = ~n3348 ;
  assign n3568 = n32847 & n3567 ;
  assign n32848 = ~n3629 ;
  assign n3689 = n3568 & n32848 ;
  assign n32849 = ~n3578 ;
  assign n3690 = n32849 & n3689 ;
  assign n3691 = n3638 | n3690 ;
  assign n3692 = x88 & n3691 ;
  assign n3693 = x88 | n3690 ;
  assign n3694 = n3638 | n3693 ;
  assign n32850 = ~n3692 ;
  assign n3695 = n32850 & n3694 ;
  assign n3696 = n3649 | n3695 ;
  assign n32851 = ~n3656 ;
  assign n3697 = n32851 & n3696 ;
  assign n32852 = ~n3697 ;
  assign n3698 = n175 & n32852 ;
  assign n3292 = n3280 | n3291 ;
  assign n32853 = ~n3292 ;
  assign n3361 = n32853 & n3355 ;
  assign n3597 = n3361 & n172 ;
  assign n3602 = n32853 & n172 ;
  assign n3603 = n3355 | n3602 ;
  assign n32854 = ~n3597 ;
  assign n3604 = n32854 & n3603 ;
  assign n3657 = n175 | n3656 ;
  assign n3660 = n174 | n3654 ;
  assign n32855 = ~n3660 ;
  assign n3661 = n3648 & n32855 ;
  assign n3704 = n3661 | n3695 ;
  assign n32856 = ~n3657 ;
  assign n3705 = n32856 & n3704 ;
  assign n3708 = n3604 | n3705 ;
  assign n32857 = ~n3698 ;
  assign n3709 = n32857 & n3708 ;
  assign n32858 = ~n3709 ;
  assign n3710 = n176 & n32858 ;
  assign n3363 = n3360 | n3362 ;
  assign n32859 = ~n3363 ;
  assign n3595 = n32859 & n172 ;
  assign n3596 = n3371 | n3595 ;
  assign n32860 = ~n3362 ;
  assign n3392 = n32860 & n3371 ;
  assign n3393 = n32718 & n3392 ;
  assign n3667 = n3393 & n3631 ;
  assign n32861 = ~n3667 ;
  assign n3668 = n3596 & n32861 ;
  assign n3700 = n2753 & n32852 ;
  assign n3701 = n2431 | n3700 ;
  assign n32862 = ~n3701 ;
  assign n3712 = n32862 & n3708 ;
  assign n3713 = n3668 | n3712 ;
  assign n32863 = ~n3710 ;
  assign n3714 = n32863 & n3713 ;
  assign n32864 = ~n3714 ;
  assign n3715 = n177 & n32864 ;
  assign n3391 = n3374 | n3377 ;
  assign n32865 = ~n3391 ;
  assign n3605 = n32865 & n172 ;
  assign n3606 = n3319 | n3605 ;
  assign n3376 = n3319 & n32706 ;
  assign n32866 = ~n3377 ;
  assign n3390 = n3376 & n32866 ;
  assign n3650 = n3390 & n3631 ;
  assign n32867 = ~n3650 ;
  assign n3651 = n3606 & n32867 ;
  assign n3711 = n177 | n3710 ;
  assign n32868 = ~n3711 ;
  assign n3718 = n32868 & n3713 ;
  assign n3719 = n3651 | n3718 ;
  assign n32869 = ~n3715 ;
  assign n3720 = n32869 & n3719 ;
  assign n32870 = ~n3720 ;
  assign n3721 = n178 & n32870 ;
  assign n3389 = n3380 | n3381 ;
  assign n32871 = ~n3389 ;
  assign n3623 = n32871 & n172 ;
  assign n3624 = n3344 | n3623 ;
  assign n32872 = ~n3381 ;
  assign n3387 = n3344 & n32872 ;
  assign n3388 = n32712 & n3387 ;
  assign n3663 = n3388 & n3631 ;
  assign n32873 = ~n3663 ;
  assign n3664 = n3624 & n32873 ;
  assign n3716 = n178 | n3715 ;
  assign n32874 = ~n3716 ;
  assign n3722 = n32874 & n3719 ;
  assign n3723 = n3664 | n3722 ;
  assign n32875 = ~n3721 ;
  assign n3724 = n32875 & n3723 ;
  assign n32876 = ~n3724 ;
  assign n3725 = n1707 & n32876 ;
  assign n3416 = n3384 | n3402 ;
  assign n32877 = ~n3416 ;
  assign n3591 = n32877 & n172 ;
  assign n3592 = n3342 | n3591 ;
  assign n3386 = n3342 & n32723 ;
  assign n32878 = ~n3402 ;
  assign n3415 = n3386 & n32878 ;
  assign n3669 = n3415 & n3631 ;
  assign n32879 = ~n3669 ;
  assign n3670 = n3592 & n32879 ;
  assign n3728 = n1707 | n3721 ;
  assign n32880 = ~n3728 ;
  assign n3729 = n3723 & n32880 ;
  assign n3730 = n3670 | n3729 ;
  assign n32881 = ~n3725 ;
  assign n3731 = n32881 & n3730 ;
  assign n32882 = ~n3731 ;
  assign n3732 = n180 & n32882 ;
  assign n3414 = n3405 | n3406 ;
  assign n32883 = ~n3414 ;
  assign n3600 = n32883 & n172 ;
  assign n3601 = n3301 | n3600 ;
  assign n32884 = ~n3406 ;
  assign n3412 = n3301 & n32884 ;
  assign n3413 = n32729 & n3412 ;
  assign n3632 = n3413 & n3631 ;
  assign n32885 = ~n3632 ;
  assign n3633 = n3601 & n32885 ;
  assign n3726 = n1487 | n3725 ;
  assign n32886 = ~n3726 ;
  assign n3733 = n32886 & n3730 ;
  assign n3734 = n3633 | n3733 ;
  assign n32887 = ~n3732 ;
  assign n3735 = n32887 & n3734 ;
  assign n32888 = ~n3735 ;
  assign n3736 = n181 & n32888 ;
  assign n3440 = n3409 | n3426 ;
  assign n32889 = ~n3440 ;
  assign n3598 = n32889 & n172 ;
  assign n3599 = n3310 | n3598 ;
  assign n3410 = n3310 & n32739 ;
  assign n32890 = ~n3426 ;
  assign n3439 = n3410 & n32890 ;
  assign n3634 = n3439 & n3631 ;
  assign n32891 = ~n3634 ;
  assign n3635 = n3599 & n32891 ;
  assign n3739 = n179 & n32876 ;
  assign n32892 = ~n3739 ;
  assign n3740 = n3730 & n32892 ;
  assign n32893 = ~n3740 ;
  assign n3741 = n1487 & n32893 ;
  assign n3742 = n181 | n3741 ;
  assign n32894 = ~n3742 ;
  assign n3743 = n3734 & n32894 ;
  assign n3744 = n3635 | n3743 ;
  assign n32895 = ~n3736 ;
  assign n3745 = n32895 & n3744 ;
  assign n32896 = ~n3745 ;
  assign n3746 = n182 & n32896 ;
  assign n3438 = n3429 | n3430 ;
  assign n32897 = ~n3438 ;
  assign n3619 = n32897 & n172 ;
  assign n3620 = n3316 | n3619 ;
  assign n32898 = ~n3430 ;
  assign n3436 = n3316 & n32898 ;
  assign n3437 = n32745 & n3436 ;
  assign n3671 = n3437 & n3631 ;
  assign n32899 = ~n3671 ;
  assign n3672 = n3620 & n32899 ;
  assign n3737 = n182 | n3736 ;
  assign n32900 = ~n3737 ;
  assign n3747 = n32900 & n3744 ;
  assign n3748 = n3672 | n3747 ;
  assign n32901 = ~n3746 ;
  assign n3749 = n32901 & n3748 ;
  assign n32902 = ~n3749 ;
  assign n3750 = n996 & n32902 ;
  assign n3464 = n3433 | n3450 ;
  assign n32903 = ~n3464 ;
  assign n3593 = n32903 & n172 ;
  assign n3594 = n3333 | n3593 ;
  assign n3435 = n3333 & n32755 ;
  assign n32904 = ~n3450 ;
  assign n3463 = n3435 & n32904 ;
  assign n3673 = n3463 & n3631 ;
  assign n32905 = ~n3673 ;
  assign n3674 = n3594 & n32905 ;
  assign n32906 = ~n3741 ;
  assign n3753 = n3734 & n32906 ;
  assign n32907 = ~n3753 ;
  assign n3754 = n181 & n32907 ;
  assign n32908 = ~n3754 ;
  assign n3755 = n3744 & n32908 ;
  assign n32909 = ~n3755 ;
  assign n3756 = n182 & n32909 ;
  assign n3757 = n183 | n3756 ;
  assign n32910 = ~n3757 ;
  assign n3758 = n3748 & n32910 ;
  assign n3759 = n3674 | n3758 ;
  assign n32911 = ~n3750 ;
  assign n3760 = n32911 & n3759 ;
  assign n32912 = ~n3760 ;
  assign n3761 = n184 & n32912 ;
  assign n3462 = n3453 | n3454 ;
  assign n32913 = ~n3462 ;
  assign n3589 = n32913 & n172 ;
  assign n3590 = n3326 | n3589 ;
  assign n32914 = ~n3454 ;
  assign n3460 = n3326 & n32914 ;
  assign n3461 = n32761 & n3460 ;
  assign n3679 = n3461 & n3631 ;
  assign n32915 = ~n3679 ;
  assign n3680 = n3590 & n32915 ;
  assign n3751 = n838 | n3750 ;
  assign n32916 = ~n3751 ;
  assign n3762 = n32916 & n3759 ;
  assign n3763 = n3680 | n3762 ;
  assign n32917 = ~n3761 ;
  assign n3764 = n32917 & n3763 ;
  assign n32918 = ~n3764 ;
  assign n3765 = n185 & n32918 ;
  assign n3488 = n3457 | n3474 ;
  assign n32919 = ~n3488 ;
  assign n3587 = n32919 & n172 ;
  assign n3588 = n3331 | n3587 ;
  assign n3459 = n3331 & n32771 ;
  assign n32920 = ~n3474 ;
  assign n3487 = n3459 & n32920 ;
  assign n3675 = n3487 & n3631 ;
  assign n32921 = ~n3675 ;
  assign n3676 = n3588 & n32921 ;
  assign n32922 = ~n3756 ;
  assign n3768 = n3748 & n32922 ;
  assign n32923 = ~n3768 ;
  assign n3769 = n183 & n32923 ;
  assign n32924 = ~n3769 ;
  assign n3772 = n3759 & n32924 ;
  assign n32925 = ~n3772 ;
  assign n3773 = n838 & n32925 ;
  assign n3774 = n185 | n3773 ;
  assign n32926 = ~n3774 ;
  assign n3775 = n3763 & n32926 ;
  assign n3776 = n3676 | n3775 ;
  assign n32927 = ~n3765 ;
  assign n3777 = n32927 & n3776 ;
  assign n32928 = ~n3777 ;
  assign n3778 = n186 & n32928 ;
  assign n3486 = n3477 | n3478 ;
  assign n32929 = ~n3486 ;
  assign n3625 = n32929 & n172 ;
  assign n3626 = n3277 | n3625 ;
  assign n32930 = ~n3478 ;
  assign n3484 = n3277 & n32930 ;
  assign n3485 = n32777 & n3484 ;
  assign n3642 = n3485 & n3631 ;
  assign n32931 = ~n3642 ;
  assign n3643 = n3626 & n32931 ;
  assign n3766 = n186 | n3765 ;
  assign n32932 = ~n3766 ;
  assign n3779 = n32932 & n3776 ;
  assign n3780 = n3643 | n3779 ;
  assign n32933 = ~n3778 ;
  assign n3781 = n32933 & n3780 ;
  assign n32934 = ~n3781 ;
  assign n3782 = n528 & n32934 ;
  assign n3512 = n3481 | n3498 ;
  assign n32935 = ~n3512 ;
  assign n3613 = n32935 & n172 ;
  assign n3614 = n3308 | n3613 ;
  assign n3482 = n3308 & n32787 ;
  assign n32936 = ~n3498 ;
  assign n3511 = n3482 & n32936 ;
  assign n3644 = n3511 & n3631 ;
  assign n32937 = ~n3644 ;
  assign n3645 = n3614 & n32937 ;
  assign n32938 = ~n3773 ;
  assign n3785 = n3763 & n32938 ;
  assign n32939 = ~n3785 ;
  assign n3786 = n185 & n32939 ;
  assign n32940 = ~n3786 ;
  assign n3787 = n3776 & n32940 ;
  assign n32941 = ~n3787 ;
  assign n3788 = n186 & n32941 ;
  assign n3789 = n528 | n3788 ;
  assign n32942 = ~n3789 ;
  assign n3790 = n3780 & n32942 ;
  assign n3791 = n3645 | n3790 ;
  assign n32943 = ~n3782 ;
  assign n3792 = n32943 & n3791 ;
  assign n32944 = ~n3792 ;
  assign n3793 = n188 & n32944 ;
  assign n3510 = n3501 | n3502 ;
  assign n32945 = ~n3510 ;
  assign n3615 = n32945 & n172 ;
  assign n3616 = n3337 | n3615 ;
  assign n32946 = ~n3502 ;
  assign n3508 = n3337 & n32946 ;
  assign n3509 = n32793 & n3508 ;
  assign n3636 = n3509 & n3631 ;
  assign n32947 = ~n3636 ;
  assign n3637 = n3616 & n32947 ;
  assign n3783 = n413 | n3782 ;
  assign n32948 = ~n3783 ;
  assign n3794 = n32948 & n3791 ;
  assign n3795 = n3637 | n3794 ;
  assign n32949 = ~n3793 ;
  assign n3796 = n32949 & n3795 ;
  assign n32950 = ~n3796 ;
  assign n3797 = n189 & n32950 ;
  assign n3534 = n3505 | n3522 ;
  assign n32951 = ~n3534 ;
  assign n3617 = n32951 & n172 ;
  assign n3618 = n3335 | n3617 ;
  assign n3507 = n3335 & n32803 ;
  assign n32952 = ~n3522 ;
  assign n3533 = n3507 & n32952 ;
  assign n3665 = n3533 & n3631 ;
  assign n32953 = ~n3665 ;
  assign n3666 = n3618 & n32953 ;
  assign n32954 = ~n3788 ;
  assign n3800 = n3780 & n32954 ;
  assign n32955 = ~n3800 ;
  assign n3801 = n187 & n32955 ;
  assign n32956 = ~n3801 ;
  assign n3802 = n3791 & n32956 ;
  assign n32957 = ~n3802 ;
  assign n3803 = n413 & n32957 ;
  assign n3804 = n189 | n3803 ;
  assign n32958 = ~n3804 ;
  assign n3805 = n3795 & n32958 ;
  assign n3806 = n3666 | n3805 ;
  assign n32959 = ~n3797 ;
  assign n3807 = n32959 & n3806 ;
  assign n32960 = ~n3807 ;
  assign n3808 = n190 & n32960 ;
  assign n3559 = n32808 & n3540 ;
  assign n3562 = n3525 | n3559 ;
  assign n32961 = ~n3562 ;
  assign n3585 = n32961 & n172 ;
  assign n3586 = n3340 | n3585 ;
  assign n32962 = ~n3559 ;
  assign n3560 = n3340 & n32962 ;
  assign n3561 = n32809 & n3560 ;
  assign n3681 = n3561 & n3631 ;
  assign n32963 = ~n3681 ;
  assign n3682 = n3586 & n32963 ;
  assign n3798 = n190 | n3797 ;
  assign n32964 = ~n3798 ;
  assign n3809 = n32964 & n3806 ;
  assign n3810 = n3682 | n3809 ;
  assign n32965 = ~n3808 ;
  assign n3811 = n32965 & n3810 ;
  assign n32966 = ~n3811 ;
  assign n3812 = n287 & n32966 ;
  assign n3549 = n3529 | n3544 ;
  assign n32967 = ~n3549 ;
  assign n3621 = n32967 & n172 ;
  assign n3622 = n3296 | n3621 ;
  assign n3531 = n3296 & n32819 ;
  assign n32968 = ~n3544 ;
  assign n3548 = n3531 & n32968 ;
  assign n3677 = n3548 & n3631 ;
  assign n32969 = ~n3677 ;
  assign n3678 = n3622 & n32969 ;
  assign n32970 = ~n3803 ;
  assign n3815 = n3795 & n32970 ;
  assign n32971 = ~n3815 ;
  assign n3816 = n189 & n32971 ;
  assign n32972 = ~n3816 ;
  assign n3817 = n3806 & n32972 ;
  assign n32973 = ~n3817 ;
  assign n3818 = n190 & n32973 ;
  assign n3819 = n287 | n3818 ;
  assign n32974 = ~n3819 ;
  assign n3820 = n3810 & n32974 ;
  assign n3821 = n3678 | n3820 ;
  assign n32975 = ~n3812 ;
  assign n3822 = n32975 & n3821 ;
  assign n3558 = n3551 | n3553 ;
  assign n32976 = ~n3558 ;
  assign n3611 = n32976 & n172 ;
  assign n3612 = n3324 | n3611 ;
  assign n32977 = ~n3553 ;
  assign n3556 = n3324 & n32977 ;
  assign n3557 = n32825 & n3556 ;
  assign n3683 = n3557 & n3631 ;
  assign n32978 = ~n3683 ;
  assign n3684 = n3612 & n32978 ;
  assign n3627 = n3552 | n3575 ;
  assign n32979 = ~n3627 ;
  assign n3685 = n32979 & n3631 ;
  assign n3871 = n3629 | n3685 ;
  assign n3872 = n3684 | n3871 ;
  assign n3875 = n3822 | n3872 ;
  assign n3876 = n31336 & n3875 ;
  assign n3813 = n3684 & n32975 ;
  assign n3823 = n3813 & n3821 ;
  assign n3628 = n192 & n3627 ;
  assign n32980 = ~n3575 ;
  assign n3686 = n32980 & n3631 ;
  assign n32981 = ~n3686 ;
  assign n3687 = n3552 & n32981 ;
  assign n32982 = ~n3687 ;
  assign n3688 = n3628 & n32982 ;
  assign n3569 = n3283 | n3565 ;
  assign n32983 = ~n3569 ;
  assign n3879 = n32983 & n3574 ;
  assign n3880 = n32847 & n3879 ;
  assign n3881 = n32848 & n3880 ;
  assign n3882 = n32849 & n3881 ;
  assign n3883 = n3688 | n3882 ;
  assign n3939 = n3823 | n3883 ;
  assign n3940 = n3876 | n3939 ;
  assign n3826 = n191 | n3818 ;
  assign n32984 = ~n3826 ;
  assign n3827 = n3810 & n32984 ;
  assign n3829 = n3812 | n3827 ;
  assign n32985 = ~n3818 ;
  assign n3830 = n3810 & n32985 ;
  assign n32986 = ~n3830 ;
  assign n3831 = n191 & n32986 ;
  assign n3832 = n3678 | n3827 ;
  assign n32987 = ~n3831 ;
  assign n3833 = n32987 & n3832 ;
  assign n3873 = n3833 | n3872 ;
  assign n3874 = n31336 & n3873 ;
  assign n3834 = n3813 & n3832 ;
  assign n3884 = n3834 | n3883 ;
  assign n171 = n3874 | n3884 ;
  assign n32988 = ~n3829 ;
  assign n3904 = n32988 & n171 ;
  assign n3905 = n3678 | n3904 ;
  assign n3814 = n3678 & n32975 ;
  assign n32989 = ~n3827 ;
  assign n3828 = n3814 & n32989 ;
  assign n3949 = n3828 & n3940 ;
  assign n32990 = ~n3949 ;
  assign n3950 = n3905 & n32990 ;
  assign n3824 = n3684 | n3822 ;
  assign n32991 = ~n3824 ;
  assign n3957 = n32991 & n3940 ;
  assign n3958 = n3823 | n3957 ;
  assign n3959 = n3950 | n3958 ;
  assign n2714 = x82 | x83 ;
  assign n32992 = ~x84 ;
  assign n3271 = n32992 & n2714 ;
  assign n32993 = ~n3940 ;
  assign n3953 = x84 & n32993 ;
  assign n3954 = n3271 | n3953 ;
  assign n32994 = ~n3954 ;
  assign n3955 = n3631 & n32994 ;
  assign n2974 = x84 | n2714 ;
  assign n3570 = n2974 & n32846 ;
  assign n3571 = n32847 & n3570 ;
  assign n3877 = n3571 & n32848 ;
  assign n3878 = n32849 & n3877 ;
  assign n3960 = x84 & n3940 ;
  assign n32995 = ~n3960 ;
  assign n3961 = n3878 & n32995 ;
  assign n3963 = n32992 & n3940 ;
  assign n32996 = ~n3963 ;
  assign n3964 = x85 & n32996 ;
  assign n32997 = ~n1906 ;
  assign n3965 = n32997 & n3940 ;
  assign n3966 = n3964 | n3965 ;
  assign n3968 = n3961 | n3966 ;
  assign n32998 = ~n3955 ;
  assign n3969 = n32998 & n3968 ;
  assign n32999 = ~n3969 ;
  assign n3970 = n173 & n32999 ;
  assign n3935 = x84 & n171 ;
  assign n33000 = ~n3935 ;
  assign n3936 = n2974 & n33000 ;
  assign n33001 = ~n3936 ;
  assign n3937 = n172 & n33001 ;
  assign n3938 = n173 | n3937 ;
  assign n33002 = ~n3938 ;
  assign n3972 = n33002 & n3968 ;
  assign n33003 = ~n3882 ;
  assign n3993 = n3631 & n33003 ;
  assign n33004 = ~n3688 ;
  assign n3994 = n33004 & n3993 ;
  assign n33005 = ~n3823 ;
  assign n3995 = n33005 & n3994 ;
  assign n33006 = ~n3876 ;
  assign n3996 = n33006 & n3995 ;
  assign n3997 = n3965 | n3996 ;
  assign n3998 = x86 & n3997 ;
  assign n3999 = x86 | n3996 ;
  assign n4000 = n3965 | n3999 ;
  assign n33007 = ~n3998 ;
  assign n4001 = n33007 & n4000 ;
  assign n4002 = n3972 | n4001 ;
  assign n33008 = ~n3970 ;
  assign n4003 = n33008 & n4002 ;
  assign n33009 = ~n4003 ;
  assign n4004 = n174 & n33009 ;
  assign n3658 = n3647 | n3654 ;
  assign n33010 = ~n3658 ;
  assign n3886 = n33010 & n171 ;
  assign n3887 = n3641 | n3886 ;
  assign n3659 = n3641 & n33010 ;
  assign n3975 = n3659 & n3940 ;
  assign n33011 = ~n3975 ;
  assign n3976 = n3887 & n33011 ;
  assign n3971 = n174 | n3970 ;
  assign n3956 = n173 | n3955 ;
  assign n33012 = ~n3956 ;
  assign n3973 = n33012 & n3968 ;
  assign n4009 = n3973 | n4001 ;
  assign n33013 = ~n3971 ;
  assign n4010 = n33013 & n4009 ;
  assign n4011 = n3976 | n4010 ;
  assign n33014 = ~n4004 ;
  assign n4012 = n33014 & n4011 ;
  assign n33015 = ~n4012 ;
  assign n4013 = n2753 & n33015 ;
  assign n3662 = n3656 | n3661 ;
  assign n33016 = ~n3662 ;
  assign n3888 = n33016 & n171 ;
  assign n3889 = n3695 | n3888 ;
  assign n33017 = ~n3661 ;
  assign n3702 = n33017 & n3695 ;
  assign n3703 = n32851 & n3702 ;
  assign n3977 = n3703 & n3940 ;
  assign n33018 = ~n3977 ;
  assign n3978 = n3889 & n33018 ;
  assign n4006 = n2753 | n4004 ;
  assign n33019 = ~n4006 ;
  assign n4015 = n33019 & n4011 ;
  assign n4016 = n3978 | n4015 ;
  assign n33020 = ~n4013 ;
  assign n4017 = n33020 & n4016 ;
  assign n33021 = ~n4017 ;
  assign n4018 = n176 & n33021 ;
  assign n3707 = n3698 | n3705 ;
  assign n33022 = ~n3707 ;
  assign n3923 = n33022 & n171 ;
  assign n3924 = n3604 | n3923 ;
  assign n3699 = n3604 & n32857 ;
  assign n33023 = ~n3705 ;
  assign n3706 = n3699 & n33023 ;
  assign n3979 = n3706 & n3940 ;
  assign n33024 = ~n3979 ;
  assign n3980 = n3924 & n33024 ;
  assign n4014 = n2431 | n4013 ;
  assign n33025 = ~n4014 ;
  assign n4019 = n33025 & n4016 ;
  assign n4020 = n3980 | n4019 ;
  assign n33026 = ~n4018 ;
  assign n4021 = n33026 & n4020 ;
  assign n33027 = ~n4021 ;
  assign n4022 = n177 & n33027 ;
  assign n3868 = n3710 | n3712 ;
  assign n33028 = ~n3868 ;
  assign n3930 = n33028 & n171 ;
  assign n3931 = n3668 | n3930 ;
  assign n33029 = ~n3712 ;
  assign n3869 = n3668 & n33029 ;
  assign n3870 = n32863 & n3869 ;
  assign n3942 = n3870 & n3940 ;
  assign n33030 = ~n3942 ;
  assign n3943 = n3931 & n33030 ;
  assign n4028 = n175 & n33015 ;
  assign n33031 = ~n4028 ;
  assign n4029 = n4016 & n33031 ;
  assign n33032 = ~n4029 ;
  assign n4030 = n2431 & n33032 ;
  assign n4031 = n177 | n4030 ;
  assign n33033 = ~n4031 ;
  assign n4032 = n4020 & n33033 ;
  assign n4033 = n3943 | n4032 ;
  assign n33034 = ~n4022 ;
  assign n4034 = n33034 & n4033 ;
  assign n33035 = ~n4034 ;
  assign n4035 = n178 & n33035 ;
  assign n3867 = n3715 | n3718 ;
  assign n33036 = ~n3867 ;
  assign n3898 = n33036 & n171 ;
  assign n3899 = n3651 | n3898 ;
  assign n3717 = n3651 & n32869 ;
  assign n33037 = ~n3718 ;
  assign n3866 = n3717 & n33037 ;
  assign n3951 = n3866 & n3940 ;
  assign n33038 = ~n3951 ;
  assign n3952 = n3899 & n33038 ;
  assign n4023 = n178 | n4022 ;
  assign n33039 = ~n4023 ;
  assign n4036 = n33039 & n4033 ;
  assign n4037 = n3952 | n4036 ;
  assign n33040 = ~n4035 ;
  assign n4038 = n33040 & n4037 ;
  assign n33041 = ~n4038 ;
  assign n4039 = n1707 & n33041 ;
  assign n3863 = n3721 | n3722 ;
  assign n33042 = ~n3863 ;
  assign n3919 = n33042 & n171 ;
  assign n3920 = n3664 | n3919 ;
  assign n33043 = ~n3722 ;
  assign n3864 = n3664 & n33043 ;
  assign n3865 = n32875 & n3864 ;
  assign n3944 = n3865 & n3940 ;
  assign n33044 = ~n3944 ;
  assign n3945 = n3920 & n33044 ;
  assign n33045 = ~n4030 ;
  assign n4047 = n4020 & n33045 ;
  assign n33046 = ~n4047 ;
  assign n4048 = n177 & n33046 ;
  assign n33047 = ~n4048 ;
  assign n4049 = n4033 & n33047 ;
  assign n33048 = ~n4049 ;
  assign n4050 = n178 & n33048 ;
  assign n4051 = n1707 | n4050 ;
  assign n33049 = ~n4051 ;
  assign n4052 = n4037 & n33049 ;
  assign n4053 = n3945 | n4052 ;
  assign n33050 = ~n4039 ;
  assign n4054 = n33050 & n4053 ;
  assign n33051 = ~n4054 ;
  assign n4055 = n180 & n33051 ;
  assign n3862 = n3729 | n3739 ;
  assign n33052 = ~n3862 ;
  assign n3908 = n33052 & n171 ;
  assign n3909 = n3670 | n3908 ;
  assign n3727 = n3670 & n32881 ;
  assign n33053 = ~n3729 ;
  assign n3861 = n3727 & n33053 ;
  assign n3981 = n3861 & n3940 ;
  assign n33054 = ~n3981 ;
  assign n3982 = n3909 & n33054 ;
  assign n4040 = n1487 | n4039 ;
  assign n33055 = ~n4040 ;
  assign n4056 = n33055 & n4053 ;
  assign n4057 = n3982 | n4056 ;
  assign n33056 = ~n4055 ;
  assign n4058 = n33056 & n4057 ;
  assign n33057 = ~n4058 ;
  assign n4059 = n181 & n33057 ;
  assign n33058 = ~n3733 ;
  assign n3858 = n3633 & n33058 ;
  assign n3859 = n32906 & n3858 ;
  assign n3890 = n3859 & n171 ;
  assign n3860 = n3733 | n3741 ;
  assign n33059 = ~n3860 ;
  assign n3891 = n33059 & n171 ;
  assign n3892 = n3633 | n3891 ;
  assign n33060 = ~n3890 ;
  assign n3893 = n33060 & n3892 ;
  assign n33061 = ~n4050 ;
  assign n4067 = n4037 & n33061 ;
  assign n33062 = ~n4067 ;
  assign n4068 = n179 & n33062 ;
  assign n33063 = ~n4068 ;
  assign n4069 = n4053 & n33063 ;
  assign n33064 = ~n4069 ;
  assign n4070 = n1487 & n33064 ;
  assign n4071 = n181 | n4070 ;
  assign n33065 = ~n4071 ;
  assign n4072 = n4057 & n33065 ;
  assign n4073 = n3893 | n4072 ;
  assign n33066 = ~n4059 ;
  assign n4074 = n33066 & n4073 ;
  assign n33067 = ~n4074 ;
  assign n4075 = n182 & n33067 ;
  assign n3857 = n3736 | n3743 ;
  assign n33068 = ~n3857 ;
  assign n3900 = n33068 & n171 ;
  assign n3901 = n3635 | n3900 ;
  assign n3738 = n3635 & n32895 ;
  assign n33069 = ~n3743 ;
  assign n3856 = n3738 & n33069 ;
  assign n3983 = n3856 & n3940 ;
  assign n33070 = ~n3983 ;
  assign n3984 = n3901 & n33070 ;
  assign n4060 = n182 | n4059 ;
  assign n33071 = ~n4060 ;
  assign n4076 = n33071 & n4073 ;
  assign n4077 = n3984 | n4076 ;
  assign n33072 = ~n4075 ;
  assign n4078 = n33072 & n4077 ;
  assign n33073 = ~n4078 ;
  assign n4079 = n996 & n33073 ;
  assign n3855 = n3747 | n3756 ;
  assign n33074 = ~n3855 ;
  assign n3896 = n33074 & n171 ;
  assign n3897 = n3672 | n3896 ;
  assign n33075 = ~n3747 ;
  assign n3853 = n3672 & n33075 ;
  assign n3854 = n32922 & n3853 ;
  assign n3906 = n3854 & n171 ;
  assign n33076 = ~n3906 ;
  assign n3907 = n3897 & n33076 ;
  assign n33077 = ~n4070 ;
  assign n4087 = n4057 & n33077 ;
  assign n33078 = ~n4087 ;
  assign n4088 = n181 & n33078 ;
  assign n33079 = ~n4088 ;
  assign n4089 = n4073 & n33079 ;
  assign n33080 = ~n4089 ;
  assign n4090 = n182 & n33080 ;
  assign n4091 = n183 | n4090 ;
  assign n33081 = ~n4091 ;
  assign n4092 = n4077 & n33081 ;
  assign n4093 = n3907 | n4092 ;
  assign n33082 = ~n4079 ;
  assign n4094 = n33082 & n4093 ;
  assign n33083 = ~n4094 ;
  assign n4095 = n184 & n33083 ;
  assign n3771 = n3750 | n3758 ;
  assign n33084 = ~n3771 ;
  assign n3902 = n33084 & n171 ;
  assign n3903 = n3674 | n3902 ;
  assign n3752 = n3674 & n32911 ;
  assign n33085 = ~n3758 ;
  assign n3770 = n3752 & n33085 ;
  assign n3985 = n3770 & n3940 ;
  assign n33086 = ~n3985 ;
  assign n3986 = n3903 & n33086 ;
  assign n4080 = n838 | n4079 ;
  assign n33087 = ~n4080 ;
  assign n4096 = n33087 & n4093 ;
  assign n4097 = n3986 | n4096 ;
  assign n33088 = ~n4095 ;
  assign n4098 = n33088 & n4097 ;
  assign n33089 = ~n4098 ;
  assign n4099 = n185 & n33089 ;
  assign n3852 = n3762 | n3773 ;
  assign n33090 = ~n3852 ;
  assign n3917 = n33090 & n171 ;
  assign n3918 = n3680 | n3917 ;
  assign n33091 = ~n3762 ;
  assign n3850 = n3680 & n33091 ;
  assign n3851 = n32938 & n3850 ;
  assign n3987 = n3851 & n3940 ;
  assign n33092 = ~n3987 ;
  assign n3988 = n3918 & n33092 ;
  assign n33093 = ~n4090 ;
  assign n4107 = n4077 & n33093 ;
  assign n33094 = ~n4107 ;
  assign n4108 = n183 & n33094 ;
  assign n33095 = ~n4108 ;
  assign n4109 = n4093 & n33095 ;
  assign n33096 = ~n4109 ;
  assign n4110 = n838 & n33096 ;
  assign n4111 = n185 | n4110 ;
  assign n33097 = ~n4111 ;
  assign n4112 = n4097 & n33097 ;
  assign n4113 = n3988 | n4112 ;
  assign n33098 = ~n4099 ;
  assign n4114 = n33098 & n4113 ;
  assign n33099 = ~n4114 ;
  assign n4115 = n186 & n33099 ;
  assign n3849 = n3765 | n3775 ;
  assign n33100 = ~n3849 ;
  assign n3910 = n33100 & n171 ;
  assign n3911 = n3676 | n3910 ;
  assign n3767 = n3676 & n32927 ;
  assign n33101 = ~n3775 ;
  assign n3848 = n3767 & n33101 ;
  assign n3989 = n3848 & n3940 ;
  assign n33102 = ~n3989 ;
  assign n3990 = n3911 & n33102 ;
  assign n4100 = n186 | n4099 ;
  assign n33103 = ~n4100 ;
  assign n4116 = n33103 & n4113 ;
  assign n4117 = n3990 | n4116 ;
  assign n33104 = ~n4115 ;
  assign n4118 = n33104 & n4117 ;
  assign n33105 = ~n4118 ;
  assign n4119 = n528 & n33105 ;
  assign n33106 = ~n3779 ;
  assign n3845 = n3643 & n33106 ;
  assign n3846 = n32954 & n3845 ;
  assign n3894 = n3846 & n171 ;
  assign n3847 = n3779 | n3788 ;
  assign n33107 = ~n3847 ;
  assign n3925 = n33107 & n171 ;
  assign n3926 = n3643 | n3925 ;
  assign n33108 = ~n3894 ;
  assign n3927 = n33108 & n3926 ;
  assign n33109 = ~n4110 ;
  assign n4127 = n4097 & n33109 ;
  assign n33110 = ~n4127 ;
  assign n4128 = n185 & n33110 ;
  assign n33111 = ~n4128 ;
  assign n4129 = n4113 & n33111 ;
  assign n33112 = ~n4129 ;
  assign n4130 = n186 & n33112 ;
  assign n4131 = n528 | n4130 ;
  assign n33113 = ~n4131 ;
  assign n4132 = n4117 & n33113 ;
  assign n4133 = n3927 | n4132 ;
  assign n33114 = ~n4119 ;
  assign n4134 = n33114 & n4133 ;
  assign n33115 = ~n4134 ;
  assign n4135 = n188 & n33115 ;
  assign n3844 = n3782 | n3790 ;
  assign n33116 = ~n3844 ;
  assign n3928 = n33116 & n171 ;
  assign n3929 = n3645 | n3928 ;
  assign n3784 = n3645 & n32943 ;
  assign n33117 = ~n3790 ;
  assign n3843 = n3784 & n33117 ;
  assign n3991 = n3843 & n3940 ;
  assign n33118 = ~n3991 ;
  assign n3992 = n3929 & n33118 ;
  assign n4120 = n413 | n4119 ;
  assign n33119 = ~n4120 ;
  assign n4136 = n33119 & n4133 ;
  assign n4137 = n3992 | n4136 ;
  assign n33120 = ~n4135 ;
  assign n4138 = n33120 & n4137 ;
  assign n33121 = ~n4138 ;
  assign n4139 = n189 & n33121 ;
  assign n33122 = ~n3794 ;
  assign n3840 = n3637 & n33122 ;
  assign n3841 = n32970 & n3840 ;
  assign n3941 = n3841 & n3940 ;
  assign n3842 = n3794 | n3803 ;
  assign n33123 = ~n3842 ;
  assign n3946 = n33123 & n3940 ;
  assign n3947 = n3637 | n3946 ;
  assign n33124 = ~n3941 ;
  assign n3948 = n33124 & n3947 ;
  assign n33125 = ~n4130 ;
  assign n4147 = n4117 & n33125 ;
  assign n33126 = ~n4147 ;
  assign n4148 = n187 & n33126 ;
  assign n33127 = ~n4148 ;
  assign n4149 = n4133 & n33127 ;
  assign n33128 = ~n4149 ;
  assign n4150 = n413 & n33128 ;
  assign n4151 = n189 | n4150 ;
  assign n33129 = ~n4151 ;
  assign n4152 = n4137 & n33129 ;
  assign n4153 = n3948 | n4152 ;
  assign n33130 = ~n4139 ;
  assign n4154 = n33130 & n4153 ;
  assign n33131 = ~n4154 ;
  assign n4155 = n190 & n33131 ;
  assign n3839 = n3797 | n3805 ;
  assign n33132 = ~n3839 ;
  assign n3912 = n33132 & n171 ;
  assign n3913 = n3666 | n3912 ;
  assign n3799 = n3666 & n32959 ;
  assign n33133 = ~n3805 ;
  assign n3838 = n3799 & n33133 ;
  assign n3921 = n3838 & n171 ;
  assign n33134 = ~n3921 ;
  assign n3922 = n3913 & n33134 ;
  assign n4140 = n190 | n4139 ;
  assign n33135 = ~n4140 ;
  assign n4156 = n33135 & n4153 ;
  assign n4157 = n3922 | n4156 ;
  assign n33136 = ~n4155 ;
  assign n4158 = n33136 & n4157 ;
  assign n33137 = ~n4158 ;
  assign n4159 = n287 & n33137 ;
  assign n33138 = ~n3809 ;
  assign n3835 = n3682 & n33138 ;
  assign n3836 = n32985 & n3835 ;
  assign n3895 = n3836 & n171 ;
  assign n3837 = n3809 | n3818 ;
  assign n33139 = ~n3837 ;
  assign n3914 = n33139 & n171 ;
  assign n3915 = n3682 | n3914 ;
  assign n33140 = ~n3895 ;
  assign n3916 = n33140 & n3915 ;
  assign n33141 = ~n4150 ;
  assign n4167 = n4137 & n33141 ;
  assign n33142 = ~n4167 ;
  assign n4168 = n189 & n33142 ;
  assign n33143 = ~n4168 ;
  assign n4169 = n4153 & n33143 ;
  assign n33144 = ~n4169 ;
  assign n4170 = n190 & n33144 ;
  assign n4171 = n287 | n4170 ;
  assign n33145 = ~n4171 ;
  assign n4172 = n4157 & n33145 ;
  assign n4176 = n3916 | n4172 ;
  assign n33146 = ~n4159 ;
  assign n4177 = n33146 & n4176 ;
  assign n4178 = n3959 | n4177 ;
  assign n4179 = n31336 & n4178 ;
  assign n4160 = n3950 & n33146 ;
  assign n4182 = n4160 & n4176 ;
  assign n3825 = n192 & n3824 ;
  assign n33147 = ~n3684 ;
  assign n3932 = n33147 & n171 ;
  assign n33148 = ~n3932 ;
  assign n3933 = n3822 & n33148 ;
  assign n33149 = ~n3933 ;
  assign n3934 = n3825 & n33149 ;
  assign n4187 = n3683 | n3882 ;
  assign n33150 = ~n4187 ;
  assign n4188 = n3612 & n33150 ;
  assign n4189 = n33004 & n4188 ;
  assign n4190 = n33005 & n4189 ;
  assign n4191 = n33006 & n4190 ;
  assign n4192 = n3934 | n4191 ;
  assign n4193 = n4182 | n4192 ;
  assign n170 = n4179 | n4193 ;
  assign n4180 = n3950 | n4177 ;
  assign n33151 = ~n4180 ;
  assign n4203 = n33151 & n170 ;
  assign n4204 = n4182 | n4203 ;
  assign n33152 = ~n4172 ;
  assign n4173 = n3916 & n33152 ;
  assign n4174 = n33146 & n4173 ;
  assign n4209 = n4174 & n170 ;
  assign n4175 = n4159 | n4172 ;
  assign n33153 = ~n4175 ;
  assign n4231 = n33153 & n170 ;
  assign n4232 = n3916 | n4231 ;
  assign n33154 = ~n4209 ;
  assign n4233 = n33154 & n4232 ;
  assign n4234 = n4204 | n4233 ;
  assign n33155 = ~n2714 ;
  assign n4202 = n33155 & n170 ;
  assign n33156 = ~n4191 ;
  assign n4293 = n3940 & n33156 ;
  assign n33157 = ~n3934 ;
  assign n4294 = n33157 & n4293 ;
  assign n33158 = ~n4182 ;
  assign n4295 = n33158 & n4294 ;
  assign n33159 = ~n4179 ;
  assign n4296 = n33159 & n4295 ;
  assign n4297 = n4202 | n4296 ;
  assign n4298 = x84 & n4297 ;
  assign n4299 = x84 | n4296 ;
  assign n4300 = n4202 | n4299 ;
  assign n33160 = ~n4298 ;
  assign n4301 = n33160 & n4300 ;
  assign n3584 = x80 | x81 ;
  assign n33161 = ~x82 ;
  assign n4194 = n33161 & n3584 ;
  assign n33162 = ~n170 ;
  assign n4197 = x82 & n33162 ;
  assign n4198 = n4194 | n4197 ;
  assign n33163 = ~n4198 ;
  assign n4199 = n3940 & n33163 ;
  assign n4200 = n3631 | n4199 ;
  assign n4290 = n33161 & n170 ;
  assign n33164 = ~n4290 ;
  assign n4291 = x83 & n33164 ;
  assign n4292 = n4202 | n4291 ;
  assign n4201 = x82 & n170 ;
  assign n3885 = x82 | n3584 ;
  assign n4319 = n3885 & n33003 ;
  assign n4320 = n33004 & n4319 ;
  assign n4321 = n33005 & n4320 ;
  assign n4322 = n33006 & n4321 ;
  assign n33165 = ~n4201 ;
  assign n4323 = n33165 & n4322 ;
  assign n4324 = n4292 | n4323 ;
  assign n33166 = ~n4200 ;
  assign n4325 = n33166 & n4324 ;
  assign n4326 = n4301 | n4325 ;
  assign n4225 = n3885 & n33165 ;
  assign n33167 = ~n4225 ;
  assign n4226 = n171 & n33167 ;
  assign n33168 = ~n4226 ;
  assign n4328 = n33168 & n4324 ;
  assign n33169 = ~n4328 ;
  assign n4329 = n3631 & n33169 ;
  assign n33170 = ~n4329 ;
  assign n4330 = n4326 & n33170 ;
  assign n33171 = ~n4330 ;
  assign n4331 = n173 & n33171 ;
  assign n3962 = n3955 | n3961 ;
  assign n33172 = ~n3962 ;
  assign n3967 = n33172 & n3966 ;
  assign n4195 = n3967 & n170 ;
  assign n4254 = n33172 & n170 ;
  assign n4255 = n3966 | n4254 ;
  assign n33173 = ~n4195 ;
  assign n4256 = n33173 & n4255 ;
  assign n4335 = n173 | n4329 ;
  assign n33174 = ~n4335 ;
  assign n4336 = n4326 & n33174 ;
  assign n4337 = n4256 | n4336 ;
  assign n33175 = ~n4331 ;
  assign n4338 = n33175 & n4337 ;
  assign n33176 = ~n4338 ;
  assign n4339 = n174 & n33176 ;
  assign n33177 = ~n3973 ;
  assign n4007 = n33177 & n4001 ;
  assign n4008 = n33008 & n4007 ;
  assign n4237 = n4008 & n170 ;
  assign n3974 = n3970 | n3973 ;
  assign n33178 = ~n3974 ;
  assign n4238 = n33178 & n170 ;
  assign n4239 = n4001 | n4238 ;
  assign n33179 = ~n4237 ;
  assign n4240 = n33179 & n4239 ;
  assign n4332 = n174 | n4331 ;
  assign n33180 = ~n4332 ;
  assign n4340 = n33180 & n4337 ;
  assign n4341 = n4240 | n4340 ;
  assign n33181 = ~n4339 ;
  assign n4342 = n33181 & n4341 ;
  assign n33182 = ~n4342 ;
  assign n4343 = n2753 & n33182 ;
  assign n4005 = n3976 & n33014 ;
  assign n33183 = ~n4010 ;
  assign n4185 = n4005 & n33183 ;
  assign n4196 = n4185 & n170 ;
  assign n4186 = n4004 | n4010 ;
  assign n33184 = ~n4186 ;
  assign n4228 = n33184 & n170 ;
  assign n4229 = n3976 | n4228 ;
  assign n33185 = ~n4196 ;
  assign n4230 = n33185 & n4229 ;
  assign n4350 = n172 & n33169 ;
  assign n4227 = n172 | n4226 ;
  assign n33186 = ~n4227 ;
  assign n4352 = n33186 & n4324 ;
  assign n4353 = n4301 | n4352 ;
  assign n33187 = ~n4350 ;
  assign n4354 = n33187 & n4353 ;
  assign n33188 = ~n4354 ;
  assign n4355 = n173 & n33188 ;
  assign n4356 = n33174 & n4353 ;
  assign n4357 = n4256 | n4356 ;
  assign n33189 = ~n4355 ;
  assign n4358 = n33189 & n4357 ;
  assign n33190 = ~n4358 ;
  assign n4359 = n174 & n33190 ;
  assign n4360 = n2753 | n4359 ;
  assign n33191 = ~n4360 ;
  assign n4361 = n4341 & n33191 ;
  assign n4362 = n4230 | n4361 ;
  assign n33192 = ~n4343 ;
  assign n4363 = n33192 & n4362 ;
  assign n33193 = ~n4363 ;
  assign n4364 = n176 & n33193 ;
  assign n4027 = n4013 | n4015 ;
  assign n33194 = ~n4027 ;
  assign n4241 = n33194 & n170 ;
  assign n4242 = n3978 | n4241 ;
  assign n33195 = ~n4015 ;
  assign n4025 = n3978 & n33195 ;
  assign n4026 = n33020 & n4025 ;
  assign n4243 = n4026 & n170 ;
  assign n33196 = ~n4243 ;
  assign n4244 = n4242 & n33196 ;
  assign n4345 = n2431 | n4343 ;
  assign n33197 = ~n4345 ;
  assign n4365 = n33197 & n4362 ;
  assign n4366 = n4244 | n4365 ;
  assign n33198 = ~n4364 ;
  assign n4367 = n33198 & n4366 ;
  assign n33199 = ~n4367 ;
  assign n4368 = n177 & n33199 ;
  assign n4024 = n4018 | n4019 ;
  assign n33200 = ~n4024 ;
  assign n4223 = n33200 & n170 ;
  assign n4224 = n3980 | n4223 ;
  assign n4045 = n3980 & n33045 ;
  assign n33201 = ~n4019 ;
  assign n4046 = n33201 & n4045 ;
  assign n4235 = n4046 & n170 ;
  assign n33202 = ~n4235 ;
  assign n4236 = n4224 & n33202 ;
  assign n4376 = n33180 & n4357 ;
  assign n4377 = n4240 | n4376 ;
  assign n33203 = ~n4359 ;
  assign n4378 = n33203 & n4377 ;
  assign n33204 = ~n4378 ;
  assign n4379 = n175 & n33204 ;
  assign n4380 = n33191 & n4377 ;
  assign n4381 = n4230 | n4380 ;
  assign n33205 = ~n4379 ;
  assign n4382 = n33205 & n4381 ;
  assign n33206 = ~n4382 ;
  assign n4383 = n2431 & n33206 ;
  assign n4384 = n177 | n4383 ;
  assign n33207 = ~n4384 ;
  assign n4385 = n4366 & n33207 ;
  assign n4386 = n4236 | n4385 ;
  assign n33208 = ~n4368 ;
  assign n4387 = n33208 & n4386 ;
  assign n33209 = ~n4387 ;
  assign n4388 = n178 & n33209 ;
  assign n4044 = n4022 | n4032 ;
  assign n33210 = ~n4044 ;
  assign n4247 = n33210 & n170 ;
  assign n4248 = n3943 | n4247 ;
  assign n33211 = ~n4032 ;
  assign n4042 = n3943 & n33211 ;
  assign n4043 = n33034 & n4042 ;
  assign n4273 = n4043 & n170 ;
  assign n33212 = ~n4273 ;
  assign n4274 = n4248 & n33212 ;
  assign n4369 = n178 | n4368 ;
  assign n33213 = ~n4369 ;
  assign n4389 = n33213 & n4386 ;
  assign n4390 = n4274 | n4389 ;
  assign n33214 = ~n4388 ;
  assign n4391 = n33214 & n4390 ;
  assign n33215 = ~n4391 ;
  assign n4392 = n1707 & n33215 ;
  assign n4041 = n4035 | n4036 ;
  assign n33216 = ~n4041 ;
  assign n4250 = n33216 & n170 ;
  assign n4251 = n3952 | n4250 ;
  assign n4065 = n3952 & n33061 ;
  assign n33217 = ~n4036 ;
  assign n4066 = n33217 & n4065 ;
  assign n4271 = n4066 & n170 ;
  assign n33218 = ~n4271 ;
  assign n4272 = n4251 & n33218 ;
  assign n4400 = n33197 & n4381 ;
  assign n4401 = n4244 | n4400 ;
  assign n33219 = ~n4383 ;
  assign n4402 = n33219 & n4401 ;
  assign n33220 = ~n4402 ;
  assign n4403 = n177 & n33220 ;
  assign n4404 = n33207 & n4401 ;
  assign n4405 = n4236 | n4404 ;
  assign n33221 = ~n4403 ;
  assign n4406 = n33221 & n4405 ;
  assign n33222 = ~n4406 ;
  assign n4407 = n178 & n33222 ;
  assign n4408 = n1707 | n4407 ;
  assign n33223 = ~n4408 ;
  assign n4409 = n4390 & n33223 ;
  assign n4410 = n4272 | n4409 ;
  assign n33224 = ~n4392 ;
  assign n4411 = n33224 & n4410 ;
  assign n33225 = ~n4411 ;
  assign n4412 = n180 & n33225 ;
  assign n4064 = n4039 | n4052 ;
  assign n33226 = ~n4064 ;
  assign n4259 = n33226 & n170 ;
  assign n4260 = n3945 | n4259 ;
  assign n33227 = ~n4052 ;
  assign n4062 = n3945 & n33227 ;
  assign n4063 = n33050 & n4062 ;
  assign n4279 = n4063 & n170 ;
  assign n33228 = ~n4279 ;
  assign n4280 = n4260 & n33228 ;
  assign n4393 = n1487 | n4392 ;
  assign n33229 = ~n4393 ;
  assign n4413 = n33229 & n4410 ;
  assign n4414 = n4280 | n4413 ;
  assign n33230 = ~n4412 ;
  assign n4415 = n33230 & n4414 ;
  assign n33231 = ~n4415 ;
  assign n4416 = n181 & n33231 ;
  assign n4085 = n3982 & n33077 ;
  assign n33232 = ~n4056 ;
  assign n4086 = n33232 & n4085 ;
  assign n4249 = n4086 & n170 ;
  assign n4061 = n4055 | n4056 ;
  assign n33233 = ~n4061 ;
  assign n4263 = n33233 & n170 ;
  assign n4264 = n3982 | n4263 ;
  assign n33234 = ~n4249 ;
  assign n4265 = n33234 & n4264 ;
  assign n4424 = n33213 & n4405 ;
  assign n4425 = n4274 | n4424 ;
  assign n33235 = ~n4407 ;
  assign n4426 = n33235 & n4425 ;
  assign n33236 = ~n4426 ;
  assign n4427 = n179 & n33236 ;
  assign n4428 = n33223 & n4425 ;
  assign n4429 = n4272 | n4428 ;
  assign n33237 = ~n4427 ;
  assign n4430 = n33237 & n4429 ;
  assign n33238 = ~n4430 ;
  assign n4431 = n1487 & n33238 ;
  assign n4432 = n181 | n4431 ;
  assign n33239 = ~n4432 ;
  assign n4433 = n4414 & n33239 ;
  assign n4434 = n4265 | n4433 ;
  assign n33240 = ~n4416 ;
  assign n4435 = n33240 & n4434 ;
  assign n33241 = ~n4435 ;
  assign n4436 = n182 & n33241 ;
  assign n4084 = n4059 | n4072 ;
  assign n33242 = ~n4084 ;
  assign n4281 = n33242 & n170 ;
  assign n4282 = n3893 | n4281 ;
  assign n33243 = ~n4072 ;
  assign n4082 = n3893 & n33243 ;
  assign n4083 = n33066 & n4082 ;
  assign n4283 = n4083 & n170 ;
  assign n33244 = ~n4283 ;
  assign n4284 = n4282 & n33244 ;
  assign n4417 = n182 | n4416 ;
  assign n33245 = ~n4417 ;
  assign n4437 = n33245 & n4434 ;
  assign n4438 = n4284 | n4437 ;
  assign n33246 = ~n4436 ;
  assign n4439 = n33246 & n4438 ;
  assign n33247 = ~n4439 ;
  assign n4440 = n996 & n33247 ;
  assign n4105 = n3984 & n33093 ;
  assign n33248 = ~n4076 ;
  assign n4106 = n33248 & n4105 ;
  assign n4208 = n4106 & n170 ;
  assign n4081 = n4075 | n4076 ;
  assign n33249 = ~n4081 ;
  assign n4285 = n33249 & n170 ;
  assign n4286 = n3984 | n4285 ;
  assign n33250 = ~n4208 ;
  assign n4287 = n33250 & n4286 ;
  assign n4448 = n33229 & n4429 ;
  assign n4449 = n4280 | n4448 ;
  assign n33251 = ~n4431 ;
  assign n4450 = n33251 & n4449 ;
  assign n33252 = ~n4450 ;
  assign n4451 = n181 & n33252 ;
  assign n4452 = n33239 & n4449 ;
  assign n4453 = n4265 | n4452 ;
  assign n33253 = ~n4451 ;
  assign n4454 = n33253 & n4453 ;
  assign n33254 = ~n4454 ;
  assign n4455 = n182 & n33254 ;
  assign n4456 = n183 | n4455 ;
  assign n33255 = ~n4456 ;
  assign n4457 = n4438 & n33255 ;
  assign n4458 = n4287 | n4457 ;
  assign n33256 = ~n4440 ;
  assign n4459 = n33256 & n4458 ;
  assign n33257 = ~n4459 ;
  assign n4460 = n184 & n33257 ;
  assign n4102 = n4079 | n4092 ;
  assign n33258 = ~n4102 ;
  assign n4277 = n33258 & n170 ;
  assign n4278 = n3907 | n4277 ;
  assign n33259 = ~n4092 ;
  assign n4103 = n3907 & n33259 ;
  assign n4104 = n33082 & n4103 ;
  assign n4288 = n4104 & n170 ;
  assign n33260 = ~n4288 ;
  assign n4289 = n4278 & n33260 ;
  assign n4441 = n838 | n4440 ;
  assign n33261 = ~n4441 ;
  assign n4461 = n33261 & n4458 ;
  assign n4462 = n4289 | n4461 ;
  assign n33262 = ~n4460 ;
  assign n4463 = n33262 & n4462 ;
  assign n33263 = ~n4463 ;
  assign n4464 = n185 & n33263 ;
  assign n4101 = n4095 | n4096 ;
  assign n33264 = ~n4101 ;
  assign n4252 = n33264 & n170 ;
  assign n4253 = n3986 | n4252 ;
  assign n4125 = n3986 & n33109 ;
  assign n33265 = ~n4096 ;
  assign n4126 = n33265 & n4125 ;
  assign n4275 = n4126 & n170 ;
  assign n33266 = ~n4275 ;
  assign n4276 = n4253 & n33266 ;
  assign n4472 = n33245 & n4453 ;
  assign n4473 = n4284 | n4472 ;
  assign n33267 = ~n4455 ;
  assign n4474 = n33267 & n4473 ;
  assign n33268 = ~n4474 ;
  assign n4475 = n183 & n33268 ;
  assign n4476 = n33255 & n4473 ;
  assign n4477 = n4287 | n4476 ;
  assign n33269 = ~n4475 ;
  assign n4478 = n33269 & n4477 ;
  assign n33270 = ~n4478 ;
  assign n4479 = n838 & n33270 ;
  assign n4480 = n185 | n4479 ;
  assign n33271 = ~n4480 ;
  assign n4481 = n4462 & n33271 ;
  assign n4482 = n4276 | n4481 ;
  assign n33272 = ~n4464 ;
  assign n4483 = n33272 & n4482 ;
  assign n33273 = ~n4483 ;
  assign n4484 = n186 & n33273 ;
  assign n4124 = n4099 | n4112 ;
  assign n33274 = ~n4124 ;
  assign n4245 = n33274 & n170 ;
  assign n4246 = n3988 | n4245 ;
  assign n33275 = ~n4112 ;
  assign n4122 = n3988 & n33275 ;
  assign n4123 = n33098 & n4122 ;
  assign n4257 = n4123 & n170 ;
  assign n33276 = ~n4257 ;
  assign n4258 = n4246 & n33276 ;
  assign n4465 = n186 | n4464 ;
  assign n33277 = ~n4465 ;
  assign n4485 = n33277 & n4482 ;
  assign n4486 = n4258 | n4485 ;
  assign n33278 = ~n4484 ;
  assign n4487 = n33278 & n4486 ;
  assign n33279 = ~n4487 ;
  assign n4488 = n528 & n33279 ;
  assign n4145 = n3990 & n33125 ;
  assign n33280 = ~n4116 ;
  assign n4146 = n33280 & n4145 ;
  assign n4219 = n4146 & n170 ;
  assign n4121 = n4115 | n4116 ;
  assign n33281 = ~n4121 ;
  assign n4220 = n33281 & n170 ;
  assign n4221 = n3990 | n4220 ;
  assign n33282 = ~n4219 ;
  assign n4222 = n33282 & n4221 ;
  assign n4496 = n33261 & n4477 ;
  assign n4497 = n4289 | n4496 ;
  assign n33283 = ~n4479 ;
  assign n4498 = n33283 & n4497 ;
  assign n33284 = ~n4498 ;
  assign n4499 = n185 & n33284 ;
  assign n4500 = n33271 & n4497 ;
  assign n4501 = n4276 | n4500 ;
  assign n33285 = ~n4499 ;
  assign n4502 = n33285 & n4501 ;
  assign n33286 = ~n4502 ;
  assign n4503 = n186 & n33286 ;
  assign n4504 = n528 | n4503 ;
  assign n33287 = ~n4504 ;
  assign n4505 = n4486 & n33287 ;
  assign n4506 = n4222 | n4505 ;
  assign n33288 = ~n4488 ;
  assign n4507 = n33288 & n4506 ;
  assign n33289 = ~n4507 ;
  assign n4508 = n188 & n33289 ;
  assign n33290 = ~n4132 ;
  assign n4142 = n3927 & n33290 ;
  assign n4143 = n33114 & n4142 ;
  assign n4215 = n4143 & n170 ;
  assign n4144 = n4119 | n4132 ;
  assign n33291 = ~n4144 ;
  assign n4216 = n33291 & n170 ;
  assign n4217 = n3927 | n4216 ;
  assign n33292 = ~n4215 ;
  assign n4218 = n33292 & n4217 ;
  assign n4489 = n413 | n4488 ;
  assign n33293 = ~n4489 ;
  assign n4509 = n33293 & n4506 ;
  assign n4510 = n4218 | n4509 ;
  assign n33294 = ~n4508 ;
  assign n4511 = n33294 & n4510 ;
  assign n33295 = ~n4511 ;
  assign n4512 = n189 & n33295 ;
  assign n4165 = n3992 & n33141 ;
  assign n33296 = ~n4136 ;
  assign n4166 = n33296 & n4165 ;
  assign n4214 = n4166 & n170 ;
  assign n4141 = n4135 | n4136 ;
  assign n33297 = ~n4141 ;
  assign n4268 = n33297 & n170 ;
  assign n4269 = n3992 | n4268 ;
  assign n33298 = ~n4214 ;
  assign n4270 = n33298 & n4269 ;
  assign n4520 = n33277 & n4501 ;
  assign n4521 = n4258 | n4520 ;
  assign n33299 = ~n4503 ;
  assign n4522 = n33299 & n4521 ;
  assign n33300 = ~n4522 ;
  assign n4523 = n187 & n33300 ;
  assign n4524 = n33287 & n4521 ;
  assign n4525 = n4222 | n4524 ;
  assign n33301 = ~n4523 ;
  assign n4526 = n33301 & n4525 ;
  assign n33302 = ~n4526 ;
  assign n4527 = n413 & n33302 ;
  assign n4528 = n189 | n4527 ;
  assign n33303 = ~n4528 ;
  assign n4529 = n4510 & n33303 ;
  assign n4530 = n4270 | n4529 ;
  assign n33304 = ~n4512 ;
  assign n4531 = n33304 & n4530 ;
  assign n33305 = ~n4531 ;
  assign n4532 = n190 & n33305 ;
  assign n4162 = n4139 | n4152 ;
  assign n33306 = ~n4162 ;
  assign n4261 = n33306 & n170 ;
  assign n4262 = n3948 | n4261 ;
  assign n33307 = ~n4152 ;
  assign n4163 = n3948 & n33307 ;
  assign n4164 = n33130 & n4163 ;
  assign n4266 = n4164 & n170 ;
  assign n33308 = ~n4266 ;
  assign n4267 = n4262 & n33308 ;
  assign n4514 = n190 | n4512 ;
  assign n33309 = ~n4514 ;
  assign n4533 = n33309 & n4530 ;
  assign n4534 = n4267 | n4533 ;
  assign n33310 = ~n4532 ;
  assign n4535 = n33310 & n4534 ;
  assign n33311 = ~n4535 ;
  assign n4536 = n287 & n33311 ;
  assign n33312 = ~n4170 ;
  assign n4183 = n3922 & n33312 ;
  assign n33313 = ~n4156 ;
  assign n4184 = n33313 & n4183 ;
  assign n4210 = n4184 & n170 ;
  assign n4161 = n4155 | n4156 ;
  assign n33314 = ~n4161 ;
  assign n4211 = n33314 & n170 ;
  assign n4212 = n3922 | n4211 ;
  assign n33315 = ~n4210 ;
  assign n4213 = n33315 & n4212 ;
  assign n4544 = n33293 & n4525 ;
  assign n4545 = n4218 | n4544 ;
  assign n33316 = ~n4527 ;
  assign n4546 = n33316 & n4545 ;
  assign n33317 = ~n4546 ;
  assign n4547 = n189 & n33317 ;
  assign n4548 = n33303 & n4545 ;
  assign n4549 = n4270 | n4548 ;
  assign n33318 = ~n4547 ;
  assign n4550 = n33318 & n4549 ;
  assign n33319 = ~n4550 ;
  assign n4551 = n190 & n33319 ;
  assign n4552 = n287 | n4551 ;
  assign n33320 = ~n4552 ;
  assign n4553 = n4534 & n33320 ;
  assign n4556 = n4213 | n4553 ;
  assign n33321 = ~n4536 ;
  assign n4557 = n33321 & n4556 ;
  assign n4560 = n4234 | n4557 ;
  assign n4561 = n31336 & n4560 ;
  assign n4181 = n192 & n4180 ;
  assign n33322 = ~n3950 ;
  assign n4205 = n33322 & n170 ;
  assign n33323 = ~n4205 ;
  assign n4206 = n4177 & n33323 ;
  assign n33324 = ~n4206 ;
  assign n4207 = n4181 & n33324 ;
  assign n4302 = n3949 | n4191 ;
  assign n33325 = ~n4302 ;
  assign n4303 = n3905 & n33325 ;
  assign n4304 = n33157 & n4303 ;
  assign n4305 = n33158 & n4304 ;
  assign n4306 = n33159 & n4305 ;
  assign n4307 = n4207 | n4306 ;
  assign n4537 = n4233 & n33321 ;
  assign n4562 = n4537 & n4556 ;
  assign n4563 = n4307 | n4562 ;
  assign n169 = n4561 | n4563 ;
  assign n4555 = n4536 | n4553 ;
  assign n33326 = ~n4555 ;
  assign n4568 = n33326 & n169 ;
  assign n4569 = n4213 | n4568 ;
  assign n4538 = n4213 & n33321 ;
  assign n33327 = ~n4553 ;
  assign n4554 = n4538 & n33327 ;
  assign n4635 = n4554 & n169 ;
  assign n33328 = ~n4635 ;
  assign n4636 = n4569 & n33328 ;
  assign n4558 = n4233 | n4557 ;
  assign n33329 = ~n4558 ;
  assign n4656 = n33329 & n169 ;
  assign n4669 = n4562 | n4656 ;
  assign n4670 = n4636 | n4669 ;
  assign n4564 = x78 | x79 ;
  assign n5012 = x80 | n4564 ;
  assign n4590 = x80 & n169 ;
  assign n33330 = ~n4590 ;
  assign n4591 = n5012 & n33330 ;
  assign n33331 = ~n4591 ;
  assign n4592 = n170 & n33331 ;
  assign n4315 = n5012 & n33156 ;
  assign n4316 = n33157 & n4315 ;
  assign n4317 = n33158 & n4316 ;
  assign n4318 = n33159 & n4317 ;
  assign n4615 = n4318 & n33330 ;
  assign n33332 = ~n3584 ;
  assign n4617 = n33332 & n169 ;
  assign n33333 = ~x80 ;
  assign n4657 = n33333 & n169 ;
  assign n33334 = ~n4657 ;
  assign n4658 = x81 & n33334 ;
  assign n4659 = n4617 | n4658 ;
  assign n4660 = n4615 | n4659 ;
  assign n33335 = ~n4592 ;
  assign n4661 = n33335 & n4660 ;
  assign n33336 = ~n4661 ;
  assign n4662 = n3940 & n33336 ;
  assign n5295 = n33333 & n4564 ;
  assign n33337 = ~n169 ;
  assign n4648 = x80 & n33337 ;
  assign n4649 = n5295 | n4648 ;
  assign n33338 = ~n4649 ;
  assign n4650 = n170 & n33338 ;
  assign n4651 = n3940 | n4650 ;
  assign n33339 = ~n4651 ;
  assign n4665 = n33339 & n4660 ;
  assign n33340 = ~n4306 ;
  assign n4308 = n170 & n33340 ;
  assign n33341 = ~n4207 ;
  assign n4309 = n33341 & n4308 ;
  assign n33342 = ~n4562 ;
  assign n4683 = n4309 & n33342 ;
  assign n33343 = ~n4561 ;
  assign n4684 = n33343 & n4683 ;
  assign n4685 = n4617 | n4684 ;
  assign n4686 = x82 & n4685 ;
  assign n4687 = x82 | n4684 ;
  assign n4688 = n4617 | n4687 ;
  assign n33344 = ~n4686 ;
  assign n4689 = n33344 & n4688 ;
  assign n4690 = n4665 | n4689 ;
  assign n33345 = ~n4662 ;
  assign n4691 = n33345 & n4690 ;
  assign n33346 = ~n4691 ;
  assign n4692 = n3631 & n33346 ;
  assign n4663 = n3631 | n4662 ;
  assign n33347 = ~n4663 ;
  assign n4694 = n33347 & n4690 ;
  assign n4706 = n4199 | n4323 ;
  assign n33348 = ~n4706 ;
  assign n4707 = n4292 & n33348 ;
  assign n4708 = n169 & n4707 ;
  assign n4709 = n169 & n33348 ;
  assign n4710 = n4292 | n4709 ;
  assign n33349 = ~n4708 ;
  assign n4711 = n33349 & n4710 ;
  assign n4714 = n4694 | n4711 ;
  assign n33350 = ~n4692 ;
  assign n4715 = n33350 & n4714 ;
  assign n33351 = ~n4715 ;
  assign n4716 = n173 & n33351 ;
  assign n4351 = n4325 | n4350 ;
  assign n33352 = ~n4351 ;
  assign n4577 = n33352 & n169 ;
  assign n4578 = n4301 | n4577 ;
  assign n33353 = ~n4325 ;
  assign n4327 = n4301 & n33353 ;
  assign n4334 = n4327 & n33170 ;
  assign n4652 = n4334 & n169 ;
  assign n33354 = ~n4652 ;
  assign n4653 = n4578 & n33354 ;
  assign n4693 = n173 | n4692 ;
  assign n33355 = ~n4693 ;
  assign n4717 = n33355 & n4714 ;
  assign n4718 = n4653 | n4717 ;
  assign n33356 = ~n4716 ;
  assign n4719 = n33356 & n4718 ;
  assign n33357 = ~n4719 ;
  assign n4720 = n174 & n33357 ;
  assign n4349 = n4331 | n4336 ;
  assign n33358 = ~n4349 ;
  assign n4611 = n33358 & n169 ;
  assign n4612 = n4256 | n4611 ;
  assign n4333 = n4256 & n33175 ;
  assign n33359 = ~n4336 ;
  assign n4348 = n4333 & n33359 ;
  assign n4654 = n4348 & n169 ;
  assign n33360 = ~n4654 ;
  assign n4655 = n4612 & n33360 ;
  assign n4664 = n171 & n33336 ;
  assign n4593 = n171 | n4592 ;
  assign n33361 = ~n4593 ;
  assign n4667 = n33361 & n4660 ;
  assign n4698 = n4667 | n4689 ;
  assign n33362 = ~n4664 ;
  assign n4699 = n33362 & n4698 ;
  assign n33363 = ~n4699 ;
  assign n4700 = n172 & n33363 ;
  assign n4701 = n33347 & n4698 ;
  assign n4726 = n4701 | n4711 ;
  assign n33364 = ~n4700 ;
  assign n4727 = n33364 & n4726 ;
  assign n33365 = ~n4727 ;
  assign n4728 = n173 & n33365 ;
  assign n4729 = n174 | n4728 ;
  assign n33366 = ~n4729 ;
  assign n4730 = n4718 & n33366 ;
  assign n4731 = n4655 | n4730 ;
  assign n33367 = ~n4720 ;
  assign n4732 = n33367 & n4731 ;
  assign n33368 = ~n4732 ;
  assign n4733 = n175 & n33368 ;
  assign n4375 = n4340 | n4359 ;
  assign n33369 = ~n4375 ;
  assign n4607 = n33369 & n169 ;
  assign n4608 = n4240 | n4607 ;
  assign n33370 = ~n4340 ;
  assign n4346 = n4240 & n33370 ;
  assign n4347 = n33181 & n4346 ;
  assign n4613 = n4347 & n169 ;
  assign n33371 = ~n4613 ;
  assign n4614 = n4608 & n33371 ;
  assign n4721 = n2753 | n4720 ;
  assign n33372 = ~n4721 ;
  assign n4734 = n33372 & n4731 ;
  assign n4735 = n4614 | n4734 ;
  assign n33373 = ~n4733 ;
  assign n4736 = n33373 & n4735 ;
  assign n33374 = ~n4736 ;
  assign n4737 = n2431 & n33374 ;
  assign n4344 = n4230 & n33192 ;
  assign n33375 = ~n4361 ;
  assign n4373 = n4344 & n33375 ;
  assign n4598 = n4373 & n169 ;
  assign n4374 = n4343 | n4361 ;
  assign n33376 = ~n4374 ;
  assign n4604 = n33376 & n169 ;
  assign n4605 = n4230 | n4604 ;
  assign n33377 = ~n4598 ;
  assign n4606 = n33377 & n4605 ;
  assign n4745 = n33355 & n4726 ;
  assign n4746 = n4653 | n4745 ;
  assign n33378 = ~n4728 ;
  assign n4747 = n33378 & n4746 ;
  assign n33379 = ~n4747 ;
  assign n4748 = n174 & n33379 ;
  assign n4749 = n33366 & n4746 ;
  assign n4750 = n4655 | n4749 ;
  assign n33380 = ~n4748 ;
  assign n4751 = n33380 & n4750 ;
  assign n33381 = ~n4751 ;
  assign n4752 = n2753 & n33381 ;
  assign n4753 = n2431 | n4752 ;
  assign n33382 = ~n4753 ;
  assign n4754 = n4735 & n33382 ;
  assign n4755 = n4606 | n4754 ;
  assign n33383 = ~n4737 ;
  assign n4756 = n33383 & n4755 ;
  assign n33384 = ~n4756 ;
  assign n4757 = n177 & n33384 ;
  assign n4399 = n4365 | n4383 ;
  assign n33385 = ~n4399 ;
  assign n4571 = n33385 & n169 ;
  assign n4572 = n4244 | n4571 ;
  assign n33386 = ~n4365 ;
  assign n4371 = n4244 & n33386 ;
  assign n4372 = n33198 & n4371 ;
  assign n4609 = n4372 & n169 ;
  assign n33387 = ~n4609 ;
  assign n4610 = n4572 & n33387 ;
  assign n4738 = n177 | n4737 ;
  assign n33388 = ~n4738 ;
  assign n4758 = n33388 & n4755 ;
  assign n4759 = n4610 | n4758 ;
  assign n33389 = ~n4757 ;
  assign n4760 = n33389 & n4759 ;
  assign n33390 = ~n4760 ;
  assign n4761 = n178 & n33390 ;
  assign n4398 = n4368 | n4385 ;
  assign n33391 = ~n4398 ;
  assign n4620 = n33391 & n169 ;
  assign n4621 = n4236 | n4620 ;
  assign n4370 = n4236 & n33208 ;
  assign n33392 = ~n4385 ;
  assign n4397 = n4370 & n33392 ;
  assign n4630 = n4397 & n169 ;
  assign n33393 = ~n4630 ;
  assign n4631 = n4621 & n33393 ;
  assign n4769 = n33372 & n4750 ;
  assign n4770 = n4614 | n4769 ;
  assign n33394 = ~n4752 ;
  assign n4771 = n33394 & n4770 ;
  assign n33395 = ~n4771 ;
  assign n4772 = n176 & n33395 ;
  assign n4773 = n33382 & n4770 ;
  assign n4774 = n4606 | n4773 ;
  assign n33396 = ~n4772 ;
  assign n4775 = n33396 & n4774 ;
  assign n33397 = ~n4775 ;
  assign n4776 = n177 & n33397 ;
  assign n4777 = n178 | n4776 ;
  assign n33398 = ~n4777 ;
  assign n4778 = n4759 & n33398 ;
  assign n4779 = n4631 | n4778 ;
  assign n33399 = ~n4761 ;
  assign n4780 = n33399 & n4779 ;
  assign n33400 = ~n4780 ;
  assign n4781 = n179 & n33400 ;
  assign n4423 = n4389 | n4407 ;
  assign n33401 = ~n4423 ;
  assign n4596 = n33401 & n169 ;
  assign n4597 = n4274 | n4596 ;
  assign n33402 = ~n4389 ;
  assign n4395 = n4274 & n33402 ;
  assign n4396 = n33214 & n4395 ;
  assign n4600 = n4396 & n169 ;
  assign n33403 = ~n4600 ;
  assign n4601 = n4597 & n33403 ;
  assign n4762 = n1707 | n4761 ;
  assign n33404 = ~n4762 ;
  assign n4782 = n33404 & n4779 ;
  assign n4783 = n4601 | n4782 ;
  assign n33405 = ~n4781 ;
  assign n4784 = n33405 & n4783 ;
  assign n33406 = ~n4784 ;
  assign n4785 = n1487 & n33406 ;
  assign n4394 = n4272 & n33224 ;
  assign n33407 = ~n4409 ;
  assign n4421 = n4394 & n33407 ;
  assign n4622 = n4421 & n169 ;
  assign n4422 = n4392 | n4409 ;
  assign n33408 = ~n4422 ;
  assign n4625 = n33408 & n169 ;
  assign n4626 = n4272 | n4625 ;
  assign n33409 = ~n4622 ;
  assign n4627 = n33409 & n4626 ;
  assign n4793 = n33388 & n4774 ;
  assign n4794 = n4610 | n4793 ;
  assign n33410 = ~n4776 ;
  assign n4795 = n33410 & n4794 ;
  assign n33411 = ~n4795 ;
  assign n4796 = n178 & n33411 ;
  assign n4797 = n33398 & n4794 ;
  assign n4798 = n4631 | n4797 ;
  assign n33412 = ~n4796 ;
  assign n4799 = n33412 & n4798 ;
  assign n33413 = ~n4799 ;
  assign n4800 = n1707 & n33413 ;
  assign n4801 = n1487 | n4800 ;
  assign n33414 = ~n4801 ;
  assign n4802 = n4783 & n33414 ;
  assign n4803 = n4627 | n4802 ;
  assign n33415 = ~n4785 ;
  assign n4804 = n33415 & n4803 ;
  assign n33416 = ~n4804 ;
  assign n4805 = n181 & n33416 ;
  assign n33417 = ~n4413 ;
  assign n4419 = n4280 & n33417 ;
  assign n4420 = n33230 & n4419 ;
  assign n4619 = n4420 & n169 ;
  assign n4447 = n4413 | n4431 ;
  assign n33418 = ~n4447 ;
  assign n4632 = n33418 & n169 ;
  assign n4633 = n4280 | n4632 ;
  assign n33419 = ~n4619 ;
  assign n4634 = n33419 & n4633 ;
  assign n4786 = n181 | n4785 ;
  assign n33420 = ~n4786 ;
  assign n4806 = n33420 & n4803 ;
  assign n4807 = n4634 | n4806 ;
  assign n33421 = ~n4805 ;
  assign n4808 = n33421 & n4807 ;
  assign n33422 = ~n4808 ;
  assign n4809 = n182 & n33422 ;
  assign n4446 = n4416 | n4433 ;
  assign n33423 = ~n4446 ;
  assign n4628 = n33423 & n169 ;
  assign n4629 = n4265 | n4628 ;
  assign n4418 = n4265 & n33240 ;
  assign n33424 = ~n4433 ;
  assign n4445 = n4418 & n33424 ;
  assign n4637 = n4445 & n169 ;
  assign n33425 = ~n4637 ;
  assign n4638 = n4629 & n33425 ;
  assign n4817 = n33404 & n4798 ;
  assign n4818 = n4601 | n4817 ;
  assign n33426 = ~n4800 ;
  assign n4819 = n33426 & n4818 ;
  assign n33427 = ~n4819 ;
  assign n4820 = n180 & n33427 ;
  assign n4821 = n33414 & n4818 ;
  assign n4822 = n4627 | n4821 ;
  assign n33428 = ~n4820 ;
  assign n4823 = n33428 & n4822 ;
  assign n33429 = ~n4823 ;
  assign n4824 = n181 & n33429 ;
  assign n4825 = n182 | n4824 ;
  assign n33430 = ~n4825 ;
  assign n4826 = n4807 & n33430 ;
  assign n4827 = n4638 | n4826 ;
  assign n33431 = ~n4809 ;
  assign n4828 = n33431 & n4827 ;
  assign n33432 = ~n4828 ;
  assign n4829 = n183 & n33432 ;
  assign n4471 = n4437 | n4455 ;
  assign n33433 = ~n4471 ;
  assign n4582 = n33433 & n169 ;
  assign n4583 = n4284 | n4582 ;
  assign n33434 = ~n4437 ;
  assign n4443 = n4284 & n33434 ;
  assign n4444 = n33246 & n4443 ;
  assign n4594 = n4444 & n169 ;
  assign n33435 = ~n4594 ;
  assign n4595 = n4583 & n33435 ;
  assign n4810 = n183 | n4809 ;
  assign n33436 = ~n4810 ;
  assign n4830 = n33436 & n4827 ;
  assign n4831 = n4595 | n4830 ;
  assign n33437 = ~n4829 ;
  assign n4832 = n33437 & n4831 ;
  assign n33438 = ~n4832 ;
  assign n4833 = n838 & n33438 ;
  assign n4442 = n4287 & n33256 ;
  assign n33439 = ~n4457 ;
  assign n4470 = n4442 & n33439 ;
  assign n4599 = n4470 & n169 ;
  assign n4469 = n4440 | n4457 ;
  assign n33440 = ~n4469 ;
  assign n4639 = n33440 & n169 ;
  assign n4640 = n4287 | n4639 ;
  assign n33441 = ~n4599 ;
  assign n4641 = n33441 & n4640 ;
  assign n4841 = n33420 & n4822 ;
  assign n4842 = n4634 | n4841 ;
  assign n33442 = ~n4824 ;
  assign n4843 = n33442 & n4842 ;
  assign n33443 = ~n4843 ;
  assign n4844 = n182 & n33443 ;
  assign n4845 = n33430 & n4842 ;
  assign n4846 = n4638 | n4845 ;
  assign n33444 = ~n4844 ;
  assign n4847 = n33444 & n4846 ;
  assign n33445 = ~n4847 ;
  assign n4848 = n996 & n33445 ;
  assign n4849 = n838 | n4848 ;
  assign n33446 = ~n4849 ;
  assign n4850 = n4831 & n33446 ;
  assign n4851 = n4641 | n4850 ;
  assign n33447 = ~n4833 ;
  assign n4852 = n33447 & n4851 ;
  assign n33448 = ~n4852 ;
  assign n4853 = n185 & n33448 ;
  assign n33449 = ~n4461 ;
  assign n4467 = n4289 & n33449 ;
  assign n4468 = n33262 & n4467 ;
  assign n4618 = n4468 & n169 ;
  assign n4495 = n4461 | n4479 ;
  assign n33450 = ~n4495 ;
  assign n4642 = n33450 & n169 ;
  assign n4643 = n4289 | n4642 ;
  assign n33451 = ~n4618 ;
  assign n4644 = n33451 & n4643 ;
  assign n4834 = n185 | n4833 ;
  assign n33452 = ~n4834 ;
  assign n4854 = n33452 & n4851 ;
  assign n4855 = n4644 | n4854 ;
  assign n33453 = ~n4853 ;
  assign n4856 = n33453 & n4855 ;
  assign n33454 = ~n4856 ;
  assign n4857 = n186 & n33454 ;
  assign n4494 = n4464 | n4481 ;
  assign n33455 = ~n4494 ;
  assign n4588 = n33455 & n169 ;
  assign n4589 = n4276 | n4588 ;
  assign n4466 = n4276 & n33272 ;
  assign n33456 = ~n4481 ;
  assign n4493 = n4466 & n33456 ;
  assign n4623 = n4493 & n169 ;
  assign n33457 = ~n4623 ;
  assign n4624 = n4589 & n33457 ;
  assign n4865 = n33436 & n4846 ;
  assign n4866 = n4595 | n4865 ;
  assign n33458 = ~n4848 ;
  assign n4867 = n33458 & n4866 ;
  assign n33459 = ~n4867 ;
  assign n4868 = n184 & n33459 ;
  assign n4869 = n33446 & n4866 ;
  assign n4870 = n4641 | n4869 ;
  assign n33460 = ~n4868 ;
  assign n4871 = n33460 & n4870 ;
  assign n33461 = ~n4871 ;
  assign n4872 = n185 & n33461 ;
  assign n4873 = n186 | n4872 ;
  assign n33462 = ~n4873 ;
  assign n4874 = n4855 & n33462 ;
  assign n4875 = n4624 | n4874 ;
  assign n33463 = ~n4857 ;
  assign n4876 = n33463 & n4875 ;
  assign n33464 = ~n4876 ;
  assign n4877 = n187 & n33464 ;
  assign n33465 = ~n4485 ;
  assign n4491 = n4258 & n33465 ;
  assign n4492 = n33278 & n4491 ;
  assign n4584 = n4492 & n169 ;
  assign n4519 = n4485 | n4503 ;
  assign n33466 = ~n4519 ;
  assign n4585 = n33466 & n169 ;
  assign n4586 = n4258 | n4585 ;
  assign n33467 = ~n4584 ;
  assign n4587 = n33467 & n4586 ;
  assign n4858 = n528 | n4857 ;
  assign n33468 = ~n4858 ;
  assign n4878 = n33468 & n4875 ;
  assign n4879 = n4587 | n4878 ;
  assign n33469 = ~n4877 ;
  assign n4880 = n33469 & n4879 ;
  assign n33470 = ~n4880 ;
  assign n4881 = n413 & n33470 ;
  assign n4490 = n4222 & n33288 ;
  assign n33471 = ~n4505 ;
  assign n4517 = n4490 & n33471 ;
  assign n4565 = n4517 & n169 ;
  assign n4518 = n4488 | n4505 ;
  assign n33472 = ~n4518 ;
  assign n4579 = n33472 & n169 ;
  assign n4580 = n4222 | n4579 ;
  assign n33473 = ~n4565 ;
  assign n4581 = n33473 & n4580 ;
  assign n4889 = n33452 & n4870 ;
  assign n4890 = n4644 | n4889 ;
  assign n33474 = ~n4872 ;
  assign n4891 = n33474 & n4890 ;
  assign n33475 = ~n4891 ;
  assign n4892 = n186 & n33475 ;
  assign n4893 = n33462 & n4890 ;
  assign n4894 = n4624 | n4893 ;
  assign n33476 = ~n4892 ;
  assign n4895 = n33476 & n4894 ;
  assign n33477 = ~n4895 ;
  assign n4896 = n528 & n33477 ;
  assign n4897 = n413 | n4896 ;
  assign n33478 = ~n4897 ;
  assign n4898 = n4879 & n33478 ;
  assign n4899 = n4581 | n4898 ;
  assign n33479 = ~n4881 ;
  assign n4900 = n33479 & n4899 ;
  assign n33480 = ~n4900 ;
  assign n4901 = n189 & n33480 ;
  assign n4543 = n4509 | n4527 ;
  assign n33481 = ~n4543 ;
  assign n4566 = n33481 & n169 ;
  assign n4567 = n4218 | n4566 ;
  assign n33482 = ~n4509 ;
  assign n4515 = n4218 & n33482 ;
  assign n4516 = n33294 & n4515 ;
  assign n4575 = n4516 & n169 ;
  assign n33483 = ~n4575 ;
  assign n4576 = n4567 & n33483 ;
  assign n4882 = n189 | n4881 ;
  assign n33484 = ~n4882 ;
  assign n4902 = n33484 & n4899 ;
  assign n4903 = n4576 | n4902 ;
  assign n33485 = ~n4901 ;
  assign n4904 = n33485 & n4903 ;
  assign n33486 = ~n4904 ;
  assign n4905 = n190 & n33486 ;
  assign n4542 = n4512 | n4529 ;
  assign n33487 = ~n4542 ;
  assign n4573 = n33487 & n169 ;
  assign n4574 = n4270 | n4573 ;
  assign n4513 = n4270 & n33304 ;
  assign n33488 = ~n4529 ;
  assign n4541 = n4513 & n33488 ;
  assign n4602 = n4541 & n169 ;
  assign n33489 = ~n4602 ;
  assign n4603 = n4574 & n33489 ;
  assign n4911 = n33468 & n4894 ;
  assign n4912 = n4587 | n4911 ;
  assign n33490 = ~n4896 ;
  assign n4913 = n33490 & n4912 ;
  assign n33491 = ~n4913 ;
  assign n4914 = n188 & n33491 ;
  assign n4915 = n33478 & n4912 ;
  assign n4916 = n4581 | n4915 ;
  assign n33492 = ~n4914 ;
  assign n4917 = n33492 & n4916 ;
  assign n33493 = ~n4917 ;
  assign n4918 = n189 & n33493 ;
  assign n4919 = n190 | n4918 ;
  assign n33494 = ~n4919 ;
  assign n4920 = n4903 & n33494 ;
  assign n4921 = n4603 | n4920 ;
  assign n33495 = ~n4905 ;
  assign n4926 = n33495 & n4921 ;
  assign n33496 = ~n4926 ;
  assign n4927 = n191 & n33496 ;
  assign n33497 = ~n4533 ;
  assign n4539 = n4267 & n33497 ;
  assign n4540 = n33310 & n4539 ;
  assign n4570 = n4540 & n169 ;
  assign n4702 = n4533 | n4551 ;
  assign n33498 = ~n4702 ;
  assign n4703 = n169 & n33498 ;
  assign n4704 = n4267 | n4703 ;
  assign n33499 = ~n4570 ;
  assign n4705 = n33499 & n4704 ;
  assign n4908 = n191 | n4905 ;
  assign n33500 = ~n4908 ;
  assign n4988 = n33500 & n4921 ;
  assign n4989 = n4705 | n4988 ;
  assign n33501 = ~n4927 ;
  assign n4990 = n33501 & n4989 ;
  assign n4991 = n4670 | n4990 ;
  assign n4992 = n31336 & n4991 ;
  assign n4559 = n192 & n4558 ;
  assign n33502 = ~n4233 ;
  assign n4645 = n33502 & n169 ;
  assign n33503 = ~n4645 ;
  assign n4646 = n4557 & n33503 ;
  assign n33504 = ~n4646 ;
  assign n4647 = n4559 & n33504 ;
  assign n4310 = n4209 | n4306 ;
  assign n33505 = ~n4310 ;
  assign n4311 = n4232 & n33505 ;
  assign n4312 = n33341 & n4311 ;
  assign n4671 = n4312 & n33342 ;
  assign n4672 = n33343 & n4671 ;
  assign n4673 = n4647 | n4672 ;
  assign n4931 = n4636 & n33501 ;
  assign n5010 = n4931 & n4989 ;
  assign n5011 = n4673 | n5010 ;
  assign n168 = n4992 | n5011 ;
  assign n4906 = n287 | n4905 ;
  assign n33506 = ~n4906 ;
  assign n4922 = n33506 & n4921 ;
  assign n4923 = n4705 | n4922 ;
  assign n4932 = n4923 & n4931 ;
  assign n4928 = n4923 & n33501 ;
  assign n4929 = n4670 | n4928 ;
  assign n4930 = n31336 & n4929 ;
  assign n4933 = n4673 | n4932 ;
  assign n4934 = n4930 | n4933 ;
  assign n4983 = n4636 | n4928 ;
  assign n33507 = ~n4983 ;
  assign n4984 = n4934 & n33507 ;
  assign n4985 = n4932 | n4984 ;
  assign n33508 = ~n4988 ;
  assign n5263 = n4705 & n33508 ;
  assign n5264 = n33501 & n5263 ;
  assign n5265 = n4934 & n5264 ;
  assign n5267 = n4927 | n4988 ;
  assign n33509 = ~n5267 ;
  assign n5268 = n168 & n33509 ;
  assign n5269 = n4705 | n5268 ;
  assign n33510 = ~n5265 ;
  assign n5270 = n33510 & n5269 ;
  assign n5271 = n4985 | n5270 ;
  assign n4883 = n4581 & n33479 ;
  assign n33511 = ~n4898 ;
  assign n4909 = n4883 & n33511 ;
  assign n4951 = n4909 & n4934 ;
  assign n4910 = n4881 | n4898 ;
  assign n33512 = ~n4910 ;
  assign n5022 = n33512 & n168 ;
  assign n5023 = n4581 | n5022 ;
  assign n33513 = ~n4951 ;
  assign n5024 = n33513 & n5023 ;
  assign n33514 = ~n4564 ;
  assign n4935 = n33514 & n4934 ;
  assign n33515 = ~x78 ;
  assign n4936 = n33515 & n4934 ;
  assign n33516 = ~n4936 ;
  assign n4937 = x79 & n33516 ;
  assign n4938 = n4935 | n4937 ;
  assign n5677 = x76 | x77 ;
  assign n6101 = x78 | n5677 ;
  assign n4313 = n6101 & n33340 ;
  assign n4314 = n33341 & n4313 ;
  assign n4681 = n4314 & n33342 ;
  assign n4682 = n33343 & n4681 ;
  assign n4939 = x78 & n4934 ;
  assign n33517 = ~n4939 ;
  assign n4940 = n4682 & n33517 ;
  assign n4941 = n4938 | n4940 ;
  assign n6542 = n33515 & n5677 ;
  assign n33518 = ~n4934 ;
  assign n4954 = x78 & n33518 ;
  assign n4955 = n6542 | n4954 ;
  assign n33519 = ~n4955 ;
  assign n4956 = n169 & n33519 ;
  assign n33520 = ~n4956 ;
  assign n4957 = n4941 & n33520 ;
  assign n33521 = ~n4957 ;
  assign n4958 = n170 & n33521 ;
  assign n4959 = n171 | n4958 ;
  assign n4962 = n170 | n4956 ;
  assign n33522 = ~n4962 ;
  assign n4963 = n4941 & n33522 ;
  assign n33523 = ~n4672 ;
  assign n4674 = n169 & n33523 ;
  assign n33524 = ~n4647 ;
  assign n4675 = n33524 & n4674 ;
  assign n33525 = ~n4932 ;
  assign n4979 = n4675 & n33525 ;
  assign n33526 = ~n4992 ;
  assign n4993 = n4979 & n33526 ;
  assign n4994 = n4935 | n4993 ;
  assign n4995 = x80 & n4994 ;
  assign n4996 = x80 | n4993 ;
  assign n4997 = n4935 | n4996 ;
  assign n33527 = ~n4995 ;
  assign n4998 = n33527 & n4997 ;
  assign n5001 = n4963 | n4998 ;
  assign n33528 = ~n4959 ;
  assign n5002 = n33528 & n5001 ;
  assign n4616 = n4592 | n4615 ;
  assign n33529 = ~n4616 ;
  assign n5037 = n33529 & n168 ;
  assign n5038 = n4659 | n5037 ;
  assign n4668 = n33529 & n4659 ;
  assign n5048 = n4668 & n168 ;
  assign n33530 = ~n5048 ;
  assign n5049 = n5038 & n33530 ;
  assign n5050 = n5002 | n5049 ;
  assign n5054 = x78 & n168 ;
  assign n33531 = ~n5054 ;
  assign n5055 = n6101 & n33531 ;
  assign n33532 = ~n5055 ;
  assign n5056 = n169 & n33532 ;
  assign n5057 = n170 | n5056 ;
  assign n33533 = ~n5057 ;
  assign n5058 = n4941 & n33533 ;
  assign n5059 = n4998 | n5058 ;
  assign n33534 = ~n4958 ;
  assign n5060 = n33534 & n5059 ;
  assign n33535 = ~n5060 ;
  assign n5061 = n171 & n33535 ;
  assign n33536 = ~n5061 ;
  assign n5062 = n5050 & n33536 ;
  assign n33537 = ~n5062 ;
  assign n5063 = n172 & n33537 ;
  assign n33538 = ~n4665 ;
  assign n4696 = n33538 & n4689 ;
  assign n4697 = n33362 & n4696 ;
  assign n4942 = n4697 & n4934 ;
  assign n4666 = n4664 | n4665 ;
  assign n33539 = ~n4666 ;
  assign n5045 = n33539 & n168 ;
  assign n5046 = n4689 | n5045 ;
  assign n33540 = ~n4942 ;
  assign n5047 = n33540 & n5046 ;
  assign n5068 = n3940 & n33535 ;
  assign n5069 = n3631 | n5068 ;
  assign n33541 = ~n5069 ;
  assign n5070 = n5050 & n33541 ;
  assign n5071 = n5047 | n5070 ;
  assign n33542 = ~n5063 ;
  assign n5072 = n33542 & n5071 ;
  assign n33543 = ~n5072 ;
  assign n5073 = n173 & n33543 ;
  assign n5064 = n173 | n5063 ;
  assign n33544 = ~n5064 ;
  assign n5075 = n33544 & n5071 ;
  assign n4712 = n33350 & n4711 ;
  assign n33545 = ~n4694 ;
  assign n4713 = n33545 & n4712 ;
  assign n4948 = n4713 & n4934 ;
  assign n4695 = n4692 | n4694 ;
  assign n33546 = ~n4695 ;
  assign n5092 = n33546 & n168 ;
  assign n5093 = n4711 | n5092 ;
  assign n33547 = ~n4948 ;
  assign n5094 = n33547 & n5093 ;
  assign n5095 = n5075 | n5094 ;
  assign n33548 = ~n5073 ;
  assign n5096 = n33548 & n5095 ;
  assign n33549 = ~n5096 ;
  assign n5097 = n174 & n33549 ;
  assign n33550 = ~n4717 ;
  assign n4723 = n4653 & n33550 ;
  assign n4724 = n33356 & n4723 ;
  assign n4968 = n4724 & n4934 ;
  assign n4725 = n4716 | n4717 ;
  assign n33551 = ~n4725 ;
  assign n5031 = n33551 & n168 ;
  assign n5032 = n4653 | n5031 ;
  assign n33552 = ~n4968 ;
  assign n5033 = n33552 & n5032 ;
  assign n5074 = n174 | n5073 ;
  assign n33553 = ~n5074 ;
  assign n5099 = n33553 & n5095 ;
  assign n5100 = n5033 | n5099 ;
  assign n33554 = ~n5097 ;
  assign n5101 = n33554 & n5100 ;
  assign n33555 = ~n5101 ;
  assign n5102 = n175 & n33555 ;
  assign n4722 = n4655 & n33367 ;
  assign n33556 = ~n4730 ;
  assign n4743 = n4722 & n33556 ;
  assign n4947 = n4743 & n4934 ;
  assign n4744 = n4720 | n4730 ;
  assign n33557 = ~n4744 ;
  assign n5042 = n33557 & n168 ;
  assign n5043 = n4655 | n5042 ;
  assign n33558 = ~n4947 ;
  assign n5044 = n33558 & n5043 ;
  assign n5098 = n2753 | n5097 ;
  assign n33559 = ~n5098 ;
  assign n5103 = n33559 & n5100 ;
  assign n5104 = n5044 | n5103 ;
  assign n33560 = ~n5102 ;
  assign n5105 = n33560 & n5104 ;
  assign n33561 = ~n5105 ;
  assign n5106 = n2431 & n33561 ;
  assign n4742 = n4733 | n4734 ;
  assign n33562 = ~n4742 ;
  assign n4952 = n33562 & n4934 ;
  assign n4953 = n4614 | n4952 ;
  assign n33563 = ~n4734 ;
  assign n4740 = n4614 & n33563 ;
  assign n4741 = n33373 & n4740 ;
  assign n4969 = n4741 & n4934 ;
  assign n33564 = ~n4969 ;
  assign n4970 = n4953 & n33564 ;
  assign n5114 = n2753 & n33555 ;
  assign n5115 = n2431 | n5114 ;
  assign n33565 = ~n5115 ;
  assign n5116 = n5104 & n33565 ;
  assign n5117 = n4970 | n5116 ;
  assign n33566 = ~n5106 ;
  assign n5118 = n33566 & n5117 ;
  assign n33567 = ~n5118 ;
  assign n5119 = n177 & n33567 ;
  assign n4739 = n4606 & n33383 ;
  assign n33568 = ~n4754 ;
  assign n4767 = n4739 & n33568 ;
  assign n4950 = n4767 & n4934 ;
  assign n4768 = n4737 | n4754 ;
  assign n33569 = ~n4768 ;
  assign n5016 = n33569 & n168 ;
  assign n5017 = n4606 | n5016 ;
  assign n33570 = ~n4950 ;
  assign n5018 = n33570 & n5017 ;
  assign n5107 = n177 | n5106 ;
  assign n33571 = ~n5107 ;
  assign n5120 = n33571 & n5117 ;
  assign n5121 = n5018 | n5120 ;
  assign n33572 = ~n5119 ;
  assign n5122 = n33572 & n5121 ;
  assign n33573 = ~n5122 ;
  assign n5123 = n178 & n33573 ;
  assign n33574 = ~n4758 ;
  assign n4764 = n4610 & n33574 ;
  assign n4765 = n33389 & n4764 ;
  assign n4971 = n4765 & n4934 ;
  assign n4766 = n4757 | n4758 ;
  assign n33575 = ~n4766 ;
  assign n5028 = n33575 & n168 ;
  assign n5029 = n4610 | n5028 ;
  assign n33576 = ~n4971 ;
  assign n5030 = n33576 & n5029 ;
  assign n33577 = ~n5114 ;
  assign n5131 = n5104 & n33577 ;
  assign n33578 = ~n5131 ;
  assign n5132 = n176 & n33578 ;
  assign n33579 = ~n5132 ;
  assign n5133 = n5117 & n33579 ;
  assign n33580 = ~n5133 ;
  assign n5134 = n177 & n33580 ;
  assign n5135 = n178 | n5134 ;
  assign n33581 = ~n5135 ;
  assign n5136 = n5121 & n33581 ;
  assign n5137 = n5030 | n5136 ;
  assign n33582 = ~n5123 ;
  assign n5138 = n33582 & n5137 ;
  assign n33583 = ~n5138 ;
  assign n5139 = n179 & n33583 ;
  assign n4763 = n4631 & n33399 ;
  assign n33584 = ~n4778 ;
  assign n4791 = n4763 & n33584 ;
  assign n4972 = n4791 & n4934 ;
  assign n4792 = n4761 | n4778 ;
  assign n33585 = ~n4792 ;
  assign n5013 = n33585 & n168 ;
  assign n5014 = n4631 | n5013 ;
  assign n33586 = ~n4972 ;
  assign n5015 = n33586 & n5014 ;
  assign n5124 = n1707 | n5123 ;
  assign n33587 = ~n5124 ;
  assign n5140 = n33587 & n5137 ;
  assign n5141 = n5015 | n5140 ;
  assign n33588 = ~n5139 ;
  assign n5142 = n33588 & n5141 ;
  assign n33589 = ~n5142 ;
  assign n5143 = n1487 & n33589 ;
  assign n33590 = ~n4782 ;
  assign n4788 = n4601 & n33590 ;
  assign n4789 = n33405 & n4788 ;
  assign n4973 = n4789 & n4934 ;
  assign n4790 = n4781 | n4782 ;
  assign n33591 = ~n4790 ;
  assign n5025 = n33591 & n168 ;
  assign n5026 = n4601 | n5025 ;
  assign n33592 = ~n4973 ;
  assign n5027 = n33592 & n5026 ;
  assign n33593 = ~n5134 ;
  assign n5151 = n5121 & n33593 ;
  assign n33594 = ~n5151 ;
  assign n5152 = n178 & n33594 ;
  assign n33595 = ~n5152 ;
  assign n5153 = n5137 & n33595 ;
  assign n33596 = ~n5153 ;
  assign n5154 = n1707 & n33596 ;
  assign n5155 = n1487 | n5154 ;
  assign n33597 = ~n5155 ;
  assign n5156 = n5141 & n33597 ;
  assign n5157 = n5027 | n5156 ;
  assign n33598 = ~n5143 ;
  assign n5158 = n33598 & n5157 ;
  assign n33599 = ~n5158 ;
  assign n5159 = n181 & n33599 ;
  assign n4787 = n4627 & n33415 ;
  assign n33600 = ~n4802 ;
  assign n4815 = n4787 & n33600 ;
  assign n4965 = n4815 & n4934 ;
  assign n4816 = n4785 | n4802 ;
  assign n33601 = ~n4816 ;
  assign n5019 = n33601 & n168 ;
  assign n5020 = n4627 | n5019 ;
  assign n33602 = ~n4965 ;
  assign n5021 = n33602 & n5020 ;
  assign n5144 = n181 | n5143 ;
  assign n33603 = ~n5144 ;
  assign n5160 = n33603 & n5157 ;
  assign n5161 = n5021 | n5160 ;
  assign n33604 = ~n5159 ;
  assign n5162 = n33604 & n5161 ;
  assign n33605 = ~n5162 ;
  assign n5163 = n182 & n33605 ;
  assign n33606 = ~n4806 ;
  assign n4812 = n4634 & n33606 ;
  assign n4813 = n33421 & n4812 ;
  assign n4974 = n4813 & n4934 ;
  assign n4814 = n4805 | n4806 ;
  assign n33607 = ~n4814 ;
  assign n5034 = n33607 & n168 ;
  assign n5035 = n4634 | n5034 ;
  assign n33608 = ~n4974 ;
  assign n5036 = n33608 & n5035 ;
  assign n33609 = ~n5154 ;
  assign n5171 = n5141 & n33609 ;
  assign n33610 = ~n5171 ;
  assign n5172 = n180 & n33610 ;
  assign n33611 = ~n5172 ;
  assign n5173 = n5157 & n33611 ;
  assign n33612 = ~n5173 ;
  assign n5174 = n181 & n33612 ;
  assign n5175 = n182 | n5174 ;
  assign n33613 = ~n5175 ;
  assign n5176 = n5161 & n33613 ;
  assign n5177 = n5036 | n5176 ;
  assign n33614 = ~n5163 ;
  assign n5178 = n33614 & n5177 ;
  assign n33615 = ~n5178 ;
  assign n5179 = n183 & n33615 ;
  assign n4811 = n4638 & n33431 ;
  assign n33616 = ~n4826 ;
  assign n4839 = n4811 & n33616 ;
  assign n4967 = n4839 & n4934 ;
  assign n4840 = n4809 | n4826 ;
  assign n33617 = ~n4840 ;
  assign n5039 = n33617 & n168 ;
  assign n5040 = n4638 | n5039 ;
  assign n33618 = ~n4967 ;
  assign n5041 = n33618 & n5040 ;
  assign n5164 = n183 | n5163 ;
  assign n33619 = ~n5164 ;
  assign n5180 = n33619 & n5177 ;
  assign n5181 = n5041 | n5180 ;
  assign n33620 = ~n5179 ;
  assign n5182 = n33620 & n5181 ;
  assign n33621 = ~n5182 ;
  assign n5183 = n838 & n33621 ;
  assign n4838 = n4829 | n4830 ;
  assign n33622 = ~n4838 ;
  assign n4945 = n33622 & n4934 ;
  assign n4946 = n4595 | n4945 ;
  assign n33623 = ~n4830 ;
  assign n4836 = n4595 & n33623 ;
  assign n4837 = n33437 & n4836 ;
  assign n4975 = n4837 & n4934 ;
  assign n33624 = ~n4975 ;
  assign n4976 = n4946 & n33624 ;
  assign n33625 = ~n5174 ;
  assign n5191 = n5161 & n33625 ;
  assign n33626 = ~n5191 ;
  assign n5192 = n182 & n33626 ;
  assign n33627 = ~n5192 ;
  assign n5193 = n5177 & n33627 ;
  assign n33628 = ~n5193 ;
  assign n5194 = n996 & n33628 ;
  assign n5195 = n838 | n5194 ;
  assign n33629 = ~n5195 ;
  assign n5196 = n5181 & n33629 ;
  assign n5197 = n4976 | n5196 ;
  assign n33630 = ~n5183 ;
  assign n5198 = n33630 & n5197 ;
  assign n33631 = ~n5198 ;
  assign n5199 = n185 & n33631 ;
  assign n4835 = n4641 & n33447 ;
  assign n33632 = ~n4850 ;
  assign n4863 = n4835 & n33632 ;
  assign n4943 = n4863 & n4934 ;
  assign n4864 = n4833 | n4850 ;
  assign n33633 = ~n4864 ;
  assign n5080 = n33633 & n168 ;
  assign n5081 = n4641 | n5080 ;
  assign n33634 = ~n4943 ;
  assign n5082 = n33634 & n5081 ;
  assign n5184 = n185 | n5183 ;
  assign n33635 = ~n5184 ;
  assign n5200 = n33635 & n5197 ;
  assign n5201 = n5082 | n5200 ;
  assign n33636 = ~n5199 ;
  assign n5202 = n33636 & n5201 ;
  assign n33637 = ~n5202 ;
  assign n5203 = n186 & n33637 ;
  assign n33638 = ~n4854 ;
  assign n4860 = n4644 & n33638 ;
  assign n4861 = n33453 & n4860 ;
  assign n4944 = n4861 & n4934 ;
  assign n4862 = n4853 | n4854 ;
  assign n33639 = ~n4862 ;
  assign n5086 = n33639 & n168 ;
  assign n5087 = n4644 | n5086 ;
  assign n33640 = ~n4944 ;
  assign n5088 = n33640 & n5087 ;
  assign n33641 = ~n5194 ;
  assign n5210 = n5181 & n33641 ;
  assign n33642 = ~n5210 ;
  assign n5211 = n184 & n33642 ;
  assign n33643 = ~n5211 ;
  assign n5212 = n5197 & n33643 ;
  assign n33644 = ~n5212 ;
  assign n5213 = n185 & n33644 ;
  assign n5214 = n186 | n5213 ;
  assign n33645 = ~n5214 ;
  assign n5215 = n5201 & n33645 ;
  assign n5216 = n5088 | n5215 ;
  assign n33646 = ~n5203 ;
  assign n5217 = n33646 & n5216 ;
  assign n33647 = ~n5217 ;
  assign n5218 = n187 & n33647 ;
  assign n4859 = n4624 & n33463 ;
  assign n33648 = ~n4874 ;
  assign n4888 = n4859 & n33648 ;
  assign n4977 = n4888 & n4934 ;
  assign n4887 = n4857 | n4874 ;
  assign n33649 = ~n4887 ;
  assign n5083 = n33649 & n168 ;
  assign n5084 = n4624 | n5083 ;
  assign n33650 = ~n4977 ;
  assign n5085 = n33650 & n5084 ;
  assign n5204 = n528 | n5203 ;
  assign n33651 = ~n5204 ;
  assign n5219 = n33651 & n5216 ;
  assign n5220 = n5085 | n5219 ;
  assign n33652 = ~n5218 ;
  assign n5221 = n33652 & n5220 ;
  assign n33653 = ~n5221 ;
  assign n5222 = n413 & n33653 ;
  assign n5223 = n189 | n5222 ;
  assign n33654 = ~n4878 ;
  assign n4884 = n4587 & n33654 ;
  assign n4885 = n33469 & n4884 ;
  assign n4966 = n4885 & n4934 ;
  assign n4886 = n4877 | n4878 ;
  assign n33655 = ~n4886 ;
  assign n5089 = n33655 & n168 ;
  assign n5090 = n4587 | n5089 ;
  assign n33656 = ~n4966 ;
  assign n5091 = n33656 & n5090 ;
  assign n33657 = ~n5213 ;
  assign n5230 = n5201 & n33657 ;
  assign n33658 = ~n5230 ;
  assign n5231 = n186 & n33658 ;
  assign n33659 = ~n5231 ;
  assign n5232 = n5216 & n33659 ;
  assign n33660 = ~n5232 ;
  assign n5233 = n528 & n33660 ;
  assign n5234 = n413 | n5233 ;
  assign n33661 = ~n5234 ;
  assign n5235 = n5220 & n33661 ;
  assign n5236 = n5091 | n5235 ;
  assign n33662 = ~n5223 ;
  assign n5239 = n33662 & n5236 ;
  assign n5240 = n5024 | n5239 ;
  assign n33663 = ~n5233 ;
  assign n5251 = n5220 & n33663 ;
  assign n33664 = ~n5251 ;
  assign n5252 = n188 & n33664 ;
  assign n33665 = ~n5252 ;
  assign n5253 = n5236 & n33665 ;
  assign n33666 = ~n5253 ;
  assign n5254 = n189 & n33666 ;
  assign n33667 = ~n5254 ;
  assign n5261 = n5240 & n33667 ;
  assign n33668 = ~n5261 ;
  assign n5262 = n190 & n33668 ;
  assign n5255 = n190 | n5254 ;
  assign n33669 = ~n5255 ;
  assign n5256 = n5240 & n33669 ;
  assign n5274 = n33484 & n4916 ;
  assign n33670 = ~n5274 ;
  assign n5275 = n4576 & n33670 ;
  assign n5276 = n33485 & n5275 ;
  assign n5277 = n4934 & n5276 ;
  assign n5278 = n4901 | n5274 ;
  assign n33671 = ~n5278 ;
  assign n5279 = n168 & n33671 ;
  assign n5280 = n4576 | n5279 ;
  assign n33672 = ~n5277 ;
  assign n5281 = n33672 & n5280 ;
  assign n5282 = n5256 | n5281 ;
  assign n33673 = ~n5262 ;
  assign n5290 = n33673 & n5282 ;
  assign n33674 = ~n5290 ;
  assign n5291 = n287 & n33674 ;
  assign n4907 = n4603 & n33495 ;
  assign n33675 = ~n4920 ;
  assign n4925 = n4907 & n33675 ;
  assign n4978 = n4925 & n4934 ;
  assign n4924 = n4905 | n4920 ;
  assign n33676 = ~n4924 ;
  assign n5051 = n33676 & n168 ;
  assign n5052 = n4603 | n5051 ;
  assign n33677 = ~n4978 ;
  assign n5053 = n33677 & n5052 ;
  assign n33678 = ~n5222 ;
  assign n5237 = n33678 & n5236 ;
  assign n33679 = ~n5237 ;
  assign n5238 = n189 & n33679 ;
  assign n33680 = ~n5238 ;
  assign n5241 = n33680 & n5240 ;
  assign n33681 = ~n5241 ;
  assign n5242 = n190 & n33681 ;
  assign n5244 = n287 | n5242 ;
  assign n33682 = ~n5244 ;
  assign n5345 = n33682 & n5282 ;
  assign n5346 = n5053 | n5345 ;
  assign n33683 = ~n5291 ;
  assign n5347 = n33683 & n5346 ;
  assign n5348 = n5271 | n5347 ;
  assign n5349 = n31336 & n5348 ;
  assign n33684 = ~n4636 ;
  assign n4949 = n33684 & n4934 ;
  assign n33685 = ~n4949 ;
  assign n4982 = n4928 & n33685 ;
  assign n4986 = n192 & n4983 ;
  assign n33686 = ~n4982 ;
  assign n4987 = n33686 & n4986 ;
  assign n4676 = n4635 | n4672 ;
  assign n33687 = ~n4676 ;
  assign n4677 = n4569 & n33687 ;
  assign n4678 = n33524 & n4677 ;
  assign n4980 = n4678 & n33525 ;
  assign n5004 = n4980 & n33526 ;
  assign n5005 = n4987 | n5004 ;
  assign n5292 = n5270 & n33683 ;
  assign n5350 = n5292 & n5346 ;
  assign n5351 = n5005 | n5350 ;
  assign n5352 = n5349 | n5351 ;
  assign n5643 = n5270 | n5347 ;
  assign n33688 = ~n5643 ;
  assign n5644 = n5352 & n33688 ;
  assign n5645 = n5350 | n5644 ;
  assign n5243 = n191 | n5242 ;
  assign n33689 = ~n5243 ;
  assign n5285 = n33689 & n5282 ;
  assign n5344 = n5053 & n33683 ;
  assign n33690 = ~n5285 ;
  assign n5651 = n33690 & n5344 ;
  assign n5652 = n5352 & n5651 ;
  assign n33691 = ~n5242 ;
  assign n5283 = n33691 & n5282 ;
  assign n33692 = ~n5283 ;
  assign n5284 = n191 & n33692 ;
  assign n5286 = n5053 | n5285 ;
  assign n33693 = ~n5284 ;
  assign n5287 = n33693 & n5286 ;
  assign n5288 = n5271 | n5287 ;
  assign n5289 = n31336 & n5288 ;
  assign n5293 = n5286 & n5292 ;
  assign n5294 = n5005 | n5293 ;
  assign n167 = n5289 | n5294 ;
  assign n5654 = n5285 | n5291 ;
  assign n33694 = ~n5654 ;
  assign n5655 = n167 & n33694 ;
  assign n5656 = n5053 | n5655 ;
  assign n33695 = ~n5652 ;
  assign n5657 = n33695 & n5656 ;
  assign n5658 = n5645 | n5657 ;
  assign n6933 = x74 | x75 ;
  assign n33696 = ~x76 ;
  assign n7878 = n33696 & n6933 ;
  assign n33697 = ~n5352 ;
  assign n5373 = x76 & n33697 ;
  assign n5374 = n7878 | n5373 ;
  assign n33698 = ~n5374 ;
  assign n5375 = n4934 & n33698 ;
  assign n7327 = x76 | n6933 ;
  assign n4679 = n7327 & n33523 ;
  assign n4680 = n33524 & n4679 ;
  assign n4981 = n4680 & n33525 ;
  assign n5003 = n4981 & n33526 ;
  assign n5363 = x76 & n5352 ;
  assign n33699 = ~n5363 ;
  assign n5364 = n5003 & n33699 ;
  assign n33700 = ~n5677 ;
  assign n5378 = n33700 & n5352 ;
  assign n5379 = n33696 & n5352 ;
  assign n33701 = ~n5379 ;
  assign n5380 = x77 & n33701 ;
  assign n5381 = n5378 | n5380 ;
  assign n5383 = n5364 | n5381 ;
  assign n33702 = ~n5375 ;
  assign n5384 = n33702 & n5383 ;
  assign n33703 = ~n5384 ;
  assign n5385 = n169 & n33703 ;
  assign n5316 = x76 & n167 ;
  assign n33704 = ~n5316 ;
  assign n5317 = n7327 & n33704 ;
  assign n33705 = ~n5317 ;
  assign n5318 = n168 & n33705 ;
  assign n5319 = n169 | n5318 ;
  assign n33706 = ~n5319 ;
  assign n5387 = n33706 & n5383 ;
  assign n33707 = ~n5004 ;
  assign n5006 = n4934 & n33707 ;
  assign n33708 = ~n4987 ;
  assign n5007 = n33708 & n5006 ;
  assign n33709 = ~n5350 ;
  assign n5414 = n5007 & n33709 ;
  assign n33710 = ~n5349 ;
  assign n5415 = n33710 & n5414 ;
  assign n5416 = n5378 | n5415 ;
  assign n5417 = x78 & n5416 ;
  assign n5418 = x78 | n5415 ;
  assign n5419 = n5378 | n5418 ;
  assign n33711 = ~n5417 ;
  assign n5420 = n33711 & n5419 ;
  assign n5421 = n5387 | n5420 ;
  assign n33712 = ~n5385 ;
  assign n5422 = n33712 & n5421 ;
  assign n33713 = ~n5422 ;
  assign n5423 = n170 & n33713 ;
  assign n4960 = n4940 | n4956 ;
  assign n33714 = ~n4960 ;
  assign n5314 = n33714 & n167 ;
  assign n5315 = n4938 | n5314 ;
  assign n4961 = n4938 & n33714 ;
  assign n5367 = n4961 & n5352 ;
  assign n33715 = ~n5367 ;
  assign n5368 = n5315 & n33715 ;
  assign n5386 = n170 | n5385 ;
  assign n5376 = n169 | n5375 ;
  assign n33716 = ~n5376 ;
  assign n5388 = n33716 & n5383 ;
  assign n5428 = n5388 | n5420 ;
  assign n33717 = ~n5386 ;
  assign n5429 = n33717 & n5428 ;
  assign n5430 = n5368 | n5429 ;
  assign n33718 = ~n5423 ;
  assign n5431 = n33718 & n5430 ;
  assign n33719 = ~n5431 ;
  assign n5432 = n3940 & n33719 ;
  assign n4964 = n4958 | n4963 ;
  assign n33720 = ~n4964 ;
  assign n5300 = n33720 & n167 ;
  assign n5301 = n4998 | n5300 ;
  assign n33721 = ~n4963 ;
  assign n4999 = n33721 & n4998 ;
  assign n5000 = n33534 & n4999 ;
  assign n5355 = n5000 & n5352 ;
  assign n33722 = ~n5355 ;
  assign n5356 = n5301 & n33722 ;
  assign n5425 = n3940 | n5423 ;
  assign n33723 = ~n5425 ;
  assign n5434 = n33723 & n5430 ;
  assign n5435 = n5356 | n5434 ;
  assign n33724 = ~n5432 ;
  assign n5436 = n33724 & n5435 ;
  assign n33725 = ~n5436 ;
  assign n5437 = n172 & n33725 ;
  assign n5067 = n5002 | n5061 ;
  assign n33726 = ~n5067 ;
  assign n5309 = n33726 & n167 ;
  assign n5310 = n5049 | n5309 ;
  assign n5065 = n5049 & n33536 ;
  assign n33727 = ~n5002 ;
  assign n5066 = n33727 & n5065 ;
  assign n5353 = n5066 & n5352 ;
  assign n33728 = ~n5353 ;
  assign n5354 = n5310 & n33728 ;
  assign n5433 = n3631 | n5432 ;
  assign n33729 = ~n5433 ;
  assign n5438 = n33729 & n5435 ;
  assign n5439 = n5354 | n5438 ;
  assign n33730 = ~n5437 ;
  assign n5440 = n33730 & n5439 ;
  assign n33731 = ~n5440 ;
  assign n5441 = n173 & n33731 ;
  assign n5079 = n5063 | n5070 ;
  assign n33732 = ~n5079 ;
  assign n5311 = n33732 & n167 ;
  assign n5312 = n5047 | n5311 ;
  assign n33733 = ~n5070 ;
  assign n5077 = n5047 & n33733 ;
  assign n5078 = n33542 & n5077 ;
  assign n5369 = n5078 & n5352 ;
  assign n33734 = ~n5369 ;
  assign n5370 = n5312 & n33734 ;
  assign n5447 = n171 & n33719 ;
  assign n33735 = ~n5447 ;
  assign n5448 = n5435 & n33735 ;
  assign n33736 = ~n5448 ;
  assign n5449 = n3631 & n33736 ;
  assign n5450 = n173 | n5449 ;
  assign n33737 = ~n5450 ;
  assign n5451 = n5439 & n33737 ;
  assign n5452 = n5370 | n5451 ;
  assign n33738 = ~n5441 ;
  assign n5453 = n33738 & n5452 ;
  assign n33739 = ~n5453 ;
  assign n5454 = n174 & n33739 ;
  assign n5112 = n33548 & n5094 ;
  assign n33740 = ~n5075 ;
  assign n5113 = n33740 & n5112 ;
  assign n5392 = n5113 & n5352 ;
  assign n5076 = n5073 | n5075 ;
  assign n33741 = ~n5076 ;
  assign n5395 = n33741 & n5352 ;
  assign n5396 = n5094 | n5395 ;
  assign n33742 = ~n5392 ;
  assign n5397 = n33742 & n5396 ;
  assign n5442 = n174 | n5441 ;
  assign n33743 = ~n5442 ;
  assign n5455 = n33743 & n5452 ;
  assign n5456 = n5397 | n5455 ;
  assign n33744 = ~n5454 ;
  assign n5457 = n33744 & n5456 ;
  assign n33745 = ~n5457 ;
  assign n5458 = n2753 & n33745 ;
  assign n5111 = n5097 | n5099 ;
  assign n33746 = ~n5111 ;
  assign n5334 = n33746 & n167 ;
  assign n5335 = n5033 | n5334 ;
  assign n33747 = ~n5099 ;
  assign n5109 = n5033 & n33747 ;
  assign n5110 = n33554 & n5109 ;
  assign n5398 = n5110 & n5352 ;
  assign n33748 = ~n5398 ;
  assign n5399 = n5335 & n33748 ;
  assign n33749 = ~n5449 ;
  assign n5466 = n5439 & n33749 ;
  assign n33750 = ~n5466 ;
  assign n5467 = n173 & n33750 ;
  assign n33751 = ~n5467 ;
  assign n5468 = n5452 & n33751 ;
  assign n33752 = ~n5468 ;
  assign n5469 = n174 & n33752 ;
  assign n5470 = n2753 | n5469 ;
  assign n33753 = ~n5470 ;
  assign n5471 = n5456 & n33753 ;
  assign n5472 = n5399 | n5471 ;
  assign n33754 = ~n5458 ;
  assign n5473 = n33754 & n5472 ;
  assign n33755 = ~n5473 ;
  assign n5474 = n176 & n33755 ;
  assign n5129 = n5044 & n33577 ;
  assign n33756 = ~n5103 ;
  assign n5130 = n33756 & n5129 ;
  assign n5304 = n5130 & n167 ;
  assign n5108 = n5102 | n5103 ;
  assign n33757 = ~n5108 ;
  assign n5341 = n33757 & n167 ;
  assign n5342 = n5044 | n5341 ;
  assign n33758 = ~n5304 ;
  assign n5343 = n33758 & n5342 ;
  assign n5459 = n2431 | n5458 ;
  assign n33759 = ~n5459 ;
  assign n5475 = n33759 & n5472 ;
  assign n5476 = n5343 | n5475 ;
  assign n33760 = ~n5474 ;
  assign n5477 = n33760 & n5476 ;
  assign n33761 = ~n5477 ;
  assign n5478 = n177 & n33761 ;
  assign n5128 = n5106 | n5116 ;
  assign n33762 = ~n5128 ;
  assign n5302 = n33762 & n167 ;
  assign n5303 = n4970 | n5302 ;
  assign n33763 = ~n5116 ;
  assign n5126 = n4970 & n33763 ;
  assign n5127 = n33566 & n5126 ;
  assign n5400 = n5127 & n5352 ;
  assign n33764 = ~n5400 ;
  assign n5401 = n5303 & n33764 ;
  assign n33765 = ~n5469 ;
  assign n5486 = n5456 & n33765 ;
  assign n33766 = ~n5486 ;
  assign n5487 = n175 & n33766 ;
  assign n33767 = ~n5487 ;
  assign n5488 = n5472 & n33767 ;
  assign n33768 = ~n5488 ;
  assign n5489 = n2431 & n33768 ;
  assign n5490 = n177 | n5489 ;
  assign n33769 = ~n5490 ;
  assign n5491 = n5476 & n33769 ;
  assign n5492 = n5401 | n5491 ;
  assign n33770 = ~n5478 ;
  assign n5493 = n33770 & n5492 ;
  assign n33771 = ~n5493 ;
  assign n5494 = n178 & n33771 ;
  assign n5125 = n5119 | n5120 ;
  assign n33772 = ~n5125 ;
  assign n5296 = n33772 & n167 ;
  assign n5297 = n5018 | n5296 ;
  assign n5149 = n5018 & n33593 ;
  assign n33773 = ~n5120 ;
  assign n5150 = n33773 & n5149 ;
  assign n5320 = n5150 & n167 ;
  assign n33774 = ~n5320 ;
  assign n5321 = n5297 & n33774 ;
  assign n5479 = n178 | n5478 ;
  assign n33775 = ~n5479 ;
  assign n5495 = n33775 & n5492 ;
  assign n5496 = n5321 | n5495 ;
  assign n33776 = ~n5494 ;
  assign n5497 = n33776 & n5496 ;
  assign n33777 = ~n5497 ;
  assign n5498 = n1707 & n33777 ;
  assign n5148 = n5123 | n5136 ;
  assign n33778 = ~n5148 ;
  assign n5298 = n33778 & n167 ;
  assign n5299 = n5030 | n5298 ;
  assign n33779 = ~n5136 ;
  assign n5146 = n5030 & n33779 ;
  assign n5147 = n33582 & n5146 ;
  assign n5390 = n5147 & n5352 ;
  assign n33780 = ~n5390 ;
  assign n5391 = n5299 & n33780 ;
  assign n33781 = ~n5489 ;
  assign n5506 = n5476 & n33781 ;
  assign n33782 = ~n5506 ;
  assign n5507 = n177 & n33782 ;
  assign n33783 = ~n5507 ;
  assign n5508 = n5492 & n33783 ;
  assign n33784 = ~n5508 ;
  assign n5509 = n178 & n33784 ;
  assign n5510 = n1707 | n5509 ;
  assign n33785 = ~n5510 ;
  assign n5511 = n5496 & n33785 ;
  assign n5512 = n5391 | n5511 ;
  assign n33786 = ~n5498 ;
  assign n5513 = n33786 & n5512 ;
  assign n33787 = ~n5513 ;
  assign n5514 = n180 & n33787 ;
  assign n5145 = n5139 | n5140 ;
  assign n33788 = ~n5145 ;
  assign n5402 = n33788 & n5352 ;
  assign n5403 = n5015 | n5402 ;
  assign n5169 = n5015 & n33609 ;
  assign n33789 = ~n5140 ;
  assign n5170 = n33789 & n5169 ;
  assign n5404 = n5170 & n5352 ;
  assign n33790 = ~n5404 ;
  assign n5405 = n5403 & n33790 ;
  assign n5499 = n1487 | n5498 ;
  assign n33791 = ~n5499 ;
  assign n5515 = n33791 & n5512 ;
  assign n5516 = n5405 | n5515 ;
  assign n33792 = ~n5514 ;
  assign n5517 = n33792 & n5516 ;
  assign n33793 = ~n5517 ;
  assign n5518 = n181 & n33793 ;
  assign n5168 = n5143 | n5156 ;
  assign n33794 = ~n5168 ;
  assign n5365 = n33794 & n5352 ;
  assign n5366 = n5027 | n5365 ;
  assign n33795 = ~n5156 ;
  assign n5166 = n5027 & n33795 ;
  assign n5167 = n33598 & n5166 ;
  assign n5406 = n5167 & n5352 ;
  assign n33796 = ~n5406 ;
  assign n5407 = n5366 & n33796 ;
  assign n33797 = ~n5509 ;
  assign n5526 = n5496 & n33797 ;
  assign n33798 = ~n5526 ;
  assign n5527 = n179 & n33798 ;
  assign n33799 = ~n5527 ;
  assign n5528 = n5512 & n33799 ;
  assign n33800 = ~n5528 ;
  assign n5529 = n1487 & n33800 ;
  assign n5530 = n181 | n5529 ;
  assign n33801 = ~n5530 ;
  assign n5531 = n5516 & n33801 ;
  assign n5532 = n5407 | n5531 ;
  assign n33802 = ~n5518 ;
  assign n5533 = n33802 & n5532 ;
  assign n33803 = ~n5533 ;
  assign n5534 = n182 & n33803 ;
  assign n5165 = n5159 | n5160 ;
  assign n33804 = ~n5165 ;
  assign n5339 = n33804 & n167 ;
  assign n5340 = n5021 | n5339 ;
  assign n5189 = n5021 & n33625 ;
  assign n33805 = ~n5160 ;
  assign n5190 = n33805 & n5189 ;
  assign n5357 = n5190 & n5352 ;
  assign n33806 = ~n5357 ;
  assign n5358 = n5340 & n33806 ;
  assign n5519 = n182 | n5518 ;
  assign n33807 = ~n5519 ;
  assign n5535 = n33807 & n5532 ;
  assign n5536 = n5358 | n5535 ;
  assign n33808 = ~n5534 ;
  assign n5537 = n33808 & n5536 ;
  assign n33809 = ~n5537 ;
  assign n5538 = n996 & n33809 ;
  assign n5188 = n5163 | n5176 ;
  assign n33810 = ~n5188 ;
  assign n5328 = n33810 & n167 ;
  assign n5329 = n5036 | n5328 ;
  assign n33811 = ~n5176 ;
  assign n5186 = n5036 & n33811 ;
  assign n5187 = n33614 & n5186 ;
  assign n5359 = n5187 & n5352 ;
  assign n33812 = ~n5359 ;
  assign n5360 = n5329 & n33812 ;
  assign n33813 = ~n5529 ;
  assign n5546 = n5516 & n33813 ;
  assign n33814 = ~n5546 ;
  assign n5547 = n181 & n33814 ;
  assign n33815 = ~n5547 ;
  assign n5548 = n5532 & n33815 ;
  assign n33816 = ~n5548 ;
  assign n5549 = n182 & n33816 ;
  assign n5550 = n183 | n5549 ;
  assign n33817 = ~n5550 ;
  assign n5551 = n5536 & n33817 ;
  assign n5552 = n5360 | n5551 ;
  assign n33818 = ~n5538 ;
  assign n5553 = n33818 & n5552 ;
  assign n33819 = ~n5553 ;
  assign n5554 = n184 & n33819 ;
  assign n5185 = n5179 | n5180 ;
  assign n33820 = ~n5185 ;
  assign n5322 = n33820 & n167 ;
  assign n5323 = n5041 | n5322 ;
  assign n5208 = n5041 & n33641 ;
  assign n33821 = ~n5180 ;
  assign n5209 = n33821 & n5208 ;
  assign n5408 = n5209 & n5352 ;
  assign n33822 = ~n5408 ;
  assign n5409 = n5323 & n33822 ;
  assign n5539 = n838 | n5538 ;
  assign n33823 = ~n5539 ;
  assign n5555 = n33823 & n5552 ;
  assign n5556 = n5409 | n5555 ;
  assign n33824 = ~n5554 ;
  assign n5557 = n33824 & n5556 ;
  assign n33825 = ~n5557 ;
  assign n5558 = n185 & n33825 ;
  assign n5207 = n5183 | n5196 ;
  assign n33826 = ~n5207 ;
  assign n5324 = n33826 & n167 ;
  assign n5325 = n4976 | n5324 ;
  assign n33827 = ~n5196 ;
  assign n5205 = n4976 & n33827 ;
  assign n5206 = n33630 & n5205 ;
  assign n5410 = n5206 & n5352 ;
  assign n33828 = ~n5410 ;
  assign n5411 = n5325 & n33828 ;
  assign n33829 = ~n5549 ;
  assign n5566 = n5536 & n33829 ;
  assign n33830 = ~n5566 ;
  assign n5567 = n183 & n33830 ;
  assign n33831 = ~n5567 ;
  assign n5568 = n5552 & n33831 ;
  assign n33832 = ~n5568 ;
  assign n5569 = n838 & n33832 ;
  assign n5570 = n185 | n5569 ;
  assign n33833 = ~n5570 ;
  assign n5571 = n5556 & n33833 ;
  assign n5572 = n5411 | n5571 ;
  assign n33834 = ~n5558 ;
  assign n5573 = n33834 & n5572 ;
  assign n33835 = ~n5573 ;
  assign n5574 = n186 & n33835 ;
  assign n5229 = n5200 | n5213 ;
  assign n33836 = ~n5229 ;
  assign n5326 = n33836 & n167 ;
  assign n5327 = n5082 | n5326 ;
  assign n5227 = n5082 & n33657 ;
  assign n33837 = ~n5200 ;
  assign n5228 = n33837 & n5227 ;
  assign n5371 = n5228 & n5352 ;
  assign n33838 = ~n5371 ;
  assign n5372 = n5327 & n33838 ;
  assign n5559 = n186 | n5558 ;
  assign n33839 = ~n5559 ;
  assign n5575 = n33839 & n5572 ;
  assign n5576 = n5372 | n5575 ;
  assign n33840 = ~n5574 ;
  assign n5577 = n33840 & n5576 ;
  assign n33841 = ~n5577 ;
  assign n5578 = n528 & n33841 ;
  assign n5226 = n5203 | n5215 ;
  assign n33842 = ~n5226 ;
  assign n5307 = n33842 & n167 ;
  assign n5308 = n5088 | n5307 ;
  assign n33843 = ~n5215 ;
  assign n5224 = n5088 & n33843 ;
  assign n5225 = n33646 & n5224 ;
  assign n5412 = n5225 & n5352 ;
  assign n33844 = ~n5412 ;
  assign n5413 = n5308 & n33844 ;
  assign n33845 = ~n5569 ;
  assign n5586 = n5556 & n33845 ;
  assign n33846 = ~n5586 ;
  assign n5587 = n185 & n33846 ;
  assign n33847 = ~n5587 ;
  assign n5588 = n5572 & n33847 ;
  assign n33848 = ~n5588 ;
  assign n5589 = n186 & n33848 ;
  assign n5590 = n528 | n5589 ;
  assign n33849 = ~n5590 ;
  assign n5591 = n5576 & n33849 ;
  assign n5592 = n5413 | n5591 ;
  assign n33850 = ~n5578 ;
  assign n5593 = n33850 & n5592 ;
  assign n33851 = ~n5593 ;
  assign n5594 = n188 & n33851 ;
  assign n5250 = n5219 | n5233 ;
  assign n33852 = ~n5250 ;
  assign n5330 = n33852 & n167 ;
  assign n5331 = n5085 | n5330 ;
  assign n5248 = n5085 & n33663 ;
  assign n33853 = ~n5219 ;
  assign n5249 = n33853 & n5248 ;
  assign n5361 = n5249 & n5352 ;
  assign n33854 = ~n5361 ;
  assign n5362 = n5331 & n33854 ;
  assign n5579 = n413 | n5578 ;
  assign n33855 = ~n5579 ;
  assign n5595 = n33855 & n5592 ;
  assign n5597 = n5362 | n5595 ;
  assign n33856 = ~n5594 ;
  assign n5598 = n33856 & n5597 ;
  assign n33857 = ~n5598 ;
  assign n5599 = n189 & n33857 ;
  assign n5247 = n5222 | n5235 ;
  assign n33858 = ~n5247 ;
  assign n5332 = n33858 & n167 ;
  assign n5333 = n5091 | n5332 ;
  assign n33859 = ~n5235 ;
  assign n5245 = n5091 & n33859 ;
  assign n5246 = n33678 & n5245 ;
  assign n5393 = n5246 & n5352 ;
  assign n33860 = ~n5393 ;
  assign n5394 = n5333 & n33860 ;
  assign n33861 = ~n5589 ;
  assign n5606 = n5576 & n33861 ;
  assign n33862 = ~n5606 ;
  assign n5607 = n187 & n33862 ;
  assign n33863 = ~n5607 ;
  assign n5608 = n5592 & n33863 ;
  assign n33864 = ~n5608 ;
  assign n5609 = n413 & n33864 ;
  assign n5610 = n189 | n5609 ;
  assign n33865 = ~n5610 ;
  assign n5611 = n5597 & n33865 ;
  assign n5612 = n5394 | n5611 ;
  assign n33866 = ~n5599 ;
  assign n5613 = n33866 & n5612 ;
  assign n33867 = ~n5613 ;
  assign n5614 = n190 & n33867 ;
  assign n5260 = n5239 | n5254 ;
  assign n33868 = ~n5260 ;
  assign n5305 = n33868 & n167 ;
  assign n5306 = n5024 | n5305 ;
  assign n5258 = n5024 & n33667 ;
  assign n33869 = ~n5239 ;
  assign n5259 = n33869 & n5258 ;
  assign n5336 = n5259 & n167 ;
  assign n33870 = ~n5336 ;
  assign n5337 = n5306 & n33870 ;
  assign n5600 = n190 | n5599 ;
  assign n33871 = ~n5600 ;
  assign n5615 = n33871 & n5612 ;
  assign n5616 = n5337 | n5615 ;
  assign n33872 = ~n5614 ;
  assign n5617 = n33872 & n5616 ;
  assign n33873 = ~n5617 ;
  assign n5618 = n287 & n33873 ;
  assign n33874 = ~n5609 ;
  assign n5625 = n5597 & n33874 ;
  assign n33875 = ~n5625 ;
  assign n5626 = n189 & n33875 ;
  assign n33876 = ~n5626 ;
  assign n5627 = n5612 & n33876 ;
  assign n33877 = ~n5627 ;
  assign n5628 = n190 & n33877 ;
  assign n5629 = n287 | n5628 ;
  assign n33878 = ~n5629 ;
  assign n5630 = n5616 & n33878 ;
  assign n33879 = ~n5256 ;
  assign n5662 = n33879 & n5281 ;
  assign n5663 = n33691 & n5662 ;
  assign n5664 = n167 & n5663 ;
  assign n5257 = n5242 | n5256 ;
  assign n33880 = ~n5257 ;
  assign n5338 = n33880 & n167 ;
  assign n5665 = n5281 | n5338 ;
  assign n33881 = ~n5664 ;
  assign n5666 = n33881 & n5665 ;
  assign n5669 = n5630 | n5666 ;
  assign n33882 = ~n5618 ;
  assign n5670 = n33882 & n5669 ;
  assign n5671 = n5658 | n5670 ;
  assign n5672 = n31336 & n5671 ;
  assign n5266 = n5004 | n5265 ;
  assign n33883 = ~n5266 ;
  assign n5272 = n33883 & n5269 ;
  assign n5273 = n33708 & n5272 ;
  assign n5638 = n5273 & n33709 ;
  assign n5639 = n33710 & n5638 ;
  assign n33884 = ~n5270 ;
  assign n5313 = n33884 & n167 ;
  assign n33885 = ~n5313 ;
  assign n5642 = n33885 & n5347 ;
  assign n5646 = n192 & n5643 ;
  assign n33886 = ~n5642 ;
  assign n5647 = n33886 & n5646 ;
  assign n5648 = n5639 | n5647 ;
  assign n5659 = n33882 & n5657 ;
  assign n5675 = n5659 & n5669 ;
  assign n5676 = n5648 | n5675 ;
  assign n166 = n5672 | n5676 ;
  assign n8390 = x72 | x73 ;
  assign n8926 = x74 | n8390 ;
  assign n5688 = x74 & n166 ;
  assign n33887 = ~n5688 ;
  assign n5752 = n8926 & n33887 ;
  assign n33888 = ~n5752 ;
  assign n5753 = n167 & n33888 ;
  assign n5008 = n8926 & n33707 ;
  assign n5009 = n33708 & n5008 ;
  assign n5636 = n5009 & n33709 ;
  assign n5637 = n33710 & n5636 ;
  assign n5689 = n5637 & n33887 ;
  assign n33889 = ~n6933 ;
  assign n5680 = n33889 & n166 ;
  assign n33890 = ~x74 ;
  assign n5787 = n33890 & n166 ;
  assign n33891 = ~n5787 ;
  assign n5788 = x75 & n33891 ;
  assign n5789 = n5680 | n5788 ;
  assign n5790 = n5689 | n5789 ;
  assign n33892 = ~n5753 ;
  assign n5793 = n33892 & n5790 ;
  assign n33893 = ~n5793 ;
  assign n5794 = n4934 & n33893 ;
  assign n9416 = n33890 & n8390 ;
  assign n33894 = ~n166 ;
  assign n5684 = x74 & n33894 ;
  assign n5685 = n9416 | n5684 ;
  assign n33895 = ~n5685 ;
  assign n5686 = n5352 & n33895 ;
  assign n5687 = n4934 | n5686 ;
  assign n33896 = ~n5687 ;
  assign n5791 = n33896 & n5790 ;
  assign n33897 = ~n5639 ;
  assign n5640 = n5352 & n33897 ;
  assign n33898 = ~n5647 ;
  assign n5649 = n5640 & n33898 ;
  assign n33899 = ~n5675 ;
  assign n5799 = n5649 & n33899 ;
  assign n33900 = ~n5672 ;
  assign n5800 = n33900 & n5799 ;
  assign n5801 = n5680 | n5800 ;
  assign n5802 = x76 & n5801 ;
  assign n5803 = x76 | n5800 ;
  assign n5804 = n5680 | n5803 ;
  assign n33901 = ~n5802 ;
  assign n5805 = n33901 & n5804 ;
  assign n5806 = n5791 | n5805 ;
  assign n33902 = ~n5794 ;
  assign n5807 = n33902 & n5806 ;
  assign n33903 = ~n5807 ;
  assign n5808 = n169 & n33903 ;
  assign n5377 = n5364 | n5375 ;
  assign n33904 = ~n5377 ;
  assign n5382 = n33904 & n5381 ;
  assign n5691 = n5382 & n166 ;
  assign n5733 = n33904 & n166 ;
  assign n5734 = n5381 | n5733 ;
  assign n33905 = ~n5691 ;
  assign n5735 = n33905 & n5734 ;
  assign n5795 = n169 | n5794 ;
  assign n33906 = ~n5795 ;
  assign n5811 = n33906 & n5806 ;
  assign n5812 = n5735 | n5811 ;
  assign n33907 = ~n5808 ;
  assign n5813 = n33907 & n5812 ;
  assign n33908 = ~n5813 ;
  assign n5814 = n170 & n33908 ;
  assign n33909 = ~n5388 ;
  assign n5426 = n33909 & n5420 ;
  assign n5427 = n33712 & n5426 ;
  assign n5731 = n5427 & n166 ;
  assign n5389 = n5385 | n5388 ;
  assign n33910 = ~n5389 ;
  assign n5761 = n33910 & n166 ;
  assign n5762 = n5420 | n5761 ;
  assign n33911 = ~n5731 ;
  assign n5763 = n33911 & n5762 ;
  assign n5809 = n170 | n5808 ;
  assign n33912 = ~n5809 ;
  assign n5815 = n33912 & n5812 ;
  assign n5816 = n5763 | n5815 ;
  assign n33913 = ~n5814 ;
  assign n5817 = n33913 & n5816 ;
  assign n33914 = ~n5817 ;
  assign n5818 = n3940 & n33914 ;
  assign n5424 = n5368 & n33718 ;
  assign n33915 = ~n5429 ;
  assign n5634 = n5424 & n33915 ;
  assign n5678 = n5634 & n166 ;
  assign n5635 = n5423 | n5429 ;
  assign n33916 = ~n5635 ;
  assign n5724 = n33916 & n166 ;
  assign n5725 = n5368 | n5724 ;
  assign n33917 = ~n5678 ;
  assign n5726 = n33917 & n5725 ;
  assign n5796 = n168 & n33893 ;
  assign n5754 = n168 | n5753 ;
  assign n33918 = ~n5754 ;
  assign n5798 = n33918 & n5790 ;
  assign n5827 = n5798 | n5805 ;
  assign n33919 = ~n5796 ;
  assign n5828 = n33919 & n5827 ;
  assign n33920 = ~n5828 ;
  assign n5829 = n169 & n33920 ;
  assign n5830 = n33906 & n5827 ;
  assign n5831 = n5735 | n5830 ;
  assign n33921 = ~n5829 ;
  assign n5832 = n33921 & n5831 ;
  assign n33922 = ~n5832 ;
  assign n5833 = n170 & n33922 ;
  assign n5834 = n3940 | n5833 ;
  assign n33923 = ~n5834 ;
  assign n5835 = n5816 & n33923 ;
  assign n5836 = n5726 | n5835 ;
  assign n33924 = ~n5818 ;
  assign n5837 = n33924 & n5836 ;
  assign n33925 = ~n5837 ;
  assign n5838 = n172 & n33925 ;
  assign n5446 = n5432 | n5434 ;
  assign n33926 = ~n5446 ;
  assign n5742 = n33926 & n166 ;
  assign n5743 = n5356 | n5742 ;
  assign n33927 = ~n5434 ;
  assign n5444 = n5356 & n33927 ;
  assign n5445 = n33724 & n5444 ;
  assign n5744 = n5445 & n166 ;
  assign n33928 = ~n5744 ;
  assign n5745 = n5743 & n33928 ;
  assign n5819 = n3631 | n5818 ;
  assign n33929 = ~n5819 ;
  assign n5839 = n33929 & n5836 ;
  assign n5840 = n5745 | n5839 ;
  assign n33930 = ~n5838 ;
  assign n5841 = n33930 & n5840 ;
  assign n33931 = ~n5841 ;
  assign n5842 = n173 & n33931 ;
  assign n5464 = n5354 & n33749 ;
  assign n33932 = ~n5438 ;
  assign n5465 = n33932 & n5464 ;
  assign n5732 = n5465 & n166 ;
  assign n5443 = n5437 | n5438 ;
  assign n33933 = ~n5443 ;
  assign n5764 = n33933 & n166 ;
  assign n5765 = n5354 | n5764 ;
  assign n33934 = ~n5732 ;
  assign n5766 = n33934 & n5765 ;
  assign n5850 = n33912 & n5831 ;
  assign n5851 = n5763 | n5850 ;
  assign n33935 = ~n5833 ;
  assign n5852 = n33935 & n5851 ;
  assign n33936 = ~n5852 ;
  assign n5853 = n171 & n33936 ;
  assign n5854 = n33923 & n5851 ;
  assign n5855 = n5726 | n5854 ;
  assign n33937 = ~n5853 ;
  assign n5856 = n33937 & n5855 ;
  assign n33938 = ~n5856 ;
  assign n5857 = n3631 & n33938 ;
  assign n5858 = n173 | n5857 ;
  assign n33939 = ~n5858 ;
  assign n5859 = n5840 & n33939 ;
  assign n5860 = n5766 | n5859 ;
  assign n33940 = ~n5842 ;
  assign n5861 = n33940 & n5860 ;
  assign n33941 = ~n5861 ;
  assign n5862 = n174 & n33941 ;
  assign n33942 = ~n5451 ;
  assign n5461 = n5370 & n33942 ;
  assign n5462 = n33738 & n5461 ;
  assign n5739 = n5462 & n166 ;
  assign n5463 = n5441 | n5451 ;
  assign n33943 = ~n5463 ;
  assign n5758 = n33943 & n166 ;
  assign n5759 = n5370 | n5758 ;
  assign n33944 = ~n5739 ;
  assign n5760 = n33944 & n5759 ;
  assign n5843 = n174 | n5842 ;
  assign n33945 = ~n5843 ;
  assign n5863 = n33945 & n5860 ;
  assign n5866 = n5760 | n5863 ;
  assign n33946 = ~n5862 ;
  assign n5867 = n33946 & n5866 ;
  assign n33947 = ~n5867 ;
  assign n5868 = n2753 & n33947 ;
  assign n5460 = n5454 | n5455 ;
  assign n33948 = ~n5460 ;
  assign n5750 = n33948 & n166 ;
  assign n5751 = n5397 | n5750 ;
  assign n5484 = n5397 & n33765 ;
  assign n33949 = ~n5455 ;
  assign n5485 = n33949 & n5484 ;
  assign n5767 = n5485 & n166 ;
  assign n33950 = ~n5767 ;
  assign n5768 = n5751 & n33950 ;
  assign n5874 = n33929 & n5855 ;
  assign n5875 = n5745 | n5874 ;
  assign n33951 = ~n5857 ;
  assign n5876 = n33951 & n5875 ;
  assign n33952 = ~n5876 ;
  assign n5877 = n173 & n33952 ;
  assign n5878 = n33939 & n5875 ;
  assign n5879 = n5766 | n5878 ;
  assign n33953 = ~n5877 ;
  assign n5880 = n33953 & n5879 ;
  assign n33954 = ~n5880 ;
  assign n5881 = n174 & n33954 ;
  assign n5882 = n2753 | n5881 ;
  assign n33955 = ~n5882 ;
  assign n5883 = n5866 & n33955 ;
  assign n5884 = n5768 | n5883 ;
  assign n33956 = ~n5868 ;
  assign n5885 = n33956 & n5884 ;
  assign n33957 = ~n5885 ;
  assign n5886 = n176 & n33957 ;
  assign n5483 = n5458 | n5471 ;
  assign n33958 = ~n5483 ;
  assign n5771 = n33958 & n166 ;
  assign n5772 = n5399 | n5771 ;
  assign n33959 = ~n5471 ;
  assign n5481 = n5399 & n33959 ;
  assign n5482 = n33754 & n5481 ;
  assign n5773 = n5482 & n166 ;
  assign n33960 = ~n5773 ;
  assign n5774 = n5772 & n33960 ;
  assign n5869 = n2431 | n5868 ;
  assign n33961 = ~n5869 ;
  assign n5887 = n33961 & n5884 ;
  assign n5888 = n5774 | n5887 ;
  assign n33962 = ~n5886 ;
  assign n5889 = n33962 & n5888 ;
  assign n33963 = ~n5889 ;
  assign n5890 = n177 & n33963 ;
  assign n5504 = n5343 & n33781 ;
  assign n33964 = ~n5475 ;
  assign n5505 = n33964 & n5504 ;
  assign n5693 = n5505 & n166 ;
  assign n5480 = n5474 | n5475 ;
  assign n33965 = ~n5480 ;
  assign n5755 = n33965 & n166 ;
  assign n5756 = n5343 | n5755 ;
  assign n33966 = ~n5693 ;
  assign n5757 = n33966 & n5756 ;
  assign n5898 = n33945 & n5879 ;
  assign n5899 = n5760 | n5898 ;
  assign n33967 = ~n5881 ;
  assign n5900 = n33967 & n5899 ;
  assign n33968 = ~n5900 ;
  assign n5901 = n175 & n33968 ;
  assign n5902 = n33955 & n5899 ;
  assign n5903 = n5768 | n5902 ;
  assign n33969 = ~n5901 ;
  assign n5904 = n33969 & n5903 ;
  assign n33970 = ~n5904 ;
  assign n5905 = n2431 & n33970 ;
  assign n5906 = n177 | n5905 ;
  assign n33971 = ~n5906 ;
  assign n5907 = n5888 & n33971 ;
  assign n5908 = n5757 | n5907 ;
  assign n33972 = ~n5890 ;
  assign n5909 = n33972 & n5908 ;
  assign n33973 = ~n5909 ;
  assign n5910 = n178 & n33973 ;
  assign n33974 = ~n5491 ;
  assign n5501 = n5401 & n33974 ;
  assign n5502 = n33770 & n5501 ;
  assign n5736 = n5502 & n166 ;
  assign n5503 = n5478 | n5491 ;
  assign n33975 = ~n5503 ;
  assign n5780 = n33975 & n166 ;
  assign n5781 = n5401 | n5780 ;
  assign n33976 = ~n5736 ;
  assign n5782 = n33976 & n5781 ;
  assign n5891 = n178 | n5890 ;
  assign n33977 = ~n5891 ;
  assign n5911 = n33977 & n5908 ;
  assign n5912 = n5782 | n5911 ;
  assign n33978 = ~n5910 ;
  assign n5913 = n33978 & n5912 ;
  assign n33979 = ~n5913 ;
  assign n5914 = n1707 & n33979 ;
  assign n5500 = n5494 | n5495 ;
  assign n33980 = ~n5500 ;
  assign n5727 = n33980 & n166 ;
  assign n5728 = n5321 | n5727 ;
  assign n5524 = n5321 & n33797 ;
  assign n33981 = ~n5495 ;
  assign n5525 = n33981 & n5524 ;
  assign n5746 = n5525 & n166 ;
  assign n33982 = ~n5746 ;
  assign n5747 = n5728 & n33982 ;
  assign n5922 = n33961 & n5903 ;
  assign n5923 = n5774 | n5922 ;
  assign n33983 = ~n5905 ;
  assign n5924 = n33983 & n5923 ;
  assign n33984 = ~n5924 ;
  assign n5925 = n177 & n33984 ;
  assign n5926 = n33971 & n5923 ;
  assign n5927 = n5757 | n5926 ;
  assign n33985 = ~n5925 ;
  assign n5928 = n33985 & n5927 ;
  assign n33986 = ~n5928 ;
  assign n5929 = n178 & n33986 ;
  assign n5930 = n1707 | n5929 ;
  assign n33987 = ~n5930 ;
  assign n5931 = n5912 & n33987 ;
  assign n5932 = n5747 | n5931 ;
  assign n33988 = ~n5914 ;
  assign n5933 = n33988 & n5932 ;
  assign n33989 = ~n5933 ;
  assign n5934 = n180 & n33989 ;
  assign n5523 = n5498 | n5511 ;
  assign n33990 = ~n5523 ;
  assign n5712 = n33990 & n166 ;
  assign n5713 = n5391 | n5712 ;
  assign n33991 = ~n5511 ;
  assign n5521 = n5391 & n33991 ;
  assign n5522 = n33786 & n5521 ;
  assign n5778 = n5522 & n166 ;
  assign n33992 = ~n5778 ;
  assign n5779 = n5713 & n33992 ;
  assign n5915 = n1487 | n5914 ;
  assign n33993 = ~n5915 ;
  assign n5935 = n33993 & n5932 ;
  assign n5936 = n5779 | n5935 ;
  assign n33994 = ~n5934 ;
  assign n5937 = n33994 & n5936 ;
  assign n33995 = ~n5937 ;
  assign n5938 = n181 & n33995 ;
  assign n5520 = n5514 | n5515 ;
  assign n33996 = ~n5520 ;
  assign n5769 = n33996 & n166 ;
  assign n5770 = n5405 | n5769 ;
  assign n5544 = n5405 & n33813 ;
  assign n33997 = ~n5515 ;
  assign n5545 = n33997 & n5544 ;
  assign n5785 = n5545 & n166 ;
  assign n33998 = ~n5785 ;
  assign n5786 = n5770 & n33998 ;
  assign n5946 = n33977 & n5927 ;
  assign n5947 = n5782 | n5946 ;
  assign n33999 = ~n5929 ;
  assign n5948 = n33999 & n5947 ;
  assign n34000 = ~n5948 ;
  assign n5949 = n179 & n34000 ;
  assign n5950 = n33987 & n5947 ;
  assign n5951 = n5747 | n5950 ;
  assign n34001 = ~n5949 ;
  assign n5952 = n34001 & n5951 ;
  assign n34002 = ~n5952 ;
  assign n5953 = n1487 & n34002 ;
  assign n5954 = n181 | n5953 ;
  assign n34003 = ~n5954 ;
  assign n5955 = n5936 & n34003 ;
  assign n5956 = n5786 | n5955 ;
  assign n34004 = ~n5938 ;
  assign n5957 = n34004 & n5956 ;
  assign n34005 = ~n5957 ;
  assign n5958 = n182 & n34005 ;
  assign n34006 = ~n5531 ;
  assign n5541 = n5407 & n34006 ;
  assign n5542 = n33802 & n5541 ;
  assign n5723 = n5542 & n166 ;
  assign n5543 = n5518 | n5531 ;
  assign n34007 = ~n5543 ;
  assign n5775 = n34007 & n166 ;
  assign n5776 = n5407 | n5775 ;
  assign n34008 = ~n5723 ;
  assign n5777 = n34008 & n5776 ;
  assign n5939 = n182 | n5938 ;
  assign n34009 = ~n5939 ;
  assign n5959 = n34009 & n5956 ;
  assign n5960 = n5777 | n5959 ;
  assign n34010 = ~n5958 ;
  assign n5961 = n34010 & n5960 ;
  assign n34011 = ~n5961 ;
  assign n5962 = n996 & n34011 ;
  assign n5564 = n5358 & n33829 ;
  assign n34012 = ~n5535 ;
  assign n5565 = n34012 & n5564 ;
  assign n5718 = n5565 & n166 ;
  assign n5540 = n5534 | n5535 ;
  assign n34013 = ~n5540 ;
  assign n5719 = n34013 & n166 ;
  assign n5720 = n5358 | n5719 ;
  assign n34014 = ~n5718 ;
  assign n5721 = n34014 & n5720 ;
  assign n5970 = n33993 & n5951 ;
  assign n5971 = n5779 | n5970 ;
  assign n34015 = ~n5953 ;
  assign n5972 = n34015 & n5971 ;
  assign n34016 = ~n5972 ;
  assign n5973 = n181 & n34016 ;
  assign n5974 = n34003 & n5971 ;
  assign n5975 = n5786 | n5974 ;
  assign n34017 = ~n5973 ;
  assign n5976 = n34017 & n5975 ;
  assign n34018 = ~n5976 ;
  assign n5977 = n182 & n34018 ;
  assign n5978 = n183 | n5977 ;
  assign n34019 = ~n5978 ;
  assign n5979 = n5960 & n34019 ;
  assign n5980 = n5721 | n5979 ;
  assign n34020 = ~n5962 ;
  assign n5981 = n34020 & n5980 ;
  assign n34021 = ~n5981 ;
  assign n5982 = n184 & n34021 ;
  assign n5561 = n5538 | n5551 ;
  assign n34022 = ~n5561 ;
  assign n5714 = n34022 & n166 ;
  assign n5715 = n5360 | n5714 ;
  assign n34023 = ~n5551 ;
  assign n5562 = n5360 & n34023 ;
  assign n5563 = n33818 & n5562 ;
  assign n5748 = n5563 & n166 ;
  assign n34024 = ~n5748 ;
  assign n5749 = n5715 & n34024 ;
  assign n5963 = n838 | n5962 ;
  assign n34025 = ~n5963 ;
  assign n5983 = n34025 & n5980 ;
  assign n5984 = n5749 | n5983 ;
  assign n34026 = ~n5982 ;
  assign n5985 = n34026 & n5984 ;
  assign n34027 = ~n5985 ;
  assign n5986 = n185 & n34027 ;
  assign n5560 = n5554 | n5555 ;
  assign n34028 = ~n5560 ;
  assign n5729 = n34028 & n166 ;
  assign n5730 = n5409 | n5729 ;
  assign n5584 = n5409 & n33845 ;
  assign n34029 = ~n5555 ;
  assign n5585 = n34029 & n5584 ;
  assign n5783 = n5585 & n166 ;
  assign n34030 = ~n5783 ;
  assign n5784 = n5730 & n34030 ;
  assign n5994 = n34009 & n5975 ;
  assign n5995 = n5777 | n5994 ;
  assign n34031 = ~n5977 ;
  assign n5996 = n34031 & n5995 ;
  assign n34032 = ~n5996 ;
  assign n5997 = n183 & n34032 ;
  assign n5998 = n34019 & n5995 ;
  assign n5999 = n5721 | n5998 ;
  assign n34033 = ~n5997 ;
  assign n6000 = n34033 & n5999 ;
  assign n34034 = ~n6000 ;
  assign n6001 = n838 & n34034 ;
  assign n6002 = n185 | n6001 ;
  assign n34035 = ~n6002 ;
  assign n6003 = n5984 & n34035 ;
  assign n6004 = n5784 | n6003 ;
  assign n34036 = ~n5986 ;
  assign n6005 = n34036 & n6004 ;
  assign n34037 = ~n6005 ;
  assign n6006 = n186 & n34037 ;
  assign n34038 = ~n5571 ;
  assign n5582 = n5411 & n34038 ;
  assign n5583 = n33834 & n5582 ;
  assign n5708 = n5583 & n166 ;
  assign n5581 = n5558 | n5571 ;
  assign n34039 = ~n5581 ;
  assign n5709 = n34039 & n166 ;
  assign n5710 = n5411 | n5709 ;
  assign n34040 = ~n5708 ;
  assign n5711 = n34040 & n5710 ;
  assign n5987 = n186 | n5986 ;
  assign n34041 = ~n5987 ;
  assign n6007 = n34041 & n6004 ;
  assign n6008 = n5711 | n6007 ;
  assign n34042 = ~n6006 ;
  assign n6009 = n34042 & n6008 ;
  assign n34043 = ~n6009 ;
  assign n6010 = n528 & n34043 ;
  assign n5580 = n5574 | n5575 ;
  assign n34044 = ~n5580 ;
  assign n5700 = n34044 & n166 ;
  assign n5701 = n5372 | n5700 ;
  assign n5604 = n5372 & n33861 ;
  assign n34045 = ~n5575 ;
  assign n5605 = n34045 & n5604 ;
  assign n5706 = n5605 & n166 ;
  assign n34046 = ~n5706 ;
  assign n5707 = n5701 & n34046 ;
  assign n6018 = n34025 & n5999 ;
  assign n6019 = n5749 | n6018 ;
  assign n34047 = ~n6001 ;
  assign n6020 = n34047 & n6019 ;
  assign n34048 = ~n6020 ;
  assign n6021 = n185 & n34048 ;
  assign n6022 = n34035 & n6019 ;
  assign n6023 = n5784 | n6022 ;
  assign n34049 = ~n6021 ;
  assign n6024 = n34049 & n6023 ;
  assign n34050 = ~n6024 ;
  assign n6025 = n186 & n34050 ;
  assign n6026 = n528 | n6025 ;
  assign n34051 = ~n6026 ;
  assign n6027 = n6008 & n34051 ;
  assign n6028 = n5707 | n6027 ;
  assign n34052 = ~n6010 ;
  assign n6029 = n34052 & n6028 ;
  assign n34053 = ~n6029 ;
  assign n6030 = n188 & n34053 ;
  assign n5603 = n5578 | n5591 ;
  assign n34054 = ~n5603 ;
  assign n5704 = n34054 & n166 ;
  assign n5705 = n5413 | n5704 ;
  assign n34055 = ~n5591 ;
  assign n5601 = n5413 & n34055 ;
  assign n5602 = n33850 & n5601 ;
  assign n5737 = n5602 & n166 ;
  assign n34056 = ~n5737 ;
  assign n5738 = n5705 & n34056 ;
  assign n6012 = n413 | n6010 ;
  assign n34057 = ~n6012 ;
  assign n6031 = n34057 & n6028 ;
  assign n6032 = n5738 | n6031 ;
  assign n34058 = ~n6030 ;
  assign n6033 = n34058 & n6032 ;
  assign n34059 = ~n6033 ;
  assign n6034 = n189 & n34059 ;
  assign n5596 = n5594 | n5595 ;
  assign n34060 = ~n5596 ;
  assign n5702 = n34060 & n166 ;
  assign n5703 = n5362 | n5702 ;
  assign n5623 = n5362 & n33874 ;
  assign n34061 = ~n5595 ;
  assign n5624 = n34061 & n5623 ;
  assign n5740 = n5624 & n166 ;
  assign n34062 = ~n5740 ;
  assign n5741 = n5703 & n34062 ;
  assign n6042 = n34041 & n6023 ;
  assign n6043 = n5711 | n6042 ;
  assign n34063 = ~n6025 ;
  assign n6044 = n34063 & n6043 ;
  assign n34064 = ~n6044 ;
  assign n6045 = n187 & n34064 ;
  assign n6046 = n34051 & n6043 ;
  assign n6047 = n5707 | n6046 ;
  assign n34065 = ~n6045 ;
  assign n6048 = n34065 & n6047 ;
  assign n34066 = ~n6048 ;
  assign n6049 = n413 & n34066 ;
  assign n6050 = n189 | n6049 ;
  assign n34067 = ~n6050 ;
  assign n6051 = n6032 & n34067 ;
  assign n6052 = n5741 | n6051 ;
  assign n34068 = ~n6034 ;
  assign n6053 = n34068 & n6052 ;
  assign n34069 = ~n6053 ;
  assign n6054 = n190 & n34069 ;
  assign n5622 = n5599 | n5611 ;
  assign n34070 = ~n5622 ;
  assign n5698 = n34070 & n166 ;
  assign n5699 = n5394 | n5698 ;
  assign n34071 = ~n5611 ;
  assign n5620 = n5394 & n34071 ;
  assign n5621 = n33866 & n5620 ;
  assign n5716 = n5621 & n166 ;
  assign n34072 = ~n5716 ;
  assign n5717 = n5699 & n34072 ;
  assign n6035 = n190 | n6034 ;
  assign n34073 = ~n6035 ;
  assign n6055 = n34073 & n6052 ;
  assign n6056 = n5717 | n6055 ;
  assign n34074 = ~n6054 ;
  assign n6057 = n34074 & n6056 ;
  assign n34075 = ~n6057 ;
  assign n6058 = n287 & n34075 ;
  assign n34076 = ~n5628 ;
  assign n5632 = n5337 & n34076 ;
  assign n34077 = ~n5615 ;
  assign n5633 = n34077 & n5632 ;
  assign n5694 = n5633 & n166 ;
  assign n5619 = n5614 | n5615 ;
  assign n34078 = ~n5619 ;
  assign n5695 = n34078 & n166 ;
  assign n5696 = n5337 | n5695 ;
  assign n34079 = ~n5694 ;
  assign n5697 = n34079 & n5696 ;
  assign n6065 = n34057 & n6047 ;
  assign n6066 = n5738 | n6065 ;
  assign n34080 = ~n6049 ;
  assign n6067 = n34080 & n6066 ;
  assign n34081 = ~n6067 ;
  assign n6068 = n189 & n34081 ;
  assign n6069 = n34067 & n6066 ;
  assign n6070 = n5741 | n6069 ;
  assign n34082 = ~n6068 ;
  assign n6071 = n34082 & n6070 ;
  assign n34083 = ~n6071 ;
  assign n6072 = n190 & n34083 ;
  assign n6073 = n287 | n6072 ;
  assign n34084 = ~n6073 ;
  assign n6074 = n6056 & n34084 ;
  assign n6077 = n5697 | n6074 ;
  assign n34085 = ~n6058 ;
  assign n6078 = n34085 & n6077 ;
  assign n5673 = n5657 | n5670 ;
  assign n34086 = ~n5673 ;
  assign n5679 = n34086 & n166 ;
  assign n6080 = n5675 | n5679 ;
  assign n34087 = ~n5630 ;
  assign n5667 = n34087 & n5666 ;
  assign n5668 = n33882 & n5667 ;
  assign n5692 = n5668 & n166 ;
  assign n5631 = n5618 | n5630 ;
  assign n34088 = ~n5631 ;
  assign n5722 = n34088 & n166 ;
  assign n6091 = n5666 | n5722 ;
  assign n34089 = ~n5692 ;
  assign n6092 = n34089 & n6091 ;
  assign n6095 = n6080 | n6092 ;
  assign n6096 = n6078 | n6095 ;
  assign n6097 = n31336 & n6096 ;
  assign n5674 = n192 & n5673 ;
  assign n34090 = ~n5657 ;
  assign n5681 = n34090 & n166 ;
  assign n34091 = ~n5681 ;
  assign n5682 = n5670 & n34091 ;
  assign n34092 = ~n5682 ;
  assign n5683 = n5674 & n34092 ;
  assign n5653 = n5639 | n5652 ;
  assign n34093 = ~n5653 ;
  assign n5660 = n34093 & n5656 ;
  assign n5661 = n33898 & n5660 ;
  assign n6081 = n5661 & n33899 ;
  assign n6082 = n33900 & n6081 ;
  assign n6083 = n5683 | n6082 ;
  assign n6098 = n34085 & n6092 ;
  assign n6099 = n6077 & n6098 ;
  assign n6100 = n6083 | n6099 ;
  assign n165 = n6097 | n6100 ;
  assign n10019 = x70 | x71 ;
  assign n10589 = x72 | n10019 ;
  assign n6180 = x72 & n165 ;
  assign n34094 = ~n6180 ;
  assign n6181 = n10589 & n34094 ;
  assign n34095 = ~n6181 ;
  assign n6182 = n166 & n34095 ;
  assign n5641 = n10589 & n33897 ;
  assign n5650 = n5641 & n33898 ;
  assign n6089 = n5650 & n33899 ;
  assign n6090 = n33900 & n6089 ;
  assign n6189 = n6090 & n34094 ;
  assign n34096 = ~n8390 ;
  assign n6166 = n34096 & n165 ;
  assign n34097 = ~x72 ;
  assign n6217 = n34097 & n165 ;
  assign n34098 = ~n6217 ;
  assign n6218 = x73 & n34098 ;
  assign n6219 = n6166 | n6218 ;
  assign n6220 = n6189 | n6219 ;
  assign n34099 = ~n6182 ;
  assign n6221 = n34099 & n6220 ;
  assign n34100 = ~n6221 ;
  assign n6222 = n5352 & n34100 ;
  assign n11144 = n34097 & n10019 ;
  assign n34101 = ~n165 ;
  assign n6207 = x72 & n34101 ;
  assign n6208 = n11144 | n6207 ;
  assign n34102 = ~n6208 ;
  assign n6209 = n166 & n34102 ;
  assign n6210 = n5352 | n6209 ;
  assign n34103 = ~n6210 ;
  assign n6225 = n34103 & n6220 ;
  assign n34104 = ~n6082 ;
  assign n6084 = n166 & n34104 ;
  assign n34105 = ~n5683 ;
  assign n6085 = n34105 & n6084 ;
  assign n34106 = ~n6099 ;
  assign n6229 = n6085 & n34106 ;
  assign n34107 = ~n6097 ;
  assign n6230 = n34107 & n6229 ;
  assign n6231 = n6166 | n6230 ;
  assign n6232 = x74 & n6231 ;
  assign n6233 = x74 | n6230 ;
  assign n6234 = n6166 | n6233 ;
  assign n34108 = ~n6232 ;
  assign n6235 = n34108 & n6234 ;
  assign n6236 = n6225 | n6235 ;
  assign n34109 = ~n6222 ;
  assign n6237 = n34109 & n6236 ;
  assign n34110 = ~n6237 ;
  assign n6238 = n4934 & n34110 ;
  assign n5690 = n5686 | n5689 ;
  assign n34111 = ~n5690 ;
  assign n5792 = n34111 & n5789 ;
  assign n6162 = n5792 & n165 ;
  assign n6163 = n34111 & n165 ;
  assign n6164 = n5789 | n6163 ;
  assign n34112 = ~n6162 ;
  assign n6165 = n34112 & n6164 ;
  assign n6223 = n4934 | n6222 ;
  assign n34113 = ~n6223 ;
  assign n6241 = n34113 & n6236 ;
  assign n6242 = n6165 | n6241 ;
  assign n34114 = ~n6238 ;
  assign n6243 = n34114 & n6242 ;
  assign n34115 = ~n6243 ;
  assign n6244 = n169 & n34115 ;
  assign n5797 = n5791 | n5796 ;
  assign n34116 = ~n5797 ;
  assign n6112 = n34116 & n165 ;
  assign n6113 = n5805 | n6112 ;
  assign n34117 = ~n5791 ;
  assign n5825 = n34117 & n5805 ;
  assign n5826 = n33902 & n5825 ;
  assign n6215 = n5826 & n165 ;
  assign n34118 = ~n6215 ;
  assign n6216 = n6113 & n34118 ;
  assign n6239 = n169 | n6238 ;
  assign n34119 = ~n6239 ;
  assign n6245 = n34119 & n6242 ;
  assign n6246 = n6216 | n6245 ;
  assign n34120 = ~n6244 ;
  assign n6247 = n34120 & n6246 ;
  assign n34121 = ~n6247 ;
  assign n6248 = n170 & n34121 ;
  assign n5824 = n5808 | n5811 ;
  assign n34122 = ~n5824 ;
  assign n6170 = n34122 & n165 ;
  assign n6171 = n5735 | n6170 ;
  assign n5810 = n5735 & n33907 ;
  assign n34123 = ~n5811 ;
  assign n5823 = n5810 & n34123 ;
  assign n6205 = n5823 & n165 ;
  assign n34124 = ~n6205 ;
  assign n6206 = n6171 & n34124 ;
  assign n6224 = n167 & n34100 ;
  assign n6183 = n167 | n6182 ;
  assign n34125 = ~n6183 ;
  assign n6227 = n34125 & n6220 ;
  assign n6258 = n6227 | n6235 ;
  assign n34126 = ~n6224 ;
  assign n6259 = n34126 & n6258 ;
  assign n34127 = ~n6259 ;
  assign n6260 = n168 & n34127 ;
  assign n6261 = n34113 & n6258 ;
  assign n6262 = n6165 | n6261 ;
  assign n34128 = ~n6260 ;
  assign n6263 = n34128 & n6262 ;
  assign n34129 = ~n6263 ;
  assign n6264 = n169 & n34129 ;
  assign n6265 = n170 | n6264 ;
  assign n34130 = ~n6265 ;
  assign n6266 = n6246 & n34130 ;
  assign n6267 = n6206 | n6266 ;
  assign n34131 = ~n6248 ;
  assign n6268 = n34131 & n6267 ;
  assign n34132 = ~n6268 ;
  assign n6269 = n171 & n34132 ;
  assign n5849 = n5815 | n5833 ;
  assign n34133 = ~n5849 ;
  assign n6142 = n34133 & n165 ;
  assign n6143 = n5763 | n6142 ;
  assign n34134 = ~n5815 ;
  assign n5821 = n5763 & n34134 ;
  assign n5822 = n33913 & n5821 ;
  assign n6195 = n5822 & n165 ;
  assign n34135 = ~n6195 ;
  assign n6196 = n6143 & n34135 ;
  assign n6249 = n3940 | n6248 ;
  assign n34136 = ~n6249 ;
  assign n6270 = n34136 & n6267 ;
  assign n6271 = n6196 | n6270 ;
  assign n34137 = ~n6269 ;
  assign n6272 = n34137 & n6271 ;
  assign n34138 = ~n6272 ;
  assign n6273 = n3631 & n34138 ;
  assign n5848 = n5818 | n5835 ;
  assign n34139 = ~n5848 ;
  assign n6146 = n34139 & n165 ;
  assign n6147 = n5726 | n6146 ;
  assign n5820 = n5726 & n33924 ;
  assign n34140 = ~n5835 ;
  assign n5847 = n5820 & n34140 ;
  assign n6157 = n5847 & n165 ;
  assign n34141 = ~n6157 ;
  assign n6158 = n6147 & n34141 ;
  assign n6281 = n34119 & n6262 ;
  assign n6282 = n6216 | n6281 ;
  assign n34142 = ~n6264 ;
  assign n6283 = n34142 & n6282 ;
  assign n34143 = ~n6283 ;
  assign n6284 = n170 & n34143 ;
  assign n6285 = n34130 & n6282 ;
  assign n6286 = n6206 | n6285 ;
  assign n34144 = ~n6284 ;
  assign n6287 = n34144 & n6286 ;
  assign n34145 = ~n6287 ;
  assign n6288 = n3940 & n34145 ;
  assign n6289 = n3631 | n6288 ;
  assign n34146 = ~n6289 ;
  assign n6290 = n6271 & n34146 ;
  assign n6291 = n6158 | n6290 ;
  assign n34147 = ~n6273 ;
  assign n6292 = n34147 & n6291 ;
  assign n34148 = ~n6292 ;
  assign n6293 = n173 & n34148 ;
  assign n5873 = n5839 | n5857 ;
  assign n34149 = ~n5873 ;
  assign n6137 = n34149 & n165 ;
  assign n6138 = n5745 | n6137 ;
  assign n34150 = ~n5839 ;
  assign n5845 = n5745 & n34150 ;
  assign n5846 = n33930 & n5845 ;
  assign n6148 = n5846 & n165 ;
  assign n34151 = ~n6148 ;
  assign n6149 = n6138 & n34151 ;
  assign n6275 = n173 | n6273 ;
  assign n34152 = ~n6275 ;
  assign n6294 = n34152 & n6291 ;
  assign n6298 = n6149 | n6294 ;
  assign n34153 = ~n6293 ;
  assign n6299 = n34153 & n6298 ;
  assign n34154 = ~n6299 ;
  assign n6300 = n174 & n34154 ;
  assign n5844 = n5766 & n33940 ;
  assign n34155 = ~n5859 ;
  assign n5871 = n5844 & n34155 ;
  assign n6159 = n5871 & n165 ;
  assign n5872 = n5842 | n5859 ;
  assign n34156 = ~n5872 ;
  assign n6167 = n34156 & n165 ;
  assign n6168 = n5766 | n6167 ;
  assign n34157 = ~n6159 ;
  assign n6169 = n34157 & n6168 ;
  assign n6305 = n34136 & n6286 ;
  assign n6306 = n6196 | n6305 ;
  assign n34158 = ~n6288 ;
  assign n6307 = n34158 & n6306 ;
  assign n34159 = ~n6307 ;
  assign n6308 = n172 & n34159 ;
  assign n6309 = n34146 & n6306 ;
  assign n6310 = n6158 | n6309 ;
  assign n34160 = ~n6308 ;
  assign n6311 = n34160 & n6310 ;
  assign n34161 = ~n6311 ;
  assign n6312 = n173 & n34161 ;
  assign n6313 = n174 | n6312 ;
  assign n34162 = ~n6313 ;
  assign n6314 = n6298 & n34162 ;
  assign n6315 = n6169 | n6314 ;
  assign n34163 = ~n6300 ;
  assign n6316 = n34163 & n6315 ;
  assign n34164 = ~n6316 ;
  assign n6317 = n175 & n34164 ;
  assign n34165 = ~n5863 ;
  assign n5864 = n5760 & n34165 ;
  assign n5865 = n33946 & n5864 ;
  assign n6114 = n5865 & n165 ;
  assign n5897 = n5863 | n5881 ;
  assign n34166 = ~n5897 ;
  assign n6197 = n34166 & n165 ;
  assign n6198 = n5760 | n6197 ;
  assign n34167 = ~n6114 ;
  assign n6199 = n34167 & n6198 ;
  assign n6301 = n2753 | n6300 ;
  assign n34168 = ~n6301 ;
  assign n6318 = n34168 & n6315 ;
  assign n6319 = n6199 | n6318 ;
  assign n34169 = ~n6317 ;
  assign n6320 = n34169 & n6319 ;
  assign n34170 = ~n6320 ;
  assign n6321 = n2431 & n34170 ;
  assign n5896 = n5868 | n5883 ;
  assign n34171 = ~n5896 ;
  assign n6121 = n34171 & n165 ;
  assign n6122 = n5768 | n6121 ;
  assign n5870 = n5768 & n33956 ;
  assign n34172 = ~n5883 ;
  assign n5895 = n5870 & n34172 ;
  assign n6174 = n5895 & n165 ;
  assign n34173 = ~n6174 ;
  assign n6175 = n6122 & n34173 ;
  assign n6329 = n34152 & n6310 ;
  assign n6330 = n6149 | n6329 ;
  assign n34174 = ~n6312 ;
  assign n6331 = n34174 & n6330 ;
  assign n34175 = ~n6331 ;
  assign n6332 = n174 & n34175 ;
  assign n6333 = n34162 & n6330 ;
  assign n6334 = n6169 | n6333 ;
  assign n34176 = ~n6332 ;
  assign n6335 = n34176 & n6334 ;
  assign n34177 = ~n6335 ;
  assign n6336 = n2753 & n34177 ;
  assign n6337 = n2431 | n6336 ;
  assign n34178 = ~n6337 ;
  assign n6338 = n6319 & n34178 ;
  assign n6339 = n6175 | n6338 ;
  assign n34179 = ~n6321 ;
  assign n6340 = n34179 & n6339 ;
  assign n34180 = ~n6340 ;
  assign n6341 = n177 & n34180 ;
  assign n34181 = ~n5887 ;
  assign n5893 = n5774 & n34181 ;
  assign n5894 = n33962 & n5893 ;
  assign n6156 = n5894 & n165 ;
  assign n5921 = n5887 | n5905 ;
  assign n34182 = ~n5921 ;
  assign n6184 = n34182 & n165 ;
  assign n6185 = n5774 | n6184 ;
  assign n34183 = ~n6156 ;
  assign n6186 = n34183 & n6185 ;
  assign n6322 = n177 | n6321 ;
  assign n34184 = ~n6322 ;
  assign n6342 = n34184 & n6339 ;
  assign n6343 = n6186 | n6342 ;
  assign n34185 = ~n6341 ;
  assign n6344 = n34185 & n6343 ;
  assign n34186 = ~n6344 ;
  assign n6345 = n178 & n34186 ;
  assign n5892 = n5757 & n33972 ;
  assign n34187 = ~n5907 ;
  assign n5919 = n5892 & n34187 ;
  assign n6191 = n5919 & n165 ;
  assign n5920 = n5890 | n5907 ;
  assign n34188 = ~n5920 ;
  assign n6192 = n34188 & n165 ;
  assign n6193 = n5757 | n6192 ;
  assign n34189 = ~n6191 ;
  assign n6194 = n34189 & n6193 ;
  assign n6353 = n34168 & n6334 ;
  assign n6354 = n6199 | n6353 ;
  assign n34190 = ~n6336 ;
  assign n6355 = n34190 & n6354 ;
  assign n34191 = ~n6355 ;
  assign n6356 = n176 & n34191 ;
  assign n6357 = n34178 & n6354 ;
  assign n6358 = n6175 | n6357 ;
  assign n34192 = ~n6356 ;
  assign n6359 = n34192 & n6358 ;
  assign n34193 = ~n6359 ;
  assign n6360 = n177 & n34193 ;
  assign n6361 = n178 | n6360 ;
  assign n34194 = ~n6361 ;
  assign n6362 = n6343 & n34194 ;
  assign n6363 = n6194 | n6362 ;
  assign n34195 = ~n6345 ;
  assign n6364 = n34195 & n6363 ;
  assign n34196 = ~n6364 ;
  assign n6365 = n179 & n34196 ;
  assign n34197 = ~n5911 ;
  assign n5917 = n5782 & n34197 ;
  assign n5918 = n33978 & n5917 ;
  assign n6179 = n5918 & n165 ;
  assign n5945 = n5911 | n5929 ;
  assign n34198 = ~n5945 ;
  assign n6202 = n34198 & n165 ;
  assign n6203 = n5782 | n6202 ;
  assign n34199 = ~n6179 ;
  assign n6204 = n34199 & n6203 ;
  assign n6346 = n1707 | n6345 ;
  assign n34200 = ~n6346 ;
  assign n6366 = n34200 & n6363 ;
  assign n6367 = n6204 | n6366 ;
  assign n34201 = ~n6365 ;
  assign n6368 = n34201 & n6367 ;
  assign n34202 = ~n6368 ;
  assign n6369 = n1487 & n34202 ;
  assign n5944 = n5914 | n5931 ;
  assign n34203 = ~n5944 ;
  assign n6160 = n34203 & n165 ;
  assign n6161 = n5747 | n6160 ;
  assign n5916 = n5747 & n33988 ;
  assign n34204 = ~n5931 ;
  assign n5943 = n5916 & n34204 ;
  assign n6200 = n5943 & n165 ;
  assign n34205 = ~n6200 ;
  assign n6201 = n6161 & n34205 ;
  assign n6377 = n34184 & n6358 ;
  assign n6378 = n6186 | n6377 ;
  assign n34206 = ~n6360 ;
  assign n6379 = n34206 & n6378 ;
  assign n34207 = ~n6379 ;
  assign n6380 = n178 & n34207 ;
  assign n6381 = n34194 & n6378 ;
  assign n6382 = n6194 | n6381 ;
  assign n34208 = ~n6380 ;
  assign n6383 = n34208 & n6382 ;
  assign n34209 = ~n6383 ;
  assign n6384 = n1707 & n34209 ;
  assign n6385 = n1487 | n6384 ;
  assign n34210 = ~n6385 ;
  assign n6386 = n6367 & n34210 ;
  assign n6387 = n6201 | n6386 ;
  assign n34211 = ~n6369 ;
  assign n6388 = n34211 & n6387 ;
  assign n34212 = ~n6388 ;
  assign n6389 = n181 & n34212 ;
  assign n5969 = n5935 | n5953 ;
  assign n34213 = ~n5969 ;
  assign n6102 = n34213 & n165 ;
  assign n6103 = n5779 | n6102 ;
  assign n34214 = ~n5935 ;
  assign n5941 = n5779 & n34214 ;
  assign n5942 = n33994 & n5941 ;
  assign n6187 = n5942 & n165 ;
  assign n34215 = ~n6187 ;
  assign n6188 = n6103 & n34215 ;
  assign n6370 = n181 | n6369 ;
  assign n34216 = ~n6370 ;
  assign n6390 = n34216 & n6387 ;
  assign n6391 = n6188 | n6390 ;
  assign n34217 = ~n6389 ;
  assign n6392 = n34217 & n6391 ;
  assign n34218 = ~n6392 ;
  assign n6393 = n182 & n34218 ;
  assign n5940 = n5786 & n34004 ;
  assign n34219 = ~n5955 ;
  assign n5967 = n5940 & n34219 ;
  assign n6133 = n5967 & n165 ;
  assign n5968 = n5938 | n5955 ;
  assign n34220 = ~n5968 ;
  assign n6134 = n34220 & n165 ;
  assign n6135 = n5786 | n6134 ;
  assign n34221 = ~n6133 ;
  assign n6136 = n34221 & n6135 ;
  assign n6401 = n34200 & n6382 ;
  assign n6402 = n6204 | n6401 ;
  assign n34222 = ~n6384 ;
  assign n6403 = n34222 & n6402 ;
  assign n34223 = ~n6403 ;
  assign n6404 = n180 & n34223 ;
  assign n6405 = n34210 & n6402 ;
  assign n6406 = n6201 | n6405 ;
  assign n34224 = ~n6404 ;
  assign n6407 = n34224 & n6406 ;
  assign n34225 = ~n6407 ;
  assign n6408 = n181 & n34225 ;
  assign n6409 = n182 | n6408 ;
  assign n34226 = ~n6409 ;
  assign n6410 = n6391 & n34226 ;
  assign n6411 = n6136 | n6410 ;
  assign n34227 = ~n6393 ;
  assign n6412 = n34227 & n6411 ;
  assign n34228 = ~n6412 ;
  assign n6413 = n183 & n34228 ;
  assign n5993 = n5959 | n5977 ;
  assign n34229 = ~n5993 ;
  assign n6131 = n34229 & n165 ;
  assign n6132 = n5777 | n6131 ;
  assign n34230 = ~n5959 ;
  assign n5965 = n5777 & n34230 ;
  assign n5966 = n34010 & n5965 ;
  assign n6152 = n5966 & n165 ;
  assign n34231 = ~n6152 ;
  assign n6153 = n6132 & n34231 ;
  assign n6394 = n183 | n6393 ;
  assign n34232 = ~n6394 ;
  assign n6414 = n34232 & n6411 ;
  assign n6415 = n6153 | n6414 ;
  assign n34233 = ~n6413 ;
  assign n6416 = n34233 & n6415 ;
  assign n34234 = ~n6416 ;
  assign n6417 = n838 & n34234 ;
  assign n5964 = n5721 & n34020 ;
  assign n34235 = ~n5979 ;
  assign n5991 = n5964 & n34235 ;
  assign n6130 = n5991 & n165 ;
  assign n5992 = n5962 | n5979 ;
  assign n34236 = ~n5992 ;
  assign n6176 = n34236 & n165 ;
  assign n6177 = n5721 | n6176 ;
  assign n34237 = ~n6130 ;
  assign n6178 = n34237 & n6177 ;
  assign n6425 = n34216 & n6406 ;
  assign n6426 = n6188 | n6425 ;
  assign n34238 = ~n6408 ;
  assign n6427 = n34238 & n6426 ;
  assign n34239 = ~n6427 ;
  assign n6428 = n182 & n34239 ;
  assign n6429 = n34226 & n6426 ;
  assign n6430 = n6136 | n6429 ;
  assign n34240 = ~n6428 ;
  assign n6431 = n34240 & n6430 ;
  assign n34241 = ~n6431 ;
  assign n6432 = n996 & n34241 ;
  assign n6433 = n838 | n6432 ;
  assign n34242 = ~n6433 ;
  assign n6434 = n6415 & n34242 ;
  assign n6435 = n6178 | n6434 ;
  assign n34243 = ~n6417 ;
  assign n6436 = n34243 & n6435 ;
  assign n34244 = ~n6436 ;
  assign n6437 = n185 & n34244 ;
  assign n34245 = ~n5983 ;
  assign n5989 = n5749 & n34245 ;
  assign n5990 = n34026 & n5989 ;
  assign n6127 = n5990 & n165 ;
  assign n6017 = n5983 | n6001 ;
  assign n34246 = ~n6017 ;
  assign n6139 = n34246 & n165 ;
  assign n6140 = n5749 | n6139 ;
  assign n34247 = ~n6127 ;
  assign n6141 = n34247 & n6140 ;
  assign n6418 = n185 | n6417 ;
  assign n34248 = ~n6418 ;
  assign n6438 = n34248 & n6435 ;
  assign n6439 = n6141 | n6438 ;
  assign n34249 = ~n6437 ;
  assign n6440 = n34249 & n6439 ;
  assign n34250 = ~n6440 ;
  assign n6441 = n186 & n34250 ;
  assign n6016 = n5986 | n6003 ;
  assign n34251 = ~n6016 ;
  assign n6125 = n34251 & n165 ;
  assign n6126 = n5784 | n6125 ;
  assign n5988 = n5784 & n34036 ;
  assign n34252 = ~n6003 ;
  assign n6015 = n5988 & n34252 ;
  assign n6154 = n6015 & n165 ;
  assign n34253 = ~n6154 ;
  assign n6155 = n6126 & n34253 ;
  assign n6449 = n34232 & n6430 ;
  assign n6450 = n6153 | n6449 ;
  assign n34254 = ~n6432 ;
  assign n6451 = n34254 & n6450 ;
  assign n34255 = ~n6451 ;
  assign n6452 = n184 & n34255 ;
  assign n6453 = n34242 & n6450 ;
  assign n6454 = n6178 | n6453 ;
  assign n34256 = ~n6452 ;
  assign n6455 = n34256 & n6454 ;
  assign n34257 = ~n6455 ;
  assign n6456 = n185 & n34257 ;
  assign n6457 = n186 | n6456 ;
  assign n34258 = ~n6457 ;
  assign n6458 = n6439 & n34258 ;
  assign n6459 = n6155 | n6458 ;
  assign n34259 = ~n6441 ;
  assign n6460 = n34259 & n6459 ;
  assign n34260 = ~n6460 ;
  assign n6461 = n187 & n34260 ;
  assign n6041 = n6007 | n6025 ;
  assign n34261 = ~n6041 ;
  assign n6119 = n34261 & n165 ;
  assign n6120 = n5711 | n6119 ;
  assign n34262 = ~n6007 ;
  assign n6013 = n5711 & n34262 ;
  assign n6014 = n34042 & n6013 ;
  assign n6128 = n6014 & n165 ;
  assign n34263 = ~n6128 ;
  assign n6129 = n6120 & n34263 ;
  assign n6442 = n528 | n6441 ;
  assign n34264 = ~n6442 ;
  assign n6462 = n34264 & n6459 ;
  assign n6466 = n6129 | n6462 ;
  assign n34265 = ~n6461 ;
  assign n6467 = n34265 & n6466 ;
  assign n34266 = ~n6467 ;
  assign n6468 = n413 & n34266 ;
  assign n6040 = n6010 | n6027 ;
  assign n34267 = ~n6040 ;
  assign n6117 = n34267 & n165 ;
  assign n6118 = n5707 | n6117 ;
  assign n6011 = n5707 & n34052 ;
  assign n34268 = ~n6027 ;
  assign n6039 = n6011 & n34268 ;
  assign n6172 = n6039 & n165 ;
  assign n34269 = ~n6172 ;
  assign n6173 = n6118 & n34269 ;
  assign n6473 = n34248 & n6454 ;
  assign n6474 = n6141 | n6473 ;
  assign n34270 = ~n6456 ;
  assign n6475 = n34270 & n6474 ;
  assign n34271 = ~n6475 ;
  assign n6476 = n186 & n34271 ;
  assign n6477 = n34258 & n6474 ;
  assign n6478 = n6155 | n6477 ;
  assign n34272 = ~n6476 ;
  assign n6479 = n34272 & n6478 ;
  assign n34273 = ~n6479 ;
  assign n6480 = n528 & n34273 ;
  assign n6481 = n413 | n6480 ;
  assign n34274 = ~n6481 ;
  assign n6482 = n6466 & n34274 ;
  assign n6483 = n6173 | n6482 ;
  assign n34275 = ~n6468 ;
  assign n6484 = n34275 & n6483 ;
  assign n34276 = ~n6484 ;
  assign n6485 = n189 & n34276 ;
  assign n6064 = n6031 | n6049 ;
  assign n34277 = ~n6064 ;
  assign n6115 = n34277 & n165 ;
  assign n6116 = n5738 | n6115 ;
  assign n34278 = ~n6031 ;
  assign n6037 = n5738 & n34278 ;
  assign n6038 = n34058 & n6037 ;
  assign n6144 = n6038 & n165 ;
  assign n34279 = ~n6144 ;
  assign n6145 = n6116 & n34279 ;
  assign n6469 = n189 | n6468 ;
  assign n34280 = ~n6469 ;
  assign n6486 = n34280 & n6483 ;
  assign n6487 = n6145 | n6486 ;
  assign n34281 = ~n6485 ;
  assign n6488 = n34281 & n6487 ;
  assign n34282 = ~n6488 ;
  assign n6489 = n190 & n34282 ;
  assign n6063 = n6034 | n6051 ;
  assign n34283 = ~n6063 ;
  assign n6108 = n34283 & n165 ;
  assign n6109 = n5741 | n6108 ;
  assign n6036 = n5741 & n34068 ;
  assign n34284 = ~n6051 ;
  assign n6062 = n6036 & n34284 ;
  assign n6110 = n6062 & n165 ;
  assign n34285 = ~n6110 ;
  assign n6111 = n6109 & n34285 ;
  assign n6495 = n34264 & n6478 ;
  assign n6496 = n6129 | n6495 ;
  assign n34286 = ~n6480 ;
  assign n6497 = n34286 & n6496 ;
  assign n34287 = ~n6497 ;
  assign n6498 = n188 & n34287 ;
  assign n6499 = n34274 & n6496 ;
  assign n6500 = n6173 | n6499 ;
  assign n34288 = ~n6498 ;
  assign n6501 = n34288 & n6500 ;
  assign n34289 = ~n6501 ;
  assign n6502 = n189 & n34289 ;
  assign n6503 = n190 | n6502 ;
  assign n34290 = ~n6503 ;
  assign n6504 = n6487 & n34290 ;
  assign n6505 = n6111 | n6504 ;
  assign n34291 = ~n6489 ;
  assign n6510 = n34291 & n6505 ;
  assign n34292 = ~n6510 ;
  assign n6511 = n191 & n34292 ;
  assign n34293 = ~n6055 ;
  assign n6060 = n5717 & n34293 ;
  assign n6061 = n34074 & n6060 ;
  assign n6104 = n6061 & n165 ;
  assign n6079 = n6055 | n6072 ;
  assign n34294 = ~n6079 ;
  assign n6105 = n34294 & n165 ;
  assign n6106 = n5717 | n6105 ;
  assign n34295 = ~n6104 ;
  assign n6107 = n34295 & n6106 ;
  assign n6491 = n191 | n6489 ;
  assign n34296 = ~n6491 ;
  assign n6517 = n34296 & n6505 ;
  assign n6521 = n6107 | n6517 ;
  assign n34297 = ~n6511 ;
  assign n6522 = n34297 & n6521 ;
  assign n6076 = n6058 | n6074 ;
  assign n34298 = ~n6076 ;
  assign n6123 = n34298 & n165 ;
  assign n6124 = n5697 | n6123 ;
  assign n6059 = n5697 & n34085 ;
  assign n34299 = ~n6074 ;
  assign n6075 = n6059 & n34299 ;
  assign n6150 = n6075 & n165 ;
  assign n34300 = ~n6150 ;
  assign n6151 = n6124 & n34300 ;
  assign n6093 = n6078 | n6092 ;
  assign n34301 = ~n6093 ;
  assign n6214 = n34301 & n165 ;
  assign n6528 = n6099 | n6214 ;
  assign n6529 = n6151 | n6528 ;
  assign n6530 = n6522 | n6529 ;
  assign n6531 = n31336 & n6530 ;
  assign n6513 = n6151 & n34297 ;
  assign n6523 = n6513 & n6521 ;
  assign n6094 = n192 & n6093 ;
  assign n34302 = ~n6092 ;
  assign n6211 = n34302 & n165 ;
  assign n34303 = ~n6211 ;
  assign n6212 = n6078 & n34303 ;
  assign n34304 = ~n6212 ;
  assign n6213 = n6094 & n34304 ;
  assign n6086 = n5692 | n6082 ;
  assign n34305 = ~n6086 ;
  assign n6536 = n34305 & n6091 ;
  assign n6537 = n34105 & n6536 ;
  assign n6538 = n34106 & n6537 ;
  assign n6539 = n34107 & n6538 ;
  assign n6540 = n6213 | n6539 ;
  assign n6541 = n6523 | n6540 ;
  assign n164 = n6531 | n6541 ;
  assign n6490 = n287 | n6489 ;
  assign n34306 = ~n6490 ;
  assign n6506 = n34306 & n6505 ;
  assign n6507 = n6107 | n6506 ;
  assign n6514 = n6507 & n6513 ;
  assign n6512 = n6507 & n34297 ;
  assign n6515 = n6151 | n6512 ;
  assign n6532 = n6512 | n6529 ;
  assign n6533 = n31336 & n6532 ;
  assign n6599 = n6514 | n6540 ;
  assign n6600 = n6533 | n6599 ;
  assign n34307 = ~n6515 ;
  assign n6612 = n34307 & n6600 ;
  assign n6613 = n6514 | n6612 ;
  assign n6520 = n6511 | n6517 ;
  assign n34308 = ~n6520 ;
  assign n6543 = n34308 & n164 ;
  assign n6544 = n6107 | n6543 ;
  assign n34309 = ~n6517 ;
  assign n6518 = n6107 & n34309 ;
  assign n6519 = n34297 & n6518 ;
  assign n6621 = n6519 & n6600 ;
  assign n34310 = ~n6621 ;
  assign n6622 = n6544 & n34310 ;
  assign n6623 = n6613 | n6622 ;
  assign n34311 = ~n10019 ;
  assign n6609 = n34311 & n6600 ;
  assign n34312 = ~x70 ;
  assign n6614 = n34312 & n6600 ;
  assign n34313 = ~n6614 ;
  assign n6615 = x71 & n34313 ;
  assign n6616 = n6609 | n6615 ;
  assign n11618 = x68 | x69 ;
  assign n12275 = x70 | n11618 ;
  assign n6087 = n12275 & n34104 ;
  assign n6088 = n34105 & n6087 ;
  assign n6534 = n6088 & n34106 ;
  assign n6535 = n34107 & n6534 ;
  assign n6617 = x70 & n6600 ;
  assign n34314 = ~n6617 ;
  assign n6618 = n6535 & n34314 ;
  assign n6619 = n6616 | n6618 ;
  assign n12914 = n34312 & n11618 ;
  assign n34315 = ~n6600 ;
  assign n6630 = x70 & n34315 ;
  assign n6631 = n12914 | n6630 ;
  assign n34316 = ~n6631 ;
  assign n6632 = n165 & n34316 ;
  assign n34317 = ~n6632 ;
  assign n6633 = n6619 & n34317 ;
  assign n34318 = ~n6633 ;
  assign n6634 = n166 & n34318 ;
  assign n6565 = x70 & n164 ;
  assign n34319 = ~n6565 ;
  assign n6566 = n12275 & n34319 ;
  assign n34320 = ~n6566 ;
  assign n6567 = n165 & n34320 ;
  assign n6568 = n166 | n6567 ;
  assign n34321 = ~n6568 ;
  assign n6620 = n34321 & n6619 ;
  assign n34322 = ~n6539 ;
  assign n6691 = n165 & n34322 ;
  assign n34323 = ~n6213 ;
  assign n6692 = n34323 & n6691 ;
  assign n34324 = ~n6514 ;
  assign n6693 = n34324 & n6692 ;
  assign n34325 = ~n6531 ;
  assign n6694 = n34325 & n6693 ;
  assign n6695 = n6609 | n6694 ;
  assign n6696 = x72 & n6695 ;
  assign n6697 = x72 | n6694 ;
  assign n6698 = n6609 | n6697 ;
  assign n34326 = ~n6696 ;
  assign n6699 = n34326 & n6698 ;
  assign n6700 = n6620 | n6699 ;
  assign n34327 = ~n6634 ;
  assign n6701 = n34327 & n6700 ;
  assign n34328 = ~n6701 ;
  assign n6702 = n167 & n34328 ;
  assign n6190 = n6182 | n6189 ;
  assign n34329 = ~n6190 ;
  assign n6555 = n34329 & n164 ;
  assign n6556 = n6219 | n6555 ;
  assign n6228 = n34329 & n6219 ;
  assign n6561 = n6228 & n164 ;
  assign n34330 = ~n6561 ;
  assign n6562 = n6556 & n34330 ;
  assign n6635 = n167 | n6634 ;
  assign n6638 = n166 | n6632 ;
  assign n34331 = ~n6638 ;
  assign n6639 = n6619 & n34331 ;
  assign n6708 = n6639 | n6699 ;
  assign n34332 = ~n6635 ;
  assign n6709 = n34332 & n6708 ;
  assign n6712 = n6562 | n6709 ;
  assign n34333 = ~n6702 ;
  assign n6713 = n34333 & n6712 ;
  assign n34334 = ~n6713 ;
  assign n6714 = n168 & n34334 ;
  assign n6226 = n6224 | n6225 ;
  assign n34335 = ~n6226 ;
  assign n6573 = n34335 & n164 ;
  assign n6574 = n6235 | n6573 ;
  assign n34336 = ~n6225 ;
  assign n6256 = n34336 & n6235 ;
  assign n6257 = n34126 & n6256 ;
  assign n6607 = n6257 & n6600 ;
  assign n34337 = ~n6607 ;
  assign n6608 = n6574 & n34337 ;
  assign n6704 = n5352 & n34328 ;
  assign n6705 = n4934 | n6704 ;
  assign n34338 = ~n6705 ;
  assign n6716 = n34338 & n6712 ;
  assign n6717 = n6608 | n6716 ;
  assign n34339 = ~n6714 ;
  assign n6718 = n34339 & n6717 ;
  assign n34340 = ~n6718 ;
  assign n6719 = n169 & n34340 ;
  assign n6255 = n6238 | n6241 ;
  assign n34341 = ~n6255 ;
  assign n6563 = n34341 & n164 ;
  assign n6564 = n6165 | n6563 ;
  assign n6240 = n6165 & n34114 ;
  assign n34342 = ~n6241 ;
  assign n6254 = n6240 & n34342 ;
  assign n6610 = n6254 & n6600 ;
  assign n34343 = ~n6610 ;
  assign n6611 = n6564 & n34343 ;
  assign n6715 = n169 | n6714 ;
  assign n34344 = ~n6715 ;
  assign n6722 = n34344 & n6717 ;
  assign n6723 = n6611 | n6722 ;
  assign n34345 = ~n6719 ;
  assign n6724 = n34345 & n6723 ;
  assign n34346 = ~n6724 ;
  assign n6725 = n170 & n34346 ;
  assign n6253 = n6244 | n6245 ;
  assign n34347 = ~n6253 ;
  assign n6545 = n34347 & n164 ;
  assign n6546 = n6216 | n6545 ;
  assign n34348 = ~n6245 ;
  assign n6251 = n6216 & n34348 ;
  assign n6252 = n34120 & n6251 ;
  assign n6626 = n6252 & n6600 ;
  assign n34349 = ~n6626 ;
  assign n6627 = n6546 & n34349 ;
  assign n6720 = n170 | n6719 ;
  assign n34350 = ~n6720 ;
  assign n6726 = n34350 & n6723 ;
  assign n6727 = n6627 | n6726 ;
  assign n34351 = ~n6725 ;
  assign n6728 = n34351 & n6727 ;
  assign n34352 = ~n6728 ;
  assign n6729 = n3940 & n34352 ;
  assign n6280 = n6248 | n6266 ;
  assign n34353 = ~n6280 ;
  assign n6559 = n34353 & n164 ;
  assign n6560 = n6206 | n6559 ;
  assign n6250 = n6206 & n34131 ;
  assign n34354 = ~n6266 ;
  assign n6279 = n6250 & n34354 ;
  assign n6605 = n6279 & n6600 ;
  assign n34355 = ~n6605 ;
  assign n6606 = n6560 & n34355 ;
  assign n6732 = n3940 | n6725 ;
  assign n34356 = ~n6732 ;
  assign n6733 = n6727 & n34356 ;
  assign n6734 = n6606 | n6733 ;
  assign n34357 = ~n6729 ;
  assign n6735 = n34357 & n6734 ;
  assign n34358 = ~n6735 ;
  assign n6736 = n172 & n34358 ;
  assign n6278 = n6269 | n6270 ;
  assign n34359 = ~n6278 ;
  assign n6557 = n34359 & n164 ;
  assign n6558 = n6196 | n6557 ;
  assign n34360 = ~n6270 ;
  assign n6276 = n6196 & n34360 ;
  assign n6277 = n34137 & n6276 ;
  assign n6628 = n6277 & n6600 ;
  assign n34361 = ~n6628 ;
  assign n6629 = n6558 & n34361 ;
  assign n6730 = n3631 | n6729 ;
  assign n34362 = ~n6730 ;
  assign n6737 = n34362 & n6734 ;
  assign n6738 = n6629 | n6737 ;
  assign n34363 = ~n6736 ;
  assign n6739 = n34363 & n6738 ;
  assign n34364 = ~n6739 ;
  assign n6740 = n173 & n34364 ;
  assign n6304 = n6273 | n6290 ;
  assign n34365 = ~n6304 ;
  assign n6547 = n34365 & n164 ;
  assign n6548 = n6158 | n6547 ;
  assign n6274 = n6158 & n34147 ;
  assign n34366 = ~n6290 ;
  assign n6303 = n6274 & n34366 ;
  assign n6603 = n6303 & n6600 ;
  assign n34367 = ~n6603 ;
  assign n6604 = n6548 & n34367 ;
  assign n6743 = n171 & n34352 ;
  assign n34368 = ~n6743 ;
  assign n6744 = n6734 & n34368 ;
  assign n34369 = ~n6744 ;
  assign n6745 = n3631 & n34369 ;
  assign n6746 = n173 | n6745 ;
  assign n34370 = ~n6746 ;
  assign n6747 = n6738 & n34370 ;
  assign n6748 = n6604 | n6747 ;
  assign n34371 = ~n6740 ;
  assign n6749 = n34371 & n6748 ;
  assign n34372 = ~n6749 ;
  assign n6750 = n174 & n34372 ;
  assign n6297 = n6293 | n6294 ;
  assign n34373 = ~n6297 ;
  assign n6571 = n34373 & n164 ;
  assign n6572 = n6149 | n6571 ;
  assign n34374 = ~n6294 ;
  assign n6295 = n6149 & n34374 ;
  assign n6296 = n34153 & n6295 ;
  assign n6601 = n6296 & n6600 ;
  assign n34375 = ~n6601 ;
  assign n6602 = n6572 & n34375 ;
  assign n6741 = n174 | n6740 ;
  assign n34376 = ~n6741 ;
  assign n6751 = n34376 & n6748 ;
  assign n6752 = n6602 | n6751 ;
  assign n34377 = ~n6750 ;
  assign n6753 = n34377 & n6752 ;
  assign n34378 = ~n6753 ;
  assign n6754 = n2753 & n34378 ;
  assign n6328 = n6300 | n6314 ;
  assign n34379 = ~n6328 ;
  assign n6551 = n34379 & n164 ;
  assign n6552 = n6169 | n6551 ;
  assign n6302 = n6169 & n34163 ;
  assign n34380 = ~n6314 ;
  assign n6327 = n6302 & n34380 ;
  assign n6646 = n6327 & n6600 ;
  assign n34381 = ~n6646 ;
  assign n6647 = n6552 & n34381 ;
  assign n34382 = ~n6745 ;
  assign n6757 = n6738 & n34382 ;
  assign n34383 = ~n6757 ;
  assign n6758 = n173 & n34383 ;
  assign n34384 = ~n6758 ;
  assign n6759 = n6748 & n34384 ;
  assign n34385 = ~n6759 ;
  assign n6760 = n174 & n34385 ;
  assign n6761 = n2753 | n6760 ;
  assign n34386 = ~n6761 ;
  assign n6762 = n6752 & n34386 ;
  assign n6763 = n6647 | n6762 ;
  assign n34387 = ~n6754 ;
  assign n6764 = n34387 & n6763 ;
  assign n34388 = ~n6764 ;
  assign n6765 = n176 & n34388 ;
  assign n6326 = n6317 | n6318 ;
  assign n34389 = ~n6326 ;
  assign n6648 = n34389 & n6600 ;
  assign n6649 = n6199 | n6648 ;
  assign n34390 = ~n6318 ;
  assign n6324 = n6199 & n34390 ;
  assign n6325 = n34169 & n6324 ;
  assign n6650 = n6325 & n6600 ;
  assign n34391 = ~n6650 ;
  assign n6651 = n6649 & n34391 ;
  assign n6755 = n2431 | n6754 ;
  assign n34392 = ~n6755 ;
  assign n6766 = n34392 & n6763 ;
  assign n6767 = n6651 | n6766 ;
  assign n34393 = ~n6765 ;
  assign n6768 = n34393 & n6767 ;
  assign n34394 = ~n6768 ;
  assign n6769 = n177 & n34394 ;
  assign n6352 = n6321 | n6338 ;
  assign n34395 = ~n6352 ;
  assign n6553 = n34395 & n164 ;
  assign n6554 = n6175 | n6553 ;
  assign n6323 = n6175 & n34179 ;
  assign n34396 = ~n6338 ;
  assign n6351 = n6323 & n34396 ;
  assign n6652 = n6351 & n6600 ;
  assign n34397 = ~n6652 ;
  assign n6653 = n6554 & n34397 ;
  assign n34398 = ~n6760 ;
  assign n6772 = n6752 & n34398 ;
  assign n34399 = ~n6772 ;
  assign n6773 = n175 & n34399 ;
  assign n34400 = ~n6773 ;
  assign n6774 = n6763 & n34400 ;
  assign n34401 = ~n6774 ;
  assign n6775 = n2431 & n34401 ;
  assign n6776 = n177 | n6775 ;
  assign n34402 = ~n6776 ;
  assign n6777 = n6767 & n34402 ;
  assign n6778 = n6653 | n6777 ;
  assign n34403 = ~n6769 ;
  assign n6779 = n34403 & n6778 ;
  assign n34404 = ~n6779 ;
  assign n6780 = n178 & n34404 ;
  assign n6350 = n6341 | n6342 ;
  assign n34405 = ~n6350 ;
  assign n6549 = n34405 & n164 ;
  assign n6550 = n6186 | n6549 ;
  assign n34406 = ~n6342 ;
  assign n6348 = n6186 & n34406 ;
  assign n6349 = n34185 & n6348 ;
  assign n6654 = n6349 & n6600 ;
  assign n34407 = ~n6654 ;
  assign n6655 = n6550 & n34407 ;
  assign n6770 = n178 | n6769 ;
  assign n34408 = ~n6770 ;
  assign n6781 = n34408 & n6778 ;
  assign n6782 = n6655 | n6781 ;
  assign n34409 = ~n6780 ;
  assign n6783 = n34409 & n6782 ;
  assign n34410 = ~n6783 ;
  assign n6784 = n1707 & n34410 ;
  assign n6376 = n6345 | n6362 ;
  assign n34411 = ~n6376 ;
  assign n6597 = n34411 & n164 ;
  assign n6598 = n6194 | n6597 ;
  assign n6347 = n6194 & n34195 ;
  assign n34412 = ~n6362 ;
  assign n6375 = n6347 & n34412 ;
  assign n6656 = n6375 & n6600 ;
  assign n34413 = ~n6656 ;
  assign n6657 = n6598 & n34413 ;
  assign n34414 = ~n6775 ;
  assign n6787 = n6767 & n34414 ;
  assign n34415 = ~n6787 ;
  assign n6788 = n177 & n34415 ;
  assign n34416 = ~n6788 ;
  assign n6789 = n6778 & n34416 ;
  assign n34417 = ~n6789 ;
  assign n6790 = n178 & n34417 ;
  assign n6791 = n1707 | n6790 ;
  assign n34418 = ~n6791 ;
  assign n6792 = n6782 & n34418 ;
  assign n6793 = n6657 | n6792 ;
  assign n34419 = ~n6784 ;
  assign n6794 = n34419 & n6793 ;
  assign n34420 = ~n6794 ;
  assign n6795 = n180 & n34420 ;
  assign n6374 = n6365 | n6366 ;
  assign n34421 = ~n6374 ;
  assign n6579 = n34421 & n164 ;
  assign n6580 = n6204 | n6579 ;
  assign n34422 = ~n6366 ;
  assign n6372 = n6204 & n34422 ;
  assign n6373 = n34201 & n6372 ;
  assign n6658 = n6373 & n6600 ;
  assign n34423 = ~n6658 ;
  assign n6659 = n6580 & n34423 ;
  assign n6785 = n1487 | n6784 ;
  assign n34424 = ~n6785 ;
  assign n6796 = n34424 & n6793 ;
  assign n6797 = n6659 | n6796 ;
  assign n34425 = ~n6795 ;
  assign n6798 = n34425 & n6797 ;
  assign n34426 = ~n6798 ;
  assign n6799 = n181 & n34426 ;
  assign n6400 = n6369 | n6386 ;
  assign n34427 = ~n6400 ;
  assign n6581 = n34427 & n164 ;
  assign n6582 = n6201 | n6581 ;
  assign n6371 = n6201 & n34211 ;
  assign n34428 = ~n6386 ;
  assign n6399 = n6371 & n34428 ;
  assign n6624 = n6399 & n6600 ;
  assign n34429 = ~n6624 ;
  assign n6625 = n6582 & n34429 ;
  assign n34430 = ~n6790 ;
  assign n6802 = n6782 & n34430 ;
  assign n34431 = ~n6802 ;
  assign n6803 = n179 & n34431 ;
  assign n34432 = ~n6803 ;
  assign n6804 = n6793 & n34432 ;
  assign n34433 = ~n6804 ;
  assign n6805 = n1487 & n34433 ;
  assign n6806 = n181 | n6805 ;
  assign n34434 = ~n6806 ;
  assign n6807 = n6797 & n34434 ;
  assign n6808 = n6625 | n6807 ;
  assign n34435 = ~n6799 ;
  assign n6809 = n34435 & n6808 ;
  assign n34436 = ~n6809 ;
  assign n6810 = n182 & n34436 ;
  assign n6398 = n6389 | n6390 ;
  assign n34437 = ~n6398 ;
  assign n6575 = n34437 & n164 ;
  assign n6576 = n6188 | n6575 ;
  assign n34438 = ~n6390 ;
  assign n6396 = n6188 & n34438 ;
  assign n6397 = n34217 & n6396 ;
  assign n6660 = n6397 & n6600 ;
  assign n34439 = ~n6660 ;
  assign n6661 = n6576 & n34439 ;
  assign n6800 = n182 | n6799 ;
  assign n34440 = ~n6800 ;
  assign n6811 = n34440 & n6808 ;
  assign n6812 = n6661 | n6811 ;
  assign n34441 = ~n6810 ;
  assign n6813 = n34441 & n6812 ;
  assign n34442 = ~n6813 ;
  assign n6814 = n996 & n34442 ;
  assign n6424 = n6393 | n6410 ;
  assign n34443 = ~n6424 ;
  assign n6583 = n34443 & n164 ;
  assign n6584 = n6136 | n6583 ;
  assign n6395 = n6136 & n34227 ;
  assign n34444 = ~n6410 ;
  assign n6423 = n6395 & n34444 ;
  assign n6662 = n6423 & n6600 ;
  assign n34445 = ~n6662 ;
  assign n6663 = n6584 & n34445 ;
  assign n34446 = ~n6805 ;
  assign n6817 = n6797 & n34446 ;
  assign n34447 = ~n6817 ;
  assign n6818 = n181 & n34447 ;
  assign n34448 = ~n6818 ;
  assign n6819 = n6808 & n34448 ;
  assign n34449 = ~n6819 ;
  assign n6820 = n182 & n34449 ;
  assign n6821 = n183 | n6820 ;
  assign n34450 = ~n6821 ;
  assign n6822 = n6812 & n34450 ;
  assign n6823 = n6663 | n6822 ;
  assign n34451 = ~n6814 ;
  assign n6824 = n34451 & n6823 ;
  assign n34452 = ~n6824 ;
  assign n6825 = n184 & n34452 ;
  assign n6422 = n6413 | n6414 ;
  assign n34453 = ~n6422 ;
  assign n6577 = n34453 & n164 ;
  assign n6578 = n6153 | n6577 ;
  assign n34454 = ~n6414 ;
  assign n6420 = n6153 & n34454 ;
  assign n6421 = n34233 & n6420 ;
  assign n6664 = n6421 & n6600 ;
  assign n34455 = ~n6664 ;
  assign n6665 = n6578 & n34455 ;
  assign n6815 = n838 | n6814 ;
  assign n34456 = ~n6815 ;
  assign n6826 = n34456 & n6823 ;
  assign n6827 = n6665 | n6826 ;
  assign n34457 = ~n6825 ;
  assign n6828 = n34457 & n6827 ;
  assign n34458 = ~n6828 ;
  assign n6829 = n185 & n34458 ;
  assign n6448 = n6417 | n6434 ;
  assign n34459 = ~n6448 ;
  assign n6591 = n34459 & n164 ;
  assign n6592 = n6178 | n6591 ;
  assign n6419 = n6178 & n34243 ;
  assign n34460 = ~n6434 ;
  assign n6447 = n6419 & n34460 ;
  assign n6666 = n6447 & n6600 ;
  assign n34461 = ~n6666 ;
  assign n6667 = n6592 & n34461 ;
  assign n34462 = ~n6820 ;
  assign n6832 = n6812 & n34462 ;
  assign n34463 = ~n6832 ;
  assign n6833 = n183 & n34463 ;
  assign n34464 = ~n6833 ;
  assign n6834 = n6823 & n34464 ;
  assign n34465 = ~n6834 ;
  assign n6835 = n838 & n34465 ;
  assign n6836 = n185 | n6835 ;
  assign n34466 = ~n6836 ;
  assign n6837 = n6827 & n34466 ;
  assign n6838 = n6667 | n6837 ;
  assign n34467 = ~n6829 ;
  assign n6839 = n34467 & n6838 ;
  assign n34468 = ~n6839 ;
  assign n6840 = n186 & n34468 ;
  assign n6446 = n6437 | n6438 ;
  assign n34469 = ~n6446 ;
  assign n6585 = n34469 & n164 ;
  assign n6586 = n6141 | n6585 ;
  assign n34470 = ~n6438 ;
  assign n6444 = n6141 & n34470 ;
  assign n6445 = n34249 & n6444 ;
  assign n6668 = n6445 & n6600 ;
  assign n34471 = ~n6668 ;
  assign n6669 = n6586 & n34471 ;
  assign n6830 = n186 | n6829 ;
  assign n34472 = ~n6830 ;
  assign n6841 = n34472 & n6838 ;
  assign n6842 = n6669 | n6841 ;
  assign n34473 = ~n6840 ;
  assign n6843 = n34473 & n6842 ;
  assign n34474 = ~n6843 ;
  assign n6844 = n528 & n34474 ;
  assign n6471 = n6441 | n6458 ;
  assign n34475 = ~n6471 ;
  assign n6587 = n34475 & n164 ;
  assign n6588 = n6155 | n6587 ;
  assign n6443 = n6155 & n34259 ;
  assign n34476 = ~n6458 ;
  assign n6472 = n6443 & n34476 ;
  assign n6644 = n6472 & n6600 ;
  assign n34477 = ~n6644 ;
  assign n6645 = n6588 & n34477 ;
  assign n34478 = ~n6835 ;
  assign n6847 = n6827 & n34478 ;
  assign n34479 = ~n6847 ;
  assign n6848 = n185 & n34479 ;
  assign n34480 = ~n6848 ;
  assign n6849 = n6838 & n34480 ;
  assign n34481 = ~n6849 ;
  assign n6850 = n186 & n34481 ;
  assign n6851 = n528 | n6850 ;
  assign n34482 = ~n6851 ;
  assign n6852 = n6842 & n34482 ;
  assign n6853 = n6645 | n6852 ;
  assign n34483 = ~n6844 ;
  assign n6854 = n34483 & n6853 ;
  assign n34484 = ~n6854 ;
  assign n6855 = n188 & n34484 ;
  assign n6465 = n6461 | n6462 ;
  assign n34485 = ~n6465 ;
  assign n6589 = n34485 & n164 ;
  assign n6590 = n6129 | n6589 ;
  assign n34486 = ~n6462 ;
  assign n6463 = n6129 & n34486 ;
  assign n6464 = n34265 & n6463 ;
  assign n6670 = n6464 & n6600 ;
  assign n34487 = ~n6670 ;
  assign n6671 = n6590 & n34487 ;
  assign n6845 = n413 | n6844 ;
  assign n34488 = ~n6845 ;
  assign n6856 = n34488 & n6853 ;
  assign n6857 = n6671 | n6856 ;
  assign n34489 = ~n6855 ;
  assign n6858 = n34489 & n6857 ;
  assign n34490 = ~n6858 ;
  assign n6859 = n189 & n34490 ;
  assign n6494 = n6468 | n6482 ;
  assign n34491 = ~n6494 ;
  assign n6593 = n34491 & n164 ;
  assign n6594 = n6173 | n6593 ;
  assign n6470 = n6173 & n34275 ;
  assign n34492 = ~n6482 ;
  assign n6493 = n6470 & n34492 ;
  assign n6674 = n6493 & n6600 ;
  assign n34493 = ~n6674 ;
  assign n6675 = n6594 & n34493 ;
  assign n34494 = ~n6850 ;
  assign n6862 = n6842 & n34494 ;
  assign n34495 = ~n6862 ;
  assign n6863 = n187 & n34495 ;
  assign n34496 = ~n6863 ;
  assign n6864 = n6853 & n34496 ;
  assign n34497 = ~n6864 ;
  assign n6865 = n413 & n34497 ;
  assign n6866 = n189 | n6865 ;
  assign n34498 = ~n6866 ;
  assign n6867 = n6857 & n34498 ;
  assign n6868 = n6675 | n6867 ;
  assign n34499 = ~n6859 ;
  assign n6869 = n34499 & n6868 ;
  assign n34500 = ~n6869 ;
  assign n6870 = n190 & n34500 ;
  assign n6524 = n34280 & n6500 ;
  assign n6527 = n6485 | n6524 ;
  assign n34501 = ~n6527 ;
  assign n6569 = n34501 & n164 ;
  assign n6570 = n6145 | n6569 ;
  assign n34502 = ~n6524 ;
  assign n6525 = n6145 & n34502 ;
  assign n6526 = n34281 & n6525 ;
  assign n6672 = n6526 & n6600 ;
  assign n34503 = ~n6672 ;
  assign n6673 = n6570 & n34503 ;
  assign n6860 = n190 | n6859 ;
  assign n34504 = ~n6860 ;
  assign n6871 = n34504 & n6868 ;
  assign n6872 = n6673 | n6871 ;
  assign n34505 = ~n6870 ;
  assign n6873 = n34505 & n6872 ;
  assign n34506 = ~n6873 ;
  assign n6874 = n287 & n34506 ;
  assign n6509 = n6489 | n6504 ;
  assign n34507 = ~n6509 ;
  assign n6595 = n34507 & n164 ;
  assign n6596 = n6111 | n6595 ;
  assign n6492 = n6111 & n34291 ;
  assign n34508 = ~n6504 ;
  assign n6508 = n6492 & n34508 ;
  assign n6676 = n6508 & n6600 ;
  assign n34509 = ~n6676 ;
  assign n6677 = n6596 & n34509 ;
  assign n34510 = ~n6865 ;
  assign n6877 = n6857 & n34510 ;
  assign n34511 = ~n6877 ;
  assign n6878 = n189 & n34511 ;
  assign n34512 = ~n6878 ;
  assign n6879 = n6868 & n34512 ;
  assign n34513 = ~n6879 ;
  assign n6880 = n190 & n34513 ;
  assign n6881 = n287 | n6880 ;
  assign n34514 = ~n6881 ;
  assign n6882 = n6872 & n34514 ;
  assign n6883 = n6677 | n6882 ;
  assign n34515 = ~n6874 ;
  assign n6884 = n34515 & n6883 ;
  assign n6885 = n6623 | n6884 ;
  assign n6886 = n31336 & n6885 ;
  assign n6516 = n192 & n6515 ;
  assign n34516 = ~n6151 ;
  assign n6641 = n34516 & n6600 ;
  assign n34517 = ~n6641 ;
  assign n6642 = n6512 & n34517 ;
  assign n34518 = ~n6642 ;
  assign n6643 = n6516 & n34518 ;
  assign n6678 = n6150 | n6539 ;
  assign n34519 = ~n6678 ;
  assign n6679 = n6124 & n34519 ;
  assign n6680 = n34323 & n6679 ;
  assign n6681 = n34324 & n6680 ;
  assign n6682 = n34325 & n6681 ;
  assign n6683 = n6643 | n6682 ;
  assign n6875 = n6622 & n34515 ;
  assign n6887 = n6875 & n6883 ;
  assign n6888 = n6683 | n6887 ;
  assign n6889 = n6886 | n6888 ;
  assign n6915 = n6622 | n6884 ;
  assign n34520 = ~n6915 ;
  assign n6916 = n6889 & n34520 ;
  assign n6917 = n6887 | n6916 ;
  assign n6876 = n6677 & n34515 ;
  assign n6919 = n191 | n6880 ;
  assign n34521 = ~n6919 ;
  assign n6920 = n6872 & n34521 ;
  assign n34522 = ~n6920 ;
  assign n6921 = n6876 & n34522 ;
  assign n6922 = n6889 & n6921 ;
  assign n6924 = n6874 | n6920 ;
  assign n34523 = ~n6880 ;
  assign n6925 = n6872 & n34523 ;
  assign n34524 = ~n6925 ;
  assign n6926 = n191 & n34524 ;
  assign n6927 = n6677 | n6920 ;
  assign n34525 = ~n6926 ;
  assign n6928 = n34525 & n6927 ;
  assign n6929 = n6623 | n6928 ;
  assign n6930 = n31336 & n6929 ;
  assign n6931 = n6875 & n6927 ;
  assign n6932 = n6683 | n6931 ;
  assign n163 = n6930 | n6932 ;
  assign n34526 = ~n6924 ;
  assign n6941 = n34526 & n163 ;
  assign n6942 = n6677 | n6941 ;
  assign n34527 = ~n6922 ;
  assign n6943 = n34527 & n6942 ;
  assign n6944 = n6917 | n6943 ;
  assign n34528 = ~n6856 ;
  assign n6970 = n6671 & n34528 ;
  assign n6971 = n34510 & n6970 ;
  assign n6972 = n6889 & n6971 ;
  assign n6973 = n6856 | n6865 ;
  assign n34529 = ~n6973 ;
  assign n6974 = n163 & n34529 ;
  assign n6975 = n6671 | n6974 ;
  assign n34530 = ~n6972 ;
  assign n6976 = n34530 & n6975 ;
  assign n13540 = x66 | x67 ;
  assign n34531 = ~x68 ;
  assign n14918 = n34531 & n13540 ;
  assign n34532 = ~n6889 ;
  assign n6898 = x68 & n34532 ;
  assign n6899 = n14918 | n6898 ;
  assign n34533 = ~n6899 ;
  assign n6900 = n6600 & n34533 ;
  assign n6890 = n34531 & n6889 ;
  assign n34534 = ~n6890 ;
  assign n6891 = x69 & n34534 ;
  assign n34535 = ~n11618 ;
  assign n6894 = n34535 & n6889 ;
  assign n6895 = n6891 | n6894 ;
  assign n6892 = x68 & n6889 ;
  assign n14207 = x68 | n13540 ;
  assign n7109 = n14207 & n34322 ;
  assign n7110 = n34323 & n7109 ;
  assign n7111 = n34324 & n7110 ;
  assign n7112 = n34325 & n7111 ;
  assign n34536 = ~n6892 ;
  assign n7113 = n34536 & n7112 ;
  assign n7114 = n6895 | n7113 ;
  assign n34537 = ~n6900 ;
  assign n7115 = n34537 & n7114 ;
  assign n34538 = ~n7115 ;
  assign n7116 = n165 & n34538 ;
  assign n34539 = ~n6682 ;
  assign n6684 = n6600 & n34539 ;
  assign n34540 = ~n6643 ;
  assign n6685 = n34540 & n6684 ;
  assign n34541 = ~n6887 ;
  assign n6902 = n6685 & n34541 ;
  assign n34542 = ~n6886 ;
  assign n6903 = n34542 & n6902 ;
  assign n6904 = n6894 | n6903 ;
  assign n6905 = x70 & n6904 ;
  assign n6906 = x70 | n6903 ;
  assign n6907 = n6894 | n6906 ;
  assign n34543 = ~n6905 ;
  assign n6908 = n34543 & n6907 ;
  assign n6934 = x68 & n163 ;
  assign n34544 = ~n6934 ;
  assign n6935 = n14207 & n34544 ;
  assign n34545 = ~n6935 ;
  assign n6936 = n164 & n34545 ;
  assign n6937 = n165 | n6936 ;
  assign n34546 = ~n6937 ;
  assign n7118 = n34546 & n7114 ;
  assign n7119 = n6908 | n7118 ;
  assign n34547 = ~n7116 ;
  assign n7120 = n34547 & n7119 ;
  assign n34548 = ~n7120 ;
  assign n7121 = n166 & n34548 ;
  assign n6636 = n6618 | n6632 ;
  assign n34549 = ~n6636 ;
  assign n6637 = n6616 & n34549 ;
  assign n6893 = n6637 & n6889 ;
  assign n6938 = n34549 & n163 ;
  assign n6939 = n6616 | n6938 ;
  assign n34550 = ~n6893 ;
  assign n6940 = n34550 & n6939 ;
  assign n7117 = n166 | n7116 ;
  assign n6901 = n165 | n6900 ;
  assign n34551 = ~n6901 ;
  assign n7126 = n34551 & n7114 ;
  assign n7127 = n6908 | n7126 ;
  assign n34552 = ~n7117 ;
  assign n7128 = n34552 & n7127 ;
  assign n7129 = n6940 | n7128 ;
  assign n34553 = ~n7121 ;
  assign n7130 = n34553 & n7129 ;
  assign n34554 = ~n7130 ;
  assign n7131 = n167 & n34554 ;
  assign n34555 = ~n6639 ;
  assign n6706 = n34555 & n6699 ;
  assign n6707 = n34327 & n6706 ;
  assign n6897 = n6707 & n6889 ;
  assign n6640 = n6634 | n6639 ;
  assign n34556 = ~n6640 ;
  assign n6946 = n34556 & n163 ;
  assign n7107 = n6699 | n6946 ;
  assign n34557 = ~n6897 ;
  assign n7108 = n34557 & n7107 ;
  assign n7123 = n5352 | n7121 ;
  assign n34558 = ~n7123 ;
  assign n7132 = n34558 & n7129 ;
  assign n7133 = n7108 | n7132 ;
  assign n34559 = ~n7131 ;
  assign n7134 = n34559 & n7133 ;
  assign n34560 = ~n7134 ;
  assign n7135 = n4934 & n34560 ;
  assign n6703 = n6562 & n34333 ;
  assign n34561 = ~n6709 ;
  assign n6710 = n6703 & n34561 ;
  assign n6896 = n6710 & n6889 ;
  assign n6711 = n6702 | n6709 ;
  assign n34562 = ~n6711 ;
  assign n6954 = n34562 & n163 ;
  assign n6955 = n6562 | n6954 ;
  assign n34563 = ~n6896 ;
  assign n6956 = n34563 & n6955 ;
  assign n7139 = n5352 & n34554 ;
  assign n7140 = n4934 | n7139 ;
  assign n34564 = ~n7140 ;
  assign n7141 = n7133 & n34564 ;
  assign n7142 = n6956 | n7141 ;
  assign n34565 = ~n7135 ;
  assign n7143 = n34565 & n7142 ;
  assign n34566 = ~n7143 ;
  assign n7144 = n169 & n34566 ;
  assign n7100 = n6714 | n6716 ;
  assign n34567 = ~n7100 ;
  assign n7101 = n163 & n34567 ;
  assign n7102 = n6608 | n7101 ;
  assign n34568 = ~n6716 ;
  assign n7103 = n6608 & n34568 ;
  assign n7104 = n34339 & n7103 ;
  assign n7105 = n6889 & n7104 ;
  assign n34569 = ~n7105 ;
  assign n7106 = n7102 & n34569 ;
  assign n7136 = n169 | n7135 ;
  assign n34570 = ~n7136 ;
  assign n7145 = n34570 & n7142 ;
  assign n7146 = n7106 | n7145 ;
  assign n34571 = ~n7144 ;
  assign n7147 = n34571 & n7146 ;
  assign n34572 = ~n7147 ;
  assign n7148 = n170 & n34572 ;
  assign n6721 = n6611 & n34345 ;
  assign n34573 = ~n6722 ;
  assign n7094 = n6721 & n34573 ;
  assign n7095 = n6889 & n7094 ;
  assign n7096 = n6719 | n6722 ;
  assign n34574 = ~n7096 ;
  assign n7097 = n163 & n34574 ;
  assign n7098 = n6611 | n7097 ;
  assign n34575 = ~n7095 ;
  assign n7099 = n34575 & n7098 ;
  assign n34576 = ~n7139 ;
  assign n7151 = n7133 & n34576 ;
  assign n34577 = ~n7151 ;
  assign n7152 = n168 & n34577 ;
  assign n34578 = ~n7152 ;
  assign n7153 = n7142 & n34578 ;
  assign n34579 = ~n7153 ;
  assign n7154 = n169 & n34579 ;
  assign n7155 = n170 | n7154 ;
  assign n34580 = ~n7155 ;
  assign n7156 = n7146 & n34580 ;
  assign n7157 = n7099 | n7156 ;
  assign n34581 = ~n7148 ;
  assign n7158 = n34581 & n7157 ;
  assign n34582 = ~n7158 ;
  assign n7159 = n171 & n34582 ;
  assign n34583 = ~n6726 ;
  assign n7087 = n6627 & n34583 ;
  assign n7088 = n34351 & n7087 ;
  assign n7089 = n6889 & n7088 ;
  assign n7090 = n6725 | n6726 ;
  assign n34584 = ~n7090 ;
  assign n7091 = n163 & n34584 ;
  assign n7092 = n6627 | n7091 ;
  assign n34585 = ~n7089 ;
  assign n7093 = n34585 & n7092 ;
  assign n7149 = n3940 | n7148 ;
  assign n34586 = ~n7149 ;
  assign n7160 = n34586 & n7157 ;
  assign n7161 = n7093 | n7160 ;
  assign n34587 = ~n7159 ;
  assign n7162 = n34587 & n7161 ;
  assign n34588 = ~n7162 ;
  assign n7163 = n3631 & n34588 ;
  assign n6731 = n6606 & n34357 ;
  assign n34589 = ~n6733 ;
  assign n7081 = n6731 & n34589 ;
  assign n7082 = n6889 & n7081 ;
  assign n7083 = n6733 | n6743 ;
  assign n34590 = ~n7083 ;
  assign n7084 = n163 & n34590 ;
  assign n7085 = n6606 | n7084 ;
  assign n34591 = ~n7082 ;
  assign n7086 = n34591 & n7085 ;
  assign n34592 = ~n7154 ;
  assign n7166 = n7146 & n34592 ;
  assign n34593 = ~n7166 ;
  assign n7167 = n170 & n34593 ;
  assign n34594 = ~n7167 ;
  assign n7170 = n7157 & n34594 ;
  assign n34595 = ~n7170 ;
  assign n7171 = n3940 & n34595 ;
  assign n7172 = n3631 | n7171 ;
  assign n34596 = ~n7172 ;
  assign n7173 = n7161 & n34596 ;
  assign n7174 = n7086 | n7173 ;
  assign n34597 = ~n7163 ;
  assign n7175 = n34597 & n7174 ;
  assign n34598 = ~n7175 ;
  assign n7176 = n173 & n34598 ;
  assign n34599 = ~n6737 ;
  assign n7074 = n6629 & n34599 ;
  assign n7075 = n34382 & n7074 ;
  assign n7076 = n6889 & n7075 ;
  assign n7077 = n6737 | n6745 ;
  assign n34600 = ~n7077 ;
  assign n7078 = n163 & n34600 ;
  assign n7079 = n6629 | n7078 ;
  assign n34601 = ~n7076 ;
  assign n7080 = n34601 & n7079 ;
  assign n7164 = n173 | n7163 ;
  assign n34602 = ~n7164 ;
  assign n7177 = n34602 & n7174 ;
  assign n7178 = n7080 | n7177 ;
  assign n34603 = ~n7176 ;
  assign n7179 = n34603 & n7178 ;
  assign n34604 = ~n7179 ;
  assign n7180 = n174 & n34604 ;
  assign n6742 = n6604 & n34371 ;
  assign n34605 = ~n6747 ;
  assign n7068 = n6742 & n34605 ;
  assign n7069 = n6889 & n7068 ;
  assign n7070 = n6740 | n6747 ;
  assign n34606 = ~n7070 ;
  assign n7071 = n163 & n34606 ;
  assign n7072 = n6604 | n7071 ;
  assign n34607 = ~n7069 ;
  assign n7073 = n34607 & n7072 ;
  assign n34608 = ~n7171 ;
  assign n7183 = n7161 & n34608 ;
  assign n34609 = ~n7183 ;
  assign n7184 = n172 & n34609 ;
  assign n34610 = ~n7184 ;
  assign n7185 = n7174 & n34610 ;
  assign n34611 = ~n7185 ;
  assign n7186 = n173 & n34611 ;
  assign n7187 = n174 | n7186 ;
  assign n34612 = ~n7187 ;
  assign n7188 = n7178 & n34612 ;
  assign n7189 = n7073 | n7188 ;
  assign n34613 = ~n7180 ;
  assign n7190 = n34613 & n7189 ;
  assign n34614 = ~n7190 ;
  assign n7191 = n175 & n34614 ;
  assign n34615 = ~n6751 ;
  assign n7061 = n6602 & n34615 ;
  assign n7062 = n34398 & n7061 ;
  assign n7063 = n6889 & n7062 ;
  assign n7064 = n6751 | n6760 ;
  assign n34616 = ~n7064 ;
  assign n7065 = n163 & n34616 ;
  assign n7066 = n6602 | n7065 ;
  assign n34617 = ~n7063 ;
  assign n7067 = n34617 & n7066 ;
  assign n7181 = n2753 | n7180 ;
  assign n34618 = ~n7181 ;
  assign n7192 = n34618 & n7189 ;
  assign n7193 = n7067 | n7192 ;
  assign n34619 = ~n7191 ;
  assign n7194 = n34619 & n7193 ;
  assign n34620 = ~n7194 ;
  assign n7195 = n2431 & n34620 ;
  assign n6756 = n6647 & n34387 ;
  assign n34621 = ~n6762 ;
  assign n7055 = n6756 & n34621 ;
  assign n7056 = n6889 & n7055 ;
  assign n7057 = n6754 | n6762 ;
  assign n34622 = ~n7057 ;
  assign n7058 = n163 & n34622 ;
  assign n7059 = n6647 | n7058 ;
  assign n34623 = ~n7056 ;
  assign n7060 = n34623 & n7059 ;
  assign n34624 = ~n7186 ;
  assign n7198 = n7178 & n34624 ;
  assign n34625 = ~n7198 ;
  assign n7199 = n174 & n34625 ;
  assign n34626 = ~n7199 ;
  assign n7200 = n7189 & n34626 ;
  assign n34627 = ~n7200 ;
  assign n7201 = n2753 & n34627 ;
  assign n7202 = n2431 | n7201 ;
  assign n34628 = ~n7202 ;
  assign n7203 = n7193 & n34628 ;
  assign n7204 = n7060 | n7203 ;
  assign n34629 = ~n7195 ;
  assign n7205 = n34629 & n7204 ;
  assign n34630 = ~n7205 ;
  assign n7206 = n177 & n34630 ;
  assign n34631 = ~n6766 ;
  assign n7048 = n6651 & n34631 ;
  assign n7049 = n34414 & n7048 ;
  assign n7050 = n6889 & n7049 ;
  assign n7051 = n6766 | n6775 ;
  assign n34632 = ~n7051 ;
  assign n7052 = n163 & n34632 ;
  assign n7053 = n6651 | n7052 ;
  assign n34633 = ~n7050 ;
  assign n7054 = n34633 & n7053 ;
  assign n7196 = n177 | n7195 ;
  assign n34634 = ~n7196 ;
  assign n7207 = n34634 & n7204 ;
  assign n7208 = n7054 | n7207 ;
  assign n34635 = ~n7206 ;
  assign n7209 = n34635 & n7208 ;
  assign n34636 = ~n7209 ;
  assign n7210 = n178 & n34636 ;
  assign n6771 = n6653 & n34403 ;
  assign n34637 = ~n6777 ;
  assign n7042 = n6771 & n34637 ;
  assign n7043 = n6889 & n7042 ;
  assign n7044 = n6769 | n6777 ;
  assign n34638 = ~n7044 ;
  assign n7045 = n163 & n34638 ;
  assign n7046 = n6653 | n7045 ;
  assign n34639 = ~n7043 ;
  assign n7047 = n34639 & n7046 ;
  assign n34640 = ~n7201 ;
  assign n7213 = n7193 & n34640 ;
  assign n34641 = ~n7213 ;
  assign n7214 = n176 & n34641 ;
  assign n34642 = ~n7214 ;
  assign n7215 = n7204 & n34642 ;
  assign n34643 = ~n7215 ;
  assign n7216 = n177 & n34643 ;
  assign n7217 = n178 | n7216 ;
  assign n34644 = ~n7217 ;
  assign n7218 = n7208 & n34644 ;
  assign n7219 = n7047 | n7218 ;
  assign n34645 = ~n7210 ;
  assign n7220 = n34645 & n7219 ;
  assign n34646 = ~n7220 ;
  assign n7221 = n179 & n34646 ;
  assign n34647 = ~n6781 ;
  assign n7035 = n6655 & n34647 ;
  assign n7036 = n34430 & n7035 ;
  assign n7037 = n6889 & n7036 ;
  assign n7038 = n6781 | n6790 ;
  assign n34648 = ~n7038 ;
  assign n7039 = n163 & n34648 ;
  assign n7040 = n6655 | n7039 ;
  assign n34649 = ~n7037 ;
  assign n7041 = n34649 & n7040 ;
  assign n7211 = n1707 | n7210 ;
  assign n34650 = ~n7211 ;
  assign n7222 = n34650 & n7219 ;
  assign n7223 = n7041 | n7222 ;
  assign n34651 = ~n7221 ;
  assign n7224 = n34651 & n7223 ;
  assign n34652 = ~n7224 ;
  assign n7225 = n1487 & n34652 ;
  assign n6786 = n6657 & n34419 ;
  assign n34653 = ~n6792 ;
  assign n7029 = n6786 & n34653 ;
  assign n7030 = n6889 & n7029 ;
  assign n7031 = n6784 | n6792 ;
  assign n34654 = ~n7031 ;
  assign n7032 = n163 & n34654 ;
  assign n7033 = n6657 | n7032 ;
  assign n34655 = ~n7030 ;
  assign n7034 = n34655 & n7033 ;
  assign n34656 = ~n7216 ;
  assign n7228 = n7208 & n34656 ;
  assign n34657 = ~n7228 ;
  assign n7229 = n178 & n34657 ;
  assign n34658 = ~n7229 ;
  assign n7230 = n7219 & n34658 ;
  assign n34659 = ~n7230 ;
  assign n7231 = n1707 & n34659 ;
  assign n7232 = n1487 | n7231 ;
  assign n34660 = ~n7232 ;
  assign n7233 = n7223 & n34660 ;
  assign n7234 = n7034 | n7233 ;
  assign n34661 = ~n7225 ;
  assign n7235 = n34661 & n7234 ;
  assign n34662 = ~n7235 ;
  assign n7236 = n181 & n34662 ;
  assign n34663 = ~n6796 ;
  assign n7022 = n6659 & n34663 ;
  assign n7023 = n34446 & n7022 ;
  assign n7024 = n6889 & n7023 ;
  assign n7025 = n6796 | n6805 ;
  assign n34664 = ~n7025 ;
  assign n7026 = n163 & n34664 ;
  assign n7027 = n6659 | n7026 ;
  assign n34665 = ~n7024 ;
  assign n7028 = n34665 & n7027 ;
  assign n7226 = n181 | n7225 ;
  assign n34666 = ~n7226 ;
  assign n7237 = n34666 & n7234 ;
  assign n7238 = n7028 | n7237 ;
  assign n34667 = ~n7236 ;
  assign n7239 = n34667 & n7238 ;
  assign n34668 = ~n7239 ;
  assign n7240 = n182 & n34668 ;
  assign n6801 = n6625 & n34435 ;
  assign n34669 = ~n6807 ;
  assign n7016 = n6801 & n34669 ;
  assign n7017 = n6889 & n7016 ;
  assign n7018 = n6799 | n6807 ;
  assign n34670 = ~n7018 ;
  assign n7019 = n163 & n34670 ;
  assign n7020 = n6625 | n7019 ;
  assign n34671 = ~n7017 ;
  assign n7021 = n34671 & n7020 ;
  assign n34672 = ~n7231 ;
  assign n7243 = n7223 & n34672 ;
  assign n34673 = ~n7243 ;
  assign n7244 = n180 & n34673 ;
  assign n34674 = ~n7244 ;
  assign n7245 = n7234 & n34674 ;
  assign n34675 = ~n7245 ;
  assign n7246 = n181 & n34675 ;
  assign n7247 = n182 | n7246 ;
  assign n34676 = ~n7247 ;
  assign n7248 = n7238 & n34676 ;
  assign n7249 = n7021 | n7248 ;
  assign n34677 = ~n7240 ;
  assign n7250 = n34677 & n7249 ;
  assign n34678 = ~n7250 ;
  assign n7251 = n183 & n34678 ;
  assign n34679 = ~n6811 ;
  assign n7009 = n6661 & n34679 ;
  assign n7010 = n34462 & n7009 ;
  assign n7011 = n6889 & n7010 ;
  assign n7012 = n6811 | n6820 ;
  assign n34680 = ~n7012 ;
  assign n7013 = n163 & n34680 ;
  assign n7014 = n6661 | n7013 ;
  assign n34681 = ~n7011 ;
  assign n7015 = n34681 & n7014 ;
  assign n7241 = n183 | n7240 ;
  assign n34682 = ~n7241 ;
  assign n7252 = n34682 & n7249 ;
  assign n7253 = n7015 | n7252 ;
  assign n34683 = ~n7251 ;
  assign n7254 = n34683 & n7253 ;
  assign n34684 = ~n7254 ;
  assign n7255 = n838 & n34684 ;
  assign n6816 = n6663 & n34451 ;
  assign n34685 = ~n6822 ;
  assign n7003 = n6816 & n34685 ;
  assign n7004 = n6889 & n7003 ;
  assign n7005 = n6814 | n6822 ;
  assign n34686 = ~n7005 ;
  assign n7006 = n163 & n34686 ;
  assign n7007 = n6663 | n7006 ;
  assign n34687 = ~n7004 ;
  assign n7008 = n34687 & n7007 ;
  assign n34688 = ~n7246 ;
  assign n7258 = n7238 & n34688 ;
  assign n34689 = ~n7258 ;
  assign n7259 = n182 & n34689 ;
  assign n34690 = ~n7259 ;
  assign n7260 = n7249 & n34690 ;
  assign n34691 = ~n7260 ;
  assign n7261 = n996 & n34691 ;
  assign n7262 = n838 | n7261 ;
  assign n34692 = ~n7262 ;
  assign n7263 = n7253 & n34692 ;
  assign n7264 = n7008 | n7263 ;
  assign n34693 = ~n7255 ;
  assign n7265 = n34693 & n7264 ;
  assign n34694 = ~n7265 ;
  assign n7266 = n185 & n34694 ;
  assign n34695 = ~n6826 ;
  assign n6996 = n6665 & n34695 ;
  assign n6997 = n34478 & n6996 ;
  assign n6998 = n6889 & n6997 ;
  assign n6999 = n6826 | n6835 ;
  assign n34696 = ~n6999 ;
  assign n7000 = n163 & n34696 ;
  assign n7001 = n6665 | n7000 ;
  assign n34697 = ~n6998 ;
  assign n7002 = n34697 & n7001 ;
  assign n7256 = n185 | n7255 ;
  assign n34698 = ~n7256 ;
  assign n7267 = n34698 & n7264 ;
  assign n7268 = n7002 | n7267 ;
  assign n34699 = ~n7266 ;
  assign n7269 = n34699 & n7268 ;
  assign n34700 = ~n7269 ;
  assign n7270 = n186 & n34700 ;
  assign n6831 = n6667 & n34467 ;
  assign n34701 = ~n6837 ;
  assign n6990 = n6831 & n34701 ;
  assign n6991 = n6889 & n6990 ;
  assign n6992 = n6829 | n6837 ;
  assign n34702 = ~n6992 ;
  assign n6993 = n163 & n34702 ;
  assign n6994 = n6667 | n6993 ;
  assign n34703 = ~n6991 ;
  assign n6995 = n34703 & n6994 ;
  assign n34704 = ~n7261 ;
  assign n7273 = n7253 & n34704 ;
  assign n34705 = ~n7273 ;
  assign n7274 = n184 & n34705 ;
  assign n34706 = ~n7274 ;
  assign n7275 = n7264 & n34706 ;
  assign n34707 = ~n7275 ;
  assign n7276 = n185 & n34707 ;
  assign n7277 = n186 | n7276 ;
  assign n34708 = ~n7277 ;
  assign n7278 = n7268 & n34708 ;
  assign n7279 = n6995 | n7278 ;
  assign n34709 = ~n7270 ;
  assign n7280 = n34709 & n7279 ;
  assign n34710 = ~n7280 ;
  assign n7281 = n187 & n34710 ;
  assign n34711 = ~n6841 ;
  assign n6983 = n6669 & n34711 ;
  assign n6984 = n34494 & n6983 ;
  assign n6985 = n6889 & n6984 ;
  assign n6986 = n6841 | n6850 ;
  assign n34712 = ~n6986 ;
  assign n6987 = n163 & n34712 ;
  assign n6988 = n6669 | n6987 ;
  assign n34713 = ~n6985 ;
  assign n6989 = n34713 & n6988 ;
  assign n7271 = n528 | n7270 ;
  assign n34714 = ~n7271 ;
  assign n7282 = n34714 & n7279 ;
  assign n7283 = n6989 | n7282 ;
  assign n34715 = ~n7281 ;
  assign n7284 = n34715 & n7283 ;
  assign n34716 = ~n7284 ;
  assign n7285 = n413 & n34716 ;
  assign n7286 = n189 | n7285 ;
  assign n6846 = n6645 & n34483 ;
  assign n34717 = ~n6852 ;
  assign n6977 = n6846 & n34717 ;
  assign n6978 = n6889 & n6977 ;
  assign n6979 = n6844 | n6852 ;
  assign n34718 = ~n6979 ;
  assign n6980 = n163 & n34718 ;
  assign n6981 = n6645 | n6980 ;
  assign n34719 = ~n6978 ;
  assign n6982 = n34719 & n6981 ;
  assign n34720 = ~n7276 ;
  assign n7288 = n7268 & n34720 ;
  assign n34721 = ~n7288 ;
  assign n7289 = n186 & n34721 ;
  assign n34722 = ~n7289 ;
  assign n7290 = n7279 & n34722 ;
  assign n34723 = ~n7290 ;
  assign n7291 = n528 & n34723 ;
  assign n7292 = n413 | n7291 ;
  assign n34724 = ~n7292 ;
  assign n7293 = n7283 & n34724 ;
  assign n7294 = n6982 | n7293 ;
  assign n34725 = ~n7286 ;
  assign n7297 = n34725 & n7294 ;
  assign n7298 = n6976 | n7297 ;
  assign n34726 = ~n7291 ;
  assign n7303 = n7283 & n34726 ;
  assign n34727 = ~n7303 ;
  assign n7304 = n188 & n34727 ;
  assign n34728 = ~n7304 ;
  assign n7305 = n7294 & n34728 ;
  assign n34729 = ~n7305 ;
  assign n7306 = n189 & n34729 ;
  assign n34730 = ~n7306 ;
  assign n7308 = n7298 & n34730 ;
  assign n34731 = ~n7308 ;
  assign n7309 = n190 & n34731 ;
  assign n6861 = n6675 & n34499 ;
  assign n34732 = ~n6867 ;
  assign n6964 = n6861 & n34732 ;
  assign n6965 = n163 & n6964 ;
  assign n6966 = n6859 | n6867 ;
  assign n34733 = ~n6966 ;
  assign n6967 = n163 & n34733 ;
  assign n6968 = n6675 | n6967 ;
  assign n34734 = ~n6965 ;
  assign n6969 = n34734 & n6968 ;
  assign n7307 = n190 | n7306 ;
  assign n34735 = ~n7307 ;
  assign n7310 = n7298 & n34735 ;
  assign n7311 = n6969 | n7310 ;
  assign n34736 = ~n7309 ;
  assign n7314 = n34736 & n7311 ;
  assign n34737 = ~n7314 ;
  assign n7315 = n287 & n34737 ;
  assign n34738 = ~n6871 ;
  assign n6957 = n6673 & n34738 ;
  assign n6958 = n34523 & n6957 ;
  assign n6959 = n163 & n6958 ;
  assign n6960 = n6871 | n6880 ;
  assign n34739 = ~n6960 ;
  assign n6961 = n163 & n34739 ;
  assign n6962 = n6673 | n6961 ;
  assign n34740 = ~n6959 ;
  assign n6963 = n34740 & n6962 ;
  assign n34741 = ~n7285 ;
  assign n7295 = n34741 & n7294 ;
  assign n34742 = ~n7295 ;
  assign n7296 = n189 & n34742 ;
  assign n34743 = ~n7296 ;
  assign n7299 = n34743 & n7298 ;
  assign n34744 = ~n7299 ;
  assign n7300 = n190 & n34744 ;
  assign n7301 = n287 | n7300 ;
  assign n34745 = ~n7301 ;
  assign n7312 = n34745 & n7311 ;
  assign n7319 = n6963 | n7312 ;
  assign n34746 = ~n7315 ;
  assign n7320 = n34746 & n7319 ;
  assign n7321 = n6944 | n7320 ;
  assign n7322 = n31336 & n7321 ;
  assign n6686 = n6621 | n6682 ;
  assign n34747 = ~n6686 ;
  assign n6687 = n6544 & n34747 ;
  assign n6688 = n34540 & n6687 ;
  assign n6909 = n6688 & n34541 ;
  assign n6910 = n34542 & n6909 ;
  assign n6918 = n192 & n6915 ;
  assign n34748 = ~n6622 ;
  assign n6947 = n34748 & n163 ;
  assign n34749 = ~n6947 ;
  assign n6948 = n6884 & n34749 ;
  assign n34750 = ~n6948 ;
  assign n6949 = n6918 & n34750 ;
  assign n6950 = n6910 | n6949 ;
  assign n7316 = n6943 & n34746 ;
  assign n7325 = n7316 & n7319 ;
  assign n7326 = n6950 | n7325 ;
  assign n162 = n7322 | n7326 ;
  assign n7318 = n7312 | n7315 ;
  assign n34751 = ~n7318 ;
  assign n7328 = n34751 & n162 ;
  assign n7329 = n6963 | n7328 ;
  assign n34752 = ~n7312 ;
  assign n7313 = n6963 & n34752 ;
  assign n7317 = n7313 & n34746 ;
  assign n7346 = n7317 & n162 ;
  assign n34753 = ~n7346 ;
  assign n7347 = n7329 & n34753 ;
  assign n7323 = n6943 | n7320 ;
  assign n34754 = ~n7323 ;
  assign n7342 = n34754 & n162 ;
  assign n7398 = n7325 | n7342 ;
  assign n7399 = n7347 | n7398 ;
  assign n15623 = x64 | x65 ;
  assign n16342 = x66 | n15623 ;
  assign n7335 = x66 & n162 ;
  assign n34755 = ~n7335 ;
  assign n7336 = n16342 & n34755 ;
  assign n34756 = ~n7336 ;
  assign n7337 = n163 & n34756 ;
  assign n6689 = n16342 & n34539 ;
  assign n6690 = n34540 & n6689 ;
  assign n6913 = n6690 & n34541 ;
  assign n6914 = n34542 & n6913 ;
  assign n7345 = n6914 & n34755 ;
  assign n34757 = ~n13540 ;
  assign n7334 = n34757 & n162 ;
  assign n34758 = ~x66 ;
  assign n7355 = n34758 & n162 ;
  assign n34759 = ~n7355 ;
  assign n7356 = x67 & n34759 ;
  assign n7357 = n7334 | n7356 ;
  assign n7358 = n7345 | n7357 ;
  assign n34760 = ~n7337 ;
  assign n7361 = n34760 & n7358 ;
  assign n34761 = ~n7361 ;
  assign n7362 = n6600 & n34761 ;
  assign n17060 = n34758 & n15623 ;
  assign n34762 = ~n162 ;
  assign n7350 = x66 & n34762 ;
  assign n7351 = n17060 | n7350 ;
  assign n34763 = ~n7351 ;
  assign n7352 = n6889 & n34763 ;
  assign n7353 = n6600 | n7352 ;
  assign n34764 = ~n7353 ;
  assign n7359 = n34764 & n7358 ;
  assign n34765 = ~n6910 ;
  assign n6911 = n6889 & n34765 ;
  assign n34766 = ~n6949 ;
  assign n6951 = n6911 & n34766 ;
  assign n34767 = ~n7325 ;
  assign n7367 = n6951 & n34767 ;
  assign n34768 = ~n7322 ;
  assign n7368 = n34768 & n7367 ;
  assign n7369 = n7334 | n7368 ;
  assign n7370 = x68 & n7369 ;
  assign n7371 = x68 | n7368 ;
  assign n7372 = n7334 | n7371 ;
  assign n34769 = ~n7370 ;
  assign n7373 = n34769 & n7372 ;
  assign n7374 = n7359 | n7373 ;
  assign n34770 = ~n7362 ;
  assign n7375 = n34770 & n7374 ;
  assign n34771 = ~n7375 ;
  assign n7376 = n165 & n34771 ;
  assign n7124 = n6900 | n7113 ;
  assign n34772 = ~n7124 ;
  assign n7343 = n34772 & n162 ;
  assign n7344 = n6895 | n7343 ;
  assign n7125 = n6895 & n34772 ;
  assign n7348 = n7125 & n162 ;
  assign n34773 = ~n7348 ;
  assign n7349 = n7344 & n34773 ;
  assign n7363 = n165 | n7362 ;
  assign n34774 = ~n7363 ;
  assign n7379 = n34774 & n7374 ;
  assign n7380 = n7349 | n7379 ;
  assign n34775 = ~n7376 ;
  assign n7381 = n34775 & n7380 ;
  assign n34776 = ~n7381 ;
  assign n7382 = n166 & n34776 ;
  assign n7377 = n166 | n7376 ;
  assign n34777 = ~n7377 ;
  assign n7383 = n34777 & n7380 ;
  assign n34778 = ~n7126 ;
  assign n7138 = n6908 & n34778 ;
  assign n7568 = n34547 & n7138 ;
  assign n7569 = n162 & n7568 ;
  assign n7570 = n7116 | n7126 ;
  assign n34779 = ~n7570 ;
  assign n7571 = n162 & n34779 ;
  assign n7572 = n6908 | n7571 ;
  assign n34780 = ~n7569 ;
  assign n7573 = n34780 & n7572 ;
  assign n7574 = n7383 | n7573 ;
  assign n34781 = ~n7382 ;
  assign n7575 = n34781 & n7574 ;
  assign n34782 = ~n7575 ;
  assign n7576 = n5352 & n34782 ;
  assign n7122 = n6940 & n34553 ;
  assign n34783 = ~n7128 ;
  assign n7562 = n7122 & n34783 ;
  assign n7563 = n162 & n7562 ;
  assign n7564 = n7121 | n7128 ;
  assign n34784 = ~n7564 ;
  assign n7565 = n162 & n34784 ;
  assign n7566 = n6940 | n7565 ;
  assign n34785 = ~n7563 ;
  assign n7567 = n34785 & n7566 ;
  assign n7364 = n164 & n34761 ;
  assign n7338 = n164 | n7337 ;
  assign n34786 = ~n7338 ;
  assign n7366 = n34786 & n7358 ;
  assign n7388 = n7366 | n7373 ;
  assign n34787 = ~n7364 ;
  assign n7389 = n34787 & n7388 ;
  assign n34788 = ~n7389 ;
  assign n7390 = n165 & n34788 ;
  assign n7391 = n34774 & n7388 ;
  assign n7392 = n7349 | n7391 ;
  assign n34789 = ~n7390 ;
  assign n7393 = n34789 & n7392 ;
  assign n34790 = ~n7393 ;
  assign n7394 = n166 & n34790 ;
  assign n7395 = n5352 | n7394 ;
  assign n34791 = ~n7395 ;
  assign n7579 = n34791 & n7574 ;
  assign n7580 = n7567 | n7579 ;
  assign n34792 = ~n7576 ;
  assign n7581 = n34792 & n7580 ;
  assign n34793 = ~n7581 ;
  assign n7582 = n168 & n34793 ;
  assign n34794 = ~n7132 ;
  assign n7555 = n7108 & n34794 ;
  assign n7556 = n34576 & n7555 ;
  assign n7557 = n162 & n7556 ;
  assign n7558 = n7132 | n7139 ;
  assign n34795 = ~n7558 ;
  assign n7559 = n162 & n34795 ;
  assign n7560 = n7108 | n7559 ;
  assign n34796 = ~n7557 ;
  assign n7561 = n34796 & n7560 ;
  assign n7577 = n4934 | n7576 ;
  assign n34797 = ~n7577 ;
  assign n7583 = n34797 & n7580 ;
  assign n7584 = n7561 | n7583 ;
  assign n34798 = ~n7582 ;
  assign n7585 = n34798 & n7584 ;
  assign n34799 = ~n7585 ;
  assign n7586 = n169 & n34799 ;
  assign n7137 = n6956 & n34565 ;
  assign n34800 = ~n7141 ;
  assign n7549 = n7137 & n34800 ;
  assign n7550 = n162 & n7549 ;
  assign n7551 = n7141 | n7152 ;
  assign n34801 = ~n7551 ;
  assign n7552 = n162 & n34801 ;
  assign n7553 = n6956 | n7552 ;
  assign n34802 = ~n7550 ;
  assign n7554 = n34802 & n7553 ;
  assign n7397 = n34777 & n7392 ;
  assign n7595 = n7397 | n7573 ;
  assign n34803 = ~n7394 ;
  assign n7596 = n34803 & n7595 ;
  assign n34804 = ~n7596 ;
  assign n7597 = n167 & n34804 ;
  assign n7598 = n34791 & n7595 ;
  assign n7599 = n7567 | n7598 ;
  assign n34805 = ~n7597 ;
  assign n7600 = n34805 & n7599 ;
  assign n34806 = ~n7600 ;
  assign n7601 = n4934 & n34806 ;
  assign n7602 = n169 | n7601 ;
  assign n34807 = ~n7602 ;
  assign n7603 = n7584 & n34807 ;
  assign n7604 = n7554 | n7603 ;
  assign n34808 = ~n7586 ;
  assign n7605 = n34808 & n7604 ;
  assign n34809 = ~n7605 ;
  assign n7606 = n170 & n34809 ;
  assign n34810 = ~n7145 ;
  assign n7542 = n7106 & n34810 ;
  assign n7543 = n34592 & n7542 ;
  assign n7544 = n162 & n7543 ;
  assign n7545 = n7145 | n7154 ;
  assign n34811 = ~n7545 ;
  assign n7546 = n162 & n34811 ;
  assign n7547 = n7106 | n7546 ;
  assign n34812 = ~n7544 ;
  assign n7548 = n34812 & n7547 ;
  assign n7587 = n170 | n7586 ;
  assign n34813 = ~n7587 ;
  assign n7607 = n34813 & n7604 ;
  assign n7608 = n7548 | n7607 ;
  assign n34814 = ~n7606 ;
  assign n7609 = n34814 & n7608 ;
  assign n34815 = ~n7609 ;
  assign n7610 = n3940 & n34815 ;
  assign n7150 = n7099 & n34581 ;
  assign n34816 = ~n7156 ;
  assign n7168 = n7150 & n34816 ;
  assign n7330 = n7168 & n162 ;
  assign n7169 = n7156 | n7167 ;
  assign n34817 = ~n7169 ;
  assign n7331 = n34817 & n162 ;
  assign n7332 = n7099 | n7331 ;
  assign n34818 = ~n7330 ;
  assign n7333 = n34818 & n7332 ;
  assign n7618 = n34797 & n7599 ;
  assign n7619 = n7561 | n7618 ;
  assign n34819 = ~n7601 ;
  assign n7620 = n34819 & n7619 ;
  assign n34820 = ~n7620 ;
  assign n7621 = n169 & n34820 ;
  assign n7622 = n34807 & n7619 ;
  assign n7623 = n7554 | n7622 ;
  assign n34821 = ~n7621 ;
  assign n7624 = n34821 & n7623 ;
  assign n34822 = ~n7624 ;
  assign n7625 = n170 & n34822 ;
  assign n7626 = n3940 | n7625 ;
  assign n34823 = ~n7626 ;
  assign n7627 = n7608 & n34823 ;
  assign n7628 = n7333 | n7627 ;
  assign n34824 = ~n7610 ;
  assign n7629 = n34824 & n7628 ;
  assign n34825 = ~n7629 ;
  assign n7630 = n172 & n34825 ;
  assign n34826 = ~n7160 ;
  assign n7535 = n7093 & n34826 ;
  assign n7536 = n34608 & n7535 ;
  assign n7537 = n162 & n7536 ;
  assign n7538 = n7160 | n7171 ;
  assign n34827 = ~n7538 ;
  assign n7539 = n162 & n34827 ;
  assign n7540 = n7093 | n7539 ;
  assign n34828 = ~n7537 ;
  assign n7541 = n34828 & n7540 ;
  assign n7612 = n3631 | n7610 ;
  assign n34829 = ~n7612 ;
  assign n7631 = n34829 & n7628 ;
  assign n7632 = n7541 | n7631 ;
  assign n34830 = ~n7630 ;
  assign n7633 = n34830 & n7632 ;
  assign n34831 = ~n7633 ;
  assign n7634 = n173 & n34831 ;
  assign n7529 = n7173 | n7184 ;
  assign n34832 = ~n7529 ;
  assign n7530 = n162 & n34832 ;
  assign n7531 = n7086 | n7530 ;
  assign n7165 = n7086 & n34597 ;
  assign n34833 = ~n7173 ;
  assign n7532 = n7165 & n34833 ;
  assign n7533 = n162 & n7532 ;
  assign n34834 = ~n7533 ;
  assign n7534 = n7531 & n34834 ;
  assign n7642 = n34813 & n7623 ;
  assign n7643 = n7548 | n7642 ;
  assign n34835 = ~n7625 ;
  assign n7644 = n34835 & n7643 ;
  assign n34836 = ~n7644 ;
  assign n7645 = n171 & n34836 ;
  assign n7646 = n34823 & n7643 ;
  assign n7647 = n7333 | n7646 ;
  assign n34837 = ~n7645 ;
  assign n7648 = n34837 & n7647 ;
  assign n34838 = ~n7648 ;
  assign n7649 = n3631 & n34838 ;
  assign n7650 = n173 | n7649 ;
  assign n34839 = ~n7650 ;
  assign n7651 = n7632 & n34839 ;
  assign n7652 = n7534 | n7651 ;
  assign n34840 = ~n7634 ;
  assign n7653 = n34840 & n7652 ;
  assign n34841 = ~n7653 ;
  assign n7654 = n174 & n34841 ;
  assign n34842 = ~n7177 ;
  assign n7522 = n7080 & n34842 ;
  assign n7523 = n34624 & n7522 ;
  assign n7524 = n162 & n7523 ;
  assign n7525 = n7177 | n7186 ;
  assign n34843 = ~n7525 ;
  assign n7526 = n162 & n34843 ;
  assign n7527 = n7080 | n7526 ;
  assign n34844 = ~n7524 ;
  assign n7528 = n34844 & n7527 ;
  assign n7635 = n174 | n7634 ;
  assign n34845 = ~n7635 ;
  assign n7655 = n34845 & n7652 ;
  assign n7656 = n7528 | n7655 ;
  assign n34846 = ~n7654 ;
  assign n7657 = n34846 & n7656 ;
  assign n34847 = ~n7657 ;
  assign n7658 = n2753 & n34847 ;
  assign n7182 = n7073 & n34613 ;
  assign n34848 = ~n7188 ;
  assign n7516 = n7182 & n34848 ;
  assign n7517 = n162 & n7516 ;
  assign n7518 = n7188 | n7199 ;
  assign n34849 = ~n7518 ;
  assign n7519 = n162 & n34849 ;
  assign n7520 = n7073 | n7519 ;
  assign n34850 = ~n7517 ;
  assign n7521 = n34850 & n7520 ;
  assign n7666 = n34829 & n7647 ;
  assign n7667 = n7541 | n7666 ;
  assign n34851 = ~n7649 ;
  assign n7668 = n34851 & n7667 ;
  assign n34852 = ~n7668 ;
  assign n7669 = n173 & n34852 ;
  assign n7670 = n34839 & n7667 ;
  assign n7671 = n7534 | n7670 ;
  assign n34853 = ~n7669 ;
  assign n7672 = n34853 & n7671 ;
  assign n34854 = ~n7672 ;
  assign n7673 = n174 & n34854 ;
  assign n7674 = n2753 | n7673 ;
  assign n34855 = ~n7674 ;
  assign n7675 = n7656 & n34855 ;
  assign n7676 = n7521 | n7675 ;
  assign n34856 = ~n7658 ;
  assign n7677 = n34856 & n7676 ;
  assign n34857 = ~n7677 ;
  assign n7678 = n176 & n34857 ;
  assign n34858 = ~n7192 ;
  assign n7509 = n7067 & n34858 ;
  assign n7510 = n34640 & n7509 ;
  assign n7511 = n162 & n7510 ;
  assign n7512 = n7192 | n7201 ;
  assign n34859 = ~n7512 ;
  assign n7513 = n162 & n34859 ;
  assign n7514 = n7067 | n7513 ;
  assign n34860 = ~n7511 ;
  assign n7515 = n34860 & n7514 ;
  assign n7659 = n2431 | n7658 ;
  assign n34861 = ~n7659 ;
  assign n7679 = n34861 & n7676 ;
  assign n7680 = n7515 | n7679 ;
  assign n34862 = ~n7678 ;
  assign n7681 = n34862 & n7680 ;
  assign n34863 = ~n7681 ;
  assign n7682 = n177 & n34863 ;
  assign n7197 = n7060 & n34629 ;
  assign n34864 = ~n7203 ;
  assign n7503 = n7197 & n34864 ;
  assign n7504 = n162 & n7503 ;
  assign n7505 = n7203 | n7214 ;
  assign n34865 = ~n7505 ;
  assign n7506 = n162 & n34865 ;
  assign n7507 = n7060 | n7506 ;
  assign n34866 = ~n7504 ;
  assign n7508 = n34866 & n7507 ;
  assign n7690 = n34845 & n7671 ;
  assign n7691 = n7528 | n7690 ;
  assign n34867 = ~n7673 ;
  assign n7692 = n34867 & n7691 ;
  assign n34868 = ~n7692 ;
  assign n7693 = n175 & n34868 ;
  assign n7694 = n34855 & n7691 ;
  assign n7695 = n7521 | n7694 ;
  assign n34869 = ~n7693 ;
  assign n7696 = n34869 & n7695 ;
  assign n34870 = ~n7696 ;
  assign n7697 = n2431 & n34870 ;
  assign n7698 = n177 | n7697 ;
  assign n34871 = ~n7698 ;
  assign n7699 = n7680 & n34871 ;
  assign n7700 = n7508 | n7699 ;
  assign n34872 = ~n7682 ;
  assign n7701 = n34872 & n7700 ;
  assign n34873 = ~n7701 ;
  assign n7702 = n178 & n34873 ;
  assign n34874 = ~n7207 ;
  assign n7496 = n7054 & n34874 ;
  assign n7497 = n34656 & n7496 ;
  assign n7498 = n162 & n7497 ;
  assign n7499 = n7207 | n7216 ;
  assign n34875 = ~n7499 ;
  assign n7500 = n162 & n34875 ;
  assign n7501 = n7054 | n7500 ;
  assign n34876 = ~n7498 ;
  assign n7502 = n34876 & n7501 ;
  assign n7683 = n178 | n7682 ;
  assign n34877 = ~n7683 ;
  assign n7703 = n34877 & n7700 ;
  assign n7706 = n7502 | n7703 ;
  assign n34878 = ~n7702 ;
  assign n7707 = n34878 & n7706 ;
  assign n34879 = ~n7707 ;
  assign n7708 = n1707 & n34879 ;
  assign n7212 = n7047 & n34645 ;
  assign n34880 = ~n7218 ;
  assign n7490 = n7212 & n34880 ;
  assign n7491 = n162 & n7490 ;
  assign n7492 = n7218 | n7229 ;
  assign n34881 = ~n7492 ;
  assign n7493 = n162 & n34881 ;
  assign n7494 = n7047 | n7493 ;
  assign n34882 = ~n7491 ;
  assign n7495 = n34882 & n7494 ;
  assign n7714 = n34861 & n7695 ;
  assign n7715 = n7515 | n7714 ;
  assign n34883 = ~n7697 ;
  assign n7716 = n34883 & n7715 ;
  assign n34884 = ~n7716 ;
  assign n7717 = n177 & n34884 ;
  assign n7718 = n34871 & n7715 ;
  assign n7719 = n7508 | n7718 ;
  assign n34885 = ~n7717 ;
  assign n7720 = n34885 & n7719 ;
  assign n34886 = ~n7720 ;
  assign n7721 = n178 & n34886 ;
  assign n7722 = n1707 | n7721 ;
  assign n34887 = ~n7722 ;
  assign n7723 = n7706 & n34887 ;
  assign n7724 = n7495 | n7723 ;
  assign n34888 = ~n7708 ;
  assign n7725 = n34888 & n7724 ;
  assign n34889 = ~n7725 ;
  assign n7726 = n180 & n34889 ;
  assign n34890 = ~n7222 ;
  assign n7483 = n7041 & n34890 ;
  assign n7484 = n34672 & n7483 ;
  assign n7485 = n162 & n7484 ;
  assign n7486 = n7222 | n7231 ;
  assign n34891 = ~n7486 ;
  assign n7487 = n162 & n34891 ;
  assign n7488 = n7041 | n7487 ;
  assign n34892 = ~n7485 ;
  assign n7489 = n34892 & n7488 ;
  assign n7709 = n1487 | n7708 ;
  assign n34893 = ~n7709 ;
  assign n7727 = n34893 & n7724 ;
  assign n7728 = n7489 | n7727 ;
  assign n34894 = ~n7726 ;
  assign n7729 = n34894 & n7728 ;
  assign n34895 = ~n7729 ;
  assign n7730 = n181 & n34895 ;
  assign n7227 = n7034 & n34661 ;
  assign n34896 = ~n7233 ;
  assign n7477 = n7227 & n34896 ;
  assign n7478 = n162 & n7477 ;
  assign n7479 = n7233 | n7244 ;
  assign n34897 = ~n7479 ;
  assign n7480 = n162 & n34897 ;
  assign n7481 = n7034 | n7480 ;
  assign n34898 = ~n7478 ;
  assign n7482 = n34898 & n7481 ;
  assign n7738 = n34877 & n7719 ;
  assign n7739 = n7502 | n7738 ;
  assign n34899 = ~n7721 ;
  assign n7740 = n34899 & n7739 ;
  assign n34900 = ~n7740 ;
  assign n7741 = n179 & n34900 ;
  assign n7742 = n34887 & n7739 ;
  assign n7743 = n7495 | n7742 ;
  assign n34901 = ~n7741 ;
  assign n7744 = n34901 & n7743 ;
  assign n34902 = ~n7744 ;
  assign n7745 = n1487 & n34902 ;
  assign n7746 = n181 | n7745 ;
  assign n34903 = ~n7746 ;
  assign n7747 = n7728 & n34903 ;
  assign n7748 = n7482 | n7747 ;
  assign n34904 = ~n7730 ;
  assign n7749 = n34904 & n7748 ;
  assign n34905 = ~n7749 ;
  assign n7750 = n182 & n34905 ;
  assign n34906 = ~n7237 ;
  assign n7470 = n7028 & n34906 ;
  assign n7471 = n34688 & n7470 ;
  assign n7472 = n162 & n7471 ;
  assign n7473 = n7237 | n7246 ;
  assign n34907 = ~n7473 ;
  assign n7474 = n162 & n34907 ;
  assign n7475 = n7028 | n7474 ;
  assign n34908 = ~n7472 ;
  assign n7476 = n34908 & n7475 ;
  assign n7731 = n182 | n7730 ;
  assign n34909 = ~n7731 ;
  assign n7751 = n34909 & n7748 ;
  assign n7752 = n7476 | n7751 ;
  assign n34910 = ~n7750 ;
  assign n7753 = n34910 & n7752 ;
  assign n34911 = ~n7753 ;
  assign n7754 = n996 & n34911 ;
  assign n7242 = n7021 & n34677 ;
  assign n34912 = ~n7248 ;
  assign n7464 = n7242 & n34912 ;
  assign n7465 = n162 & n7464 ;
  assign n7466 = n7248 | n7259 ;
  assign n34913 = ~n7466 ;
  assign n7467 = n162 & n34913 ;
  assign n7468 = n7021 | n7467 ;
  assign n34914 = ~n7465 ;
  assign n7469 = n34914 & n7468 ;
  assign n7762 = n34893 & n7743 ;
  assign n7763 = n7489 | n7762 ;
  assign n34915 = ~n7745 ;
  assign n7764 = n34915 & n7763 ;
  assign n34916 = ~n7764 ;
  assign n7765 = n181 & n34916 ;
  assign n7766 = n34903 & n7763 ;
  assign n7767 = n7482 | n7766 ;
  assign n34917 = ~n7765 ;
  assign n7768 = n34917 & n7767 ;
  assign n34918 = ~n7768 ;
  assign n7769 = n182 & n34918 ;
  assign n7770 = n183 | n7769 ;
  assign n34919 = ~n7770 ;
  assign n7771 = n7752 & n34919 ;
  assign n7772 = n7469 | n7771 ;
  assign n34920 = ~n7754 ;
  assign n7773 = n34920 & n7772 ;
  assign n34921 = ~n7773 ;
  assign n7774 = n184 & n34921 ;
  assign n34922 = ~n7252 ;
  assign n7457 = n7015 & n34922 ;
  assign n7458 = n34704 & n7457 ;
  assign n7459 = n162 & n7458 ;
  assign n7460 = n7252 | n7261 ;
  assign n34923 = ~n7460 ;
  assign n7461 = n162 & n34923 ;
  assign n7462 = n7015 | n7461 ;
  assign n34924 = ~n7459 ;
  assign n7463 = n34924 & n7462 ;
  assign n7755 = n838 | n7754 ;
  assign n34925 = ~n7755 ;
  assign n7775 = n34925 & n7772 ;
  assign n7776 = n7463 | n7775 ;
  assign n34926 = ~n7774 ;
  assign n7777 = n34926 & n7776 ;
  assign n34927 = ~n7777 ;
  assign n7778 = n185 & n34927 ;
  assign n7257 = n7008 & n34693 ;
  assign n34928 = ~n7263 ;
  assign n7451 = n7257 & n34928 ;
  assign n7452 = n162 & n7451 ;
  assign n7453 = n7263 | n7274 ;
  assign n34929 = ~n7453 ;
  assign n7454 = n162 & n34929 ;
  assign n7455 = n7008 | n7454 ;
  assign n34930 = ~n7452 ;
  assign n7456 = n34930 & n7455 ;
  assign n7786 = n34909 & n7767 ;
  assign n7787 = n7476 | n7786 ;
  assign n34931 = ~n7769 ;
  assign n7788 = n34931 & n7787 ;
  assign n34932 = ~n7788 ;
  assign n7789 = n183 & n34932 ;
  assign n7790 = n34919 & n7787 ;
  assign n7791 = n7469 | n7790 ;
  assign n34933 = ~n7789 ;
  assign n7792 = n34933 & n7791 ;
  assign n34934 = ~n7792 ;
  assign n7793 = n838 & n34934 ;
  assign n7794 = n185 | n7793 ;
  assign n34935 = ~n7794 ;
  assign n7795 = n7776 & n34935 ;
  assign n7796 = n7456 | n7795 ;
  assign n34936 = ~n7778 ;
  assign n7797 = n34936 & n7796 ;
  assign n34937 = ~n7797 ;
  assign n7798 = n186 & n34937 ;
  assign n34938 = ~n7267 ;
  assign n7444 = n7002 & n34938 ;
  assign n7445 = n34720 & n7444 ;
  assign n7446 = n162 & n7445 ;
  assign n7447 = n7267 | n7276 ;
  assign n34939 = ~n7447 ;
  assign n7448 = n162 & n34939 ;
  assign n7449 = n7002 | n7448 ;
  assign n34940 = ~n7446 ;
  assign n7450 = n34940 & n7449 ;
  assign n7779 = n186 | n7778 ;
  assign n34941 = ~n7779 ;
  assign n7799 = n34941 & n7796 ;
  assign n7800 = n7450 | n7799 ;
  assign n34942 = ~n7798 ;
  assign n7801 = n34942 & n7800 ;
  assign n34943 = ~n7801 ;
  assign n7802 = n528 & n34943 ;
  assign n7272 = n6995 & n34709 ;
  assign n34944 = ~n7278 ;
  assign n7438 = n7272 & n34944 ;
  assign n7439 = n162 & n7438 ;
  assign n7440 = n7278 | n7289 ;
  assign n34945 = ~n7440 ;
  assign n7441 = n162 & n34945 ;
  assign n7442 = n6995 | n7441 ;
  assign n34946 = ~n7439 ;
  assign n7443 = n34946 & n7442 ;
  assign n7810 = n34925 & n7791 ;
  assign n7811 = n7463 | n7810 ;
  assign n34947 = ~n7793 ;
  assign n7812 = n34947 & n7811 ;
  assign n34948 = ~n7812 ;
  assign n7813 = n185 & n34948 ;
  assign n7814 = n34935 & n7811 ;
  assign n7815 = n7456 | n7814 ;
  assign n34949 = ~n7813 ;
  assign n7816 = n34949 & n7815 ;
  assign n34950 = ~n7816 ;
  assign n7817 = n186 & n34950 ;
  assign n7818 = n528 | n7817 ;
  assign n34951 = ~n7818 ;
  assign n7819 = n7800 & n34951 ;
  assign n7820 = n7443 | n7819 ;
  assign n34952 = ~n7802 ;
  assign n7821 = n34952 & n7820 ;
  assign n34953 = ~n7821 ;
  assign n7822 = n188 & n34953 ;
  assign n34954 = ~n7282 ;
  assign n7431 = n6989 & n34954 ;
  assign n7432 = n34726 & n7431 ;
  assign n7433 = n162 & n7432 ;
  assign n7434 = n7282 | n7291 ;
  assign n34955 = ~n7434 ;
  assign n7435 = n162 & n34955 ;
  assign n7436 = n6989 | n7435 ;
  assign n34956 = ~n7433 ;
  assign n7437 = n34956 & n7436 ;
  assign n7803 = n413 | n7802 ;
  assign n34957 = ~n7803 ;
  assign n7823 = n34957 & n7820 ;
  assign n7824 = n7437 | n7823 ;
  assign n34958 = ~n7822 ;
  assign n7825 = n34958 & n7824 ;
  assign n34959 = ~n7825 ;
  assign n7826 = n189 & n34959 ;
  assign n7287 = n6982 & n34741 ;
  assign n34960 = ~n7293 ;
  assign n7425 = n7287 & n34960 ;
  assign n7426 = n162 & n7425 ;
  assign n7427 = n7293 | n7304 ;
  assign n34961 = ~n7427 ;
  assign n7428 = n162 & n34961 ;
  assign n7429 = n6982 | n7428 ;
  assign n34962 = ~n7426 ;
  assign n7430 = n34962 & n7429 ;
  assign n7834 = n34941 & n7815 ;
  assign n7835 = n7450 | n7834 ;
  assign n34963 = ~n7817 ;
  assign n7836 = n34963 & n7835 ;
  assign n34964 = ~n7836 ;
  assign n7837 = n187 & n34964 ;
  assign n7838 = n34951 & n7835 ;
  assign n7839 = n7443 | n7838 ;
  assign n34965 = ~n7837 ;
  assign n7840 = n34965 & n7839 ;
  assign n34966 = ~n7840 ;
  assign n7841 = n413 & n34966 ;
  assign n7842 = n189 | n7841 ;
  assign n34967 = ~n7842 ;
  assign n7843 = n7824 & n34967 ;
  assign n7844 = n7430 | n7843 ;
  assign n34968 = ~n7826 ;
  assign n7845 = n34968 & n7844 ;
  assign n34969 = ~n7845 ;
  assign n7846 = n190 & n34969 ;
  assign n34970 = ~n7297 ;
  assign n7418 = n6976 & n34970 ;
  assign n7419 = n34730 & n7418 ;
  assign n7420 = n162 & n7419 ;
  assign n7421 = n7297 | n7306 ;
  assign n34971 = ~n7421 ;
  assign n7422 = n162 & n34971 ;
  assign n7423 = n6976 | n7422 ;
  assign n34972 = ~n7420 ;
  assign n7424 = n34972 & n7423 ;
  assign n7827 = n190 | n7826 ;
  assign n34973 = ~n7827 ;
  assign n7847 = n34973 & n7844 ;
  assign n7848 = n7424 | n7847 ;
  assign n34974 = ~n7846 ;
  assign n7849 = n34974 & n7848 ;
  assign n34975 = ~n7849 ;
  assign n7850 = n287 & n34975 ;
  assign n34976 = ~n7300 ;
  assign n7302 = n6969 & n34976 ;
  assign n34977 = ~n7310 ;
  assign n7412 = n7302 & n34977 ;
  assign n7413 = n162 & n7412 ;
  assign n7414 = n7309 | n7310 ;
  assign n34978 = ~n7414 ;
  assign n7415 = n162 & n34978 ;
  assign n7416 = n6969 | n7415 ;
  assign n34979 = ~n7413 ;
  assign n7417 = n34979 & n7416 ;
  assign n7858 = n34957 & n7839 ;
  assign n7859 = n7437 | n7858 ;
  assign n34980 = ~n7841 ;
  assign n7860 = n34980 & n7859 ;
  assign n34981 = ~n7860 ;
  assign n7861 = n189 & n34981 ;
  assign n7862 = n34967 & n7859 ;
  assign n7863 = n7430 | n7862 ;
  assign n34982 = ~n7861 ;
  assign n7864 = n34982 & n7863 ;
  assign n34983 = ~n7864 ;
  assign n7865 = n190 & n34983 ;
  assign n7866 = n287 | n7865 ;
  assign n34984 = ~n7866 ;
  assign n7867 = n7848 & n34984 ;
  assign n7870 = n7417 | n7867 ;
  assign n34985 = ~n7850 ;
  assign n7871 = n34985 & n7870 ;
  assign n7874 = n7399 | n7871 ;
  assign n7875 = n31336 & n7874 ;
  assign n7324 = n192 & n7323 ;
  assign n34986 = ~n6943 ;
  assign n7339 = n34986 & n162 ;
  assign n34987 = ~n7339 ;
  assign n7340 = n7320 & n34987 ;
  assign n34988 = ~n7340 ;
  assign n7341 = n7324 & n34988 ;
  assign n6923 = n6910 | n6922 ;
  assign n34989 = ~n6923 ;
  assign n6945 = n34989 & n6942 ;
  assign n6952 = n6945 & n34766 ;
  assign n7400 = n6952 & n34767 ;
  assign n7401 = n34768 & n7400 ;
  assign n7402 = n7341 | n7401 ;
  assign n7851 = n7347 & n34985 ;
  assign n7876 = n7851 & n7870 ;
  assign n7877 = n7402 | n7876 ;
  assign n161 = n7875 | n7877 ;
  assign n7852 = n7417 & n34985 ;
  assign n34990 = ~n7867 ;
  assign n7868 = n7852 & n34990 ;
  assign n7879 = n7868 & n161 ;
  assign n7869 = n7850 | n7867 ;
  assign n34991 = ~n7869 ;
  assign n7989 = n34991 & n161 ;
  assign n7990 = n7417 | n7989 ;
  assign n34992 = ~n7879 ;
  assign n7991 = n34992 & n7990 ;
  assign n7872 = n7347 | n7871 ;
  assign n34993 = ~n7872 ;
  assign n8017 = n34993 & n161 ;
  assign n8073 = n7876 | n8017 ;
  assign n8074 = n7991 | n8073 ;
  assign n17827 = x62 | x63 ;
  assign n18594 = x64 | n17827 ;
  assign n7930 = x64 & n161 ;
  assign n34994 = ~n7930 ;
  assign n7931 = n18594 & n34994 ;
  assign n34995 = ~n7931 ;
  assign n7932 = n162 & n34995 ;
  assign n6912 = n18594 & n34765 ;
  assign n6953 = n6912 & n34766 ;
  assign n7410 = n6953 & n34767 ;
  assign n7411 = n34768 & n7410 ;
  assign n7986 = n7411 & n34994 ;
  assign n34996 = ~n15623 ;
  assign n7899 = n34996 & n161 ;
  assign n34997 = ~x64 ;
  assign n7992 = n34997 & n161 ;
  assign n34998 = ~n7992 ;
  assign n7993 = x65 & n34998 ;
  assign n7994 = n7899 | n7993 ;
  assign n7995 = n7986 | n7994 ;
  assign n34999 = ~n7932 ;
  assign n7997 = n34999 & n7995 ;
  assign n35000 = ~n7997 ;
  assign n7998 = n6889 & n35000 ;
  assign n19398 = n34997 & n17827 ;
  assign n35001 = ~n161 ;
  assign n8004 = x64 & n35001 ;
  assign n8005 = n19398 | n8004 ;
  assign n35002 = ~n8005 ;
  assign n8006 = n162 & n35002 ;
  assign n8007 = n6889 | n8006 ;
  assign n35003 = ~n8007 ;
  assign n8008 = n7995 & n35003 ;
  assign n35004 = ~n7401 ;
  assign n7403 = n162 & n35004 ;
  assign n35005 = ~n7341 ;
  assign n7404 = n35005 & n7403 ;
  assign n35006 = ~n7876 ;
  assign n8018 = n7404 & n35006 ;
  assign n35007 = ~n7875 ;
  assign n8019 = n35007 & n8018 ;
  assign n8020 = n7899 | n8019 ;
  assign n8021 = x66 & n8020 ;
  assign n8022 = x66 | n8019 ;
  assign n8023 = n7899 | n8022 ;
  assign n35008 = ~n8021 ;
  assign n8024 = n35008 & n8023 ;
  assign n8025 = n8008 | n8024 ;
  assign n35009 = ~n7998 ;
  assign n8026 = n35009 & n8025 ;
  assign n35010 = ~n8026 ;
  assign n8027 = n6600 & n35010 ;
  assign n7354 = n7345 | n7352 ;
  assign n35011 = ~n7354 ;
  assign n7947 = n35011 & n161 ;
  assign n7948 = n7357 | n7947 ;
  assign n7360 = n35011 & n7357 ;
  assign n7962 = n7360 & n161 ;
  assign n35012 = ~n7962 ;
  assign n7963 = n7948 & n35012 ;
  assign n7999 = n6600 | n7998 ;
  assign n35013 = ~n7999 ;
  assign n8030 = n35013 & n8025 ;
  assign n8031 = n7963 | n8030 ;
  assign n35014 = ~n8027 ;
  assign n8032 = n35014 & n8031 ;
  assign n35015 = ~n8032 ;
  assign n8033 = n165 & n35015 ;
  assign n7365 = n7359 | n7364 ;
  assign n35016 = ~n7365 ;
  assign n7941 = n35016 & n161 ;
  assign n7942 = n7373 | n7941 ;
  assign n35017 = ~n7359 ;
  assign n7386 = n35017 & n7373 ;
  assign n7387 = n34770 & n7386 ;
  assign n8012 = n7387 & n161 ;
  assign n35018 = ~n8012 ;
  assign n8013 = n7942 & n35018 ;
  assign n8028 = n165 | n8027 ;
  assign n35019 = ~n8028 ;
  assign n8034 = n35019 & n8031 ;
  assign n8038 = n8013 | n8034 ;
  assign n35020 = ~n8033 ;
  assign n8039 = n35020 & n8038 ;
  assign n35021 = ~n8039 ;
  assign n8040 = n166 & n35021 ;
  assign n7385 = n7376 | n7379 ;
  assign n35022 = ~n7385 ;
  assign n7949 = n35022 & n161 ;
  assign n7950 = n7349 | n7949 ;
  assign n7378 = n7349 & n34775 ;
  assign n35023 = ~n7379 ;
  assign n7384 = n7378 & n35023 ;
  assign n8002 = n7384 & n161 ;
  assign n35024 = ~n8002 ;
  assign n8003 = n7950 & n35024 ;
  assign n8000 = n163 & n35000 ;
  assign n7933 = n163 | n7932 ;
  assign n35025 = ~n7933 ;
  assign n7996 = n35025 & n7995 ;
  assign n8047 = n7996 | n8024 ;
  assign n35026 = ~n8000 ;
  assign n8048 = n35026 & n8047 ;
  assign n35027 = ~n8048 ;
  assign n8049 = n164 & n35027 ;
  assign n8050 = n35013 & n8047 ;
  assign n8051 = n7963 | n8050 ;
  assign n35028 = ~n8049 ;
  assign n8052 = n35028 & n8051 ;
  assign n35029 = ~n8052 ;
  assign n8053 = n165 & n35029 ;
  assign n8054 = n166 | n8053 ;
  assign n35030 = ~n8054 ;
  assign n8055 = n8038 & n35030 ;
  assign n8056 = n8003 | n8055 ;
  assign n35031 = ~n8040 ;
  assign n8057 = n35031 & n8056 ;
  assign n35032 = ~n8057 ;
  assign n8058 = n167 & n35032 ;
  assign n8041 = n5352 | n8040 ;
  assign n35033 = ~n8041 ;
  assign n8059 = n35033 & n8056 ;
  assign n35034 = ~n7383 ;
  assign n7593 = n35034 & n7573 ;
  assign n7594 = n34781 & n7593 ;
  assign n7934 = n7594 & n161 ;
  assign n7396 = n7383 | n7394 ;
  assign n35035 = ~n7396 ;
  assign n7937 = n35035 & n161 ;
  assign n8091 = n7573 | n7937 ;
  assign n35036 = ~n7934 ;
  assign n8092 = n35036 & n8091 ;
  assign n8093 = n8059 | n8092 ;
  assign n35037 = ~n8058 ;
  assign n8094 = n35037 & n8093 ;
  assign n35038 = ~n8094 ;
  assign n8095 = n4934 & n35038 ;
  assign n7578 = n7567 & n34792 ;
  assign n35039 = ~n7579 ;
  assign n7591 = n7578 & n35039 ;
  assign n7918 = n7591 & n161 ;
  assign n7592 = n7576 | n7579 ;
  assign n35040 = ~n7592 ;
  assign n7951 = n35040 & n161 ;
  assign n7952 = n7567 | n7951 ;
  assign n35041 = ~n7918 ;
  assign n7953 = n35041 & n7952 ;
  assign n8063 = n35019 & n8051 ;
  assign n8064 = n8013 | n8063 ;
  assign n35042 = ~n8053 ;
  assign n8065 = n35042 & n8064 ;
  assign n35043 = ~n8065 ;
  assign n8066 = n166 & n35043 ;
  assign n8067 = n35030 & n8064 ;
  assign n8068 = n8003 | n8067 ;
  assign n35044 = ~n8066 ;
  assign n8069 = n35044 & n8068 ;
  assign n35045 = ~n8069 ;
  assign n8070 = n5352 & n35045 ;
  assign n8071 = n4934 | n8070 ;
  assign n35046 = ~n8071 ;
  assign n8098 = n35046 & n8093 ;
  assign n8099 = n7953 | n8098 ;
  assign n35047 = ~n8095 ;
  assign n8100 = n35047 & n8099 ;
  assign n35048 = ~n8100 ;
  assign n8101 = n169 & n35048 ;
  assign n7617 = n7583 | n7601 ;
  assign n35049 = ~n7617 ;
  assign n7928 = n35049 & n161 ;
  assign n7929 = n7561 | n7928 ;
  assign n35050 = ~n7583 ;
  assign n7589 = n7561 & n35050 ;
  assign n7590 = n34798 & n7589 ;
  assign n7958 = n7590 & n161 ;
  assign n35051 = ~n7958 ;
  assign n7959 = n7929 & n35051 ;
  assign n8096 = n169 | n8095 ;
  assign n35052 = ~n8096 ;
  assign n8102 = n35052 & n8099 ;
  assign n8103 = n7959 | n8102 ;
  assign n35053 = ~n8101 ;
  assign n8104 = n35053 & n8103 ;
  assign n35054 = ~n8104 ;
  assign n8105 = n170 & n35054 ;
  assign n7588 = n7554 & n34808 ;
  assign n35055 = ~n7603 ;
  assign n7615 = n7588 & n35055 ;
  assign n7886 = n7615 & n161 ;
  assign n7616 = n7586 | n7603 ;
  assign n35056 = ~n7616 ;
  assign n7977 = n35056 & n161 ;
  assign n7978 = n7554 | n7977 ;
  assign n35057 = ~n7886 ;
  assign n7979 = n35057 & n7978 ;
  assign n8072 = n35033 & n8068 ;
  assign n8115 = n8072 | n8092 ;
  assign n35058 = ~n8070 ;
  assign n8116 = n35058 & n8115 ;
  assign n35059 = ~n8116 ;
  assign n8117 = n168 & n35059 ;
  assign n8118 = n35046 & n8115 ;
  assign n8119 = n7953 | n8118 ;
  assign n35060 = ~n8117 ;
  assign n8120 = n35060 & n8119 ;
  assign n35061 = ~n8120 ;
  assign n8121 = n169 & n35061 ;
  assign n8122 = n170 | n8121 ;
  assign n35062 = ~n8122 ;
  assign n8123 = n8103 & n35062 ;
  assign n8124 = n7979 | n8123 ;
  assign n35063 = ~n8105 ;
  assign n8125 = n35063 & n8124 ;
  assign n35064 = ~n8125 ;
  assign n8126 = n171 & n35064 ;
  assign n35065 = ~n7607 ;
  assign n7613 = n7548 & n35065 ;
  assign n7614 = n34814 & n7613 ;
  assign n7912 = n7614 & n161 ;
  assign n7641 = n7607 | n7625 ;
  assign n35066 = ~n7641 ;
  assign n7964 = n35066 & n161 ;
  assign n7965 = n7548 | n7964 ;
  assign n35067 = ~n7912 ;
  assign n7966 = n35067 & n7965 ;
  assign n8106 = n3940 | n8105 ;
  assign n35068 = ~n8106 ;
  assign n8127 = n35068 & n8124 ;
  assign n8128 = n7966 | n8127 ;
  assign n35069 = ~n8126 ;
  assign n8129 = n35069 & n8128 ;
  assign n35070 = ~n8129 ;
  assign n8130 = n3631 & n35070 ;
  assign n7640 = n7610 | n7627 ;
  assign n35071 = ~n7640 ;
  assign n7967 = n35071 & n161 ;
  assign n7968 = n7333 | n7967 ;
  assign n7611 = n7333 & n34824 ;
  assign n35072 = ~n7627 ;
  assign n7639 = n7611 & n35072 ;
  assign n7969 = n7639 & n161 ;
  assign n35073 = ~n7969 ;
  assign n7970 = n7968 & n35073 ;
  assign n8138 = n35052 & n8119 ;
  assign n8139 = n7959 | n8138 ;
  assign n35074 = ~n8121 ;
  assign n8140 = n35074 & n8139 ;
  assign n35075 = ~n8140 ;
  assign n8141 = n170 & n35075 ;
  assign n8142 = n35062 & n8139 ;
  assign n8143 = n7979 | n8142 ;
  assign n35076 = ~n8141 ;
  assign n8144 = n35076 & n8143 ;
  assign n35077 = ~n8144 ;
  assign n8145 = n3940 & n35077 ;
  assign n8146 = n3631 | n8145 ;
  assign n35078 = ~n8146 ;
  assign n8147 = n8128 & n35078 ;
  assign n8148 = n7970 | n8147 ;
  assign n35079 = ~n8130 ;
  assign n8149 = n35079 & n8148 ;
  assign n35080 = ~n8149 ;
  assign n8150 = n173 & n35080 ;
  assign n35081 = ~n7631 ;
  assign n7637 = n7541 & n35081 ;
  assign n7638 = n34830 & n7637 ;
  assign n7945 = n7638 & n161 ;
  assign n7665 = n7631 | n7649 ;
  assign n35082 = ~n7665 ;
  assign n7971 = n35082 & n161 ;
  assign n7972 = n7541 | n7971 ;
  assign n35083 = ~n7945 ;
  assign n7973 = n35083 & n7972 ;
  assign n8132 = n173 | n8130 ;
  assign n35084 = ~n8132 ;
  assign n8151 = n35084 & n8148 ;
  assign n8152 = n7973 | n8151 ;
  assign n35085 = ~n8150 ;
  assign n8153 = n35085 & n8152 ;
  assign n35086 = ~n8153 ;
  assign n8154 = n174 & n35086 ;
  assign n7636 = n7534 & n34840 ;
  assign n35087 = ~n7651 ;
  assign n7664 = n7636 & n35087 ;
  assign n7946 = n7664 & n161 ;
  assign n7663 = n7634 | n7651 ;
  assign n35088 = ~n7663 ;
  assign n7974 = n35088 & n161 ;
  assign n7975 = n7534 | n7974 ;
  assign n35089 = ~n7946 ;
  assign n7976 = n35089 & n7975 ;
  assign n8162 = n35068 & n8143 ;
  assign n8163 = n7966 | n8162 ;
  assign n35090 = ~n8145 ;
  assign n8164 = n35090 & n8163 ;
  assign n35091 = ~n8164 ;
  assign n8165 = n172 & n35091 ;
  assign n8166 = n35078 & n8163 ;
  assign n8167 = n7970 | n8166 ;
  assign n35092 = ~n8165 ;
  assign n8168 = n35092 & n8167 ;
  assign n35093 = ~n8168 ;
  assign n8169 = n173 & n35093 ;
  assign n8170 = n174 | n8169 ;
  assign n35094 = ~n8170 ;
  assign n8171 = n8152 & n35094 ;
  assign n8172 = n7976 | n8171 ;
  assign n35095 = ~n8154 ;
  assign n8173 = n35095 & n8172 ;
  assign n35096 = ~n8173 ;
  assign n8174 = n175 & n35096 ;
  assign n7689 = n7655 | n7673 ;
  assign n35097 = ~n7689 ;
  assign n7980 = n35097 & n161 ;
  assign n7981 = n7528 | n7980 ;
  assign n35098 = ~n7655 ;
  assign n7661 = n7528 & n35098 ;
  assign n7662 = n34846 & n7661 ;
  assign n7982 = n7662 & n161 ;
  assign n35099 = ~n7982 ;
  assign n7983 = n7981 & n35099 ;
  assign n8155 = n2753 | n8154 ;
  assign n35100 = ~n8155 ;
  assign n8175 = n35100 & n8172 ;
  assign n8179 = n7983 | n8175 ;
  assign n35101 = ~n8174 ;
  assign n8180 = n35101 & n8179 ;
  assign n35102 = ~n8180 ;
  assign n8181 = n2431 & n35102 ;
  assign n7688 = n7658 | n7675 ;
  assign n35103 = ~n7688 ;
  assign n7984 = n35103 & n161 ;
  assign n7985 = n7521 | n7984 ;
  assign n7660 = n7521 & n34856 ;
  assign n35104 = ~n7675 ;
  assign n7687 = n7660 & n35104 ;
  assign n7987 = n7687 & n161 ;
  assign n35105 = ~n7987 ;
  assign n7988 = n7985 & n35105 ;
  assign n8186 = n35084 & n8167 ;
  assign n8187 = n7973 | n8186 ;
  assign n35106 = ~n8169 ;
  assign n8188 = n35106 & n8187 ;
  assign n35107 = ~n8188 ;
  assign n8189 = n174 & n35107 ;
  assign n8190 = n35094 & n8187 ;
  assign n8191 = n7976 | n8190 ;
  assign n35108 = ~n8189 ;
  assign n8192 = n35108 & n8191 ;
  assign n35109 = ~n8192 ;
  assign n8193 = n2753 & n35109 ;
  assign n8194 = n2431 | n8193 ;
  assign n35110 = ~n8194 ;
  assign n8195 = n8179 & n35110 ;
  assign n8196 = n7988 | n8195 ;
  assign n35111 = ~n8181 ;
  assign n8197 = n35111 & n8196 ;
  assign n35112 = ~n8197 ;
  assign n8198 = n177 & n35112 ;
  assign n7713 = n7679 | n7697 ;
  assign n35113 = ~n7713 ;
  assign n7890 = n35113 & n161 ;
  assign n7891 = n7515 | n7890 ;
  assign n35114 = ~n7679 ;
  assign n7685 = n7515 & n35114 ;
  assign n7686 = n34862 & n7685 ;
  assign n7922 = n7686 & n161 ;
  assign n35115 = ~n7922 ;
  assign n7923 = n7891 & n35115 ;
  assign n8182 = n177 | n8181 ;
  assign n35116 = ~n8182 ;
  assign n8199 = n35116 & n8196 ;
  assign n8200 = n7923 | n8199 ;
  assign n35117 = ~n8198 ;
  assign n8201 = n35117 & n8200 ;
  assign n35118 = ~n8201 ;
  assign n8202 = n178 & n35118 ;
  assign n7684 = n7508 & n34872 ;
  assign n35119 = ~n7699 ;
  assign n7711 = n7684 & n35119 ;
  assign n7917 = n7711 & n161 ;
  assign n7712 = n7682 | n7699 ;
  assign n35120 = ~n7712 ;
  assign n7919 = n35120 & n161 ;
  assign n7920 = n7508 | n7919 ;
  assign n35121 = ~n7917 ;
  assign n7921 = n35121 & n7920 ;
  assign n8210 = n35100 & n8191 ;
  assign n8211 = n7983 | n8210 ;
  assign n35122 = ~n8193 ;
  assign n8212 = n35122 & n8211 ;
  assign n35123 = ~n8212 ;
  assign n8213 = n176 & n35123 ;
  assign n8214 = n35110 & n8211 ;
  assign n8215 = n7988 | n8214 ;
  assign n35124 = ~n8213 ;
  assign n8216 = n35124 & n8215 ;
  assign n35125 = ~n8216 ;
  assign n8217 = n177 & n35125 ;
  assign n8218 = n178 | n8217 ;
  assign n35126 = ~n8218 ;
  assign n8219 = n8200 & n35126 ;
  assign n8220 = n7921 | n8219 ;
  assign n35127 = ~n8202 ;
  assign n8221 = n35127 & n8220 ;
  assign n35128 = ~n8221 ;
  assign n8222 = n179 & n35128 ;
  assign n35129 = ~n7703 ;
  assign n7704 = n7502 & n35129 ;
  assign n7705 = n34878 & n7704 ;
  assign n7913 = n7705 & n161 ;
  assign n7737 = n7703 | n7721 ;
  assign n35130 = ~n7737 ;
  assign n7914 = n35130 & n161 ;
  assign n7915 = n7502 | n7914 ;
  assign n35131 = ~n7913 ;
  assign n7916 = n35131 & n7915 ;
  assign n8203 = n1707 | n8202 ;
  assign n35132 = ~n8203 ;
  assign n8223 = n35132 & n8220 ;
  assign n8224 = n7916 | n8223 ;
  assign n35133 = ~n8222 ;
  assign n8225 = n35133 & n8224 ;
  assign n35134 = ~n8225 ;
  assign n8226 = n1487 & n35134 ;
  assign n7710 = n7495 & n34888 ;
  assign n35135 = ~n7723 ;
  assign n7735 = n7710 & n35135 ;
  assign n7906 = n7735 & n161 ;
  assign n7736 = n7708 | n7723 ;
  assign n35136 = ~n7736 ;
  assign n7909 = n35136 & n161 ;
  assign n7910 = n7495 | n7909 ;
  assign n35137 = ~n7906 ;
  assign n7911 = n35137 & n7910 ;
  assign n8234 = n35116 & n8215 ;
  assign n8235 = n7923 | n8234 ;
  assign n35138 = ~n8217 ;
  assign n8236 = n35138 & n8235 ;
  assign n35139 = ~n8236 ;
  assign n8237 = n178 & n35139 ;
  assign n8238 = n35126 & n8235 ;
  assign n8239 = n7921 | n8238 ;
  assign n35140 = ~n8237 ;
  assign n8240 = n35140 & n8239 ;
  assign n35141 = ~n8240 ;
  assign n8241 = n1707 & n35141 ;
  assign n8242 = n1487 | n8241 ;
  assign n35142 = ~n8242 ;
  assign n8243 = n8224 & n35142 ;
  assign n8244 = n7911 | n8243 ;
  assign n35143 = ~n8226 ;
  assign n8245 = n35143 & n8244 ;
  assign n35144 = ~n8245 ;
  assign n8246 = n181 & n35144 ;
  assign n7761 = n7727 | n7745 ;
  assign n35145 = ~n7761 ;
  assign n7924 = n35145 & n161 ;
  assign n7925 = n7489 | n7924 ;
  assign n35146 = ~n7727 ;
  assign n7733 = n7489 & n35146 ;
  assign n7734 = n34894 & n7733 ;
  assign n7954 = n7734 & n161 ;
  assign n35147 = ~n7954 ;
  assign n7955 = n7925 & n35147 ;
  assign n8227 = n181 | n8226 ;
  assign n35148 = ~n8227 ;
  assign n8247 = n35148 & n8244 ;
  assign n8248 = n7955 | n8247 ;
  assign n35149 = ~n8246 ;
  assign n8249 = n35149 & n8248 ;
  assign n35150 = ~n8249 ;
  assign n8250 = n182 & n35150 ;
  assign n7732 = n7482 & n34904 ;
  assign n35151 = ~n7747 ;
  assign n7759 = n7732 & n35151 ;
  assign n7894 = n7759 & n161 ;
  assign n7760 = n7730 | n7747 ;
  assign n35152 = ~n7760 ;
  assign n7938 = n35152 & n161 ;
  assign n7939 = n7482 | n7938 ;
  assign n35153 = ~n7894 ;
  assign n7940 = n35153 & n7939 ;
  assign n8258 = n35132 & n8239 ;
  assign n8259 = n7916 | n8258 ;
  assign n35154 = ~n8241 ;
  assign n8260 = n35154 & n8259 ;
  assign n35155 = ~n8260 ;
  assign n8261 = n180 & n35155 ;
  assign n8262 = n35142 & n8259 ;
  assign n8263 = n7911 | n8262 ;
  assign n35156 = ~n8261 ;
  assign n8264 = n35156 & n8263 ;
  assign n35157 = ~n8264 ;
  assign n8265 = n181 & n35157 ;
  assign n8266 = n182 | n8265 ;
  assign n35158 = ~n8266 ;
  assign n8267 = n8248 & n35158 ;
  assign n8268 = n7940 | n8267 ;
  assign n35159 = ~n8250 ;
  assign n8269 = n35159 & n8268 ;
  assign n35160 = ~n8269 ;
  assign n8270 = n183 & n35160 ;
  assign n7785 = n7751 | n7769 ;
  assign n35161 = ~n7785 ;
  assign n7907 = n35161 & n161 ;
  assign n7908 = n7476 | n7907 ;
  assign n35162 = ~n7751 ;
  assign n7757 = n7476 & n35162 ;
  assign n7758 = n34910 & n7757 ;
  assign n7935 = n7758 & n161 ;
  assign n35163 = ~n7935 ;
  assign n7936 = n7908 & n35163 ;
  assign n8251 = n183 | n8250 ;
  assign n35164 = ~n8251 ;
  assign n8271 = n35164 & n8268 ;
  assign n8272 = n7936 | n8271 ;
  assign n35165 = ~n8270 ;
  assign n8273 = n35165 & n8272 ;
  assign n35166 = ~n8273 ;
  assign n8274 = n838 & n35166 ;
  assign n7756 = n7469 & n34920 ;
  assign n35167 = ~n7771 ;
  assign n7783 = n7756 & n35167 ;
  assign n7881 = n7783 & n161 ;
  assign n7784 = n7754 | n7771 ;
  assign n35168 = ~n7784 ;
  assign n7900 = n35168 & n161 ;
  assign n7901 = n7469 | n7900 ;
  assign n35169 = ~n7881 ;
  assign n7902 = n35169 & n7901 ;
  assign n8282 = n35148 & n8263 ;
  assign n8283 = n7955 | n8282 ;
  assign n35170 = ~n8265 ;
  assign n8284 = n35170 & n8283 ;
  assign n35171 = ~n8284 ;
  assign n8285 = n182 & n35171 ;
  assign n8286 = n35158 & n8283 ;
  assign n8287 = n7940 | n8286 ;
  assign n35172 = ~n8285 ;
  assign n8288 = n35172 & n8287 ;
  assign n35173 = ~n8288 ;
  assign n8289 = n996 & n35173 ;
  assign n8290 = n838 | n8289 ;
  assign n35174 = ~n8290 ;
  assign n8291 = n8272 & n35174 ;
  assign n8292 = n7902 | n8291 ;
  assign n35175 = ~n8274 ;
  assign n8293 = n35175 & n8292 ;
  assign n35176 = ~n8293 ;
  assign n8294 = n185 & n35176 ;
  assign n35177 = ~n7775 ;
  assign n7781 = n7463 & n35177 ;
  assign n7782 = n34926 & n7781 ;
  assign n7895 = n7782 & n161 ;
  assign n7809 = n7775 | n7793 ;
  assign n35178 = ~n7809 ;
  assign n7903 = n35178 & n161 ;
  assign n7904 = n7463 | n7903 ;
  assign n35179 = ~n7895 ;
  assign n7905 = n35179 & n7904 ;
  assign n8275 = n185 | n8274 ;
  assign n35180 = ~n8275 ;
  assign n8295 = n35180 & n8292 ;
  assign n8296 = n7905 | n8295 ;
  assign n35181 = ~n8294 ;
  assign n8297 = n35181 & n8296 ;
  assign n35182 = ~n8297 ;
  assign n8298 = n186 & n35182 ;
  assign n7808 = n7778 | n7795 ;
  assign n35183 = ~n7808 ;
  assign n7892 = n35183 & n161 ;
  assign n7893 = n7456 | n7892 ;
  assign n7780 = n7456 & n34936 ;
  assign n35184 = ~n7795 ;
  assign n7807 = n7780 & n35184 ;
  assign n7956 = n7807 & n161 ;
  assign n35185 = ~n7956 ;
  assign n7957 = n7893 & n35185 ;
  assign n8306 = n35164 & n8287 ;
  assign n8307 = n7936 | n8306 ;
  assign n35186 = ~n8289 ;
  assign n8308 = n35186 & n8307 ;
  assign n35187 = ~n8308 ;
  assign n8309 = n184 & n35187 ;
  assign n8310 = n35174 & n8307 ;
  assign n8311 = n7902 | n8310 ;
  assign n35188 = ~n8309 ;
  assign n8312 = n35188 & n8311 ;
  assign n35189 = ~n8312 ;
  assign n8313 = n185 & n35189 ;
  assign n8314 = n186 | n8313 ;
  assign n35190 = ~n8314 ;
  assign n8315 = n8296 & n35190 ;
  assign n8316 = n7957 | n8315 ;
  assign n35191 = ~n8298 ;
  assign n8317 = n35191 & n8316 ;
  assign n35192 = ~n8317 ;
  assign n8318 = n187 & n35192 ;
  assign n35193 = ~n7799 ;
  assign n7805 = n7450 & n35193 ;
  assign n7806 = n34942 & n7805 ;
  assign n7887 = n7806 & n161 ;
  assign n7833 = n7799 | n7817 ;
  assign n35194 = ~n7833 ;
  assign n7896 = n35194 & n161 ;
  assign n7897 = n7450 | n7896 ;
  assign n35195 = ~n7887 ;
  assign n7898 = n35195 & n7897 ;
  assign n8299 = n528 | n8298 ;
  assign n35196 = ~n8299 ;
  assign n8319 = n35196 & n8316 ;
  assign n8320 = n7898 | n8319 ;
  assign n35197 = ~n8318 ;
  assign n8321 = n35197 & n8320 ;
  assign n35198 = ~n8321 ;
  assign n8322 = n413 & n35198 ;
  assign n7832 = n7802 | n7819 ;
  assign n35199 = ~n7832 ;
  assign n7888 = n35199 & n161 ;
  assign n7889 = n7443 | n7888 ;
  assign n7804 = n7443 & n34952 ;
  assign n35200 = ~n7819 ;
  assign n7831 = n7804 & n35200 ;
  assign n7960 = n7831 & n161 ;
  assign n35201 = ~n7960 ;
  assign n7961 = n7889 & n35201 ;
  assign n8330 = n35180 & n8311 ;
  assign n8331 = n7905 | n8330 ;
  assign n35202 = ~n8313 ;
  assign n8332 = n35202 & n8331 ;
  assign n35203 = ~n8332 ;
  assign n8333 = n186 & n35203 ;
  assign n8334 = n35190 & n8331 ;
  assign n8335 = n7957 | n8334 ;
  assign n35204 = ~n8333 ;
  assign n8336 = n35204 & n8335 ;
  assign n35205 = ~n8336 ;
  assign n8337 = n528 & n35205 ;
  assign n8338 = n413 | n8337 ;
  assign n35206 = ~n8338 ;
  assign n8339 = n8320 & n35206 ;
  assign n8340 = n7961 | n8339 ;
  assign n35207 = ~n8322 ;
  assign n8341 = n35207 & n8340 ;
  assign n35208 = ~n8341 ;
  assign n8342 = n189 & n35208 ;
  assign n7857 = n7823 | n7841 ;
  assign n35209 = ~n7857 ;
  assign n7884 = n35209 & n161 ;
  assign n7885 = n7437 | n7884 ;
  assign n35210 = ~n7823 ;
  assign n7829 = n7437 & n35210 ;
  assign n7830 = n34958 & n7829 ;
  assign n7926 = n7830 & n161 ;
  assign n35211 = ~n7926 ;
  assign n7927 = n7885 & n35211 ;
  assign n8323 = n189 | n8322 ;
  assign n35212 = ~n8323 ;
  assign n8343 = n35212 & n8340 ;
  assign n8344 = n7927 | n8343 ;
  assign n35213 = ~n8342 ;
  assign n8345 = n35213 & n8344 ;
  assign n35214 = ~n8345 ;
  assign n8346 = n190 & n35214 ;
  assign n7856 = n7826 | n7843 ;
  assign n35215 = ~n7856 ;
  assign n7882 = n35215 & n161 ;
  assign n7883 = n7430 | n7882 ;
  assign n7828 = n7430 & n34968 ;
  assign n35216 = ~n7843 ;
  assign n7855 = n7828 & n35216 ;
  assign n7943 = n7855 & n161 ;
  assign n35217 = ~n7943 ;
  assign n7944 = n7883 & n35217 ;
  assign n8352 = n35196 & n8335 ;
  assign n8353 = n7898 | n8352 ;
  assign n35218 = ~n8337 ;
  assign n8354 = n35218 & n8353 ;
  assign n35219 = ~n8354 ;
  assign n8355 = n188 & n35219 ;
  assign n8356 = n35206 & n8353 ;
  assign n8357 = n7961 | n8356 ;
  assign n35220 = ~n8355 ;
  assign n8358 = n35220 & n8357 ;
  assign n35221 = ~n8358 ;
  assign n8359 = n189 & n35221 ;
  assign n8360 = n190 | n8359 ;
  assign n35222 = ~n8360 ;
  assign n8361 = n8344 & n35222 ;
  assign n8362 = n7944 | n8361 ;
  assign n35223 = ~n8346 ;
  assign n8367 = n35223 & n8362 ;
  assign n35224 = ~n8367 ;
  assign n8368 = n191 & n35224 ;
  assign n35225 = ~n7847 ;
  assign n7853 = n7424 & n35225 ;
  assign n7854 = n34974 & n7853 ;
  assign n7880 = n7854 & n161 ;
  assign n8087 = n7847 | n7865 ;
  assign n35226 = ~n8087 ;
  assign n8088 = n161 & n35226 ;
  assign n8089 = n7424 | n8088 ;
  assign n35227 = ~n7880 ;
  assign n8090 = n35227 & n8089 ;
  assign n8348 = n191 | n8346 ;
  assign n35228 = ~n8348 ;
  assign n8378 = n35228 & n8362 ;
  assign n8379 = n8090 | n8378 ;
  assign n35229 = ~n8368 ;
  assign n8380 = n35229 & n8379 ;
  assign n8381 = n8074 | n8380 ;
  assign n8382 = n31336 & n8381 ;
  assign n7873 = n192 & n7872 ;
  assign n35230 = ~n7347 ;
  assign n8014 = n35230 & n161 ;
  assign n35231 = ~n8014 ;
  assign n8015 = n7871 & n35231 ;
  assign n35232 = ~n8015 ;
  assign n8016 = n7873 & n35232 ;
  assign n7405 = n7346 | n7401 ;
  assign n35233 = ~n7405 ;
  assign n7406 = n7329 & n35233 ;
  assign n7407 = n35005 & n7406 ;
  assign n8075 = n7407 & n35006 ;
  assign n8076 = n35007 & n8075 ;
  assign n8077 = n8016 | n8076 ;
  assign n8369 = n7991 & n35229 ;
  assign n8388 = n8369 & n8379 ;
  assign n8389 = n8077 | n8388 ;
  assign n160 = n8382 | n8389 ;
  assign n8349 = n287 | n8346 ;
  assign n35234 = ~n8349 ;
  assign n8363 = n35234 & n8362 ;
  assign n8364 = n8090 | n8363 ;
  assign n8370 = n8364 & n8369 ;
  assign n8375 = n8364 & n35229 ;
  assign n8376 = n7991 | n8375 ;
  assign n35235 = ~n8376 ;
  assign n8463 = n35235 & n160 ;
  assign n8464 = n8370 | n8463 ;
  assign n35236 = ~n8378 ;
  assign n8610 = n8090 & n35236 ;
  assign n8611 = n35229 & n8610 ;
  assign n8612 = n160 & n8611 ;
  assign n8614 = n8368 | n8378 ;
  assign n35237 = ~n8614 ;
  assign n8615 = n160 & n35237 ;
  assign n8616 = n8090 | n8615 ;
  assign n35238 = ~n8612 ;
  assign n8617 = n35238 & n8616 ;
  assign n8618 = n8464 | n8617 ;
  assign n20170 = x60 | x61 ;
  assign n20991 = x62 | n20170 ;
  assign n8402 = x62 & n160 ;
  assign n35239 = ~n8402 ;
  assign n8403 = n20991 & n35239 ;
  assign n35240 = ~n8403 ;
  assign n8404 = n161 & n35240 ;
  assign n8405 = n162 | n8404 ;
  assign n7408 = n20991 & n35004 ;
  assign n7409 = n35005 & n7408 ;
  assign n8085 = n7409 & n35006 ;
  assign n8086 = n35007 & n8085 ;
  assign n8415 = n8086 & n35239 ;
  assign n35241 = ~n17827 ;
  assign n8412 = n35241 & n160 ;
  assign n35242 = ~x62 ;
  assign n8472 = n35242 & n160 ;
  assign n35243 = ~n8472 ;
  assign n8473 = x63 & n35243 ;
  assign n8476 = n8412 | n8473 ;
  assign n8477 = n8415 | n8476 ;
  assign n35244 = ~n8405 ;
  assign n8478 = n35244 & n8477 ;
  assign n35245 = ~n8076 ;
  assign n8078 = n161 & n35245 ;
  assign n35246 = ~n8016 ;
  assign n8079 = n35246 & n8078 ;
  assign n35247 = ~n8370 ;
  assign n8372 = n8079 & n35247 ;
  assign n35248 = ~n8382 ;
  assign n8383 = n8372 & n35248 ;
  assign n8384 = x64 | n8383 ;
  assign n8413 = n8384 | n8412 ;
  assign n8479 = n8383 | n8412 ;
  assign n8480 = x64 & n8479 ;
  assign n35249 = ~n8480 ;
  assign n8485 = n8413 & n35249 ;
  assign n8486 = n8478 | n8485 ;
  assign n21824 = n35242 & n20170 ;
  assign n8371 = n8077 | n8370 ;
  assign n8532 = n8074 | n8375 ;
  assign n8533 = n31336 & n8532 ;
  assign n8534 = n8371 | n8533 ;
  assign n35250 = ~n8534 ;
  assign n8537 = x62 & n35250 ;
  assign n8538 = n21824 | n8537 ;
  assign n35251 = ~n8538 ;
  assign n8539 = n161 & n35251 ;
  assign n35252 = ~n8539 ;
  assign n8540 = n8477 & n35252 ;
  assign n35253 = ~n8540 ;
  assign n8541 = n162 & n35253 ;
  assign n35254 = ~n8541 ;
  assign n8542 = n8486 & n35254 ;
  assign n35255 = ~n8542 ;
  assign n8564 = n163 & n35255 ;
  assign n8011 = n7986 | n8006 ;
  assign n35256 = ~n8011 ;
  assign n8393 = n35256 & n160 ;
  assign n8394 = n7994 | n8393 ;
  assign n35257 = ~n7986 ;
  assign n8001 = n35257 & n7994 ;
  assign n35258 = ~n8006 ;
  assign n8010 = n8001 & n35258 ;
  assign n8474 = n8010 & n160 ;
  assign n35259 = ~n8474 ;
  assign n8475 = n8394 & n35259 ;
  assign n8565 = n163 | n8541 ;
  assign n35260 = ~n8565 ;
  assign n8566 = n8486 & n35260 ;
  assign n8567 = n8475 | n8566 ;
  assign n35261 = ~n8564 ;
  assign n8568 = n35261 & n8567 ;
  assign n35262 = ~n8568 ;
  assign n8569 = n164 & n35262 ;
  assign n8009 = n8000 | n8008 ;
  assign n35263 = ~n8009 ;
  assign n8468 = n35263 & n160 ;
  assign n8469 = n8024 | n8468 ;
  assign n35264 = ~n8008 ;
  assign n8045 = n35264 & n8024 ;
  assign n8046 = n35026 & n8045 ;
  assign n8494 = n8046 & n160 ;
  assign n35265 = ~n8494 ;
  assign n8495 = n8469 & n35265 ;
  assign n8543 = n6889 & n35255 ;
  assign n8550 = n6600 | n8543 ;
  assign n35266 = ~n8550 ;
  assign n8570 = n35266 & n8567 ;
  assign n8571 = n8495 | n8570 ;
  assign n35267 = ~n8569 ;
  assign n8572 = n35267 & n8571 ;
  assign n35268 = ~n8572 ;
  assign n8573 = n165 & n35268 ;
  assign n8044 = n8027 | n8030 ;
  assign n35269 = ~n8044 ;
  assign n8457 = n35269 & n160 ;
  assign n8458 = n7963 | n8457 ;
  assign n8029 = n7963 & n35014 ;
  assign n35270 = ~n8030 ;
  assign n8043 = n8029 & n35270 ;
  assign n8510 = n8043 & n160 ;
  assign n35271 = ~n8510 ;
  assign n8511 = n8458 & n35271 ;
  assign n35272 = ~n8404 ;
  assign n8481 = n35272 & n8477 ;
  assign n35273 = ~n8481 ;
  assign n8482 = n162 & n35273 ;
  assign n8483 = n6889 | n8482 ;
  assign n35274 = ~n8483 ;
  assign n8489 = n35274 & n8486 ;
  assign n8490 = n8475 | n8489 ;
  assign n35275 = ~n8543 ;
  assign n8544 = n8490 & n35275 ;
  assign n35276 = ~n8544 ;
  assign n8545 = n6600 & n35276 ;
  assign n8546 = n165 | n8545 ;
  assign n35277 = ~n8546 ;
  assign n8590 = n35277 & n8571 ;
  assign n8591 = n8511 | n8590 ;
  assign n35278 = ~n8573 ;
  assign n8592 = n35278 & n8591 ;
  assign n35279 = ~n8592 ;
  assign n8593 = n166 & n35279 ;
  assign n8037 = n8033 | n8034 ;
  assign n35280 = ~n8037 ;
  assign n8391 = n35280 & n160 ;
  assign n8392 = n8013 | n8391 ;
  assign n35281 = ~n8034 ;
  assign n8035 = n8013 & n35281 ;
  assign n8036 = n35020 & n8035 ;
  assign n8459 = n8036 & n160 ;
  assign n35282 = ~n8459 ;
  assign n8460 = n8392 & n35282 ;
  assign n8574 = n166 | n8573 ;
  assign n35283 = ~n8574 ;
  assign n8594 = n35283 & n8591 ;
  assign n8595 = n8460 | n8594 ;
  assign n35284 = ~n8593 ;
  assign n8596 = n35284 & n8595 ;
  assign n35285 = ~n8596 ;
  assign n8597 = n5352 & n35285 ;
  assign n8062 = n8040 | n8055 ;
  assign n35286 = ~n8062 ;
  assign n8400 = n35286 & n160 ;
  assign n8401 = n8003 | n8400 ;
  assign n8042 = n8003 & n35031 ;
  assign n35287 = ~n8055 ;
  assign n8061 = n8042 & n35287 ;
  assign n8450 = n8061 & n160 ;
  assign n35288 = ~n8450 ;
  assign n8451 = n8401 & n35288 ;
  assign n8551 = n8490 & n35266 ;
  assign n8552 = n8495 | n8551 ;
  assign n35289 = ~n8545 ;
  assign n8553 = n35289 & n8552 ;
  assign n35290 = ~n8553 ;
  assign n8554 = n165 & n35290 ;
  assign n8555 = n35277 & n8552 ;
  assign n8556 = n8511 | n8555 ;
  assign n35291 = ~n8554 ;
  assign n8557 = n35291 & n8556 ;
  assign n35292 = ~n8557 ;
  assign n8558 = n166 & n35292 ;
  assign n8559 = n5352 | n8558 ;
  assign n35293 = ~n8559 ;
  assign n8603 = n35293 & n8595 ;
  assign n8604 = n8451 | n8603 ;
  assign n35294 = ~n8597 ;
  assign n8605 = n35294 & n8604 ;
  assign n35295 = ~n8605 ;
  assign n8606 = n168 & n35295 ;
  assign n8598 = n4934 | n8597 ;
  assign n35296 = ~n8598 ;
  assign n8607 = n35296 & n8604 ;
  assign n35297 = ~n8059 ;
  assign n8113 = n35297 & n8092 ;
  assign n8114 = n35037 & n8113 ;
  assign n8439 = n8114 & n160 ;
  assign n8060 = n8058 | n8059 ;
  assign n35298 = ~n8060 ;
  assign n8436 = n35298 & n160 ;
  assign n8629 = n8092 | n8436 ;
  assign n35299 = ~n8439 ;
  assign n8630 = n35299 & n8629 ;
  assign n8631 = n8607 | n8630 ;
  assign n35300 = ~n8606 ;
  assign n8632 = n35300 & n8631 ;
  assign n35301 = ~n8632 ;
  assign n8633 = n169 & n35301 ;
  assign n8112 = n8095 | n8098 ;
  assign n35302 = ~n8112 ;
  assign n8433 = n35302 & n160 ;
  assign n8434 = n7953 | n8433 ;
  assign n8097 = n7953 & n35047 ;
  assign n35303 = ~n8098 ;
  assign n8111 = n8097 & n35303 ;
  assign n8522 = n8111 & n160 ;
  assign n35304 = ~n8522 ;
  assign n8523 = n8434 & n35304 ;
  assign n8575 = n8556 & n35283 ;
  assign n8576 = n8460 | n8575 ;
  assign n35305 = ~n8558 ;
  assign n8577 = n35305 & n8576 ;
  assign n35306 = ~n8577 ;
  assign n8578 = n167 & n35306 ;
  assign n8579 = n35293 & n8576 ;
  assign n8580 = n8451 | n8579 ;
  assign n35307 = ~n8578 ;
  assign n8581 = n35307 & n8580 ;
  assign n35308 = ~n8581 ;
  assign n8582 = n4934 & n35308 ;
  assign n8583 = n169 | n8582 ;
  assign n35309 = ~n8583 ;
  assign n8636 = n35309 & n8631 ;
  assign n8637 = n8523 | n8636 ;
  assign n35310 = ~n8633 ;
  assign n8638 = n35310 & n8637 ;
  assign n35311 = ~n8638 ;
  assign n8639 = n170 & n35311 ;
  assign n8110 = n8101 | n8102 ;
  assign n35312 = ~n8110 ;
  assign n8410 = n35312 & n160 ;
  assign n8411 = n7959 | n8410 ;
  assign n35313 = ~n8102 ;
  assign n8108 = n7959 & n35313 ;
  assign n8109 = n35053 & n8108 ;
  assign n8498 = n8109 & n160 ;
  assign n35314 = ~n8498 ;
  assign n8499 = n8411 & n35314 ;
  assign n8634 = n170 | n8633 ;
  assign n35315 = ~n8634 ;
  assign n8640 = n35315 & n8637 ;
  assign n8641 = n8499 | n8640 ;
  assign n35316 = ~n8639 ;
  assign n8642 = n35316 & n8641 ;
  assign n35317 = ~n8642 ;
  assign n8643 = n3940 & n35317 ;
  assign n8107 = n7979 & n35063 ;
  assign n35318 = ~n8123 ;
  assign n8136 = n8107 & n35318 ;
  assign n8467 = n8136 & n160 ;
  assign n8137 = n8105 | n8123 ;
  assign n35319 = ~n8137 ;
  assign n8506 = n35319 & n160 ;
  assign n8507 = n7979 | n8506 ;
  assign n35320 = ~n8467 ;
  assign n8508 = n35320 & n8507 ;
  assign n8599 = n8580 & n35296 ;
  assign n8648 = n8599 | n8630 ;
  assign n35321 = ~n8582 ;
  assign n8649 = n35321 & n8648 ;
  assign n35322 = ~n8649 ;
  assign n8650 = n169 & n35322 ;
  assign n8651 = n35309 & n8648 ;
  assign n8652 = n8523 | n8651 ;
  assign n35323 = ~n8650 ;
  assign n8653 = n35323 & n8652 ;
  assign n35324 = ~n8653 ;
  assign n8654 = n170 & n35324 ;
  assign n8655 = n3940 | n8654 ;
  assign n35325 = ~n8655 ;
  assign n8656 = n8641 & n35325 ;
  assign n8657 = n8508 | n8656 ;
  assign n35326 = ~n8643 ;
  assign n8658 = n35326 & n8657 ;
  assign n35327 = ~n8658 ;
  assign n8659 = n172 & n35327 ;
  assign n35328 = ~n8127 ;
  assign n8133 = n7966 & n35328 ;
  assign n8134 = n35069 & n8133 ;
  assign n8414 = n8134 & n160 ;
  assign n8135 = n8126 | n8127 ;
  assign n35329 = ~n8135 ;
  assign n8445 = n35329 & n160 ;
  assign n8446 = n7966 | n8445 ;
  assign n35330 = ~n8414 ;
  assign n8447 = n35330 & n8446 ;
  assign n8644 = n3631 | n8643 ;
  assign n35331 = ~n8644 ;
  assign n8660 = n35331 & n8657 ;
  assign n8661 = n8447 | n8660 ;
  assign n35332 = ~n8659 ;
  assign n8662 = n35332 & n8661 ;
  assign n35333 = ~n8662 ;
  assign n8663 = n173 & n35333 ;
  assign n8161 = n8130 | n8147 ;
  assign n35334 = ~n8161 ;
  assign n8416 = n35334 & n160 ;
  assign n8417 = n7970 | n8416 ;
  assign n8131 = n7970 & n35079 ;
  assign n35335 = ~n8147 ;
  assign n8160 = n8131 & n35335 ;
  assign n8452 = n8160 & n160 ;
  assign n35336 = ~n8452 ;
  assign n8453 = n8417 & n35336 ;
  assign n8666 = n35315 & n8652 ;
  assign n8667 = n8499 | n8666 ;
  assign n35337 = ~n8654 ;
  assign n8668 = n35337 & n8667 ;
  assign n35338 = ~n8668 ;
  assign n8669 = n171 & n35338 ;
  assign n8670 = n35325 & n8667 ;
  assign n8671 = n8508 | n8670 ;
  assign n35339 = ~n8669 ;
  assign n8672 = n35339 & n8671 ;
  assign n35340 = ~n8672 ;
  assign n8673 = n3631 & n35340 ;
  assign n8674 = n173 | n8673 ;
  assign n35341 = ~n8674 ;
  assign n8675 = n8661 & n35341 ;
  assign n8676 = n8453 | n8675 ;
  assign n35342 = ~n8663 ;
  assign n8677 = n35342 & n8676 ;
  assign n35343 = ~n8677 ;
  assign n8678 = n174 & n35343 ;
  assign n35344 = ~n8151 ;
  assign n8157 = n7973 & n35344 ;
  assign n8158 = n35085 & n8157 ;
  assign n8432 = n8158 & n160 ;
  assign n8159 = n8150 | n8151 ;
  assign n35345 = ~n8159 ;
  assign n8454 = n35345 & n160 ;
  assign n8455 = n7973 | n8454 ;
  assign n35346 = ~n8432 ;
  assign n8456 = n35346 & n8455 ;
  assign n8664 = n174 | n8663 ;
  assign n35347 = ~n8664 ;
  assign n8679 = n35347 & n8676 ;
  assign n8680 = n8456 | n8679 ;
  assign n35348 = ~n8678 ;
  assign n8681 = n35348 & n8680 ;
  assign n35349 = ~n8681 ;
  assign n8682 = n2753 & n35349 ;
  assign n8156 = n7976 & n35095 ;
  assign n35350 = ~n8171 ;
  assign n8184 = n8156 & n35350 ;
  assign n8406 = n8184 & n160 ;
  assign n8185 = n8154 | n8171 ;
  assign n35351 = ~n8185 ;
  assign n8512 = n35351 & n160 ;
  assign n8513 = n7976 | n8512 ;
  assign n35352 = ~n8406 ;
  assign n8514 = n35352 & n8513 ;
  assign n8685 = n35331 & n8671 ;
  assign n8686 = n8447 | n8685 ;
  assign n35353 = ~n8673 ;
  assign n8687 = n35353 & n8686 ;
  assign n35354 = ~n8687 ;
  assign n8688 = n173 & n35354 ;
  assign n8689 = n35341 & n8686 ;
  assign n8690 = n8453 | n8689 ;
  assign n35355 = ~n8688 ;
  assign n8691 = n35355 & n8690 ;
  assign n35356 = ~n8691 ;
  assign n8692 = n174 & n35356 ;
  assign n8693 = n2753 | n8692 ;
  assign n35357 = ~n8693 ;
  assign n8694 = n8680 & n35357 ;
  assign n8695 = n8514 | n8694 ;
  assign n35358 = ~n8682 ;
  assign n8696 = n35358 & n8695 ;
  assign n35359 = ~n8696 ;
  assign n8697 = n176 & n35359 ;
  assign n8178 = n8174 | n8175 ;
  assign n35360 = ~n8178 ;
  assign n8448 = n35360 & n160 ;
  assign n8449 = n7983 | n8448 ;
  assign n35361 = ~n8175 ;
  assign n8176 = n7983 & n35361 ;
  assign n8177 = n35101 & n8176 ;
  assign n8515 = n8177 & n160 ;
  assign n35362 = ~n8515 ;
  assign n8516 = n8449 & n35362 ;
  assign n8683 = n2431 | n8682 ;
  assign n35363 = ~n8683 ;
  assign n8698 = n35363 & n8695 ;
  assign n8699 = n8516 | n8698 ;
  assign n35364 = ~n8697 ;
  assign n8700 = n35364 & n8699 ;
  assign n35365 = ~n8700 ;
  assign n8701 = n177 & n35365 ;
  assign n8209 = n8181 | n8195 ;
  assign n35366 = ~n8209 ;
  assign n8470 = n35366 & n160 ;
  assign n8471 = n7988 | n8470 ;
  assign n8183 = n7988 & n35111 ;
  assign n35367 = ~n8195 ;
  assign n8208 = n8183 & n35367 ;
  assign n8496 = n8208 & n160 ;
  assign n35368 = ~n8496 ;
  assign n8497 = n8471 & n35368 ;
  assign n8704 = n35347 & n8690 ;
  assign n8705 = n8456 | n8704 ;
  assign n35369 = ~n8692 ;
  assign n8706 = n35369 & n8705 ;
  assign n35370 = ~n8706 ;
  assign n8707 = n175 & n35370 ;
  assign n8708 = n35357 & n8705 ;
  assign n8709 = n8514 | n8708 ;
  assign n35371 = ~n8707 ;
  assign n8710 = n35371 & n8709 ;
  assign n35372 = ~n8710 ;
  assign n8711 = n2431 & n35372 ;
  assign n8712 = n177 | n8711 ;
  assign n35373 = ~n8712 ;
  assign n8713 = n8699 & n35373 ;
  assign n8714 = n8497 | n8713 ;
  assign n35374 = ~n8701 ;
  assign n8715 = n35374 & n8714 ;
  assign n35375 = ~n8715 ;
  assign n8716 = n178 & n35375 ;
  assign n35376 = ~n8199 ;
  assign n8205 = n7923 & n35376 ;
  assign n8206 = n35117 & n8205 ;
  assign n8435 = n8206 & n160 ;
  assign n8207 = n8198 | n8199 ;
  assign n35377 = ~n8207 ;
  assign n8491 = n35377 & n160 ;
  assign n8492 = n7923 | n8491 ;
  assign n35378 = ~n8435 ;
  assign n8493 = n35378 & n8492 ;
  assign n8702 = n178 | n8701 ;
  assign n35379 = ~n8702 ;
  assign n8717 = n35379 & n8714 ;
  assign n8718 = n8493 | n8717 ;
  assign n35380 = ~n8716 ;
  assign n8719 = n35380 & n8718 ;
  assign n35381 = ~n8719 ;
  assign n8720 = n1707 & n35381 ;
  assign n8233 = n8202 | n8219 ;
  assign n35382 = ~n8233 ;
  assign n8500 = n35382 & n160 ;
  assign n8501 = n7921 | n8500 ;
  assign n8204 = n7921 & n35127 ;
  assign n35383 = ~n8219 ;
  assign n8232 = n8204 & n35383 ;
  assign n8517 = n8232 & n160 ;
  assign n35384 = ~n8517 ;
  assign n8518 = n8501 & n35384 ;
  assign n8723 = n35363 & n8709 ;
  assign n8724 = n8516 | n8723 ;
  assign n35385 = ~n8711 ;
  assign n8725 = n35385 & n8724 ;
  assign n35386 = ~n8725 ;
  assign n8726 = n177 & n35386 ;
  assign n8727 = n35373 & n8724 ;
  assign n8728 = n8497 | n8727 ;
  assign n35387 = ~n8726 ;
  assign n8729 = n35387 & n8728 ;
  assign n35388 = ~n8729 ;
  assign n8730 = n178 & n35388 ;
  assign n8731 = n1707 | n8730 ;
  assign n35389 = ~n8731 ;
  assign n8732 = n8718 & n35389 ;
  assign n8733 = n8518 | n8732 ;
  assign n35390 = ~n8720 ;
  assign n8734 = n35390 & n8733 ;
  assign n35391 = ~n8734 ;
  assign n8735 = n180 & n35391 ;
  assign n35392 = ~n8223 ;
  assign n8229 = n7916 & n35392 ;
  assign n8230 = n35133 & n8229 ;
  assign n8398 = n8230 & n160 ;
  assign n8231 = n8222 | n8223 ;
  assign n35393 = ~n8231 ;
  assign n8519 = n35393 & n160 ;
  assign n8520 = n7916 | n8519 ;
  assign n35394 = ~n8398 ;
  assign n8521 = n35394 & n8520 ;
  assign n8721 = n1487 | n8720 ;
  assign n35395 = ~n8721 ;
  assign n8736 = n35395 & n8733 ;
  assign n8737 = n8521 | n8736 ;
  assign n35396 = ~n8735 ;
  assign n8738 = n35396 & n8737 ;
  assign n35397 = ~n8738 ;
  assign n8739 = n181 & n35397 ;
  assign n8257 = n8226 | n8243 ;
  assign n35398 = ~n8257 ;
  assign n8437 = n35398 & n160 ;
  assign n8438 = n7911 | n8437 ;
  assign n8228 = n7911 & n35143 ;
  assign n35399 = ~n8243 ;
  assign n8256 = n8228 & n35399 ;
  assign n8443 = n8256 & n160 ;
  assign n35400 = ~n8443 ;
  assign n8444 = n8438 & n35400 ;
  assign n8742 = n35379 & n8728 ;
  assign n8743 = n8493 | n8742 ;
  assign n35401 = ~n8730 ;
  assign n8744 = n35401 & n8743 ;
  assign n35402 = ~n8744 ;
  assign n8745 = n179 & n35402 ;
  assign n8746 = n35389 & n8743 ;
  assign n8747 = n8518 | n8746 ;
  assign n35403 = ~n8745 ;
  assign n8748 = n35403 & n8747 ;
  assign n35404 = ~n8748 ;
  assign n8749 = n1487 & n35404 ;
  assign n8750 = n181 | n8749 ;
  assign n35405 = ~n8750 ;
  assign n8751 = n8737 & n35405 ;
  assign n8752 = n8444 | n8751 ;
  assign n35406 = ~n8739 ;
  assign n8753 = n35406 & n8752 ;
  assign n35407 = ~n8753 ;
  assign n8754 = n182 & n35407 ;
  assign n35408 = ~n8247 ;
  assign n8253 = n7955 & n35408 ;
  assign n8254 = n35149 & n8253 ;
  assign n8397 = n8254 & n160 ;
  assign n8255 = n8246 | n8247 ;
  assign n35409 = ~n8255 ;
  assign n8426 = n35409 & n160 ;
  assign n8427 = n7955 | n8426 ;
  assign n35410 = ~n8397 ;
  assign n8428 = n35410 & n8427 ;
  assign n8740 = n182 | n8739 ;
  assign n35411 = ~n8740 ;
  assign n8755 = n35411 & n8752 ;
  assign n8756 = n8428 | n8755 ;
  assign n35412 = ~n8754 ;
  assign n8757 = n35412 & n8756 ;
  assign n35413 = ~n8757 ;
  assign n8758 = n996 & n35413 ;
  assign n8281 = n8250 | n8267 ;
  assign n35414 = ~n8281 ;
  assign n8524 = n35414 & n160 ;
  assign n8525 = n7940 | n8524 ;
  assign n8252 = n7940 & n35159 ;
  assign n35415 = ~n8267 ;
  assign n8280 = n8252 & n35415 ;
  assign n8535 = n8280 & n8534 ;
  assign n35416 = ~n8535 ;
  assign n8536 = n8525 & n35416 ;
  assign n8761 = n35395 & n8747 ;
  assign n8762 = n8521 | n8761 ;
  assign n35417 = ~n8749 ;
  assign n8763 = n35417 & n8762 ;
  assign n35418 = ~n8763 ;
  assign n8764 = n181 & n35418 ;
  assign n8765 = n35405 & n8762 ;
  assign n8766 = n8444 | n8765 ;
  assign n35419 = ~n8764 ;
  assign n8767 = n35419 & n8766 ;
  assign n35420 = ~n8767 ;
  assign n8768 = n182 & n35420 ;
  assign n8769 = n183 | n8768 ;
  assign n35421 = ~n8769 ;
  assign n8770 = n8756 & n35421 ;
  assign n8771 = n8536 | n8770 ;
  assign n35422 = ~n8758 ;
  assign n8772 = n35422 & n8771 ;
  assign n35423 = ~n8772 ;
  assign n8773 = n184 & n35423 ;
  assign n35424 = ~n8271 ;
  assign n8277 = n7936 & n35424 ;
  assign n8278 = n35165 & n8277 ;
  assign n8429 = n8278 & n160 ;
  assign n8279 = n8270 | n8271 ;
  assign n35425 = ~n8279 ;
  assign n8526 = n35425 & n160 ;
  assign n8527 = n7936 | n8526 ;
  assign n35426 = ~n8429 ;
  assign n8528 = n35426 & n8527 ;
  assign n8759 = n838 | n8758 ;
  assign n35427 = ~n8759 ;
  assign n8774 = n35427 & n8771 ;
  assign n8775 = n8528 | n8774 ;
  assign n35428 = ~n8773 ;
  assign n8776 = n35428 & n8775 ;
  assign n35429 = ~n8776 ;
  assign n8777 = n185 & n35429 ;
  assign n8305 = n8274 | n8291 ;
  assign n35430 = ~n8305 ;
  assign n8395 = n35430 & n160 ;
  assign n8396 = n7902 | n8395 ;
  assign n8276 = n7902 & n35175 ;
  assign n35431 = ~n8291 ;
  assign n8304 = n8276 & n35431 ;
  assign n8502 = n8304 & n160 ;
  assign n35432 = ~n8502 ;
  assign n8503 = n8396 & n35432 ;
  assign n8780 = n35411 & n8766 ;
  assign n8781 = n8428 | n8780 ;
  assign n35433 = ~n8768 ;
  assign n8782 = n35433 & n8781 ;
  assign n35434 = ~n8782 ;
  assign n8783 = n183 & n35434 ;
  assign n8784 = n35421 & n8781 ;
  assign n8785 = n8536 | n8784 ;
  assign n35435 = ~n8783 ;
  assign n8786 = n35435 & n8785 ;
  assign n35436 = ~n8786 ;
  assign n8787 = n838 & n35436 ;
  assign n8788 = n185 | n8787 ;
  assign n35437 = ~n8788 ;
  assign n8789 = n8775 & n35437 ;
  assign n8790 = n8503 | n8789 ;
  assign n35438 = ~n8777 ;
  assign n8791 = n35438 & n8790 ;
  assign n35439 = ~n8791 ;
  assign n8792 = n186 & n35439 ;
  assign n35440 = ~n8295 ;
  assign n8301 = n7905 & n35440 ;
  assign n8302 = n35181 & n8301 ;
  assign n8418 = n8302 & n160 ;
  assign n8303 = n8294 | n8295 ;
  assign n35441 = ~n8303 ;
  assign n8440 = n35441 & n160 ;
  assign n8441 = n7905 | n8440 ;
  assign n35442 = ~n8418 ;
  assign n8442 = n35442 & n8441 ;
  assign n8778 = n186 | n8777 ;
  assign n35443 = ~n8778 ;
  assign n8793 = n35443 & n8790 ;
  assign n8794 = n8442 | n8793 ;
  assign n35444 = ~n8792 ;
  assign n8795 = n35444 & n8794 ;
  assign n35445 = ~n8795 ;
  assign n8796 = n528 & n35445 ;
  assign n8300 = n7957 & n35191 ;
  assign n35446 = ~n8315 ;
  assign n8328 = n8300 & n35446 ;
  assign n8399 = n8328 & n160 ;
  assign n8329 = n8298 | n8315 ;
  assign n35447 = ~n8329 ;
  assign n8407 = n35447 & n160 ;
  assign n8408 = n7957 | n8407 ;
  assign n35448 = ~n8399 ;
  assign n8409 = n35448 & n8408 ;
  assign n8799 = n35427 & n8785 ;
  assign n8800 = n8528 | n8799 ;
  assign n35449 = ~n8787 ;
  assign n8801 = n35449 & n8800 ;
  assign n35450 = ~n8801 ;
  assign n8802 = n185 & n35450 ;
  assign n8803 = n35437 & n8800 ;
  assign n8804 = n8503 | n8803 ;
  assign n35451 = ~n8802 ;
  assign n8805 = n35451 & n8804 ;
  assign n35452 = ~n8805 ;
  assign n8806 = n186 & n35452 ;
  assign n8807 = n528 | n8806 ;
  assign n35453 = ~n8807 ;
  assign n8808 = n8794 & n35453 ;
  assign n8809 = n8409 | n8808 ;
  assign n35454 = ~n8796 ;
  assign n8810 = n35454 & n8809 ;
  assign n35455 = ~n8810 ;
  assign n8811 = n188 & n35455 ;
  assign n8327 = n8318 | n8319 ;
  assign n35456 = ~n8327 ;
  assign n8461 = n35456 & n160 ;
  assign n8462 = n7898 | n8461 ;
  assign n35457 = ~n8319 ;
  assign n8325 = n7898 & n35457 ;
  assign n8326 = n35197 & n8325 ;
  assign n8465 = n8326 & n160 ;
  assign n35458 = ~n8465 ;
  assign n8466 = n8462 & n35458 ;
  assign n8797 = n413 | n8796 ;
  assign n35459 = ~n8797 ;
  assign n8812 = n35459 & n8809 ;
  assign n8813 = n8466 | n8812 ;
  assign n35460 = ~n8811 ;
  assign n8814 = n35460 & n8813 ;
  assign n35461 = ~n8814 ;
  assign n8815 = n189 & n35461 ;
  assign n8324 = n7961 & n35207 ;
  assign n35462 = ~n8339 ;
  assign n8350 = n8324 & n35462 ;
  assign n8509 = n8350 & n160 ;
  assign n8351 = n8322 | n8339 ;
  assign n35463 = ~n8351 ;
  assign n8529 = n35463 & n160 ;
  assign n8530 = n7961 | n8529 ;
  assign n35464 = ~n8509 ;
  assign n8531 = n35464 & n8530 ;
  assign n8818 = n35443 & n8804 ;
  assign n8819 = n8442 | n8818 ;
  assign n35465 = ~n8806 ;
  assign n8820 = n35465 & n8819 ;
  assign n35466 = ~n8820 ;
  assign n8821 = n187 & n35466 ;
  assign n8822 = n35453 & n8819 ;
  assign n8823 = n8409 | n8822 ;
  assign n35467 = ~n8821 ;
  assign n8824 = n35467 & n8823 ;
  assign n35468 = ~n8824 ;
  assign n8825 = n413 & n35468 ;
  assign n8826 = n189 | n8825 ;
  assign n35469 = ~n8826 ;
  assign n8827 = n8813 & n35469 ;
  assign n8828 = n8531 | n8827 ;
  assign n35470 = ~n8815 ;
  assign n8829 = n35470 & n8828 ;
  assign n35471 = ~n8829 ;
  assign n8830 = n190 & n35471 ;
  assign n8621 = n35212 & n8357 ;
  assign n35472 = ~n8621 ;
  assign n8622 = n7927 & n35472 ;
  assign n8623 = n35213 & n8622 ;
  assign n8624 = n160 & n8623 ;
  assign n8625 = n8342 | n8621 ;
  assign n35473 = ~n8625 ;
  assign n8626 = n160 & n35473 ;
  assign n8627 = n7927 | n8626 ;
  assign n35474 = ~n8624 ;
  assign n8628 = n35474 & n8627 ;
  assign n8816 = n190 | n8815 ;
  assign n35475 = ~n8816 ;
  assign n8831 = n35475 & n8828 ;
  assign n8832 = n8628 | n8831 ;
  assign n35476 = ~n8830 ;
  assign n8833 = n35476 & n8832 ;
  assign n35477 = ~n8833 ;
  assign n8834 = n287 & n35477 ;
  assign n8366 = n8346 | n8361 ;
  assign n35478 = ~n8366 ;
  assign n8424 = n35478 & n160 ;
  assign n8425 = n7944 | n8424 ;
  assign n8347 = n7944 & n35223 ;
  assign n35479 = ~n8361 ;
  assign n8365 = n8347 & n35479 ;
  assign n8430 = n8365 & n160 ;
  assign n35480 = ~n8430 ;
  assign n8431 = n8425 & n35480 ;
  assign n8837 = n35459 & n8823 ;
  assign n8838 = n8466 | n8837 ;
  assign n35481 = ~n8825 ;
  assign n8839 = n35481 & n8838 ;
  assign n35482 = ~n8839 ;
  assign n8840 = n189 & n35482 ;
  assign n8841 = n35469 & n8838 ;
  assign n8842 = n8531 | n8841 ;
  assign n35483 = ~n8840 ;
  assign n8843 = n35483 & n8842 ;
  assign n35484 = ~n8843 ;
  assign n8844 = n190 & n35484 ;
  assign n8849 = n287 | n8844 ;
  assign n35485 = ~n8849 ;
  assign n8850 = n8832 & n35485 ;
  assign n8851 = n8431 | n8850 ;
  assign n35486 = ~n8834 ;
  assign n8852 = n35486 & n8851 ;
  assign n8853 = n8618 | n8852 ;
  assign n8854 = n31336 & n8853 ;
  assign n8080 = n7879 | n8076 ;
  assign n35487 = ~n8080 ;
  assign n8081 = n7990 & n35487 ;
  assign n8082 = n35246 & n8081 ;
  assign n8373 = n8082 & n35247 ;
  assign n8385 = n8373 & n35248 ;
  assign n8377 = n192 & n8376 ;
  assign n35488 = ~n7991 ;
  assign n8419 = n35488 & n160 ;
  assign n35489 = ~n8419 ;
  assign n8420 = n8375 & n35489 ;
  assign n35490 = ~n8420 ;
  assign n8421 = n8377 & n35490 ;
  assign n8422 = n8385 | n8421 ;
  assign n8835 = n8617 & n35486 ;
  assign n8855 = n8835 & n8851 ;
  assign n8856 = n8422 | n8855 ;
  assign n8857 = n8854 | n8856 ;
  assign n8911 = n8617 | n8852 ;
  assign n35491 = ~n8911 ;
  assign n8912 = n8857 & n35491 ;
  assign n8913 = n8855 | n8912 ;
  assign n8836 = n8431 & n35486 ;
  assign n8845 = n191 | n8844 ;
  assign n35492 = ~n8845 ;
  assign n8846 = n8832 & n35492 ;
  assign n35493 = ~n8846 ;
  assign n8847 = n8836 & n35493 ;
  assign n8865 = n8847 & n8857 ;
  assign n8848 = n8834 | n8846 ;
  assign n8915 = n35475 & n8842 ;
  assign n8916 = n8628 | n8915 ;
  assign n35494 = ~n8844 ;
  assign n8917 = n35494 & n8916 ;
  assign n35495 = ~n8917 ;
  assign n8918 = n191 & n35495 ;
  assign n8919 = n35492 & n8916 ;
  assign n8920 = n8431 | n8919 ;
  assign n35496 = ~n8918 ;
  assign n8921 = n35496 & n8920 ;
  assign n8922 = n8618 | n8921 ;
  assign n8923 = n31336 & n8922 ;
  assign n8924 = n8835 & n8920 ;
  assign n8925 = n8422 | n8924 ;
  assign n159 = n8923 | n8925 ;
  assign n35497 = ~n8848 ;
  assign n8936 = n35497 & n159 ;
  assign n8937 = n8431 | n8936 ;
  assign n35498 = ~n8865 ;
  assign n8938 = n35498 & n8937 ;
  assign n8939 = n8913 | n8938 ;
  assign n22692 = x58 | x59 ;
  assign n23545 = x60 | n22692 ;
  assign n8083 = n23545 & n35245 ;
  assign n8084 = n35246 & n8083 ;
  assign n8374 = n8084 & n35247 ;
  assign n8387 = n8374 & n35248 ;
  assign n8866 = x60 & n8857 ;
  assign n35499 = ~n8866 ;
  assign n8867 = n8387 & n35499 ;
  assign n35500 = ~n20170 ;
  assign n8864 = n35500 & n8857 ;
  assign n35501 = ~x60 ;
  assign n8869 = n35501 & n8857 ;
  assign n35502 = ~n8869 ;
  assign n8870 = x61 & n35502 ;
  assign n8871 = n8864 | n8870 ;
  assign n8872 = n8867 | n8871 ;
  assign n24413 = n35501 & n22692 ;
  assign n35503 = ~n8857 ;
  assign n8873 = x60 & n35503 ;
  assign n8874 = n24413 | n8873 ;
  assign n35504 = ~n8874 ;
  assign n8881 = n160 & n35504 ;
  assign n35505 = ~n8881 ;
  assign n8882 = n8872 & n35505 ;
  assign n35506 = ~n8882 ;
  assign n8883 = n161 & n35506 ;
  assign n8884 = n162 | n8883 ;
  assign n8875 = n8534 & n35504 ;
  assign n8879 = n161 | n8875 ;
  assign n35507 = ~n8879 ;
  assign n8880 = n8872 & n35507 ;
  assign n35508 = ~n8385 ;
  assign n8504 = n35508 & n160 ;
  assign n35509 = ~n8421 ;
  assign n8505 = n35509 & n8504 ;
  assign n35510 = ~n8855 ;
  assign n8892 = n8505 & n35510 ;
  assign n35511 = ~n8854 ;
  assign n8893 = n35511 & n8892 ;
  assign n8894 = n8864 | n8893 ;
  assign n8895 = x62 & n8894 ;
  assign n8896 = x62 | n8893 ;
  assign n8897 = n8864 | n8896 ;
  assign n35512 = ~n8895 ;
  assign n8898 = n35512 & n8897 ;
  assign n8901 = n8880 | n8898 ;
  assign n35513 = ~n8884 ;
  assign n8902 = n35513 & n8901 ;
  assign n8608 = n8415 | n8539 ;
  assign n35514 = ~n8608 ;
  assign n8609 = n8476 & n35514 ;
  assign n8858 = n8609 & n8857 ;
  assign n8942 = n35514 & n159 ;
  assign n8943 = n8476 | n8942 ;
  assign n35515 = ~n8858 ;
  assign n8944 = n35515 & n8943 ;
  assign n8945 = n8902 | n8944 ;
  assign n35516 = ~n8875 ;
  assign n8876 = n8872 & n35516 ;
  assign n35517 = ~n8876 ;
  assign n8877 = n161 & n35517 ;
  assign n8954 = x60 & n159 ;
  assign n35518 = ~n8954 ;
  assign n8955 = n23545 & n35518 ;
  assign n35519 = ~n8955 ;
  assign n8956 = n160 & n35519 ;
  assign n8957 = n161 | n8956 ;
  assign n35520 = ~n8957 ;
  assign n8958 = n8872 & n35520 ;
  assign n8959 = n8898 | n8958 ;
  assign n35521 = ~n8877 ;
  assign n8960 = n35521 & n8959 ;
  assign n35522 = ~n8960 ;
  assign n8961 = n162 & n35522 ;
  assign n35523 = ~n8961 ;
  assign n8962 = n8945 & n35523 ;
  assign n35524 = ~n8962 ;
  assign n8963 = n6889 & n35524 ;
  assign n8967 = n6889 | n8961 ;
  assign n35525 = ~n8967 ;
  assign n8968 = n8945 & n35525 ;
  assign n35526 = ~n8478 ;
  assign n8487 = n35526 & n8485 ;
  assign n35527 = ~n8482 ;
  assign n8488 = n35527 & n8487 ;
  assign n8863 = n8488 & n8857 ;
  assign n8484 = n8478 | n8482 ;
  assign n35528 = ~n8484 ;
  assign n8977 = n35528 & n159 ;
  assign n8978 = n8485 | n8977 ;
  assign n35529 = ~n8863 ;
  assign n8979 = n35529 & n8978 ;
  assign n8980 = n8968 | n8979 ;
  assign n35530 = ~n8963 ;
  assign n8981 = n35530 & n8980 ;
  assign n35531 = ~n8981 ;
  assign n8982 = n164 & n35531 ;
  assign n8547 = n8475 & n35275 ;
  assign n35532 = ~n8489 ;
  assign n8548 = n35532 & n8547 ;
  assign n8861 = n8548 & n8857 ;
  assign n8549 = n8489 | n8543 ;
  assign n35533 = ~n8549 ;
  assign n8888 = n35533 & n8857 ;
  assign n8889 = n8475 | n8888 ;
  assign n35534 = ~n8861 ;
  assign n8890 = n35534 & n8889 ;
  assign n8964 = n6600 | n8963 ;
  assign n35535 = ~n8964 ;
  assign n8983 = n35535 & n8980 ;
  assign n8984 = n8890 | n8983 ;
  assign n35536 = ~n8982 ;
  assign n8985 = n35536 & n8984 ;
  assign n35537 = ~n8985 ;
  assign n8986 = n165 & n35537 ;
  assign n35538 = ~n8551 ;
  assign n8561 = n8495 & n35538 ;
  assign n8562 = n35289 & n8561 ;
  assign n8891 = n8562 & n8857 ;
  assign n8563 = n8545 | n8551 ;
  assign n35539 = ~n8563 ;
  assign n8948 = n35539 & n159 ;
  assign n8949 = n8495 | n8948 ;
  assign n35540 = ~n8891 ;
  assign n8950 = n35540 & n8949 ;
  assign n8878 = n162 | n8877 ;
  assign n35541 = ~n8878 ;
  assign n8903 = n35541 & n8901 ;
  assign n8946 = n8903 | n8944 ;
  assign n8971 = n8946 & n35523 ;
  assign n35542 = ~n8971 ;
  assign n8972 = n163 & n35542 ;
  assign n8970 = n8946 & n35525 ;
  assign n8989 = n8970 | n8979 ;
  assign n35543 = ~n8972 ;
  assign n8990 = n35543 & n8989 ;
  assign n35544 = ~n8990 ;
  assign n8991 = n6600 & n35544 ;
  assign n8992 = n165 | n8991 ;
  assign n35545 = ~n8992 ;
  assign n8993 = n8984 & n35545 ;
  assign n8994 = n8950 | n8993 ;
  assign n35546 = ~n8986 ;
  assign n8995 = n35546 & n8994 ;
  assign n35547 = ~n8995 ;
  assign n8996 = n166 & n35547 ;
  assign n8588 = n8511 & n35278 ;
  assign n35548 = ~n8555 ;
  assign n8589 = n35548 & n8588 ;
  assign n8868 = n8589 & n8857 ;
  assign n8560 = n8554 | n8555 ;
  assign n35549 = ~n8560 ;
  assign n8933 = n35549 & n159 ;
  assign n8934 = n8511 | n8933 ;
  assign n35550 = ~n8868 ;
  assign n8935 = n35550 & n8934 ;
  assign n8987 = n166 | n8986 ;
  assign n35551 = ~n8987 ;
  assign n8997 = n35551 & n8994 ;
  assign n8998 = n8935 | n8997 ;
  assign n35552 = ~n8996 ;
  assign n8999 = n35552 & n8998 ;
  assign n35553 = ~n8999 ;
  assign n9000 = n5352 & n35553 ;
  assign n35554 = ~n8575 ;
  assign n8585 = n8460 & n35554 ;
  assign n8586 = n35305 & n8585 ;
  assign n8862 = n8586 & n8857 ;
  assign n8587 = n8558 | n8575 ;
  assign n35555 = ~n8587 ;
  assign n8974 = n35555 & n159 ;
  assign n8975 = n8460 | n8974 ;
  assign n35556 = ~n8862 ;
  assign n8976 = n35556 & n8975 ;
  assign n9008 = n35535 & n8989 ;
  assign n9009 = n8890 | n9008 ;
  assign n35557 = ~n8991 ;
  assign n9010 = n35557 & n9009 ;
  assign n35558 = ~n9010 ;
  assign n9011 = n165 & n35558 ;
  assign n9012 = n35545 & n9009 ;
  assign n9013 = n8950 | n9012 ;
  assign n35559 = ~n9011 ;
  assign n9014 = n35559 & n9013 ;
  assign n35560 = ~n9014 ;
  assign n9015 = n166 & n35560 ;
  assign n9016 = n5352 | n9015 ;
  assign n35561 = ~n9016 ;
  assign n9017 = n8998 & n35561 ;
  assign n9018 = n8976 | n9017 ;
  assign n35562 = ~n9000 ;
  assign n9019 = n35562 & n9018 ;
  assign n35563 = ~n9019 ;
  assign n9020 = n168 & n35563 ;
  assign n8601 = n8451 & n35294 ;
  assign n35564 = ~n8579 ;
  assign n8602 = n35564 & n8601 ;
  assign n8860 = n8602 & n8857 ;
  assign n8584 = n8578 | n8579 ;
  assign n35565 = ~n8584 ;
  assign n8951 = n35565 & n159 ;
  assign n8952 = n8451 | n8951 ;
  assign n35566 = ~n8860 ;
  assign n8953 = n35566 & n8952 ;
  assign n9001 = n4934 | n9000 ;
  assign n35567 = ~n9001 ;
  assign n9021 = n35567 & n9018 ;
  assign n9023 = n8953 | n9021 ;
  assign n35568 = ~n9020 ;
  assign n9024 = n35568 & n9023 ;
  assign n35569 = ~n9024 ;
  assign n9025 = n169 & n35569 ;
  assign n9032 = n35551 & n9013 ;
  assign n9033 = n8935 | n9032 ;
  assign n35570 = ~n9015 ;
  assign n9034 = n35570 & n9033 ;
  assign n35571 = ~n9034 ;
  assign n9035 = n167 & n35571 ;
  assign n9036 = n35561 & n9033 ;
  assign n9037 = n8976 | n9036 ;
  assign n35572 = ~n9035 ;
  assign n9038 = n35572 & n9037 ;
  assign n35573 = ~n9038 ;
  assign n9039 = n4934 & n35573 ;
  assign n9040 = n169 | n9039 ;
  assign n35574 = ~n9040 ;
  assign n9041 = n9023 & n35574 ;
  assign n35575 = ~n8599 ;
  assign n8646 = n35575 & n8630 ;
  assign n8647 = n35321 & n8646 ;
  assign n8859 = n8647 & n8857 ;
  assign n8600 = n8582 | n8599 ;
  assign n35576 = ~n8600 ;
  assign n8947 = n35576 & n159 ;
  assign n9195 = n8630 | n8947 ;
  assign n35577 = ~n8859 ;
  assign n9196 = n35577 & n9195 ;
  assign n9212 = n9041 | n9196 ;
  assign n35578 = ~n9025 ;
  assign n9213 = n35578 & n9212 ;
  assign n35579 = ~n9213 ;
  assign n9214 = n170 & n35579 ;
  assign n8635 = n8523 & n35310 ;
  assign n35580 = ~n8651 ;
  assign n9189 = n8635 & n35580 ;
  assign n9190 = n8857 & n9189 ;
  assign n9191 = n8633 | n8651 ;
  assign n35581 = ~n9191 ;
  assign n9192 = n159 & n35581 ;
  assign n9193 = n8523 | n9192 ;
  assign n35582 = ~n9190 ;
  assign n9194 = n35582 & n9193 ;
  assign n9026 = n170 | n9025 ;
  assign n35583 = ~n9026 ;
  assign n9215 = n35583 & n9212 ;
  assign n9216 = n9194 | n9215 ;
  assign n35584 = ~n9214 ;
  assign n9217 = n35584 & n9216 ;
  assign n35585 = ~n9217 ;
  assign n9218 = n3940 & n35585 ;
  assign n35586 = ~n8666 ;
  assign n9182 = n8499 & n35586 ;
  assign n9183 = n35337 & n9182 ;
  assign n9184 = n8857 & n9183 ;
  assign n9185 = n8654 | n8666 ;
  assign n35587 = ~n9185 ;
  assign n9186 = n159 & n35587 ;
  assign n9187 = n8499 | n9186 ;
  assign n35588 = ~n9184 ;
  assign n9188 = n35588 & n9187 ;
  assign n9045 = n35567 & n9037 ;
  assign n9046 = n8953 | n9045 ;
  assign n35589 = ~n9039 ;
  assign n9047 = n35589 & n9046 ;
  assign n35590 = ~n9047 ;
  assign n9048 = n169 & n35590 ;
  assign n9049 = n35574 & n9046 ;
  assign n9197 = n9049 | n9196 ;
  assign n35591 = ~n9048 ;
  assign n9198 = n35591 & n9197 ;
  assign n35592 = ~n9198 ;
  assign n9199 = n170 & n35592 ;
  assign n9200 = n3940 | n9199 ;
  assign n35593 = ~n9200 ;
  assign n9230 = n35593 & n9216 ;
  assign n9231 = n9188 | n9230 ;
  assign n35594 = ~n9218 ;
  assign n9232 = n35594 & n9231 ;
  assign n35595 = ~n9232 ;
  assign n9233 = n172 & n35595 ;
  assign n8645 = n8508 & n35326 ;
  assign n35596 = ~n8670 ;
  assign n9176 = n8645 & n35596 ;
  assign n9177 = n8857 & n9176 ;
  assign n9178 = n8643 | n8670 ;
  assign n35597 = ~n9178 ;
  assign n9179 = n159 & n35597 ;
  assign n9180 = n8508 | n9179 ;
  assign n35598 = ~n9177 ;
  assign n9181 = n35598 & n9180 ;
  assign n9219 = n3631 | n9218 ;
  assign n35599 = ~n9219 ;
  assign n9234 = n35599 & n9231 ;
  assign n9237 = n9181 | n9234 ;
  assign n35600 = ~n9233 ;
  assign n9238 = n35600 & n9237 ;
  assign n35601 = ~n9238 ;
  assign n9239 = n173 & n35601 ;
  assign n35602 = ~n8685 ;
  assign n9169 = n8447 & n35602 ;
  assign n9170 = n35353 & n9169 ;
  assign n9171 = n8857 & n9170 ;
  assign n9172 = n8673 | n8685 ;
  assign n35603 = ~n9172 ;
  assign n9173 = n159 & n35603 ;
  assign n9174 = n8447 | n9173 ;
  assign n35604 = ~n9171 ;
  assign n9175 = n35604 & n9174 ;
  assign n9202 = n35583 & n9197 ;
  assign n9203 = n9194 | n9202 ;
  assign n35605 = ~n9199 ;
  assign n9204 = n35605 & n9203 ;
  assign n35606 = ~n9204 ;
  assign n9205 = n171 & n35606 ;
  assign n9206 = n35593 & n9203 ;
  assign n9207 = n9188 | n9206 ;
  assign n35607 = ~n9205 ;
  assign n9208 = n35607 & n9207 ;
  assign n35608 = ~n9208 ;
  assign n9209 = n3631 & n35608 ;
  assign n9210 = n173 | n9209 ;
  assign n35609 = ~n9210 ;
  assign n9251 = n35609 & n9237 ;
  assign n9252 = n9175 | n9251 ;
  assign n35610 = ~n9239 ;
  assign n9253 = n35610 & n9252 ;
  assign n35611 = ~n9253 ;
  assign n9254 = n174 & n35611 ;
  assign n8665 = n8453 & n35342 ;
  assign n35612 = ~n8689 ;
  assign n9163 = n8665 & n35612 ;
  assign n9164 = n159 & n9163 ;
  assign n9165 = n8688 | n8689 ;
  assign n35613 = ~n9165 ;
  assign n9166 = n159 & n35613 ;
  assign n9167 = n8453 | n9166 ;
  assign n35614 = ~n9164 ;
  assign n9168 = n35614 & n9167 ;
  assign n9240 = n174 | n9239 ;
  assign n35615 = ~n9240 ;
  assign n9255 = n35615 & n9252 ;
  assign n9256 = n9168 | n9255 ;
  assign n35616 = ~n9254 ;
  assign n9257 = n35616 & n9256 ;
  assign n35617 = ~n9257 ;
  assign n9258 = n2753 & n35617 ;
  assign n35618 = ~n8704 ;
  assign n9156 = n8456 & n35618 ;
  assign n9157 = n35369 & n9156 ;
  assign n9158 = n8857 & n9157 ;
  assign n9159 = n8692 | n8704 ;
  assign n35619 = ~n9159 ;
  assign n9160 = n159 & n35619 ;
  assign n9161 = n8456 | n9160 ;
  assign n35620 = ~n9158 ;
  assign n9162 = n35620 & n9161 ;
  assign n9220 = n9207 & n35599 ;
  assign n9221 = n9181 | n9220 ;
  assign n35621 = ~n9209 ;
  assign n9222 = n35621 & n9221 ;
  assign n35622 = ~n9222 ;
  assign n9223 = n173 & n35622 ;
  assign n9224 = n35609 & n9221 ;
  assign n9225 = n9175 | n9224 ;
  assign n35623 = ~n9223 ;
  assign n9226 = n35623 & n9225 ;
  assign n35624 = ~n9226 ;
  assign n9227 = n174 & n35624 ;
  assign n9228 = n2753 | n9227 ;
  assign n35625 = ~n9228 ;
  assign n9270 = n35625 & n9256 ;
  assign n9271 = n9162 | n9270 ;
  assign n35626 = ~n9258 ;
  assign n9272 = n35626 & n9271 ;
  assign n35627 = ~n9272 ;
  assign n9273 = n176 & n35627 ;
  assign n8684 = n8514 & n35358 ;
  assign n35628 = ~n8708 ;
  assign n9150 = n8684 & n35628 ;
  assign n9151 = n8857 & n9150 ;
  assign n9152 = n8707 | n8708 ;
  assign n35629 = ~n9152 ;
  assign n9153 = n159 & n35629 ;
  assign n9154 = n8514 | n9153 ;
  assign n35630 = ~n9151 ;
  assign n9155 = n35630 & n9154 ;
  assign n9259 = n2431 | n9258 ;
  assign n35631 = ~n9259 ;
  assign n9274 = n35631 & n9271 ;
  assign n9275 = n9155 | n9274 ;
  assign n35632 = ~n9273 ;
  assign n9276 = n35632 & n9275 ;
  assign n35633 = ~n9276 ;
  assign n9277 = n177 & n35633 ;
  assign n35634 = ~n8723 ;
  assign n9143 = n8516 & n35634 ;
  assign n9144 = n35385 & n9143 ;
  assign n9145 = n8857 & n9144 ;
  assign n9146 = n8711 | n8723 ;
  assign n35635 = ~n9146 ;
  assign n9147 = n159 & n35635 ;
  assign n9148 = n8516 | n9147 ;
  assign n35636 = ~n9145 ;
  assign n9149 = n35636 & n9148 ;
  assign n9241 = n9225 & n35615 ;
  assign n9242 = n9168 | n9241 ;
  assign n35637 = ~n9227 ;
  assign n9243 = n35637 & n9242 ;
  assign n35638 = ~n9243 ;
  assign n9244 = n175 & n35638 ;
  assign n9245 = n35625 & n9242 ;
  assign n9246 = n9162 | n9245 ;
  assign n35639 = ~n9244 ;
  assign n9247 = n35639 & n9246 ;
  assign n35640 = ~n9247 ;
  assign n9248 = n2431 & n35640 ;
  assign n9249 = n177 | n9248 ;
  assign n35641 = ~n9249 ;
  assign n9289 = n35641 & n9275 ;
  assign n9290 = n9149 | n9289 ;
  assign n35642 = ~n9277 ;
  assign n9291 = n35642 & n9290 ;
  assign n35643 = ~n9291 ;
  assign n9292 = n178 & n35643 ;
  assign n8703 = n8497 & n35374 ;
  assign n35644 = ~n8727 ;
  assign n9137 = n8703 & n35644 ;
  assign n9138 = n8857 & n9137 ;
  assign n9139 = n8726 | n8727 ;
  assign n35645 = ~n9139 ;
  assign n9140 = n159 & n35645 ;
  assign n9141 = n8497 | n9140 ;
  assign n35646 = ~n9138 ;
  assign n9142 = n35646 & n9141 ;
  assign n9278 = n178 | n9277 ;
  assign n35647 = ~n9278 ;
  assign n9293 = n35647 & n9290 ;
  assign n9294 = n9142 | n9293 ;
  assign n35648 = ~n9292 ;
  assign n9295 = n35648 & n9294 ;
  assign n35649 = ~n9295 ;
  assign n9296 = n1707 & n35649 ;
  assign n35650 = ~n8742 ;
  assign n9130 = n8493 & n35650 ;
  assign n9131 = n35401 & n9130 ;
  assign n9132 = n8857 & n9131 ;
  assign n9133 = n8730 | n8742 ;
  assign n35651 = ~n9133 ;
  assign n9134 = n159 & n35651 ;
  assign n9135 = n8493 | n9134 ;
  assign n35652 = ~n9132 ;
  assign n9136 = n35652 & n9135 ;
  assign n9260 = n9246 & n35631 ;
  assign n9261 = n9155 | n9260 ;
  assign n35653 = ~n9248 ;
  assign n9262 = n35653 & n9261 ;
  assign n35654 = ~n9262 ;
  assign n9263 = n177 & n35654 ;
  assign n9264 = n35641 & n9261 ;
  assign n9265 = n9149 | n9264 ;
  assign n35655 = ~n9263 ;
  assign n9266 = n35655 & n9265 ;
  assign n35656 = ~n9266 ;
  assign n9267 = n178 & n35656 ;
  assign n9268 = n1707 | n9267 ;
  assign n35657 = ~n9268 ;
  assign n9308 = n35657 & n9294 ;
  assign n9309 = n9136 | n9308 ;
  assign n35658 = ~n9296 ;
  assign n9310 = n35658 & n9309 ;
  assign n35659 = ~n9310 ;
  assign n9311 = n180 & n35659 ;
  assign n8722 = n8518 & n35390 ;
  assign n35660 = ~n8746 ;
  assign n9124 = n8722 & n35660 ;
  assign n9125 = n8857 & n9124 ;
  assign n9126 = n8720 | n8746 ;
  assign n35661 = ~n9126 ;
  assign n9127 = n159 & n35661 ;
  assign n9128 = n8518 | n9127 ;
  assign n35662 = ~n9125 ;
  assign n9129 = n35662 & n9128 ;
  assign n9297 = n1487 | n9296 ;
  assign n35663 = ~n9297 ;
  assign n9312 = n35663 & n9309 ;
  assign n9313 = n9129 | n9312 ;
  assign n35664 = ~n9311 ;
  assign n9314 = n35664 & n9313 ;
  assign n35665 = ~n9314 ;
  assign n9315 = n181 & n35665 ;
  assign n35666 = ~n8761 ;
  assign n9117 = n8521 & n35666 ;
  assign n9118 = n35417 & n9117 ;
  assign n9119 = n8857 & n9118 ;
  assign n9120 = n8749 | n8761 ;
  assign n35667 = ~n9120 ;
  assign n9121 = n8857 & n35667 ;
  assign n9122 = n8521 | n9121 ;
  assign n35668 = ~n9119 ;
  assign n9123 = n35668 & n9122 ;
  assign n9279 = n9265 & n35647 ;
  assign n9280 = n9142 | n9279 ;
  assign n35669 = ~n9267 ;
  assign n9281 = n35669 & n9280 ;
  assign n35670 = ~n9281 ;
  assign n9282 = n179 & n35670 ;
  assign n9283 = n35657 & n9280 ;
  assign n9284 = n9136 | n9283 ;
  assign n35671 = ~n9282 ;
  assign n9285 = n35671 & n9284 ;
  assign n35672 = ~n9285 ;
  assign n9286 = n1487 & n35672 ;
  assign n9287 = n181 | n9286 ;
  assign n35673 = ~n9287 ;
  assign n9327 = n35673 & n9313 ;
  assign n9328 = n9123 | n9327 ;
  assign n35674 = ~n9315 ;
  assign n9329 = n35674 & n9328 ;
  assign n35675 = ~n9329 ;
  assign n9330 = n182 & n35675 ;
  assign n8741 = n8444 & n35406 ;
  assign n35676 = ~n8765 ;
  assign n9111 = n8741 & n35676 ;
  assign n9112 = n8857 & n9111 ;
  assign n9113 = n8764 | n8765 ;
  assign n35677 = ~n9113 ;
  assign n9114 = n159 & n35677 ;
  assign n9115 = n8444 | n9114 ;
  assign n35678 = ~n9112 ;
  assign n9116 = n35678 & n9115 ;
  assign n9316 = n182 | n9315 ;
  assign n35679 = ~n9316 ;
  assign n9331 = n35679 & n9328 ;
  assign n9334 = n9116 | n9331 ;
  assign n35680 = ~n9330 ;
  assign n9335 = n35680 & n9334 ;
  assign n35681 = ~n9335 ;
  assign n9336 = n996 & n35681 ;
  assign n35682 = ~n8780 ;
  assign n9104 = n8428 & n35682 ;
  assign n9105 = n35433 & n9104 ;
  assign n9106 = n8857 & n9105 ;
  assign n9107 = n8768 | n8780 ;
  assign n35683 = ~n9107 ;
  assign n9108 = n159 & n35683 ;
  assign n9109 = n8428 | n9108 ;
  assign n35684 = ~n9106 ;
  assign n9110 = n35684 & n9109 ;
  assign n9298 = n9284 & n35663 ;
  assign n9299 = n9129 | n9298 ;
  assign n35685 = ~n9286 ;
  assign n9300 = n35685 & n9299 ;
  assign n35686 = ~n9300 ;
  assign n9301 = n181 & n35686 ;
  assign n9302 = n35673 & n9299 ;
  assign n9303 = n9123 | n9302 ;
  assign n35687 = ~n9301 ;
  assign n9304 = n35687 & n9303 ;
  assign n35688 = ~n9304 ;
  assign n9305 = n182 & n35688 ;
  assign n9306 = n183 | n9305 ;
  assign n35689 = ~n9306 ;
  assign n9348 = n35689 & n9334 ;
  assign n9349 = n9110 | n9348 ;
  assign n35690 = ~n9336 ;
  assign n9350 = n35690 & n9349 ;
  assign n35691 = ~n9350 ;
  assign n9351 = n184 & n35691 ;
  assign n8760 = n8536 & n35422 ;
  assign n35692 = ~n8784 ;
  assign n9098 = n8760 & n35692 ;
  assign n9099 = n8857 & n9098 ;
  assign n9100 = n8758 | n8784 ;
  assign n35693 = ~n9100 ;
  assign n9101 = n159 & n35693 ;
  assign n9102 = n8536 | n9101 ;
  assign n35694 = ~n9099 ;
  assign n9103 = n35694 & n9102 ;
  assign n9337 = n838 | n9336 ;
  assign n35695 = ~n9337 ;
  assign n9352 = n35695 & n9349 ;
  assign n9353 = n9103 | n9352 ;
  assign n35696 = ~n9351 ;
  assign n9354 = n35696 & n9353 ;
  assign n35697 = ~n9354 ;
  assign n9355 = n185 & n35697 ;
  assign n35698 = ~n8799 ;
  assign n9091 = n8528 & n35698 ;
  assign n9092 = n35449 & n9091 ;
  assign n9093 = n8857 & n9092 ;
  assign n9094 = n8787 | n8799 ;
  assign n35699 = ~n9094 ;
  assign n9095 = n159 & n35699 ;
  assign n9096 = n8528 | n9095 ;
  assign n35700 = ~n9093 ;
  assign n9097 = n35700 & n9096 ;
  assign n9317 = n9303 & n35679 ;
  assign n9318 = n9116 | n9317 ;
  assign n35701 = ~n9305 ;
  assign n9319 = n35701 & n9318 ;
  assign n35702 = ~n9319 ;
  assign n9320 = n183 & n35702 ;
  assign n9321 = n35689 & n9318 ;
  assign n9322 = n9110 | n9321 ;
  assign n35703 = ~n9320 ;
  assign n9323 = n35703 & n9322 ;
  assign n35704 = ~n9323 ;
  assign n9324 = n838 & n35704 ;
  assign n9325 = n185 | n9324 ;
  assign n35705 = ~n9325 ;
  assign n9367 = n35705 & n9353 ;
  assign n9368 = n9097 | n9367 ;
  assign n35706 = ~n9355 ;
  assign n9369 = n35706 & n9368 ;
  assign n35707 = ~n9369 ;
  assign n9370 = n186 & n35707 ;
  assign n8779 = n8503 & n35438 ;
  assign n35708 = ~n8803 ;
  assign n9085 = n8779 & n35708 ;
  assign n9086 = n8857 & n9085 ;
  assign n9087 = n8777 | n8803 ;
  assign n35709 = ~n9087 ;
  assign n9088 = n159 & n35709 ;
  assign n9089 = n8503 | n9088 ;
  assign n35710 = ~n9086 ;
  assign n9090 = n35710 & n9089 ;
  assign n9356 = n186 | n9355 ;
  assign n35711 = ~n9356 ;
  assign n9371 = n35711 & n9368 ;
  assign n9372 = n9090 | n9371 ;
  assign n35712 = ~n9370 ;
  assign n9373 = n35712 & n9372 ;
  assign n35713 = ~n9373 ;
  assign n9374 = n528 & n35713 ;
  assign n35714 = ~n8818 ;
  assign n9078 = n8442 & n35714 ;
  assign n9079 = n35465 & n9078 ;
  assign n9080 = n8857 & n9079 ;
  assign n9081 = n8806 | n8818 ;
  assign n35715 = ~n9081 ;
  assign n9082 = n159 & n35715 ;
  assign n9083 = n8442 | n9082 ;
  assign n35716 = ~n9080 ;
  assign n9084 = n35716 & n9083 ;
  assign n9338 = n9322 & n35695 ;
  assign n9339 = n9103 | n9338 ;
  assign n35717 = ~n9324 ;
  assign n9340 = n35717 & n9339 ;
  assign n35718 = ~n9340 ;
  assign n9341 = n185 & n35718 ;
  assign n9342 = n35705 & n9339 ;
  assign n9343 = n9097 | n9342 ;
  assign n35719 = ~n9341 ;
  assign n9344 = n35719 & n9343 ;
  assign n35720 = ~n9344 ;
  assign n9345 = n186 & n35720 ;
  assign n9346 = n528 | n9345 ;
  assign n35721 = ~n9346 ;
  assign n9386 = n35721 & n9372 ;
  assign n9387 = n9084 | n9386 ;
  assign n35722 = ~n9374 ;
  assign n9388 = n35722 & n9387 ;
  assign n35723 = ~n9388 ;
  assign n9389 = n188 & n35723 ;
  assign n8798 = n8409 & n35454 ;
  assign n35724 = ~n8822 ;
  assign n9072 = n8798 & n35724 ;
  assign n9073 = n8857 & n9072 ;
  assign n9074 = n8796 | n8822 ;
  assign n35725 = ~n9074 ;
  assign n9075 = n159 & n35725 ;
  assign n9076 = n8409 | n9075 ;
  assign n35726 = ~n9073 ;
  assign n9077 = n35726 & n9076 ;
  assign n9375 = n413 | n9374 ;
  assign n35727 = ~n9375 ;
  assign n9390 = n35727 & n9387 ;
  assign n9391 = n9077 | n9390 ;
  assign n35728 = ~n9389 ;
  assign n9392 = n35728 & n9391 ;
  assign n35729 = ~n9392 ;
  assign n9393 = n189 & n35729 ;
  assign n35730 = ~n8837 ;
  assign n9065 = n8466 & n35730 ;
  assign n9066 = n35481 & n9065 ;
  assign n9067 = n8857 & n9066 ;
  assign n9068 = n8825 | n8837 ;
  assign n35731 = ~n9068 ;
  assign n9069 = n159 & n35731 ;
  assign n9070 = n8466 | n9069 ;
  assign n35732 = ~n9067 ;
  assign n9071 = n35732 & n9070 ;
  assign n9357 = n9343 & n35711 ;
  assign n9358 = n9090 | n9357 ;
  assign n35733 = ~n9345 ;
  assign n9359 = n35733 & n9358 ;
  assign n35734 = ~n9359 ;
  assign n9360 = n187 & n35734 ;
  assign n9361 = n35721 & n9358 ;
  assign n9362 = n9084 | n9361 ;
  assign n35735 = ~n9360 ;
  assign n9363 = n35735 & n9362 ;
  assign n35736 = ~n9363 ;
  assign n9364 = n413 & n35736 ;
  assign n9365 = n189 | n9364 ;
  assign n35737 = ~n9365 ;
  assign n9395 = n35737 & n9391 ;
  assign n9396 = n9071 | n9395 ;
  assign n35738 = ~n9393 ;
  assign n9397 = n35738 & n9396 ;
  assign n35739 = ~n9397 ;
  assign n9398 = n190 & n35739 ;
  assign n8817 = n8531 & n35470 ;
  assign n35740 = ~n8841 ;
  assign n9059 = n8817 & n35740 ;
  assign n9060 = n159 & n9059 ;
  assign n9061 = n8815 | n8841 ;
  assign n35741 = ~n9061 ;
  assign n9062 = n159 & n35741 ;
  assign n9063 = n8531 | n9062 ;
  assign n35742 = ~n9060 ;
  assign n9064 = n35742 & n9063 ;
  assign n9394 = n190 | n9393 ;
  assign n35743 = ~n9394 ;
  assign n9399 = n35743 & n9396 ;
  assign n9400 = n9064 | n9399 ;
  assign n35744 = ~n9398 ;
  assign n9403 = n35744 & n9400 ;
  assign n35745 = ~n9403 ;
  assign n9404 = n287 & n35745 ;
  assign n35746 = ~n8915 ;
  assign n9052 = n8628 & n35746 ;
  assign n9053 = n35494 & n9052 ;
  assign n9054 = n159 & n9053 ;
  assign n9055 = n8844 | n8915 ;
  assign n35747 = ~n9055 ;
  assign n9056 = n159 & n35747 ;
  assign n9057 = n8628 | n9056 ;
  assign n35748 = ~n9054 ;
  assign n9058 = n35748 & n9057 ;
  assign n9376 = n9362 & n35727 ;
  assign n9377 = n9077 | n9376 ;
  assign n35749 = ~n9364 ;
  assign n9378 = n35749 & n9377 ;
  assign n35750 = ~n9378 ;
  assign n9379 = n189 & n35750 ;
  assign n9380 = n35737 & n9377 ;
  assign n9381 = n9071 | n9380 ;
  assign n35751 = ~n9379 ;
  assign n9382 = n35751 & n9381 ;
  assign n35752 = ~n9382 ;
  assign n9383 = n190 & n35752 ;
  assign n9384 = n287 | n9383 ;
  assign n35753 = ~n9384 ;
  assign n9401 = n35753 & n9400 ;
  assign n9408 = n9058 | n9401 ;
  assign n35754 = ~n9404 ;
  assign n9409 = n35754 & n9408 ;
  assign n9410 = n8939 | n9409 ;
  assign n9411 = n31336 & n9410 ;
  assign n8613 = n8385 | n8612 ;
  assign n35755 = ~n8613 ;
  assign n8619 = n35755 & n8616 ;
  assign n8620 = n35509 & n8619 ;
  assign n8906 = n8620 & n35510 ;
  assign n8907 = n35511 & n8906 ;
  assign n8914 = n192 & n8911 ;
  assign n35756 = ~n8617 ;
  assign n8927 = n35756 & n159 ;
  assign n35757 = ~n8927 ;
  assign n8928 = n8852 & n35757 ;
  assign n35758 = ~n8928 ;
  assign n8929 = n8914 & n35758 ;
  assign n8930 = n8907 | n8929 ;
  assign n9405 = n8938 & n35754 ;
  assign n9414 = n9405 & n9408 ;
  assign n9415 = n8930 | n9414 ;
  assign n158 = n9411 | n9415 ;
  assign n35759 = ~n9401 ;
  assign n9402 = n9058 & n35759 ;
  assign n9406 = n9402 & n35754 ;
  assign n9463 = n9406 & n158 ;
  assign n9407 = n9401 | n9404 ;
  assign n35760 = ~n9407 ;
  assign n9464 = n35760 & n158 ;
  assign n9465 = n9058 | n9464 ;
  assign n35761 = ~n9463 ;
  assign n9466 = n35761 & n9465 ;
  assign n9412 = n8938 | n9409 ;
  assign n35762 = ~n9412 ;
  assign n9474 = n35762 & n158 ;
  assign n9620 = n9414 | n9474 ;
  assign n9621 = n9466 | n9620 ;
  assign n25304 = x56 | x57 ;
  assign n26221 = x58 | n25304 ;
  assign n9425 = x58 & n158 ;
  assign n35763 = ~n9425 ;
  assign n9426 = n26221 & n35763 ;
  assign n35764 = ~n9426 ;
  assign n9427 = n159 & n35764 ;
  assign n8386 = n26221 & n35508 ;
  assign n8423 = n8386 & n35509 ;
  assign n8904 = n8423 & n35510 ;
  assign n8905 = n35511 & n8904 ;
  assign n9477 = n8905 & n35763 ;
  assign n35765 = ~n22692 ;
  assign n9443 = n35765 & n158 ;
  assign n35766 = ~x58 ;
  assign n9481 = n35766 & n158 ;
  assign n35767 = ~n9481 ;
  assign n9482 = x59 & n35767 ;
  assign n9483 = n9443 | n9482 ;
  assign n9484 = n9477 | n9483 ;
  assign n35768 = ~n9427 ;
  assign n9487 = n35768 & n9484 ;
  assign n35769 = ~n9487 ;
  assign n9488 = n8534 & n35769 ;
  assign n27031 = n35766 & n25304 ;
  assign n35770 = ~n158 ;
  assign n9470 = x58 & n35770 ;
  assign n9471 = n27031 | n9470 ;
  assign n35771 = ~n9471 ;
  assign n9472 = n8857 & n35771 ;
  assign n9473 = n8534 | n9472 ;
  assign n35772 = ~n9473 ;
  assign n9485 = n35772 & n9484 ;
  assign n35773 = ~n8907 ;
  assign n8908 = n8857 & n35773 ;
  assign n35774 = ~n8929 ;
  assign n8931 = n8908 & n35774 ;
  assign n35775 = ~n9414 ;
  assign n9493 = n8931 & n35775 ;
  assign n35776 = ~n9411 ;
  assign n9494 = n35776 & n9493 ;
  assign n9495 = n9443 | n9494 ;
  assign n9496 = x60 & n9495 ;
  assign n9497 = x60 | n9494 ;
  assign n9498 = n9443 | n9497 ;
  assign n35777 = ~n9496 ;
  assign n9499 = n35777 & n9498 ;
  assign n9500 = n9485 | n9499 ;
  assign n35778 = ~n9488 ;
  assign n9501 = n35778 & n9500 ;
  assign n35779 = ~n9501 ;
  assign n9502 = n161 & n35779 ;
  assign n8886 = n8867 | n8881 ;
  assign n35780 = ~n8886 ;
  assign n9423 = n35780 & n158 ;
  assign n9424 = n8871 | n9423 ;
  assign n8887 = n8871 & n35780 ;
  assign n9475 = n8887 & n158 ;
  assign n35781 = ~n9475 ;
  assign n9476 = n9424 & n35781 ;
  assign n9489 = n161 | n9488 ;
  assign n35782 = ~n9489 ;
  assign n9505 = n35782 & n9500 ;
  assign n9506 = n9476 | n9505 ;
  assign n35783 = ~n9502 ;
  assign n9507 = n35783 & n9506 ;
  assign n35784 = ~n9507 ;
  assign n9508 = n162 & n35784 ;
  assign n35785 = ~n8880 ;
  assign n8899 = n35785 & n8898 ;
  assign n35786 = ~n8883 ;
  assign n8900 = n35786 & n8899 ;
  assign n9435 = n8900 & n158 ;
  assign n8885 = n8880 | n8883 ;
  assign n35787 = ~n8885 ;
  assign n9438 = n35787 & n158 ;
  assign n9439 = n8898 | n9438 ;
  assign n35788 = ~n9435 ;
  assign n9440 = n35788 & n9439 ;
  assign n9503 = n162 | n9502 ;
  assign n35789 = ~n9503 ;
  assign n9509 = n35789 & n9506 ;
  assign n9510 = n9440 | n9509 ;
  assign n35790 = ~n9508 ;
  assign n9511 = n35790 & n9510 ;
  assign n35791 = ~n9511 ;
  assign n9512 = n6889 & n35791 ;
  assign n8973 = n8902 | n8961 ;
  assign n35792 = ~n8973 ;
  assign n9461 = n35792 & n158 ;
  assign n9462 = n8944 | n9461 ;
  assign n8965 = n8944 & n35523 ;
  assign n35793 = ~n8902 ;
  assign n8966 = n35793 & n8965 ;
  assign n9479 = n8966 & n158 ;
  assign n35794 = ~n9479 ;
  assign n9480 = n9462 & n35794 ;
  assign n9490 = n160 & n35769 ;
  assign n9428 = n160 | n9427 ;
  assign n35795 = ~n9428 ;
  assign n9492 = n35795 & n9484 ;
  assign n9521 = n9492 | n9499 ;
  assign n35796 = ~n9490 ;
  assign n9522 = n35796 & n9521 ;
  assign n35797 = ~n9522 ;
  assign n9523 = n161 & n35797 ;
  assign n9524 = n35782 & n9521 ;
  assign n9525 = n9476 | n9524 ;
  assign n35798 = ~n9523 ;
  assign n9526 = n35798 & n9525 ;
  assign n35799 = ~n9526 ;
  assign n9527 = n162 & n35799 ;
  assign n9528 = n6889 | n9527 ;
  assign n35800 = ~n9528 ;
  assign n9529 = n9510 & n35800 ;
  assign n9530 = n9480 | n9529 ;
  assign n35801 = ~n9512 ;
  assign n9531 = n35801 & n9530 ;
  assign n35802 = ~n9531 ;
  assign n9532 = n164 & n35802 ;
  assign n8969 = n8963 | n8968 ;
  assign n35803 = ~n8969 ;
  assign n9421 = n35803 & n158 ;
  assign n9422 = n8979 | n9421 ;
  assign n35804 = ~n8968 ;
  assign n9050 = n35804 & n8979 ;
  assign n9051 = n35530 & n9050 ;
  assign n9441 = n9051 & n158 ;
  assign n35805 = ~n9441 ;
  assign n9442 = n9422 & n35805 ;
  assign n9513 = n6600 | n9512 ;
  assign n35806 = ~n9513 ;
  assign n9533 = n35806 & n9530 ;
  assign n9534 = n9442 | n9533 ;
  assign n35807 = ~n9532 ;
  assign n9535 = n35807 & n9534 ;
  assign n35808 = ~n9535 ;
  assign n9536 = n165 & n35808 ;
  assign n8988 = n8982 | n8983 ;
  assign n35809 = ~n8988 ;
  assign n9431 = n35809 & n158 ;
  assign n9432 = n8890 | n9431 ;
  assign n9006 = n8890 & n35557 ;
  assign n35810 = ~n8983 ;
  assign n9007 = n35810 & n9006 ;
  assign n9436 = n9007 & n158 ;
  assign n35811 = ~n9436 ;
  assign n9437 = n9432 & n35811 ;
  assign n9544 = n35789 & n9525 ;
  assign n9545 = n9440 | n9544 ;
  assign n35812 = ~n9527 ;
  assign n9546 = n35812 & n9545 ;
  assign n35813 = ~n9546 ;
  assign n9547 = n163 & n35813 ;
  assign n9548 = n35800 & n9545 ;
  assign n9549 = n9480 | n9548 ;
  assign n35814 = ~n9547 ;
  assign n9550 = n35814 & n9549 ;
  assign n35815 = ~n9550 ;
  assign n9551 = n6600 & n35815 ;
  assign n9552 = n165 | n9551 ;
  assign n35816 = ~n9552 ;
  assign n9553 = n9534 & n35816 ;
  assign n9554 = n9437 | n9553 ;
  assign n35817 = ~n9536 ;
  assign n9555 = n35817 & n9554 ;
  assign n35818 = ~n9555 ;
  assign n9556 = n166 & n35818 ;
  assign n9005 = n8986 | n8993 ;
  assign n35819 = ~n9005 ;
  assign n9433 = n35819 & n158 ;
  assign n9434 = n8950 | n9433 ;
  assign n35820 = ~n8993 ;
  assign n9003 = n8950 & n35820 ;
  assign n9004 = n35546 & n9003 ;
  assign n9450 = n9004 & n158 ;
  assign n35821 = ~n9450 ;
  assign n9451 = n9434 & n35821 ;
  assign n9537 = n166 | n9536 ;
  assign n35822 = ~n9537 ;
  assign n9557 = n35822 & n9554 ;
  assign n9558 = n9451 | n9557 ;
  assign n35823 = ~n9556 ;
  assign n9559 = n35823 & n9558 ;
  assign n35824 = ~n9559 ;
  assign n9560 = n5352 & n35824 ;
  assign n9002 = n8996 | n8997 ;
  assign n35825 = ~n9002 ;
  assign n9452 = n35825 & n158 ;
  assign n9453 = n8935 | n9452 ;
  assign n9030 = n8935 & n35570 ;
  assign n35826 = ~n8997 ;
  assign n9031 = n35826 & n9030 ;
  assign n9454 = n9031 & n158 ;
  assign n35827 = ~n9454 ;
  assign n9455 = n9453 & n35827 ;
  assign n9568 = n35806 & n9549 ;
  assign n9569 = n9442 | n9568 ;
  assign n35828 = ~n9551 ;
  assign n9570 = n35828 & n9569 ;
  assign n35829 = ~n9570 ;
  assign n9571 = n165 & n35829 ;
  assign n9572 = n35816 & n9569 ;
  assign n9573 = n9437 | n9572 ;
  assign n35830 = ~n9571 ;
  assign n9574 = n35830 & n9573 ;
  assign n35831 = ~n9574 ;
  assign n9575 = n166 & n35831 ;
  assign n9576 = n5352 | n9575 ;
  assign n35832 = ~n9576 ;
  assign n9577 = n9558 & n35832 ;
  assign n9578 = n9455 | n9577 ;
  assign n35833 = ~n9560 ;
  assign n9579 = n35833 & n9578 ;
  assign n35834 = ~n9579 ;
  assign n9580 = n168 & n35834 ;
  assign n35835 = ~n9017 ;
  assign n9027 = n8976 & n35835 ;
  assign n9028 = n35562 & n9027 ;
  assign n9445 = n9028 & n158 ;
  assign n9029 = n9000 | n9017 ;
  assign n35836 = ~n9029 ;
  assign n9456 = n35836 & n158 ;
  assign n9457 = n8976 | n9456 ;
  assign n35837 = ~n9445 ;
  assign n9458 = n35837 & n9457 ;
  assign n9561 = n4934 | n9560 ;
  assign n35838 = ~n9561 ;
  assign n9581 = n35838 & n9578 ;
  assign n9582 = n9458 | n9581 ;
  assign n35839 = ~n9580 ;
  assign n9583 = n35839 & n9582 ;
  assign n35840 = ~n9583 ;
  assign n9584 = n169 & n35840 ;
  assign n9022 = n9020 | n9021 ;
  assign n35841 = ~n9022 ;
  assign n9417 = n35841 & n158 ;
  assign n9418 = n8953 | n9417 ;
  assign n9043 = n8953 & n35589 ;
  assign n35842 = ~n9021 ;
  assign n9044 = n35842 & n9043 ;
  assign n9459 = n9044 & n158 ;
  assign n35843 = ~n9459 ;
  assign n9460 = n9418 & n35843 ;
  assign n9592 = n35822 & n9573 ;
  assign n9593 = n9451 | n9592 ;
  assign n35844 = ~n9575 ;
  assign n9594 = n35844 & n9593 ;
  assign n35845 = ~n9594 ;
  assign n9595 = n167 & n35845 ;
  assign n9596 = n35832 & n9593 ;
  assign n9597 = n9455 | n9596 ;
  assign n35846 = ~n9595 ;
  assign n9598 = n35846 & n9597 ;
  assign n35847 = ~n9598 ;
  assign n9599 = n4934 & n35847 ;
  assign n9600 = n169 | n9599 ;
  assign n35848 = ~n9600 ;
  assign n9601 = n9582 & n35848 ;
  assign n9602 = n9460 | n9601 ;
  assign n35849 = ~n9584 ;
  assign n9603 = n35849 & n9602 ;
  assign n35850 = ~n9603 ;
  assign n9604 = n170 & n35850 ;
  assign n9585 = n170 | n9584 ;
  assign n35851 = ~n9585 ;
  assign n9605 = n35851 & n9602 ;
  assign n35852 = ~n9041 ;
  assign n9758 = n35852 & n9196 ;
  assign n9759 = n35578 & n9758 ;
  assign n9760 = n158 & n9759 ;
  assign n9042 = n9025 | n9041 ;
  assign n35853 = ~n9042 ;
  assign n9444 = n35853 & n158 ;
  assign n9761 = n9196 | n9444 ;
  assign n35854 = ~n9760 ;
  assign n9762 = n35854 & n9761 ;
  assign n9763 = n9605 | n9762 ;
  assign n35855 = ~n9604 ;
  assign n9764 = n35855 & n9763 ;
  assign n35856 = ~n9764 ;
  assign n9765 = n3940 & n35856 ;
  assign n9201 = n9194 & n35605 ;
  assign n35857 = ~n9215 ;
  assign n9752 = n9201 & n35857 ;
  assign n9753 = n158 & n9752 ;
  assign n9754 = n9214 | n9215 ;
  assign n35858 = ~n9754 ;
  assign n9755 = n158 & n35858 ;
  assign n9756 = n9194 | n9755 ;
  assign n35859 = ~n9753 ;
  assign n9757 = n35859 & n9756 ;
  assign n9609 = n35838 & n9597 ;
  assign n9610 = n9458 | n9609 ;
  assign n35860 = ~n9599 ;
  assign n9611 = n35860 & n9610 ;
  assign n35861 = ~n9611 ;
  assign n9612 = n169 & n35861 ;
  assign n9613 = n35848 & n9610 ;
  assign n9614 = n9460 | n9613 ;
  assign n35862 = ~n9612 ;
  assign n9615 = n35862 & n9614 ;
  assign n35863 = ~n9615 ;
  assign n9616 = n170 & n35863 ;
  assign n9617 = n3940 | n9616 ;
  assign n35864 = ~n9617 ;
  assign n9768 = n35864 & n9763 ;
  assign n9769 = n9757 | n9768 ;
  assign n35865 = ~n9765 ;
  assign n9770 = n35865 & n9769 ;
  assign n35866 = ~n9770 ;
  assign n9771 = n172 & n35866 ;
  assign n35867 = ~n9230 ;
  assign n9745 = n9188 & n35867 ;
  assign n9746 = n35594 & n9745 ;
  assign n9747 = n158 & n9746 ;
  assign n9748 = n9218 | n9230 ;
  assign n35868 = ~n9748 ;
  assign n9749 = n158 & n35868 ;
  assign n9750 = n9188 | n9749 ;
  assign n35869 = ~n9747 ;
  assign n9751 = n35869 & n9750 ;
  assign n9766 = n3631 | n9765 ;
  assign n35870 = ~n9766 ;
  assign n9772 = n35870 & n9769 ;
  assign n9773 = n9751 | n9772 ;
  assign n35871 = ~n9771 ;
  assign n9774 = n35871 & n9773 ;
  assign n35872 = ~n9774 ;
  assign n9775 = n173 & n35872 ;
  assign n9211 = n9181 & n35621 ;
  assign n35873 = ~n9234 ;
  assign n9235 = n9211 & n35873 ;
  assign n9446 = n9235 & n158 ;
  assign n9236 = n9233 | n9234 ;
  assign n35874 = ~n9236 ;
  assign n9447 = n35874 & n158 ;
  assign n9448 = n9181 | n9447 ;
  assign n35875 = ~n9446 ;
  assign n9449 = n35875 & n9448 ;
  assign n9619 = n35851 & n9614 ;
  assign n9784 = n9619 | n9762 ;
  assign n35876 = ~n9616 ;
  assign n9785 = n35876 & n9784 ;
  assign n35877 = ~n9785 ;
  assign n9786 = n171 & n35877 ;
  assign n9787 = n35864 & n9784 ;
  assign n9788 = n9757 | n9787 ;
  assign n35878 = ~n9786 ;
  assign n9789 = n35878 & n9788 ;
  assign n35879 = ~n9789 ;
  assign n9790 = n3631 & n35879 ;
  assign n9791 = n173 | n9790 ;
  assign n35880 = ~n9791 ;
  assign n9792 = n9773 & n35880 ;
  assign n9793 = n9449 | n9792 ;
  assign n35881 = ~n9775 ;
  assign n9794 = n35881 & n9793 ;
  assign n35882 = ~n9794 ;
  assign n9795 = n174 & n35882 ;
  assign n35883 = ~n9251 ;
  assign n9738 = n9175 & n35883 ;
  assign n9739 = n35610 & n9738 ;
  assign n9740 = n158 & n9739 ;
  assign n9741 = n9239 | n9251 ;
  assign n35884 = ~n9741 ;
  assign n9742 = n158 & n35884 ;
  assign n9743 = n9175 | n9742 ;
  assign n35885 = ~n9740 ;
  assign n9744 = n35885 & n9743 ;
  assign n9776 = n174 | n9775 ;
  assign n35886 = ~n9776 ;
  assign n9796 = n35886 & n9793 ;
  assign n9797 = n9744 | n9796 ;
  assign n35887 = ~n9795 ;
  assign n9798 = n35887 & n9797 ;
  assign n35888 = ~n9798 ;
  assign n9799 = n2753 & n35888 ;
  assign n9229 = n9168 & n35637 ;
  assign n35889 = ~n9255 ;
  assign n9732 = n9229 & n35889 ;
  assign n9733 = n158 & n9732 ;
  assign n9734 = n9254 | n9255 ;
  assign n35890 = ~n9734 ;
  assign n9735 = n158 & n35890 ;
  assign n9736 = n9168 | n9735 ;
  assign n35891 = ~n9733 ;
  assign n9737 = n35891 & n9736 ;
  assign n9807 = n35870 & n9788 ;
  assign n9808 = n9751 | n9807 ;
  assign n35892 = ~n9790 ;
  assign n9809 = n35892 & n9808 ;
  assign n35893 = ~n9809 ;
  assign n9810 = n173 & n35893 ;
  assign n9811 = n35880 & n9808 ;
  assign n9812 = n9449 | n9811 ;
  assign n35894 = ~n9810 ;
  assign n9813 = n35894 & n9812 ;
  assign n35895 = ~n9813 ;
  assign n9814 = n174 & n35895 ;
  assign n9815 = n2753 | n9814 ;
  assign n35896 = ~n9815 ;
  assign n9816 = n9797 & n35896 ;
  assign n9817 = n9737 | n9816 ;
  assign n35897 = ~n9799 ;
  assign n9818 = n35897 & n9817 ;
  assign n35898 = ~n9818 ;
  assign n9819 = n176 & n35898 ;
  assign n35899 = ~n9270 ;
  assign n9725 = n9162 & n35899 ;
  assign n9726 = n35626 & n9725 ;
  assign n9727 = n158 & n9726 ;
  assign n9728 = n9258 | n9270 ;
  assign n35900 = ~n9728 ;
  assign n9729 = n158 & n35900 ;
  assign n9730 = n9162 | n9729 ;
  assign n35901 = ~n9727 ;
  assign n9731 = n35901 & n9730 ;
  assign n9800 = n2431 | n9799 ;
  assign n35902 = ~n9800 ;
  assign n9820 = n35902 & n9817 ;
  assign n9821 = n9731 | n9820 ;
  assign n35903 = ~n9819 ;
  assign n9822 = n35903 & n9821 ;
  assign n35904 = ~n9822 ;
  assign n9823 = n177 & n35904 ;
  assign n9250 = n9155 & n35653 ;
  assign n35905 = ~n9274 ;
  assign n9719 = n9250 & n35905 ;
  assign n9720 = n158 & n9719 ;
  assign n9721 = n9273 | n9274 ;
  assign n35906 = ~n9721 ;
  assign n9722 = n158 & n35906 ;
  assign n9723 = n9155 | n9722 ;
  assign n35907 = ~n9720 ;
  assign n9724 = n35907 & n9723 ;
  assign n9831 = n35886 & n9812 ;
  assign n9832 = n9744 | n9831 ;
  assign n35908 = ~n9814 ;
  assign n9833 = n35908 & n9832 ;
  assign n35909 = ~n9833 ;
  assign n9834 = n175 & n35909 ;
  assign n9835 = n35896 & n9832 ;
  assign n9836 = n9737 | n9835 ;
  assign n35910 = ~n9834 ;
  assign n9837 = n35910 & n9836 ;
  assign n35911 = ~n9837 ;
  assign n9838 = n2431 & n35911 ;
  assign n9839 = n177 | n9838 ;
  assign n35912 = ~n9839 ;
  assign n9840 = n9821 & n35912 ;
  assign n9841 = n9724 | n9840 ;
  assign n35913 = ~n9823 ;
  assign n9842 = n35913 & n9841 ;
  assign n35914 = ~n9842 ;
  assign n9843 = n178 & n35914 ;
  assign n35915 = ~n9289 ;
  assign n9712 = n9149 & n35915 ;
  assign n9713 = n35642 & n9712 ;
  assign n9714 = n158 & n9713 ;
  assign n9715 = n9277 | n9289 ;
  assign n35916 = ~n9715 ;
  assign n9716 = n158 & n35916 ;
  assign n9717 = n9149 | n9716 ;
  assign n35917 = ~n9714 ;
  assign n9718 = n35917 & n9717 ;
  assign n9824 = n178 | n9823 ;
  assign n35918 = ~n9824 ;
  assign n9844 = n35918 & n9841 ;
  assign n9845 = n9718 | n9844 ;
  assign n35919 = ~n9843 ;
  assign n9846 = n35919 & n9845 ;
  assign n35920 = ~n9846 ;
  assign n9847 = n1707 & n35920 ;
  assign n9269 = n9142 & n35669 ;
  assign n35921 = ~n9293 ;
  assign n9706 = n9269 & n35921 ;
  assign n9707 = n158 & n9706 ;
  assign n9708 = n9292 | n9293 ;
  assign n35922 = ~n9708 ;
  assign n9709 = n158 & n35922 ;
  assign n9710 = n9142 | n9709 ;
  assign n35923 = ~n9707 ;
  assign n9711 = n35923 & n9710 ;
  assign n9855 = n35902 & n9836 ;
  assign n9856 = n9731 | n9855 ;
  assign n35924 = ~n9838 ;
  assign n9857 = n35924 & n9856 ;
  assign n35925 = ~n9857 ;
  assign n9858 = n177 & n35925 ;
  assign n9859 = n35912 & n9856 ;
  assign n9860 = n9724 | n9859 ;
  assign n35926 = ~n9858 ;
  assign n9861 = n35926 & n9860 ;
  assign n35927 = ~n9861 ;
  assign n9862 = n178 & n35927 ;
  assign n9863 = n1707 | n9862 ;
  assign n35928 = ~n9863 ;
  assign n9864 = n9845 & n35928 ;
  assign n9865 = n9711 | n9864 ;
  assign n35929 = ~n9847 ;
  assign n9866 = n35929 & n9865 ;
  assign n35930 = ~n9866 ;
  assign n9867 = n180 & n35930 ;
  assign n35931 = ~n9308 ;
  assign n9699 = n9136 & n35931 ;
  assign n9700 = n35658 & n9699 ;
  assign n9701 = n158 & n9700 ;
  assign n9702 = n9296 | n9308 ;
  assign n35932 = ~n9702 ;
  assign n9703 = n158 & n35932 ;
  assign n9704 = n9136 | n9703 ;
  assign n35933 = ~n9701 ;
  assign n9705 = n35933 & n9704 ;
  assign n9848 = n1487 | n9847 ;
  assign n35934 = ~n9848 ;
  assign n9868 = n35934 & n9865 ;
  assign n9869 = n9705 | n9868 ;
  assign n35935 = ~n9867 ;
  assign n9870 = n35935 & n9869 ;
  assign n35936 = ~n9870 ;
  assign n9871 = n181 & n35936 ;
  assign n9288 = n9129 & n35685 ;
  assign n35937 = ~n9312 ;
  assign n9693 = n9288 & n35937 ;
  assign n9694 = n158 & n9693 ;
  assign n9695 = n9311 | n9312 ;
  assign n35938 = ~n9695 ;
  assign n9696 = n158 & n35938 ;
  assign n9697 = n9129 | n9696 ;
  assign n35939 = ~n9694 ;
  assign n9698 = n35939 & n9697 ;
  assign n9879 = n35918 & n9860 ;
  assign n9880 = n9718 | n9879 ;
  assign n35940 = ~n9862 ;
  assign n9881 = n35940 & n9880 ;
  assign n35941 = ~n9881 ;
  assign n9882 = n179 & n35941 ;
  assign n9883 = n35928 & n9880 ;
  assign n9884 = n9711 | n9883 ;
  assign n35942 = ~n9882 ;
  assign n9885 = n35942 & n9884 ;
  assign n35943 = ~n9885 ;
  assign n9886 = n1487 & n35943 ;
  assign n9887 = n181 | n9886 ;
  assign n35944 = ~n9887 ;
  assign n9888 = n9869 & n35944 ;
  assign n9889 = n9698 | n9888 ;
  assign n35945 = ~n9871 ;
  assign n9890 = n35945 & n9889 ;
  assign n35946 = ~n9890 ;
  assign n9891 = n182 & n35946 ;
  assign n35947 = ~n9327 ;
  assign n9686 = n9123 & n35947 ;
  assign n9687 = n35674 & n9686 ;
  assign n9688 = n158 & n9687 ;
  assign n9689 = n9315 | n9327 ;
  assign n35948 = ~n9689 ;
  assign n9690 = n158 & n35948 ;
  assign n9691 = n9123 | n9690 ;
  assign n35949 = ~n9688 ;
  assign n9692 = n35949 & n9691 ;
  assign n9872 = n182 | n9871 ;
  assign n35950 = ~n9872 ;
  assign n9892 = n35950 & n9889 ;
  assign n9893 = n9692 | n9892 ;
  assign n35951 = ~n9891 ;
  assign n9894 = n35951 & n9893 ;
  assign n35952 = ~n9894 ;
  assign n9895 = n996 & n35952 ;
  assign n9333 = n9330 | n9331 ;
  assign n35953 = ~n9333 ;
  assign n9419 = n35953 & n158 ;
  assign n9420 = n9116 | n9419 ;
  assign n9307 = n9116 & n35701 ;
  assign n35954 = ~n9331 ;
  assign n9332 = n9307 & n35954 ;
  assign n9429 = n9332 & n158 ;
  assign n35955 = ~n9429 ;
  assign n9430 = n9420 & n35955 ;
  assign n9903 = n35934 & n9884 ;
  assign n9904 = n9705 | n9903 ;
  assign n35956 = ~n9886 ;
  assign n9905 = n35956 & n9904 ;
  assign n35957 = ~n9905 ;
  assign n9906 = n181 & n35957 ;
  assign n9907 = n35944 & n9904 ;
  assign n9908 = n9698 | n9907 ;
  assign n35958 = ~n9906 ;
  assign n9909 = n35958 & n9908 ;
  assign n35959 = ~n9909 ;
  assign n9910 = n182 & n35959 ;
  assign n9911 = n183 | n9910 ;
  assign n35960 = ~n9911 ;
  assign n9912 = n9893 & n35960 ;
  assign n9913 = n9430 | n9912 ;
  assign n35961 = ~n9895 ;
  assign n9914 = n35961 & n9913 ;
  assign n35962 = ~n9914 ;
  assign n9915 = n184 & n35962 ;
  assign n35963 = ~n9348 ;
  assign n9679 = n9110 & n35963 ;
  assign n9680 = n35690 & n9679 ;
  assign n9681 = n158 & n9680 ;
  assign n9682 = n9336 | n9348 ;
  assign n35964 = ~n9682 ;
  assign n9683 = n158 & n35964 ;
  assign n9684 = n9110 | n9683 ;
  assign n35965 = ~n9681 ;
  assign n9685 = n35965 & n9684 ;
  assign n9896 = n838 | n9895 ;
  assign n35966 = ~n9896 ;
  assign n9916 = n35966 & n9913 ;
  assign n9917 = n9685 | n9916 ;
  assign n35967 = ~n9915 ;
  assign n9918 = n35967 & n9917 ;
  assign n35968 = ~n9918 ;
  assign n9919 = n185 & n35968 ;
  assign n9326 = n9103 & n35717 ;
  assign n35969 = ~n9352 ;
  assign n9673 = n9326 & n35969 ;
  assign n9674 = n158 & n9673 ;
  assign n9675 = n9351 | n9352 ;
  assign n35970 = ~n9675 ;
  assign n9676 = n158 & n35970 ;
  assign n9677 = n9103 | n9676 ;
  assign n35971 = ~n9674 ;
  assign n9678 = n35971 & n9677 ;
  assign n9927 = n35950 & n9908 ;
  assign n9928 = n9692 | n9927 ;
  assign n35972 = ~n9910 ;
  assign n9929 = n35972 & n9928 ;
  assign n35973 = ~n9929 ;
  assign n9930 = n183 & n35973 ;
  assign n9931 = n35960 & n9928 ;
  assign n9932 = n9430 | n9931 ;
  assign n35974 = ~n9930 ;
  assign n9933 = n35974 & n9932 ;
  assign n35975 = ~n9933 ;
  assign n9934 = n838 & n35975 ;
  assign n9935 = n185 | n9934 ;
  assign n35976 = ~n9935 ;
  assign n9936 = n9917 & n35976 ;
  assign n9937 = n9678 | n9936 ;
  assign n35977 = ~n9919 ;
  assign n9938 = n35977 & n9937 ;
  assign n35978 = ~n9938 ;
  assign n9939 = n186 & n35978 ;
  assign n35979 = ~n9367 ;
  assign n9666 = n9097 & n35979 ;
  assign n9667 = n35706 & n9666 ;
  assign n9668 = n158 & n9667 ;
  assign n9669 = n9355 | n9367 ;
  assign n35980 = ~n9669 ;
  assign n9670 = n158 & n35980 ;
  assign n9671 = n9097 | n9670 ;
  assign n35981 = ~n9668 ;
  assign n9672 = n35981 & n9671 ;
  assign n9920 = n186 | n9919 ;
  assign n35982 = ~n9920 ;
  assign n9940 = n35982 & n9937 ;
  assign n9941 = n9672 | n9940 ;
  assign n35983 = ~n9939 ;
  assign n9942 = n35983 & n9941 ;
  assign n35984 = ~n9942 ;
  assign n9943 = n528 & n35984 ;
  assign n9347 = n9090 & n35733 ;
  assign n35985 = ~n9371 ;
  assign n9660 = n9347 & n35985 ;
  assign n9661 = n158 & n9660 ;
  assign n9662 = n9370 | n9371 ;
  assign n35986 = ~n9662 ;
  assign n9663 = n158 & n35986 ;
  assign n9664 = n9090 | n9663 ;
  assign n35987 = ~n9661 ;
  assign n9665 = n35987 & n9664 ;
  assign n9951 = n35966 & n9932 ;
  assign n9952 = n9685 | n9951 ;
  assign n35988 = ~n9934 ;
  assign n9953 = n35988 & n9952 ;
  assign n35989 = ~n9953 ;
  assign n9954 = n185 & n35989 ;
  assign n9955 = n35976 & n9952 ;
  assign n9956 = n9678 | n9955 ;
  assign n35990 = ~n9954 ;
  assign n9957 = n35990 & n9956 ;
  assign n35991 = ~n9957 ;
  assign n9958 = n186 & n35991 ;
  assign n9959 = n528 | n9958 ;
  assign n35992 = ~n9959 ;
  assign n9960 = n9941 & n35992 ;
  assign n9961 = n9665 | n9960 ;
  assign n35993 = ~n9943 ;
  assign n9962 = n35993 & n9961 ;
  assign n35994 = ~n9962 ;
  assign n9963 = n188 & n35994 ;
  assign n35995 = ~n9386 ;
  assign n9653 = n9084 & n35995 ;
  assign n9654 = n35722 & n9653 ;
  assign n9655 = n158 & n9654 ;
  assign n9656 = n9374 | n9386 ;
  assign n35996 = ~n9656 ;
  assign n9657 = n158 & n35996 ;
  assign n9658 = n9084 | n9657 ;
  assign n35997 = ~n9655 ;
  assign n9659 = n35997 & n9658 ;
  assign n9944 = n413 | n9943 ;
  assign n35998 = ~n9944 ;
  assign n9964 = n35998 & n9961 ;
  assign n9965 = n9659 | n9964 ;
  assign n35999 = ~n9963 ;
  assign n9966 = n35999 & n9965 ;
  assign n36000 = ~n9966 ;
  assign n9967 = n189 & n36000 ;
  assign n9366 = n9077 & n35749 ;
  assign n36001 = ~n9390 ;
  assign n9647 = n9366 & n36001 ;
  assign n9648 = n158 & n9647 ;
  assign n9649 = n9389 | n9390 ;
  assign n36002 = ~n9649 ;
  assign n9650 = n158 & n36002 ;
  assign n9651 = n9077 | n9650 ;
  assign n36003 = ~n9648 ;
  assign n9652 = n36003 & n9651 ;
  assign n9975 = n35982 & n9956 ;
  assign n9976 = n9672 | n9975 ;
  assign n36004 = ~n9958 ;
  assign n9977 = n36004 & n9976 ;
  assign n36005 = ~n9977 ;
  assign n9978 = n187 & n36005 ;
  assign n9979 = n35992 & n9976 ;
  assign n9980 = n9665 | n9979 ;
  assign n36006 = ~n9978 ;
  assign n9981 = n36006 & n9980 ;
  assign n36007 = ~n9981 ;
  assign n9982 = n413 & n36007 ;
  assign n9983 = n189 | n9982 ;
  assign n36008 = ~n9983 ;
  assign n9984 = n9965 & n36008 ;
  assign n9985 = n9652 | n9984 ;
  assign n36009 = ~n9967 ;
  assign n9986 = n36009 & n9985 ;
  assign n36010 = ~n9986 ;
  assign n9987 = n190 & n36010 ;
  assign n36011 = ~n9395 ;
  assign n9640 = n9071 & n36011 ;
  assign n9641 = n35738 & n9640 ;
  assign n9642 = n158 & n9641 ;
  assign n9643 = n9393 | n9395 ;
  assign n36012 = ~n9643 ;
  assign n9644 = n158 & n36012 ;
  assign n9645 = n9071 | n9644 ;
  assign n36013 = ~n9642 ;
  assign n9646 = n36013 & n9645 ;
  assign n9968 = n190 | n9967 ;
  assign n36014 = ~n9968 ;
  assign n9988 = n36014 & n9985 ;
  assign n9989 = n9646 | n9988 ;
  assign n36015 = ~n9987 ;
  assign n9990 = n36015 & n9989 ;
  assign n36016 = ~n9990 ;
  assign n9991 = n287 & n36016 ;
  assign n36017 = ~n9383 ;
  assign n9385 = n9064 & n36017 ;
  assign n36018 = ~n9399 ;
  assign n9634 = n9385 & n36018 ;
  assign n9635 = n158 & n9634 ;
  assign n9636 = n9398 | n9399 ;
  assign n36019 = ~n9636 ;
  assign n9637 = n158 & n36019 ;
  assign n9638 = n9064 | n9637 ;
  assign n36020 = ~n9635 ;
  assign n9639 = n36020 & n9638 ;
  assign n9999 = n35998 & n9980 ;
  assign n10000 = n9659 | n9999 ;
  assign n36021 = ~n9982 ;
  assign n10001 = n36021 & n10000 ;
  assign n36022 = ~n10001 ;
  assign n10002 = n189 & n36022 ;
  assign n10003 = n36008 & n10000 ;
  assign n10004 = n9652 | n10003 ;
  assign n36023 = ~n10002 ;
  assign n10005 = n36023 & n10004 ;
  assign n36024 = ~n10005 ;
  assign n10006 = n190 & n36024 ;
  assign n10007 = n287 | n10006 ;
  assign n36025 = ~n10007 ;
  assign n10008 = n9989 & n36025 ;
  assign n10011 = n9639 | n10008 ;
  assign n36026 = ~n9991 ;
  assign n10012 = n36026 & n10011 ;
  assign n10015 = n9621 | n10012 ;
  assign n10016 = n31336 & n10015 ;
  assign n9413 = n192 & n9412 ;
  assign n36027 = ~n8938 ;
  assign n9467 = n36027 & n158 ;
  assign n36028 = ~n9467 ;
  assign n9468 = n9409 & n36028 ;
  assign n36029 = ~n9468 ;
  assign n9469 = n9413 & n36029 ;
  assign n8909 = n8865 | n8907 ;
  assign n36030 = ~n8909 ;
  assign n8940 = n36030 & n8937 ;
  assign n8941 = n35774 & n8940 ;
  assign n9622 = n8941 & n35775 ;
  assign n9623 = n35776 & n9622 ;
  assign n9624 = n9469 | n9623 ;
  assign n9992 = n9466 & n36026 ;
  assign n10017 = n9992 & n10011 ;
  assign n10018 = n9624 | n10017 ;
  assign n157 = n10016 | n10018 ;
  assign n9993 = n9639 & n36026 ;
  assign n36031 = ~n10008 ;
  assign n10009 = n9993 & n36031 ;
  assign n10146 = n10009 & n157 ;
  assign n10010 = n9991 | n10008 ;
  assign n36032 = ~n10010 ;
  assign n10147 = n36032 & n157 ;
  assign n10148 = n9639 | n10147 ;
  assign n36033 = ~n10146 ;
  assign n10149 = n36033 & n10148 ;
  assign n10013 = n9466 | n10012 ;
  assign n36034 = ~n10013 ;
  assign n10153 = n36034 & n157 ;
  assign n10174 = n10017 | n10153 ;
  assign n10175 = n10149 | n10174 ;
  assign n27977 = x54 | x55 ;
  assign n28941 = x56 | n27977 ;
  assign n10074 = x56 & n157 ;
  assign n36035 = ~n10074 ;
  assign n10097 = n28941 & n36035 ;
  assign n36036 = ~n10097 ;
  assign n10098 = n158 & n36036 ;
  assign n8910 = n28941 & n35773 ;
  assign n8932 = n8910 & n35774 ;
  assign n9632 = n8932 & n35775 ;
  assign n9633 = n35776 & n9632 ;
  assign n10075 = n9633 & n36035 ;
  assign n36037 = ~n25304 ;
  assign n10048 = n36037 & n157 ;
  assign n36038 = ~x56 ;
  assign n10162 = n36038 & n157 ;
  assign n36039 = ~n10162 ;
  assign n10163 = x57 & n36039 ;
  assign n10164 = n10048 | n10163 ;
  assign n10165 = n10075 | n10164 ;
  assign n36040 = ~n10098 ;
  assign n10166 = n36040 & n10165 ;
  assign n36041 = ~n10166 ;
  assign n10167 = n8857 & n36041 ;
  assign n29770 = n36038 & n27977 ;
  assign n36042 = ~n157 ;
  assign n10156 = x56 & n36042 ;
  assign n10157 = n29770 | n10156 ;
  assign n36043 = ~n10157 ;
  assign n10158 = n158 & n36043 ;
  assign n10159 = n8857 | n10158 ;
  assign n36044 = ~n10159 ;
  assign n10170 = n36044 & n10165 ;
  assign n36045 = ~n9623 ;
  assign n9625 = n158 & n36045 ;
  assign n36046 = ~n9469 ;
  assign n9626 = n36046 & n9625 ;
  assign n36047 = ~n10017 ;
  assign n10188 = n9626 & n36047 ;
  assign n36048 = ~n10016 ;
  assign n10189 = n36048 & n10188 ;
  assign n10190 = n10048 | n10189 ;
  assign n10191 = x58 & n10190 ;
  assign n10192 = x58 | n10189 ;
  assign n10193 = n10048 | n10192 ;
  assign n36049 = ~n10191 ;
  assign n10194 = n36049 & n10193 ;
  assign n10195 = n10170 | n10194 ;
  assign n36050 = ~n10167 ;
  assign n10196 = n36050 & n10195 ;
  assign n36051 = ~n10196 ;
  assign n10197 = n8534 & n36051 ;
  assign n9478 = n9472 | n9477 ;
  assign n36052 = ~n9478 ;
  assign n10069 = n36052 & n157 ;
  assign n10070 = n9483 | n10069 ;
  assign n9486 = n36052 & n9483 ;
  assign n10076 = n9486 & n157 ;
  assign n36053 = ~n10076 ;
  assign n10077 = n10070 & n36053 ;
  assign n10168 = n8534 | n10167 ;
  assign n36054 = ~n10168 ;
  assign n10200 = n36054 & n10195 ;
  assign n10201 = n10077 | n10200 ;
  assign n36055 = ~n10197 ;
  assign n10202 = n36055 & n10201 ;
  assign n36056 = ~n10202 ;
  assign n10203 = n161 & n36056 ;
  assign n9491 = n9485 | n9490 ;
  assign n36057 = ~n9491 ;
  assign n10063 = n36057 & n157 ;
  assign n10064 = n9499 | n10063 ;
  assign n36058 = ~n9485 ;
  assign n9519 = n36058 & n9499 ;
  assign n9520 = n35778 & n9519 ;
  assign n10160 = n9520 & n157 ;
  assign n36059 = ~n10160 ;
  assign n10161 = n10064 & n36059 ;
  assign n10198 = n161 | n10197 ;
  assign n36060 = ~n10198 ;
  assign n10204 = n36060 & n10201 ;
  assign n10205 = n10161 | n10204 ;
  assign n36061 = ~n10203 ;
  assign n10206 = n36061 & n10205 ;
  assign n36062 = ~n10206 ;
  assign n10207 = n162 & n36062 ;
  assign n9518 = n9502 | n9505 ;
  assign n36063 = ~n9518 ;
  assign n10059 = n36063 & n157 ;
  assign n10060 = n9476 | n10059 ;
  assign n9504 = n9476 & n35783 ;
  assign n36064 = ~n9505 ;
  assign n9517 = n9504 & n36064 ;
  assign n10154 = n9517 & n157 ;
  assign n36065 = ~n10154 ;
  assign n10155 = n10060 & n36065 ;
  assign n10169 = n159 & n36041 ;
  assign n10099 = n159 | n10098 ;
  assign n36066 = ~n10099 ;
  assign n10172 = n36066 & n10165 ;
  assign n10217 = n10172 | n10194 ;
  assign n36067 = ~n10169 ;
  assign n10218 = n36067 & n10217 ;
  assign n36068 = ~n10218 ;
  assign n10219 = n160 & n36068 ;
  assign n10220 = n36054 & n10217 ;
  assign n10221 = n10077 | n10220 ;
  assign n36069 = ~n10219 ;
  assign n10222 = n36069 & n10221 ;
  assign n36070 = ~n10222 ;
  assign n10223 = n161 & n36070 ;
  assign n10224 = n162 | n10223 ;
  assign n36071 = ~n10224 ;
  assign n10225 = n10205 & n36071 ;
  assign n10226 = n10155 | n10225 ;
  assign n36072 = ~n10207 ;
  assign n10227 = n36072 & n10226 ;
  assign n36073 = ~n10227 ;
  assign n10228 = n163 & n36073 ;
  assign n36074 = ~n9509 ;
  assign n9515 = n9440 & n36074 ;
  assign n9516 = n35790 & n9515 ;
  assign n10039 = n9516 & n157 ;
  assign n9543 = n9509 | n9527 ;
  assign n36075 = ~n9543 ;
  assign n10049 = n36075 & n157 ;
  assign n10050 = n9440 | n10049 ;
  assign n36076 = ~n10039 ;
  assign n10051 = n36076 & n10050 ;
  assign n10209 = n6889 | n10207 ;
  assign n36077 = ~n10209 ;
  assign n10229 = n36077 & n10226 ;
  assign n10230 = n10051 | n10229 ;
  assign n36078 = ~n10228 ;
  assign n10231 = n36078 & n10230 ;
  assign n36079 = ~n10231 ;
  assign n10232 = n6600 & n36079 ;
  assign n9514 = n9480 & n35801 ;
  assign n36080 = ~n9529 ;
  assign n9542 = n9514 & n36080 ;
  assign n10047 = n9542 & n157 ;
  assign n9541 = n9512 | n9529 ;
  assign n36081 = ~n9541 ;
  assign n10071 = n36081 & n157 ;
  assign n10072 = n9480 | n10071 ;
  assign n36082 = ~n10047 ;
  assign n10073 = n36082 & n10072 ;
  assign n10240 = n36060 & n10221 ;
  assign n10241 = n10161 | n10240 ;
  assign n36083 = ~n10223 ;
  assign n10242 = n36083 & n10241 ;
  assign n36084 = ~n10242 ;
  assign n10243 = n162 & n36084 ;
  assign n10244 = n36071 & n10241 ;
  assign n10245 = n10155 | n10244 ;
  assign n36085 = ~n10243 ;
  assign n10246 = n36085 & n10245 ;
  assign n36086 = ~n10246 ;
  assign n10247 = n6889 & n36086 ;
  assign n10248 = n6600 | n10247 ;
  assign n36087 = ~n10248 ;
  assign n10249 = n10230 & n36087 ;
  assign n10250 = n10073 | n10249 ;
  assign n36088 = ~n10232 ;
  assign n10251 = n36088 & n10250 ;
  assign n36089 = ~n10251 ;
  assign n10252 = n165 & n36089 ;
  assign n9567 = n9533 | n9551 ;
  assign n36090 = ~n9567 ;
  assign n10056 = n36090 & n157 ;
  assign n10057 = n9442 | n10056 ;
  assign n36091 = ~n9533 ;
  assign n9539 = n9442 & n36091 ;
  assign n9540 = n35807 & n9539 ;
  assign n10104 = n9540 & n157 ;
  assign n36092 = ~n10104 ;
  assign n10105 = n10057 & n36092 ;
  assign n10233 = n165 | n10232 ;
  assign n36093 = ~n10233 ;
  assign n10253 = n36093 & n10250 ;
  assign n10254 = n10105 | n10253 ;
  assign n36094 = ~n10252 ;
  assign n10255 = n36094 & n10254 ;
  assign n36095 = ~n10255 ;
  assign n10256 = n166 & n36095 ;
  assign n9566 = n9536 | n9553 ;
  assign n36096 = ~n9566 ;
  assign n10095 = n36096 & n157 ;
  assign n10096 = n9437 | n10095 ;
  assign n9538 = n9437 & n35817 ;
  assign n36097 = ~n9553 ;
  assign n9565 = n9538 & n36097 ;
  assign n10106 = n9565 & n157 ;
  assign n36098 = ~n10106 ;
  assign n10107 = n10096 & n36098 ;
  assign n10264 = n36077 & n10245 ;
  assign n10265 = n10051 | n10264 ;
  assign n36099 = ~n10247 ;
  assign n10266 = n36099 & n10265 ;
  assign n36100 = ~n10266 ;
  assign n10267 = n164 & n36100 ;
  assign n10268 = n36087 & n10265 ;
  assign n10269 = n10073 | n10268 ;
  assign n36101 = ~n10267 ;
  assign n10270 = n36101 & n10269 ;
  assign n36102 = ~n10270 ;
  assign n10271 = n165 & n36102 ;
  assign n10272 = n166 | n10271 ;
  assign n36103 = ~n10272 ;
  assign n10273 = n10254 & n36103 ;
  assign n10274 = n10107 | n10273 ;
  assign n36104 = ~n10256 ;
  assign n10275 = n36104 & n10274 ;
  assign n36105 = ~n10275 ;
  assign n10276 = n167 & n36105 ;
  assign n36106 = ~n9557 ;
  assign n9563 = n9451 & n36106 ;
  assign n9564 = n35823 & n9563 ;
  assign n10079 = n9564 & n157 ;
  assign n9591 = n9557 | n9575 ;
  assign n36107 = ~n9591 ;
  assign n10108 = n36107 & n157 ;
  assign n10109 = n9451 | n10108 ;
  assign n36108 = ~n10079 ;
  assign n10110 = n36108 & n10109 ;
  assign n10257 = n5352 | n10256 ;
  assign n36109 = ~n10257 ;
  assign n10277 = n36109 & n10274 ;
  assign n10278 = n10110 | n10277 ;
  assign n36110 = ~n10276 ;
  assign n10279 = n36110 & n10278 ;
  assign n36111 = ~n10279 ;
  assign n10280 = n4934 & n36111 ;
  assign n9562 = n9455 & n35833 ;
  assign n36112 = ~n9577 ;
  assign n9589 = n9562 & n36112 ;
  assign n10058 = n9589 & n157 ;
  assign n9590 = n9560 | n9577 ;
  assign n36113 = ~n9590 ;
  assign n10065 = n36113 & n157 ;
  assign n10066 = n9455 | n10065 ;
  assign n36114 = ~n10058 ;
  assign n10067 = n36114 & n10066 ;
  assign n10288 = n36093 & n10269 ;
  assign n10289 = n10105 | n10288 ;
  assign n36115 = ~n10271 ;
  assign n10290 = n36115 & n10289 ;
  assign n36116 = ~n10290 ;
  assign n10291 = n166 & n36116 ;
  assign n10292 = n36103 & n10289 ;
  assign n10293 = n10107 | n10292 ;
  assign n36117 = ~n10291 ;
  assign n10294 = n36117 & n10293 ;
  assign n36118 = ~n10294 ;
  assign n10295 = n5352 & n36118 ;
  assign n10296 = n4934 | n10295 ;
  assign n36119 = ~n10296 ;
  assign n10297 = n10278 & n36119 ;
  assign n10298 = n10067 | n10297 ;
  assign n36120 = ~n10280 ;
  assign n10299 = n36120 & n10298 ;
  assign n36121 = ~n10299 ;
  assign n10300 = n169 & n36121 ;
  assign n9608 = n9581 | n9599 ;
  assign n36122 = ~n9608 ;
  assign n10125 = n36122 & n157 ;
  assign n10126 = n9458 | n10125 ;
  assign n36123 = ~n9581 ;
  assign n9587 = n9458 & n36123 ;
  assign n9588 = n35839 & n9587 ;
  assign n10129 = n9588 & n157 ;
  assign n36124 = ~n10129 ;
  assign n10130 = n10126 & n36124 ;
  assign n10281 = n169 | n10280 ;
  assign n36125 = ~n10281 ;
  assign n10301 = n36125 & n10298 ;
  assign n10302 = n10130 | n10301 ;
  assign n36126 = ~n10300 ;
  assign n10303 = n36126 & n10302 ;
  assign n36127 = ~n10303 ;
  assign n10304 = n170 & n36127 ;
  assign n9607 = n9584 | n9601 ;
  assign n36128 = ~n9607 ;
  assign n10082 = n36128 & n157 ;
  assign n10083 = n9460 | n10082 ;
  assign n9586 = n9460 & n35849 ;
  assign n36129 = ~n9601 ;
  assign n9606 = n9586 & n36129 ;
  assign n10088 = n9606 & n157 ;
  assign n36130 = ~n10088 ;
  assign n10089 = n10083 & n36130 ;
  assign n10312 = n36109 & n10293 ;
  assign n10313 = n10110 | n10312 ;
  assign n36131 = ~n10295 ;
  assign n10314 = n36131 & n10313 ;
  assign n36132 = ~n10314 ;
  assign n10315 = n168 & n36132 ;
  assign n10316 = n36119 & n10313 ;
  assign n10317 = n10067 | n10316 ;
  assign n36133 = ~n10315 ;
  assign n10318 = n36133 & n10317 ;
  assign n36134 = ~n10318 ;
  assign n10319 = n169 & n36134 ;
  assign n10320 = n170 | n10319 ;
  assign n36135 = ~n10320 ;
  assign n10321 = n10302 & n36135 ;
  assign n10322 = n10089 | n10321 ;
  assign n36136 = ~n10304 ;
  assign n10323 = n36136 & n10322 ;
  assign n36137 = ~n10323 ;
  assign n10324 = n171 & n36137 ;
  assign n10305 = n3940 | n10304 ;
  assign n36138 = ~n10305 ;
  assign n10325 = n36138 & n10322 ;
  assign n36139 = ~n9605 ;
  assign n9782 = n36139 & n9762 ;
  assign n9783 = n35855 & n9782 ;
  assign n10116 = n9783 & n157 ;
  assign n9618 = n9605 | n9616 ;
  assign n36140 = ~n9618 ;
  assign n10136 = n36140 & n157 ;
  assign n10343 = n9762 | n10136 ;
  assign n36141 = ~n10116 ;
  assign n10344 = n36141 & n10343 ;
  assign n10345 = n10325 | n10344 ;
  assign n36142 = ~n10324 ;
  assign n10346 = n36142 & n10345 ;
  assign n36143 = ~n10346 ;
  assign n10347 = n3631 & n36143 ;
  assign n9781 = n9765 | n9768 ;
  assign n36144 = ~n9781 ;
  assign n10032 = n36144 & n157 ;
  assign n10033 = n9757 | n10032 ;
  assign n9767 = n9757 & n35865 ;
  assign n36145 = ~n9768 ;
  assign n9780 = n9767 & n36145 ;
  assign n10117 = n9780 & n157 ;
  assign n36146 = ~n10117 ;
  assign n10118 = n10033 & n36146 ;
  assign n10329 = n36125 & n10317 ;
  assign n10330 = n10130 | n10329 ;
  assign n36147 = ~n10319 ;
  assign n10331 = n36147 & n10330 ;
  assign n36148 = ~n10331 ;
  assign n10332 = n170 & n36148 ;
  assign n10333 = n36135 & n10330 ;
  assign n10334 = n10089 | n10333 ;
  assign n36149 = ~n10332 ;
  assign n10335 = n36149 & n10334 ;
  assign n36150 = ~n10335 ;
  assign n10336 = n3940 & n36150 ;
  assign n10337 = n3631 | n10336 ;
  assign n36151 = ~n10337 ;
  assign n10350 = n36151 & n10345 ;
  assign n10351 = n10118 | n10350 ;
  assign n36152 = ~n10347 ;
  assign n10352 = n36152 & n10351 ;
  assign n36153 = ~n10352 ;
  assign n10353 = n173 & n36153 ;
  assign n9806 = n9772 | n9790 ;
  assign n36154 = ~n9806 ;
  assign n10080 = n36154 & n157 ;
  assign n10081 = n9751 | n10080 ;
  assign n36155 = ~n9772 ;
  assign n9778 = n9751 & n36155 ;
  assign n9779 = n35871 & n9778 ;
  assign n10127 = n9779 & n157 ;
  assign n36156 = ~n10127 ;
  assign n10128 = n10081 & n36156 ;
  assign n10348 = n173 | n10347 ;
  assign n36157 = ~n10348 ;
  assign n10354 = n36157 & n10351 ;
  assign n10355 = n10128 | n10354 ;
  assign n36158 = ~n10353 ;
  assign n10356 = n36158 & n10355 ;
  assign n36159 = ~n10356 ;
  assign n10357 = n174 & n36159 ;
  assign n9777 = n9449 & n35881 ;
  assign n36160 = ~n9792 ;
  assign n9804 = n9777 & n36160 ;
  assign n10046 = n9804 & n157 ;
  assign n9805 = n9775 | n9792 ;
  assign n36161 = ~n9805 ;
  assign n10113 = n36161 & n157 ;
  assign n10114 = n9449 | n10113 ;
  assign n36162 = ~n10046 ;
  assign n10115 = n36162 & n10114 ;
  assign n10338 = n36138 & n10334 ;
  assign n10367 = n10338 | n10344 ;
  assign n36163 = ~n10336 ;
  assign n10368 = n36163 & n10367 ;
  assign n36164 = ~n10368 ;
  assign n10369 = n172 & n36164 ;
  assign n10370 = n36151 & n10367 ;
  assign n10371 = n10118 | n10370 ;
  assign n36165 = ~n10369 ;
  assign n10372 = n36165 & n10371 ;
  assign n36166 = ~n10372 ;
  assign n10373 = n173 & n36166 ;
  assign n10374 = n174 | n10373 ;
  assign n36167 = ~n10374 ;
  assign n10375 = n10355 & n36167 ;
  assign n10376 = n10115 | n10375 ;
  assign n36168 = ~n10357 ;
  assign n10377 = n36168 & n10376 ;
  assign n36169 = ~n10377 ;
  assign n10378 = n175 & n36169 ;
  assign n36170 = ~n9796 ;
  assign n9802 = n9744 & n36170 ;
  assign n9803 = n35887 & n9802 ;
  assign n10042 = n9803 & n157 ;
  assign n9830 = n9796 | n9814 ;
  assign n36171 = ~n9830 ;
  assign n10043 = n36171 & n157 ;
  assign n10044 = n9744 | n10043 ;
  assign n36172 = ~n10042 ;
  assign n10045 = n36172 & n10044 ;
  assign n10358 = n2753 | n10357 ;
  assign n36173 = ~n10358 ;
  assign n10379 = n36173 & n10376 ;
  assign n10380 = n10045 | n10379 ;
  assign n36174 = ~n10378 ;
  assign n10381 = n36174 & n10380 ;
  assign n36175 = ~n10381 ;
  assign n10382 = n2431 & n36175 ;
  assign n9829 = n9799 | n9816 ;
  assign n36176 = ~n9829 ;
  assign n10040 = n36176 & n157 ;
  assign n10041 = n9737 | n10040 ;
  assign n9801 = n9737 & n35897 ;
  assign n36177 = ~n9816 ;
  assign n9828 = n9801 & n36177 ;
  assign n10086 = n9828 & n157 ;
  assign n36178 = ~n10086 ;
  assign n10087 = n10041 & n36178 ;
  assign n10390 = n36157 & n10371 ;
  assign n10391 = n10128 | n10390 ;
  assign n36179 = ~n10373 ;
  assign n10392 = n36179 & n10391 ;
  assign n36180 = ~n10392 ;
  assign n10393 = n174 & n36180 ;
  assign n10394 = n36167 & n10391 ;
  assign n10395 = n10115 | n10394 ;
  assign n36181 = ~n10393 ;
  assign n10396 = n36181 & n10395 ;
  assign n36182 = ~n10396 ;
  assign n10397 = n2753 & n36182 ;
  assign n10398 = n2431 | n10397 ;
  assign n36183 = ~n10398 ;
  assign n10399 = n10380 & n36183 ;
  assign n10400 = n10087 | n10399 ;
  assign n36184 = ~n10382 ;
  assign n10401 = n36184 & n10400 ;
  assign n36185 = ~n10401 ;
  assign n10402 = n177 & n36185 ;
  assign n36186 = ~n9820 ;
  assign n9826 = n9731 & n36186 ;
  assign n9827 = n35903 & n9826 ;
  assign n10094 = n9827 & n157 ;
  assign n9854 = n9820 | n9838 ;
  assign n36187 = ~n9854 ;
  assign n10122 = n36187 & n157 ;
  assign n10123 = n9731 | n10122 ;
  assign n36188 = ~n10094 ;
  assign n10124 = n36188 & n10123 ;
  assign n10383 = n177 | n10382 ;
  assign n36189 = ~n10383 ;
  assign n10403 = n36189 & n10400 ;
  assign n10404 = n10124 | n10403 ;
  assign n36190 = ~n10402 ;
  assign n10405 = n36190 & n10404 ;
  assign n36191 = ~n10405 ;
  assign n10406 = n178 & n36191 ;
  assign n9825 = n9724 & n35913 ;
  assign n36192 = ~n9840 ;
  assign n9852 = n9825 & n36192 ;
  assign n10093 = n9852 & n157 ;
  assign n9853 = n9823 | n9840 ;
  assign n36193 = ~n9853 ;
  assign n10119 = n36193 & n157 ;
  assign n10120 = n9724 | n10119 ;
  assign n36194 = ~n10093 ;
  assign n10121 = n36194 & n10120 ;
  assign n10414 = n36173 & n10395 ;
  assign n10415 = n10045 | n10414 ;
  assign n36195 = ~n10397 ;
  assign n10416 = n36195 & n10415 ;
  assign n36196 = ~n10416 ;
  assign n10417 = n176 & n36196 ;
  assign n10418 = n36183 & n10415 ;
  assign n10419 = n10087 | n10418 ;
  assign n36197 = ~n10417 ;
  assign n10420 = n36197 & n10419 ;
  assign n36198 = ~n10420 ;
  assign n10421 = n177 & n36198 ;
  assign n10422 = n178 | n10421 ;
  assign n36199 = ~n10422 ;
  assign n10423 = n10404 & n36199 ;
  assign n10424 = n10121 | n10423 ;
  assign n36200 = ~n10406 ;
  assign n10425 = n36200 & n10424 ;
  assign n36201 = ~n10425 ;
  assign n10426 = n179 & n36201 ;
  assign n36202 = ~n9844 ;
  assign n9850 = n9718 & n36202 ;
  assign n9851 = n35919 & n9850 ;
  assign n10038 = n9851 & n157 ;
  assign n9878 = n9844 | n9862 ;
  assign n36203 = ~n9878 ;
  assign n10133 = n36203 & n157 ;
  assign n10134 = n9718 | n10133 ;
  assign n36204 = ~n10038 ;
  assign n10135 = n36204 & n10134 ;
  assign n10407 = n1707 | n10406 ;
  assign n36205 = ~n10407 ;
  assign n10427 = n36205 & n10424 ;
  assign n10428 = n10135 | n10427 ;
  assign n36206 = ~n10426 ;
  assign n10429 = n36206 & n10428 ;
  assign n36207 = ~n10429 ;
  assign n10430 = n1487 & n36207 ;
  assign n9877 = n9847 | n9864 ;
  assign n36208 = ~n9877 ;
  assign n10034 = n36208 & n157 ;
  assign n10035 = n9711 | n10034 ;
  assign n9849 = n9711 & n35929 ;
  assign n36209 = ~n9864 ;
  assign n9876 = n9849 & n36209 ;
  assign n10054 = n9876 & n157 ;
  assign n36210 = ~n10054 ;
  assign n10055 = n10035 & n36210 ;
  assign n10436 = n36189 & n10419 ;
  assign n10437 = n10124 | n10436 ;
  assign n36211 = ~n10421 ;
  assign n10438 = n36211 & n10437 ;
  assign n36212 = ~n10438 ;
  assign n10439 = n178 & n36212 ;
  assign n10440 = n36199 & n10437 ;
  assign n10441 = n10121 | n10440 ;
  assign n36213 = ~n10439 ;
  assign n10442 = n36213 & n10441 ;
  assign n36214 = ~n10442 ;
  assign n10443 = n1707 & n36214 ;
  assign n10444 = n1487 | n10443 ;
  assign n36215 = ~n10444 ;
  assign n10445 = n10428 & n36215 ;
  assign n10446 = n10055 | n10445 ;
  assign n36216 = ~n10430 ;
  assign n10447 = n36216 & n10446 ;
  assign n36217 = ~n10447 ;
  assign n10448 = n181 & n36217 ;
  assign n9902 = n9868 | n9886 ;
  assign n36218 = ~n9902 ;
  assign n10026 = n36218 & n157 ;
  assign n10027 = n9705 | n10026 ;
  assign n36219 = ~n9868 ;
  assign n9874 = n9705 & n36219 ;
  assign n9875 = n35935 & n9874 ;
  assign n10030 = n9875 & n157 ;
  assign n36220 = ~n10030 ;
  assign n10031 = n10027 & n36220 ;
  assign n10432 = n181 | n10430 ;
  assign n36221 = ~n10432 ;
  assign n10449 = n36221 & n10446 ;
  assign n10450 = n10031 | n10449 ;
  assign n36222 = ~n10448 ;
  assign n10451 = n36222 & n10450 ;
  assign n36223 = ~n10451 ;
  assign n10452 = n182 & n36223 ;
  assign n9901 = n9871 | n9888 ;
  assign n36224 = ~n9901 ;
  assign n10028 = n36224 & n157 ;
  assign n10029 = n9698 | n10028 ;
  assign n9873 = n9698 & n35945 ;
  assign n36225 = ~n9888 ;
  assign n9900 = n9873 & n36225 ;
  assign n10131 = n9900 & n157 ;
  assign n36226 = ~n10131 ;
  assign n10132 = n10029 & n36226 ;
  assign n10462 = n36205 & n10441 ;
  assign n10463 = n10135 | n10462 ;
  assign n36227 = ~n10443 ;
  assign n10464 = n36227 & n10463 ;
  assign n36228 = ~n10464 ;
  assign n10465 = n180 & n36228 ;
  assign n10466 = n36215 & n10463 ;
  assign n10467 = n10055 | n10466 ;
  assign n36229 = ~n10465 ;
  assign n10468 = n36229 & n10467 ;
  assign n36230 = ~n10468 ;
  assign n10469 = n181 & n36230 ;
  assign n10470 = n182 | n10469 ;
  assign n36231 = ~n10470 ;
  assign n10471 = n10450 & n36231 ;
  assign n10472 = n10132 | n10471 ;
  assign n36232 = ~n10452 ;
  assign n10473 = n36232 & n10472 ;
  assign n36233 = ~n10473 ;
  assign n10474 = n183 & n36233 ;
  assign n9926 = n9892 | n9910 ;
  assign n36234 = ~n9926 ;
  assign n10024 = n36234 & n157 ;
  assign n10025 = n9692 | n10024 ;
  assign n36235 = ~n9892 ;
  assign n9898 = n9692 & n36235 ;
  assign n9899 = n35951 & n9898 ;
  assign n10052 = n9899 & n157 ;
  assign n36236 = ~n10052 ;
  assign n10053 = n10025 & n36236 ;
  assign n10453 = n183 | n10452 ;
  assign n36237 = ~n10453 ;
  assign n10475 = n36237 & n10472 ;
  assign n10476 = n10053 | n10475 ;
  assign n36238 = ~n10474 ;
  assign n10477 = n36238 & n10476 ;
  assign n36239 = ~n10477 ;
  assign n10478 = n838 & n36239 ;
  assign n9897 = n9430 & n35961 ;
  assign n36240 = ~n9912 ;
  assign n9924 = n9897 & n36240 ;
  assign n10068 = n9924 & n157 ;
  assign n9925 = n9895 | n9912 ;
  assign n36241 = ~n9925 ;
  assign n10101 = n36241 & n157 ;
  assign n10102 = n9430 | n10101 ;
  assign n36242 = ~n10068 ;
  assign n10103 = n36242 & n10102 ;
  assign n10486 = n36221 & n10467 ;
  assign n10487 = n10031 | n10486 ;
  assign n36243 = ~n10469 ;
  assign n10488 = n36243 & n10487 ;
  assign n36244 = ~n10488 ;
  assign n10489 = n182 & n36244 ;
  assign n10490 = n36231 & n10487 ;
  assign n10491 = n10132 | n10490 ;
  assign n36245 = ~n10489 ;
  assign n10492 = n36245 & n10491 ;
  assign n36246 = ~n10492 ;
  assign n10493 = n996 & n36246 ;
  assign n10494 = n838 | n10493 ;
  assign n36247 = ~n10494 ;
  assign n10495 = n10476 & n36247 ;
  assign n10496 = n10103 | n10495 ;
  assign n36248 = ~n10478 ;
  assign n10497 = n36248 & n10496 ;
  assign n36249 = ~n10497 ;
  assign n10498 = n185 & n36249 ;
  assign n9950 = n9916 | n9934 ;
  assign n36250 = ~n9950 ;
  assign n10022 = n36250 & n157 ;
  assign n10023 = n9685 | n10022 ;
  assign n36251 = ~n9916 ;
  assign n9922 = n9685 & n36251 ;
  assign n9923 = n35967 & n9922 ;
  assign n10111 = n9923 & n157 ;
  assign n36252 = ~n10111 ;
  assign n10112 = n10023 & n36252 ;
  assign n10479 = n185 | n10478 ;
  assign n36253 = ~n10479 ;
  assign n10499 = n36253 & n10496 ;
  assign n10500 = n10112 | n10499 ;
  assign n36254 = ~n10498 ;
  assign n10501 = n36254 & n10500 ;
  assign n36255 = ~n10501 ;
  assign n10502 = n186 & n36255 ;
  assign n9949 = n9919 | n9936 ;
  assign n36256 = ~n9949 ;
  assign n10020 = n36256 & n157 ;
  assign n10021 = n9678 | n10020 ;
  assign n9921 = n9678 & n35977 ;
  assign n36257 = ~n9936 ;
  assign n9948 = n9921 & n36257 ;
  assign n10036 = n9948 & n157 ;
  assign n36258 = ~n10036 ;
  assign n10037 = n10021 & n36258 ;
  assign n10510 = n36237 & n10491 ;
  assign n10511 = n10053 | n10510 ;
  assign n36259 = ~n10493 ;
  assign n10512 = n36259 & n10511 ;
  assign n36260 = ~n10512 ;
  assign n10513 = n184 & n36260 ;
  assign n10514 = n36247 & n10511 ;
  assign n10515 = n10103 | n10514 ;
  assign n36261 = ~n10513 ;
  assign n10516 = n36261 & n10515 ;
  assign n36262 = ~n10516 ;
  assign n10517 = n185 & n36262 ;
  assign n10518 = n186 | n10517 ;
  assign n36263 = ~n10518 ;
  assign n10519 = n10500 & n36263 ;
  assign n10520 = n10037 | n10519 ;
  assign n36264 = ~n10502 ;
  assign n10521 = n36264 & n10520 ;
  assign n36265 = ~n10521 ;
  assign n10522 = n187 & n36265 ;
  assign n9974 = n9940 | n9958 ;
  assign n36266 = ~n9974 ;
  assign n10061 = n36266 & n157 ;
  assign n10062 = n9672 | n10061 ;
  assign n36267 = ~n9940 ;
  assign n9946 = n9672 & n36267 ;
  assign n9947 = n35983 & n9946 ;
  assign n10090 = n9947 & n157 ;
  assign n36268 = ~n10090 ;
  assign n10091 = n10062 & n36268 ;
  assign n10503 = n528 | n10502 ;
  assign n36269 = ~n10503 ;
  assign n10523 = n36269 & n10520 ;
  assign n10524 = n10091 | n10523 ;
  assign n36270 = ~n10522 ;
  assign n10525 = n36270 & n10524 ;
  assign n36271 = ~n10525 ;
  assign n10526 = n413 & n36271 ;
  assign n9973 = n9943 | n9960 ;
  assign n36272 = ~n9973 ;
  assign n10137 = n36272 & n157 ;
  assign n10138 = n9665 | n10137 ;
  assign n9945 = n9665 & n35993 ;
  assign n36273 = ~n9960 ;
  assign n9972 = n9945 & n36273 ;
  assign n10141 = n9972 & n157 ;
  assign n36274 = ~n10141 ;
  assign n10142 = n10138 & n36274 ;
  assign n10533 = n36253 & n10515 ;
  assign n10534 = n10112 | n10533 ;
  assign n36275 = ~n10517 ;
  assign n10535 = n36275 & n10534 ;
  assign n36276 = ~n10535 ;
  assign n10536 = n186 & n36276 ;
  assign n10537 = n36263 & n10534 ;
  assign n10538 = n10037 | n10537 ;
  assign n36277 = ~n10536 ;
  assign n10539 = n36277 & n10538 ;
  assign n36278 = ~n10539 ;
  assign n10540 = n528 & n36278 ;
  assign n10541 = n413 | n10540 ;
  assign n36279 = ~n10541 ;
  assign n10542 = n10524 & n36279 ;
  assign n10543 = n10142 | n10542 ;
  assign n36280 = ~n10526 ;
  assign n10544 = n36280 & n10543 ;
  assign n36281 = ~n10544 ;
  assign n10545 = n189 & n36281 ;
  assign n9998 = n9964 | n9982 ;
  assign n36282 = ~n9998 ;
  assign n10084 = n36282 & n157 ;
  assign n10085 = n9659 | n10084 ;
  assign n36283 = ~n9964 ;
  assign n9970 = n9659 & n36283 ;
  assign n9971 = n35999 & n9970 ;
  assign n10139 = n9971 & n157 ;
  assign n36284 = ~n10139 ;
  assign n10140 = n10085 & n36284 ;
  assign n10527 = n189 | n10526 ;
  assign n36285 = ~n10527 ;
  assign n10546 = n36285 & n10543 ;
  assign n10547 = n10140 | n10546 ;
  assign n36286 = ~n10545 ;
  assign n10548 = n36286 & n10547 ;
  assign n36287 = ~n10548 ;
  assign n10549 = n190 & n36287 ;
  assign n9969 = n9652 & n36009 ;
  assign n36288 = ~n9984 ;
  assign n9996 = n9969 & n36288 ;
  assign n10092 = n9996 & n157 ;
  assign n9997 = n9967 | n9984 ;
  assign n36289 = ~n9997 ;
  assign n10143 = n36289 & n157 ;
  assign n10144 = n9652 | n10143 ;
  assign n36290 = ~n10092 ;
  assign n10145 = n36290 & n10144 ;
  assign n10556 = n36269 & n10538 ;
  assign n10557 = n10091 | n10556 ;
  assign n36291 = ~n10540 ;
  assign n10558 = n36291 & n10557 ;
  assign n36292 = ~n10558 ;
  assign n10559 = n188 & n36292 ;
  assign n10560 = n36279 & n10557 ;
  assign n10561 = n10142 | n10560 ;
  assign n36293 = ~n10559 ;
  assign n10562 = n36293 & n10561 ;
  assign n36294 = ~n10562 ;
  assign n10563 = n189 & n36294 ;
  assign n10564 = n190 | n10563 ;
  assign n36295 = ~n10564 ;
  assign n10565 = n10547 & n36295 ;
  assign n10566 = n10145 | n10565 ;
  assign n36296 = ~n10549 ;
  assign n10571 = n36296 & n10566 ;
  assign n36297 = ~n10571 ;
  assign n10572 = n191 & n36297 ;
  assign n36298 = ~n9988 ;
  assign n9994 = n9646 & n36298 ;
  assign n9995 = n36015 & n9994 ;
  assign n10078 = n9995 & n157 ;
  assign n10339 = n9988 | n10006 ;
  assign n36299 = ~n10339 ;
  assign n10340 = n157 & n36299 ;
  assign n10341 = n9646 | n10340 ;
  assign n36300 = ~n10078 ;
  assign n10342 = n36300 & n10341 ;
  assign n10550 = n191 | n10549 ;
  assign n36301 = ~n10550 ;
  assign n10582 = n36301 & n10566 ;
  assign n10583 = n10342 | n10582 ;
  assign n36302 = ~n10572 ;
  assign n10584 = n36302 & n10583 ;
  assign n10585 = n10175 | n10584 ;
  assign n10586 = n31336 & n10585 ;
  assign n10014 = n192 & n10013 ;
  assign n36303 = ~n9466 ;
  assign n10150 = n36303 & n157 ;
  assign n36304 = ~n10150 ;
  assign n10151 = n10012 & n36304 ;
  assign n36305 = ~n10151 ;
  assign n10152 = n10014 & n36305 ;
  assign n9627 = n9463 | n9623 ;
  assign n36306 = ~n9627 ;
  assign n9628 = n9465 & n36306 ;
  assign n9629 = n36046 & n9628 ;
  assign n10176 = n9629 & n36047 ;
  assign n10177 = n36048 & n10176 ;
  assign n10178 = n10152 | n10177 ;
  assign n10573 = n10149 & n36302 ;
  assign n10587 = n10573 & n10583 ;
  assign n10588 = n10178 | n10587 ;
  assign n156 = n10586 | n10588 ;
  assign n10551 = n287 | n10549 ;
  assign n36307 = ~n10551 ;
  assign n10567 = n36307 & n10566 ;
  assign n10568 = n10342 | n10567 ;
  assign n10574 = n10568 & n10573 ;
  assign n10579 = n10568 & n36302 ;
  assign n10580 = n10149 | n10579 ;
  assign n10575 = n10178 | n10574 ;
  assign n10655 = n10175 | n10579 ;
  assign n10656 = n31336 & n10655 ;
  assign n10657 = n10575 | n10656 ;
  assign n36308 = ~n10580 ;
  assign n10742 = n36308 & n10657 ;
  assign n10743 = n10574 | n10742 ;
  assign n36309 = ~n10582 ;
  assign n10893 = n10342 & n36309 ;
  assign n10894 = n36302 & n10893 ;
  assign n10895 = n10657 & n10894 ;
  assign n10897 = n10572 | n10582 ;
  assign n36310 = ~n10897 ;
  assign n10898 = n156 & n36310 ;
  assign n10899 = n10342 | n10898 ;
  assign n36311 = ~n10895 ;
  assign n10900 = n36311 & n10899 ;
  assign n10901 = n10743 | n10900 ;
  assign n30758 = x52 | x53 ;
  assign n31330 = x54 | n30758 ;
  assign n9630 = n31330 & n36045 ;
  assign n9631 = n36046 & n9630 ;
  assign n10186 = n9631 & n36047 ;
  assign n10187 = n36048 & n10186 ;
  assign n10683 = x54 & n10657 ;
  assign n36312 = ~n10683 ;
  assign n10684 = n10187 & n36312 ;
  assign n36313 = ~x54 ;
  assign n10679 = n36313 & n10657 ;
  assign n36314 = ~n10679 ;
  assign n10680 = x55 & n36314 ;
  assign n36315 = ~n27977 ;
  assign n10694 = n36315 & n10657 ;
  assign n10695 = n10680 | n10694 ;
  assign n10696 = n10684 | n10695 ;
  assign n193 = n36313 & n30758 ;
  assign n36316 = ~n10657 ;
  assign n10700 = x54 & n36316 ;
  assign n10701 = n193 | n10700 ;
  assign n36317 = ~n10701 ;
  assign n10702 = n157 & n36317 ;
  assign n36318 = ~n10702 ;
  assign n10703 = n10696 & n36318 ;
  assign n36319 = ~n10703 ;
  assign n10704 = n158 & n36319 ;
  assign n10629 = x54 & n156 ;
  assign n36320 = ~n10629 ;
  assign n10630 = n31330 & n36320 ;
  assign n36321 = ~n10630 ;
  assign n10631 = n157 & n36321 ;
  assign n10632 = n158 | n10631 ;
  assign n36322 = ~n10632 ;
  assign n10697 = n36322 & n10696 ;
  assign n36323 = ~n10177 ;
  assign n10179 = n157 & n36323 ;
  assign n36324 = ~n10152 ;
  assign n10180 = n36324 & n10179 ;
  assign n36325 = ~n10574 ;
  assign n10576 = n10180 & n36325 ;
  assign n36326 = ~n10656 ;
  assign n10747 = n10576 & n36326 ;
  assign n10748 = n10694 | n10747 ;
  assign n10749 = x56 & n10748 ;
  assign n10750 = x56 | n10747 ;
  assign n10751 = n10694 | n10750 ;
  assign n36327 = ~n10749 ;
  assign n10752 = n36327 & n10751 ;
  assign n10753 = n10697 | n10752 ;
  assign n36328 = ~n10704 ;
  assign n10754 = n36328 & n10753 ;
  assign n36329 = ~n10754 ;
  assign n10755 = n159 & n36329 ;
  assign n10100 = n10075 | n10098 ;
  assign n36330 = ~n10100 ;
  assign n10173 = n36330 & n10164 ;
  assign n10607 = n10173 & n156 ;
  assign n10626 = n36330 & n156 ;
  assign n10627 = n10164 | n10626 ;
  assign n36331 = ~n10607 ;
  assign n10628 = n36331 & n10627 ;
  assign n10705 = n159 | n10704 ;
  assign n10708 = n158 | n10702 ;
  assign n36332 = ~n10708 ;
  assign n10709 = n10696 & n36332 ;
  assign n10761 = n10709 | n10752 ;
  assign n36333 = ~n10705 ;
  assign n10762 = n36333 & n10761 ;
  assign n10765 = n10628 | n10762 ;
  assign n36334 = ~n10755 ;
  assign n10766 = n36334 & n10765 ;
  assign n36335 = ~n10766 ;
  assign n10767 = n160 & n36335 ;
  assign n10171 = n10169 | n10170 ;
  assign n36336 = ~n10171 ;
  assign n10624 = n36336 & n156 ;
  assign n10625 = n10194 | n10624 ;
  assign n36337 = ~n10170 ;
  assign n10215 = n36337 & n10194 ;
  assign n10216 = n36050 & n10215 ;
  assign n10673 = n10216 & n10657 ;
  assign n36338 = ~n10673 ;
  assign n10674 = n10625 & n36338 ;
  assign n10757 = n8857 & n36329 ;
  assign n10758 = n8534 | n10757 ;
  assign n36339 = ~n10758 ;
  assign n10769 = n36339 & n10765 ;
  assign n10770 = n10674 | n10769 ;
  assign n36340 = ~n10767 ;
  assign n10771 = n36340 & n10770 ;
  assign n36341 = ~n10771 ;
  assign n10772 = n161 & n36341 ;
  assign n10214 = n10197 | n10200 ;
  assign n36342 = ~n10214 ;
  assign n10616 = n36342 & n156 ;
  assign n10617 = n10077 | n10616 ;
  assign n10199 = n10077 & n36055 ;
  assign n36343 = ~n10200 ;
  assign n10213 = n10199 & n36343 ;
  assign n10692 = n10213 & n10657 ;
  assign n36344 = ~n10692 ;
  assign n10693 = n10617 & n36344 ;
  assign n10768 = n161 | n10767 ;
  assign n36345 = ~n10768 ;
  assign n10775 = n36345 & n10770 ;
  assign n10776 = n10693 | n10775 ;
  assign n36346 = ~n10772 ;
  assign n10777 = n36346 & n10776 ;
  assign n36347 = ~n10777 ;
  assign n10778 = n162 & n36347 ;
  assign n10212 = n10203 | n10204 ;
  assign n36348 = ~n10212 ;
  assign n10612 = n36348 & n156 ;
  assign n10613 = n10161 | n10612 ;
  assign n36349 = ~n10204 ;
  assign n10210 = n10161 & n36349 ;
  assign n10211 = n36061 & n10210 ;
  assign n10687 = n10211 & n10657 ;
  assign n36350 = ~n10687 ;
  assign n10688 = n10613 & n36350 ;
  assign n10773 = n162 | n10772 ;
  assign n36351 = ~n10773 ;
  assign n10779 = n36351 & n10776 ;
  assign n10780 = n10688 | n10779 ;
  assign n36352 = ~n10778 ;
  assign n10781 = n36352 & n10780 ;
  assign n36353 = ~n10781 ;
  assign n10782 = n6889 & n36353 ;
  assign n10239 = n10207 | n10225 ;
  assign n36354 = ~n10239 ;
  assign n10614 = n36354 & n156 ;
  assign n10615 = n10155 | n10614 ;
  assign n10208 = n10155 & n36072 ;
  assign n36355 = ~n10225 ;
  assign n10238 = n10208 & n36355 ;
  assign n10671 = n10238 & n10657 ;
  assign n36356 = ~n10671 ;
  assign n10672 = n10615 & n36356 ;
  assign n10785 = n6889 | n10778 ;
  assign n36357 = ~n10785 ;
  assign n10786 = n10780 & n36357 ;
  assign n10787 = n10672 | n10786 ;
  assign n36358 = ~n10782 ;
  assign n10788 = n36358 & n10787 ;
  assign n36359 = ~n10788 ;
  assign n10789 = n164 & n36359 ;
  assign n10237 = n10228 | n10229 ;
  assign n36360 = ~n10237 ;
  assign n10605 = n36360 & n156 ;
  assign n10606 = n10051 | n10605 ;
  assign n36361 = ~n10229 ;
  assign n10235 = n10051 & n36361 ;
  assign n10236 = n36078 & n10235 ;
  assign n10669 = n10236 & n10657 ;
  assign n36362 = ~n10669 ;
  assign n10670 = n10606 & n36362 ;
  assign n10783 = n6600 | n10782 ;
  assign n36363 = ~n10783 ;
  assign n10790 = n36363 & n10787 ;
  assign n10791 = n10670 | n10790 ;
  assign n36364 = ~n10789 ;
  assign n10792 = n36364 & n10791 ;
  assign n36365 = ~n10792 ;
  assign n10793 = n165 & n36365 ;
  assign n10263 = n10232 | n10249 ;
  assign n36366 = ~n10263 ;
  assign n10599 = n36366 & n156 ;
  assign n10600 = n10073 | n10599 ;
  assign n10234 = n10073 & n36088 ;
  assign n36367 = ~n10249 ;
  assign n10262 = n10234 & n36367 ;
  assign n10716 = n10262 & n10657 ;
  assign n36368 = ~n10716 ;
  assign n10717 = n10600 & n36368 ;
  assign n10796 = n163 & n36353 ;
  assign n36369 = ~n10796 ;
  assign n10799 = n10787 & n36369 ;
  assign n36370 = ~n10799 ;
  assign n10800 = n6600 & n36370 ;
  assign n10801 = n165 | n10800 ;
  assign n36371 = ~n10801 ;
  assign n10802 = n10791 & n36371 ;
  assign n10803 = n10717 | n10802 ;
  assign n36372 = ~n10793 ;
  assign n10804 = n36372 & n10803 ;
  assign n36373 = ~n10804 ;
  assign n10805 = n166 & n36373 ;
  assign n10261 = n10252 | n10253 ;
  assign n36374 = ~n10261 ;
  assign n10592 = n36374 & n156 ;
  assign n10593 = n10105 | n10592 ;
  assign n36375 = ~n10253 ;
  assign n10259 = n10105 & n36375 ;
  assign n10260 = n36094 & n10259 ;
  assign n10665 = n10260 & n10657 ;
  assign n36376 = ~n10665 ;
  assign n10666 = n10593 & n36376 ;
  assign n10794 = n166 | n10793 ;
  assign n36377 = ~n10794 ;
  assign n10806 = n36377 & n10803 ;
  assign n10807 = n10666 | n10806 ;
  assign n36378 = ~n10805 ;
  assign n10808 = n36378 & n10807 ;
  assign n36379 = ~n10808 ;
  assign n10809 = n5352 & n36379 ;
  assign n10287 = n10256 | n10273 ;
  assign n36380 = ~n10287 ;
  assign n10622 = n36380 & n156 ;
  assign n10623 = n10107 | n10622 ;
  assign n10258 = n10107 & n36104 ;
  assign n36381 = ~n10273 ;
  assign n10286 = n10258 & n36381 ;
  assign n10661 = n10286 & n10657 ;
  assign n36382 = ~n10661 ;
  assign n10662 = n10623 & n36382 ;
  assign n36383 = ~n10800 ;
  assign n10812 = n10791 & n36383 ;
  assign n36384 = ~n10812 ;
  assign n10813 = n165 & n36384 ;
  assign n36385 = ~n10813 ;
  assign n10814 = n10803 & n36385 ;
  assign n36386 = ~n10814 ;
  assign n10815 = n166 & n36386 ;
  assign n10816 = n5352 | n10815 ;
  assign n36387 = ~n10816 ;
  assign n10817 = n10807 & n36387 ;
  assign n10818 = n10662 | n10817 ;
  assign n36388 = ~n10809 ;
  assign n10819 = n36388 & n10818 ;
  assign n36389 = ~n10819 ;
  assign n10820 = n168 & n36389 ;
  assign n10285 = n10276 | n10277 ;
  assign n36390 = ~n10285 ;
  assign n10601 = n36390 & n156 ;
  assign n10602 = n10110 | n10601 ;
  assign n36391 = ~n10277 ;
  assign n10283 = n10110 & n36391 ;
  assign n10284 = n36110 & n10283 ;
  assign n10685 = n10284 & n10657 ;
  assign n36392 = ~n10685 ;
  assign n10686 = n10602 & n36392 ;
  assign n10810 = n4934 | n10809 ;
  assign n36393 = ~n10810 ;
  assign n10821 = n36393 & n10818 ;
  assign n10822 = n10686 | n10821 ;
  assign n36394 = ~n10820 ;
  assign n10823 = n36394 & n10822 ;
  assign n36395 = ~n10823 ;
  assign n10824 = n169 & n36395 ;
  assign n10311 = n10280 | n10297 ;
  assign n36396 = ~n10311 ;
  assign n10608 = n36396 & n156 ;
  assign n10609 = n10067 | n10608 ;
  assign n10282 = n10067 & n36120 ;
  assign n36397 = ~n10297 ;
  assign n10310 = n10282 & n36397 ;
  assign n10667 = n10310 & n10657 ;
  assign n36398 = ~n10667 ;
  assign n10668 = n10609 & n36398 ;
  assign n36399 = ~n10815 ;
  assign n10827 = n10807 & n36399 ;
  assign n36400 = ~n10827 ;
  assign n10828 = n167 & n36400 ;
  assign n36401 = ~n10828 ;
  assign n10829 = n10818 & n36401 ;
  assign n36402 = ~n10829 ;
  assign n10830 = n4934 & n36402 ;
  assign n10831 = n169 | n10830 ;
  assign n36403 = ~n10831 ;
  assign n10832 = n10822 & n36403 ;
  assign n10833 = n10668 | n10832 ;
  assign n36404 = ~n10824 ;
  assign n10834 = n36404 & n10833 ;
  assign n36405 = ~n10834 ;
  assign n10835 = n170 & n36405 ;
  assign n10309 = n10300 | n10301 ;
  assign n36406 = ~n10309 ;
  assign n10610 = n36406 & n156 ;
  assign n10611 = n10130 | n10610 ;
  assign n36407 = ~n10301 ;
  assign n10307 = n10130 & n36407 ;
  assign n10308 = n36126 & n10307 ;
  assign n10663 = n10308 & n10657 ;
  assign n36408 = ~n10663 ;
  assign n10664 = n10611 & n36408 ;
  assign n10825 = n170 | n10824 ;
  assign n36409 = ~n10825 ;
  assign n10836 = n36409 & n10833 ;
  assign n10837 = n10664 | n10836 ;
  assign n36410 = ~n10835 ;
  assign n10838 = n36410 & n10837 ;
  assign n36411 = ~n10838 ;
  assign n10839 = n3940 & n36411 ;
  assign n10306 = n10089 & n36136 ;
  assign n36412 = ~n10321 ;
  assign n10327 = n10306 & n36412 ;
  assign n10660 = n10327 & n10657 ;
  assign n10328 = n10304 | n10321 ;
  assign n36413 = ~n10328 ;
  assign n10689 = n36413 & n10657 ;
  assign n10690 = n10089 | n10689 ;
  assign n36414 = ~n10660 ;
  assign n10691 = n36414 & n10690 ;
  assign n36415 = ~n10830 ;
  assign n10842 = n10822 & n36415 ;
  assign n36416 = ~n10842 ;
  assign n10843 = n169 & n36416 ;
  assign n36417 = ~n10843 ;
  assign n10844 = n10833 & n36417 ;
  assign n36418 = ~n10844 ;
  assign n10845 = n170 & n36418 ;
  assign n10846 = n3940 | n10845 ;
  assign n36419 = ~n10846 ;
  assign n10847 = n10837 & n36419 ;
  assign n10848 = n10691 | n10847 ;
  assign n36420 = ~n10839 ;
  assign n10849 = n36420 & n10848 ;
  assign n36421 = ~n10849 ;
  assign n10850 = n172 & n36421 ;
  assign n10840 = n3631 | n10839 ;
  assign n36422 = ~n10840 ;
  assign n10851 = n36422 & n10848 ;
  assign n36423 = ~n10325 ;
  assign n10365 = n36423 & n10344 ;
  assign n10366 = n36142 & n10365 ;
  assign n10715 = n10366 & n10657 ;
  assign n10326 = n10324 | n10325 ;
  assign n36424 = ~n10326 ;
  assign n10635 = n36424 & n156 ;
  assign n10912 = n10344 | n10635 ;
  assign n36425 = ~n10715 ;
  assign n10913 = n36425 & n10912 ;
  assign n10914 = n10851 | n10913 ;
  assign n36426 = ~n10850 ;
  assign n10915 = n36426 & n10914 ;
  assign n36427 = ~n10915 ;
  assign n10916 = n173 & n36427 ;
  assign n10364 = n10347 | n10350 ;
  assign n36428 = ~n10364 ;
  assign n10675 = n36428 & n10657 ;
  assign n10676 = n10118 | n10675 ;
  assign n10349 = n10118 & n36152 ;
  assign n36429 = ~n10350 ;
  assign n10363 = n10349 & n36429 ;
  assign n10681 = n10363 & n10657 ;
  assign n36430 = ~n10681 ;
  assign n10682 = n10676 & n36430 ;
  assign n36431 = ~n10845 ;
  assign n10852 = n10837 & n36431 ;
  assign n36432 = ~n10852 ;
  assign n10853 = n171 & n36432 ;
  assign n36433 = ~n10853 ;
  assign n10854 = n10848 & n36433 ;
  assign n36434 = ~n10854 ;
  assign n10855 = n3631 & n36434 ;
  assign n10856 = n173 | n10855 ;
  assign n36435 = ~n10856 ;
  assign n10919 = n36435 & n10914 ;
  assign n10920 = n10682 | n10919 ;
  assign n36436 = ~n10916 ;
  assign n10921 = n36436 & n10920 ;
  assign n36437 = ~n10921 ;
  assign n10922 = n174 & n36437 ;
  assign n10362 = n10353 | n10354 ;
  assign n36438 = ~n10362 ;
  assign n10636 = n36438 & n156 ;
  assign n10637 = n10128 | n10636 ;
  assign n36439 = ~n10354 ;
  assign n10360 = n10128 & n36439 ;
  assign n10361 = n36158 & n10360 ;
  assign n10658 = n10361 & n10657 ;
  assign n36440 = ~n10658 ;
  assign n10659 = n10637 & n36440 ;
  assign n10917 = n174 | n10916 ;
  assign n36441 = ~n10917 ;
  assign n10923 = n36441 & n10920 ;
  assign n10924 = n10659 | n10923 ;
  assign n36442 = ~n10922 ;
  assign n10925 = n36442 & n10924 ;
  assign n36443 = ~n10925 ;
  assign n10926 = n2753 & n36443 ;
  assign n10389 = n10357 | n10375 ;
  assign n36444 = ~n10389 ;
  assign n10642 = n36444 & n156 ;
  assign n10643 = n10115 | n10642 ;
  assign n10359 = n10115 & n36168 ;
  assign n36445 = ~n10375 ;
  assign n10388 = n10359 & n36445 ;
  assign n10713 = n10388 & n10657 ;
  assign n36446 = ~n10713 ;
  assign n10714 = n10643 & n36446 ;
  assign n36447 = ~n10855 ;
  assign n10931 = n36447 & n10914 ;
  assign n36448 = ~n10931 ;
  assign n10932 = n173 & n36448 ;
  assign n36449 = ~n10932 ;
  assign n10933 = n10920 & n36449 ;
  assign n36450 = ~n10933 ;
  assign n10934 = n174 & n36450 ;
  assign n10935 = n2753 | n10934 ;
  assign n36451 = ~n10935 ;
  assign n10936 = n10924 & n36451 ;
  assign n10937 = n10714 | n10936 ;
  assign n36452 = ~n10926 ;
  assign n10938 = n36452 & n10937 ;
  assign n36453 = ~n10938 ;
  assign n10939 = n176 & n36453 ;
  assign n10387 = n10378 | n10379 ;
  assign n36454 = ~n10387 ;
  assign n10618 = n36454 & n156 ;
  assign n10619 = n10045 | n10618 ;
  assign n36455 = ~n10379 ;
  assign n10385 = n10045 & n36455 ;
  assign n10386 = n36174 & n10385 ;
  assign n10728 = n10386 & n10657 ;
  assign n36456 = ~n10728 ;
  assign n10729 = n10619 & n36456 ;
  assign n10927 = n2431 | n10926 ;
  assign n36457 = ~n10927 ;
  assign n10940 = n36457 & n10937 ;
  assign n10941 = n10729 | n10940 ;
  assign n36458 = ~n10939 ;
  assign n10942 = n36458 & n10941 ;
  assign n36459 = ~n10942 ;
  assign n10943 = n177 & n36459 ;
  assign n10413 = n10382 | n10399 ;
  assign n36460 = ~n10413 ;
  assign n10720 = n36460 & n10657 ;
  assign n10721 = n10087 | n10720 ;
  assign n10384 = n10087 & n36184 ;
  assign n36461 = ~n10399 ;
  assign n10412 = n10384 & n36461 ;
  assign n10730 = n10412 & n10657 ;
  assign n36462 = ~n10730 ;
  assign n10731 = n10721 & n36462 ;
  assign n36463 = ~n10934 ;
  assign n10946 = n10924 & n36463 ;
  assign n36464 = ~n10946 ;
  assign n10947 = n175 & n36464 ;
  assign n36465 = ~n10947 ;
  assign n10948 = n10937 & n36465 ;
  assign n36466 = ~n10948 ;
  assign n10949 = n2431 & n36466 ;
  assign n10950 = n177 | n10949 ;
  assign n36467 = ~n10950 ;
  assign n10951 = n10941 & n36467 ;
  assign n10952 = n10731 | n10951 ;
  assign n36468 = ~n10943 ;
  assign n10953 = n36468 & n10952 ;
  assign n36469 = ~n10953 ;
  assign n10954 = n178 & n36469 ;
  assign n10411 = n10402 | n10403 ;
  assign n36470 = ~n10411 ;
  assign n10640 = n36470 & n156 ;
  assign n10641 = n10124 | n10640 ;
  assign n36471 = ~n10403 ;
  assign n10409 = n10124 & n36471 ;
  assign n10410 = n36190 & n10409 ;
  assign n10732 = n10410 & n10657 ;
  assign n36472 = ~n10732 ;
  assign n10733 = n10641 & n36472 ;
  assign n10944 = n178 | n10943 ;
  assign n36473 = ~n10944 ;
  assign n10955 = n36473 & n10952 ;
  assign n10956 = n10733 | n10955 ;
  assign n36474 = ~n10954 ;
  assign n10957 = n36474 & n10956 ;
  assign n36475 = ~n10957 ;
  assign n10958 = n1707 & n36475 ;
  assign n10435 = n10406 | n10423 ;
  assign n36476 = ~n10435 ;
  assign n10646 = n36476 & n156 ;
  assign n10647 = n10121 | n10646 ;
  assign n10408 = n10121 & n36200 ;
  assign n36477 = ~n10423 ;
  assign n10434 = n10408 & n36477 ;
  assign n10711 = n10434 & n10657 ;
  assign n36478 = ~n10711 ;
  assign n10712 = n10647 & n36478 ;
  assign n36479 = ~n10949 ;
  assign n10961 = n10941 & n36479 ;
  assign n36480 = ~n10961 ;
  assign n10962 = n177 & n36480 ;
  assign n36481 = ~n10962 ;
  assign n10965 = n10952 & n36481 ;
  assign n36482 = ~n10965 ;
  assign n10966 = n178 & n36482 ;
  assign n10967 = n1707 | n10966 ;
  assign n36483 = ~n10967 ;
  assign n10968 = n10956 & n36483 ;
  assign n10969 = n10712 | n10968 ;
  assign n36484 = ~n10958 ;
  assign n10970 = n36484 & n10969 ;
  assign n36485 = ~n10970 ;
  assign n10971 = n180 & n36485 ;
  assign n10461 = n10427 | n10443 ;
  assign n36486 = ~n10461 ;
  assign n10597 = n36486 & n156 ;
  assign n10598 = n10135 | n10597 ;
  assign n36487 = ~n10427 ;
  assign n10433 = n10135 & n36487 ;
  assign n10460 = n10433 & n36227 ;
  assign n10734 = n10460 & n10657 ;
  assign n36488 = ~n10734 ;
  assign n10735 = n10598 & n36488 ;
  assign n10959 = n1487 | n10958 ;
  assign n36489 = ~n10959 ;
  assign n10972 = n36489 & n10969 ;
  assign n10973 = n10735 | n10972 ;
  assign n36490 = ~n10971 ;
  assign n10974 = n36490 & n10973 ;
  assign n36491 = ~n10974 ;
  assign n10975 = n181 & n36491 ;
  assign n10459 = n10430 | n10445 ;
  assign n36492 = ~n10459 ;
  assign n10644 = n36492 & n156 ;
  assign n10645 = n10055 | n10644 ;
  assign n10431 = n10055 & n36216 ;
  assign n36493 = ~n10445 ;
  assign n10458 = n10431 & n36493 ;
  assign n10736 = n10458 & n10657 ;
  assign n36494 = ~n10736 ;
  assign n10737 = n10645 & n36494 ;
  assign n36495 = ~n10966 ;
  assign n10978 = n10956 & n36495 ;
  assign n36496 = ~n10978 ;
  assign n10979 = n179 & n36496 ;
  assign n36497 = ~n10979 ;
  assign n10980 = n10969 & n36497 ;
  assign n36498 = ~n10980 ;
  assign n10981 = n1487 & n36498 ;
  assign n10982 = n181 | n10981 ;
  assign n36499 = ~n10982 ;
  assign n10983 = n10973 & n36499 ;
  assign n10984 = n10737 | n10983 ;
  assign n36500 = ~n10975 ;
  assign n10985 = n36500 & n10984 ;
  assign n36501 = ~n10985 ;
  assign n10986 = n182 & n36501 ;
  assign n10457 = n10448 | n10449 ;
  assign n36502 = ~n10457 ;
  assign n10648 = n36502 & n156 ;
  assign n10649 = n10031 | n10648 ;
  assign n36503 = ~n10449 ;
  assign n10455 = n10031 & n36503 ;
  assign n10456 = n36222 & n10455 ;
  assign n10738 = n10456 & n10657 ;
  assign n36504 = ~n10738 ;
  assign n10739 = n10649 & n36504 ;
  assign n10976 = n182 | n10975 ;
  assign n36505 = ~n10976 ;
  assign n10987 = n36505 & n10984 ;
  assign n10988 = n10739 | n10987 ;
  assign n36506 = ~n10986 ;
  assign n10989 = n36506 & n10988 ;
  assign n36507 = ~n10989 ;
  assign n10990 = n996 & n36507 ;
  assign n10485 = n10452 | n10471 ;
  assign n36508 = ~n10485 ;
  assign n10650 = n36508 & n156 ;
  assign n10651 = n10132 | n10650 ;
  assign n10454 = n10132 & n36232 ;
  assign n36509 = ~n10471 ;
  assign n10484 = n10454 & n36509 ;
  assign n10740 = n10484 & n10657 ;
  assign n36510 = ~n10740 ;
  assign n10741 = n10651 & n36510 ;
  assign n36511 = ~n10981 ;
  assign n10993 = n10973 & n36511 ;
  assign n36512 = ~n10993 ;
  assign n10994 = n181 & n36512 ;
  assign n36513 = ~n10994 ;
  assign n10995 = n10984 & n36513 ;
  assign n36514 = ~n10995 ;
  assign n10996 = n182 & n36514 ;
  assign n10997 = n183 | n10996 ;
  assign n36515 = ~n10997 ;
  assign n10998 = n10988 & n36515 ;
  assign n10999 = n10741 | n10998 ;
  assign n36516 = ~n10990 ;
  assign n11000 = n36516 & n10999 ;
  assign n36517 = ~n11000 ;
  assign n11001 = n184 & n36517 ;
  assign n10483 = n10474 | n10475 ;
  assign n36518 = ~n10483 ;
  assign n10638 = n36518 & n156 ;
  assign n10639 = n10053 | n10638 ;
  assign n36519 = ~n10475 ;
  assign n10481 = n10053 & n36519 ;
  assign n10482 = n36238 & n10481 ;
  assign n10698 = n10482 & n10657 ;
  assign n36520 = ~n10698 ;
  assign n10699 = n10639 & n36520 ;
  assign n10991 = n838 | n10990 ;
  assign n36521 = ~n10991 ;
  assign n11002 = n36521 & n10999 ;
  assign n11003 = n10699 | n11002 ;
  assign n36522 = ~n11001 ;
  assign n11004 = n36522 & n11003 ;
  assign n36523 = ~n11004 ;
  assign n11005 = n185 & n36523 ;
  assign n10509 = n10478 | n10495 ;
  assign n36524 = ~n10509 ;
  assign n10620 = n36524 & n156 ;
  assign n10621 = n10103 | n10620 ;
  assign n10480 = n10103 & n36248 ;
  assign n36525 = ~n10495 ;
  assign n10508 = n10480 & n36525 ;
  assign n10726 = n10508 & n10657 ;
  assign n36526 = ~n10726 ;
  assign n10727 = n10621 & n36526 ;
  assign n36527 = ~n10996 ;
  assign n11008 = n10988 & n36527 ;
  assign n36528 = ~n11008 ;
  assign n11009 = n183 & n36528 ;
  assign n36529 = ~n11009 ;
  assign n11010 = n10999 & n36529 ;
  assign n36530 = ~n11010 ;
  assign n11011 = n838 & n36530 ;
  assign n11012 = n185 | n11011 ;
  assign n36531 = ~n11012 ;
  assign n11013 = n11003 & n36531 ;
  assign n11014 = n10727 | n11013 ;
  assign n36532 = ~n11005 ;
  assign n11015 = n36532 & n11014 ;
  assign n36533 = ~n11015 ;
  assign n11016 = n186 & n36533 ;
  assign n10507 = n10498 | n10499 ;
  assign n36534 = ~n10507 ;
  assign n10590 = n36534 & n156 ;
  assign n10591 = n10112 | n10590 ;
  assign n36535 = ~n10499 ;
  assign n10505 = n10112 & n36535 ;
  assign n10506 = n36254 & n10505 ;
  assign n10677 = n10506 & n10657 ;
  assign n36536 = ~n10677 ;
  assign n10678 = n10591 & n36536 ;
  assign n11006 = n186 | n11005 ;
  assign n36537 = ~n11006 ;
  assign n11017 = n36537 & n11014 ;
  assign n11018 = n10678 | n11017 ;
  assign n36538 = ~n11016 ;
  assign n11019 = n36538 & n11018 ;
  assign n36539 = ~n11019 ;
  assign n11020 = n528 & n36539 ;
  assign n10532 = n10502 | n10519 ;
  assign n36540 = ~n10532 ;
  assign n10633 = n36540 & n156 ;
  assign n10634 = n10037 | n10633 ;
  assign n10504 = n10037 & n36264 ;
  assign n36541 = ~n10519 ;
  assign n10531 = n10504 & n36541 ;
  assign n10724 = n10531 & n10657 ;
  assign n36542 = ~n10724 ;
  assign n10725 = n10634 & n36542 ;
  assign n36543 = ~n11011 ;
  assign n11023 = n11003 & n36543 ;
  assign n36544 = ~n11023 ;
  assign n11024 = n185 & n36544 ;
  assign n36545 = ~n11024 ;
  assign n11025 = n11014 & n36545 ;
  assign n36546 = ~n11025 ;
  assign n11026 = n186 & n36546 ;
  assign n11027 = n528 | n11026 ;
  assign n36547 = ~n11027 ;
  assign n11028 = n11018 & n36547 ;
  assign n11029 = n10725 | n11028 ;
  assign n36548 = ~n11020 ;
  assign n11030 = n36548 & n11029 ;
  assign n36549 = ~n11030 ;
  assign n11031 = n188 & n36549 ;
  assign n36550 = ~n10523 ;
  assign n10529 = n10091 & n36550 ;
  assign n10530 = n36270 & n10529 ;
  assign n10596 = n10530 & n156 ;
  assign n10555 = n10523 | n10540 ;
  assign n36551 = ~n10555 ;
  assign n10652 = n36551 & n156 ;
  assign n10653 = n10091 | n10652 ;
  assign n36552 = ~n10596 ;
  assign n10654 = n36552 & n10653 ;
  assign n11021 = n413 | n11020 ;
  assign n36553 = ~n11021 ;
  assign n11032 = n36553 & n11029 ;
  assign n11033 = n10654 | n11032 ;
  assign n36554 = ~n11031 ;
  assign n11034 = n36554 & n11033 ;
  assign n36555 = ~n11034 ;
  assign n11035 = n189 & n36555 ;
  assign n10554 = n10526 | n10542 ;
  assign n36556 = ~n10554 ;
  assign n10603 = n36556 & n156 ;
  assign n10604 = n10142 | n10603 ;
  assign n10528 = n10142 & n36280 ;
  assign n36557 = ~n10542 ;
  assign n10553 = n10528 & n36557 ;
  assign n10722 = n10553 & n10657 ;
  assign n36558 = ~n10722 ;
  assign n10723 = n10604 & n36558 ;
  assign n36559 = ~n11026 ;
  assign n11038 = n11018 & n36559 ;
  assign n36560 = ~n11038 ;
  assign n11039 = n187 & n36560 ;
  assign n36561 = ~n11039 ;
  assign n11042 = n11029 & n36561 ;
  assign n36562 = ~n11042 ;
  assign n11043 = n413 & n36562 ;
  assign n11044 = n189 | n11043 ;
  assign n36563 = ~n11044 ;
  assign n11045 = n11033 & n36563 ;
  assign n11046 = n10723 | n11045 ;
  assign n36564 = ~n11035 ;
  assign n11047 = n36564 & n11046 ;
  assign n36565 = ~n11047 ;
  assign n11048 = n190 & n36565 ;
  assign n10904 = n36285 & n10561 ;
  assign n36566 = ~n10904 ;
  assign n10905 = n10140 & n36566 ;
  assign n10906 = n36286 & n10905 ;
  assign n10907 = n10657 & n10906 ;
  assign n10908 = n10545 | n10904 ;
  assign n36567 = ~n10908 ;
  assign n10909 = n156 & n36567 ;
  assign n10910 = n10140 | n10909 ;
  assign n36568 = ~n10907 ;
  assign n10911 = n36568 & n10910 ;
  assign n11036 = n190 | n11035 ;
  assign n36569 = ~n11036 ;
  assign n11049 = n36569 & n11046 ;
  assign n11050 = n10911 | n11049 ;
  assign n36570 = ~n11048 ;
  assign n11051 = n36570 & n11050 ;
  assign n36571 = ~n11051 ;
  assign n11052 = n287 & n36571 ;
  assign n10569 = n10549 | n10565 ;
  assign n36572 = ~n10569 ;
  assign n10594 = n36572 & n156 ;
  assign n10595 = n10145 | n10594 ;
  assign n10552 = n10145 & n36296 ;
  assign n36573 = ~n10565 ;
  assign n10570 = n10552 & n36573 ;
  assign n10718 = n10570 & n10657 ;
  assign n36574 = ~n10718 ;
  assign n10719 = n10595 & n36574 ;
  assign n36575 = ~n11043 ;
  assign n11055 = n11033 & n36575 ;
  assign n36576 = ~n11055 ;
  assign n11056 = n189 & n36576 ;
  assign n36577 = ~n11056 ;
  assign n11057 = n11046 & n36577 ;
  assign n36578 = ~n11057 ;
  assign n11058 = n190 & n36578 ;
  assign n11059 = n287 | n11058 ;
  assign n36579 = ~n11059 ;
  assign n11060 = n11050 & n36579 ;
  assign n11061 = n10719 | n11060 ;
  assign n36580 = ~n11052 ;
  assign n11062 = n36580 & n11061 ;
  assign n11063 = n10901 | n11062 ;
  assign n11064 = n31336 & n11063 ;
  assign n10581 = n192 & n10580 ;
  assign n36581 = ~n10149 ;
  assign n10744 = n36581 & n10657 ;
  assign n36582 = ~n10744 ;
  assign n10745 = n10579 & n36582 ;
  assign n36583 = ~n10745 ;
  assign n10746 = n10581 & n36583 ;
  assign n10183 = n10146 | n10177 ;
  assign n36584 = ~n10183 ;
  assign n10184 = n10148 & n36584 ;
  assign n10185 = n36324 & n10184 ;
  assign n10577 = n10185 & n36325 ;
  assign n10886 = n10577 & n36326 ;
  assign n10887 = n10746 | n10886 ;
  assign n11053 = n10900 & n36580 ;
  assign n11065 = n11053 & n11061 ;
  assign n11066 = n10887 | n11065 ;
  assign n11067 = n11064 | n11066 ;
  assign n11126 = n10900 | n11062 ;
  assign n36585 = ~n11126 ;
  assign n11127 = n11067 & n36585 ;
  assign n11128 = n11065 | n11127 ;
  assign n11054 = n10719 & n36580 ;
  assign n11130 = n191 | n11058 ;
  assign n36586 = ~n11130 ;
  assign n11131 = n11050 & n36586 ;
  assign n36587 = ~n11131 ;
  assign n11132 = n11054 & n36587 ;
  assign n11133 = n11067 & n11132 ;
  assign n11135 = n11052 | n11131 ;
  assign n36588 = ~n11058 ;
  assign n11136 = n11050 & n36588 ;
  assign n36589 = ~n11136 ;
  assign n11137 = n191 & n36589 ;
  assign n11138 = n10719 | n11131 ;
  assign n36590 = ~n11137 ;
  assign n11139 = n36590 & n11138 ;
  assign n11140 = n10901 | n11139 ;
  assign n11141 = n31336 & n11140 ;
  assign n11142 = n11053 & n11138 ;
  assign n11143 = n10887 | n11142 ;
  assign n155 = n11141 | n11143 ;
  assign n36591 = ~n11135 ;
  assign n11148 = n36591 & n155 ;
  assign n11149 = n10719 | n11148 ;
  assign n36592 = ~n11133 ;
  assign n11150 = n36592 & n11149 ;
  assign n11151 = n11128 | n11150 ;
  assign n11376 = n11032 | n11043 ;
  assign n36593 = ~n11376 ;
  assign n11377 = n155 & n36593 ;
  assign n11378 = n10654 | n11377 ;
  assign n36594 = ~n11032 ;
  assign n11379 = n10654 & n36594 ;
  assign n11380 = n36575 & n11379 ;
  assign n11381 = n11067 & n11380 ;
  assign n36595 = ~n11381 ;
  assign n11382 = n11378 & n36595 ;
  assign n10841 = n10691 & n36420 ;
  assign n36596 = ~n10847 ;
  assign n10858 = n10841 & n36596 ;
  assign n11073 = n10858 & n11067 ;
  assign n10859 = n10839 | n10847 ;
  assign n36597 = ~n10859 ;
  assign n11160 = n36597 & n155 ;
  assign n11161 = n10691 | n11160 ;
  assign n36598 = ~n11073 ;
  assign n11162 = n36598 & n11161 ;
  assign n194 = x50 | x51 ;
  assign n36599 = ~x52 ;
  assign n196 = n36599 & n194 ;
  assign n36600 = ~n11067 ;
  assign n11069 = x52 & n36600 ;
  assign n11070 = n196 | n11069 ;
  assign n36601 = ~n11070 ;
  assign n11071 = n10657 & n36601 ;
  assign n195 = x52 | n194 ;
  assign n10181 = n195 & n36323 ;
  assign n10182 = n36324 & n10181 ;
  assign n10578 = n10182 & n36325 ;
  assign n10892 = n10578 & n36326 ;
  assign n11085 = x52 & n11067 ;
  assign n36602 = ~n11085 ;
  assign n11086 = n10892 & n36602 ;
  assign n36603 = ~n30758 ;
  assign n11083 = n36603 & n11067 ;
  assign n11090 = n36599 & n11067 ;
  assign n36604 = ~n11090 ;
  assign n11091 = x53 & n36604 ;
  assign n11092 = n11083 | n11091 ;
  assign n11094 = n11086 | n11092 ;
  assign n36605 = ~n11071 ;
  assign n11095 = n36605 & n11094 ;
  assign n36606 = ~n11095 ;
  assign n11096 = n157 & n36606 ;
  assign n36607 = ~n10886 ;
  assign n10888 = n10657 & n36607 ;
  assign n36608 = ~n10746 ;
  assign n10889 = n36608 & n10888 ;
  assign n36609 = ~n11065 ;
  assign n11109 = n10889 & n36609 ;
  assign n36610 = ~n11064 ;
  assign n11110 = n36610 & n11109 ;
  assign n11111 = n11083 | n11110 ;
  assign n11112 = x54 & n11111 ;
  assign n11113 = x54 | n11110 ;
  assign n11114 = n11083 | n11113 ;
  assign n36611 = ~n11112 ;
  assign n11115 = n36611 & n11114 ;
  assign n11184 = x52 & n155 ;
  assign n36612 = ~n11184 ;
  assign n11185 = n195 & n36612 ;
  assign n36613 = ~n11185 ;
  assign n11186 = n156 & n36613 ;
  assign n11187 = n157 | n11186 ;
  assign n36614 = ~n11187 ;
  assign n11188 = n11094 & n36614 ;
  assign n11189 = n11115 | n11188 ;
  assign n36615 = ~n11096 ;
  assign n11190 = n36615 & n11189 ;
  assign n36616 = ~n11190 ;
  assign n11191 = n158 & n36616 ;
  assign n11097 = n158 | n11096 ;
  assign n11072 = n157 | n11071 ;
  assign n36617 = ~n11072 ;
  assign n11098 = n36617 & n11094 ;
  assign n11118 = n11098 | n11115 ;
  assign n36618 = ~n11097 ;
  assign n11119 = n36618 & n11118 ;
  assign n10706 = n10684 | n10702 ;
  assign n36619 = ~n10706 ;
  assign n10707 = n10695 & n36619 ;
  assign n11082 = n10707 & n11067 ;
  assign n11197 = n36619 & n155 ;
  assign n11198 = n10695 | n11197 ;
  assign n36620 = ~n11082 ;
  assign n11199 = n36620 & n11198 ;
  assign n11200 = n11119 | n11199 ;
  assign n36621 = ~n11191 ;
  assign n11201 = n36621 & n11200 ;
  assign n36622 = ~n11201 ;
  assign n11202 = n8857 & n36622 ;
  assign n36623 = ~n10709 ;
  assign n10759 = n36623 & n10752 ;
  assign n10760 = n36328 & n10759 ;
  assign n11106 = n10760 & n11067 ;
  assign n10710 = n10704 | n10709 ;
  assign n36624 = ~n10710 ;
  assign n11194 = n36624 & n155 ;
  assign n11195 = n10752 | n11194 ;
  assign n36625 = ~n11106 ;
  assign n11196 = n36625 & n11195 ;
  assign n11193 = n8857 | n11191 ;
  assign n36626 = ~n11193 ;
  assign n11204 = n36626 & n11200 ;
  assign n11205 = n11196 | n11204 ;
  assign n36627 = ~n11202 ;
  assign n11206 = n36627 & n11205 ;
  assign n36628 = ~n11206 ;
  assign n11207 = n160 & n36628 ;
  assign n10756 = n10628 & n36334 ;
  assign n36629 = ~n10762 ;
  assign n10763 = n10756 & n36629 ;
  assign n11088 = n10763 & n11067 ;
  assign n10764 = n10755 | n10762 ;
  assign n36630 = ~n10764 ;
  assign n11175 = n36630 & n155 ;
  assign n11176 = n10628 | n11175 ;
  assign n36631 = ~n11088 ;
  assign n11177 = n36631 & n11176 ;
  assign n11203 = n160 | n11202 ;
  assign n36632 = ~n11203 ;
  assign n11208 = n36632 & n11205 ;
  assign n11209 = n11177 | n11208 ;
  assign n36633 = ~n11207 ;
  assign n11210 = n36633 & n11209 ;
  assign n36634 = ~n11210 ;
  assign n11211 = n161 & n36634 ;
  assign n36635 = ~n10769 ;
  assign n10883 = n10674 & n36635 ;
  assign n10884 = n36340 & n10883 ;
  assign n11075 = n10884 & n11067 ;
  assign n10885 = n10767 | n10769 ;
  assign n36636 = ~n10885 ;
  assign n11169 = n36636 & n155 ;
  assign n11170 = n10674 | n11169 ;
  assign n36637 = ~n11075 ;
  assign n11171 = n36637 & n11170 ;
  assign n11219 = n159 & n36622 ;
  assign n36638 = ~n11219 ;
  assign n11220 = n11205 & n36638 ;
  assign n36639 = ~n11220 ;
  assign n11221 = n8534 & n36639 ;
  assign n11222 = n161 | n11221 ;
  assign n36640 = ~n11222 ;
  assign n11223 = n11209 & n36640 ;
  assign n11224 = n11171 | n11223 ;
  assign n36641 = ~n11211 ;
  assign n11225 = n36641 & n11224 ;
  assign n36642 = ~n11225 ;
  assign n11226 = n162 & n36642 ;
  assign n10882 = n10772 | n10775 ;
  assign n36643 = ~n10882 ;
  assign n11080 = n36643 & n11067 ;
  assign n11081 = n10693 | n11080 ;
  assign n10774 = n10693 & n36346 ;
  assign n36644 = ~n10775 ;
  assign n10881 = n10774 & n36644 ;
  assign n11104 = n10881 & n11067 ;
  assign n36645 = ~n11104 ;
  assign n11105 = n11081 & n36645 ;
  assign n11212 = n162 | n11211 ;
  assign n36646 = ~n11212 ;
  assign n11227 = n36646 & n11224 ;
  assign n11228 = n11105 | n11227 ;
  assign n36647 = ~n11226 ;
  assign n11229 = n36647 & n11228 ;
  assign n36648 = ~n11229 ;
  assign n11230 = n6889 & n36648 ;
  assign n36649 = ~n10779 ;
  assign n10878 = n10688 & n36649 ;
  assign n10879 = n36352 & n10878 ;
  assign n11089 = n10879 & n11067 ;
  assign n10880 = n10778 | n10779 ;
  assign n36650 = ~n10880 ;
  assign n11172 = n36650 & n155 ;
  assign n11173 = n10688 | n11172 ;
  assign n36651 = ~n11089 ;
  assign n11174 = n36651 & n11173 ;
  assign n36652 = ~n11221 ;
  assign n11238 = n11209 & n36652 ;
  assign n36653 = ~n11238 ;
  assign n11239 = n161 & n36653 ;
  assign n36654 = ~n11239 ;
  assign n11240 = n11224 & n36654 ;
  assign n36655 = ~n11240 ;
  assign n11241 = n162 & n36655 ;
  assign n11242 = n6889 | n11241 ;
  assign n36656 = ~n11242 ;
  assign n11243 = n11228 & n36656 ;
  assign n11244 = n11174 | n11243 ;
  assign n36657 = ~n11230 ;
  assign n11245 = n36657 & n11244 ;
  assign n36658 = ~n11245 ;
  assign n11246 = n164 & n36658 ;
  assign n10798 = n10782 | n10786 ;
  assign n36659 = ~n10798 ;
  assign n11078 = n36659 & n11067 ;
  assign n11079 = n10672 | n11078 ;
  assign n10784 = n10672 & n36358 ;
  assign n36660 = ~n10786 ;
  assign n10797 = n10784 & n36660 ;
  assign n11101 = n10797 & n11067 ;
  assign n36661 = ~n11101 ;
  assign n11102 = n11079 & n36661 ;
  assign n11231 = n6600 | n11230 ;
  assign n36662 = ~n11231 ;
  assign n11247 = n36662 & n11244 ;
  assign n11248 = n11102 | n11247 ;
  assign n36663 = ~n11246 ;
  assign n11249 = n36663 & n11248 ;
  assign n36664 = ~n11249 ;
  assign n11250 = n165 & n36664 ;
  assign n36665 = ~n10790 ;
  assign n10875 = n10670 & n36665 ;
  assign n10876 = n36383 & n10875 ;
  assign n11103 = n10876 & n11067 ;
  assign n10877 = n10790 | n10800 ;
  assign n36666 = ~n10877 ;
  assign n11166 = n36666 & n155 ;
  assign n11167 = n10670 | n11166 ;
  assign n36667 = ~n11103 ;
  assign n11168 = n36667 & n11167 ;
  assign n36668 = ~n11241 ;
  assign n11258 = n11228 & n36668 ;
  assign n36669 = ~n11258 ;
  assign n11259 = n163 & n36669 ;
  assign n36670 = ~n11259 ;
  assign n11260 = n11244 & n36670 ;
  assign n36671 = ~n11260 ;
  assign n11261 = n6600 & n36671 ;
  assign n11262 = n165 | n11261 ;
  assign n36672 = ~n11262 ;
  assign n11263 = n11248 & n36672 ;
  assign n11264 = n11168 | n11263 ;
  assign n36673 = ~n11250 ;
  assign n11265 = n36673 & n11264 ;
  assign n36674 = ~n11265 ;
  assign n11266 = n166 & n36674 ;
  assign n10795 = n10717 & n36372 ;
  assign n36675 = ~n10802 ;
  assign n10873 = n10795 & n36675 ;
  assign n11159 = n10873 & n155 ;
  assign n10874 = n10802 | n10813 ;
  assign n36676 = ~n10874 ;
  assign n11181 = n36676 & n155 ;
  assign n11182 = n10717 | n11181 ;
  assign n36677 = ~n11159 ;
  assign n11183 = n36677 & n11182 ;
  assign n11251 = n166 | n11250 ;
  assign n36678 = ~n11251 ;
  assign n11267 = n36678 & n11264 ;
  assign n11268 = n11183 | n11267 ;
  assign n36679 = ~n11266 ;
  assign n11269 = n36679 & n11268 ;
  assign n36680 = ~n11269 ;
  assign n11270 = n5352 & n36680 ;
  assign n36681 = ~n10806 ;
  assign n10871 = n10666 & n36681 ;
  assign n10872 = n36399 & n10871 ;
  assign n11077 = n10872 & n11067 ;
  assign n10870 = n10806 | n10815 ;
  assign n36682 = ~n10870 ;
  assign n11178 = n36682 & n155 ;
  assign n11179 = n10666 | n11178 ;
  assign n36683 = ~n11077 ;
  assign n11180 = n36683 & n11179 ;
  assign n36684 = ~n11261 ;
  assign n11278 = n11248 & n36684 ;
  assign n36685 = ~n11278 ;
  assign n11279 = n165 & n36685 ;
  assign n36686 = ~n11279 ;
  assign n11280 = n11264 & n36686 ;
  assign n36687 = ~n11280 ;
  assign n11281 = n166 & n36687 ;
  assign n11282 = n5352 | n11281 ;
  assign n36688 = ~n11282 ;
  assign n11283 = n11268 & n36688 ;
  assign n11284 = n11180 | n11283 ;
  assign n36689 = ~n11270 ;
  assign n11285 = n36689 & n11284 ;
  assign n36690 = ~n11285 ;
  assign n11286 = n168 & n36690 ;
  assign n11271 = n4934 | n11270 ;
  assign n36691 = ~n11271 ;
  assign n11287 = n36691 & n11284 ;
  assign n10811 = n10662 & n36388 ;
  assign n36692 = ~n10817 ;
  assign n10868 = n10811 & n36692 ;
  assign n11076 = n10868 & n11067 ;
  assign n10869 = n10817 | n10828 ;
  assign n36693 = ~n10869 ;
  assign n11310 = n36693 & n155 ;
  assign n11311 = n10662 | n11310 ;
  assign n36694 = ~n11076 ;
  assign n11312 = n36694 & n11311 ;
  assign n11313 = n11287 | n11312 ;
  assign n36695 = ~n11286 ;
  assign n11314 = n36695 & n11313 ;
  assign n36696 = ~n11314 ;
  assign n11315 = n169 & n36696 ;
  assign n36697 = ~n10821 ;
  assign n10865 = n10686 & n36697 ;
  assign n10866 = n36415 & n10865 ;
  assign n11074 = n10866 & n11067 ;
  assign n10867 = n10821 | n10830 ;
  assign n36698 = ~n10867 ;
  assign n11145 = n36698 & n155 ;
  assign n11146 = n10686 | n11145 ;
  assign n36699 = ~n11074 ;
  assign n11147 = n36699 & n11146 ;
  assign n36700 = ~n11281 ;
  assign n11294 = n11268 & n36700 ;
  assign n36701 = ~n11294 ;
  assign n11295 = n167 & n36701 ;
  assign n36702 = ~n11295 ;
  assign n11296 = n11284 & n36702 ;
  assign n36703 = ~n11296 ;
  assign n11297 = n4934 & n36703 ;
  assign n11298 = n169 | n11297 ;
  assign n36704 = ~n11298 ;
  assign n11317 = n36704 & n11313 ;
  assign n11318 = n11147 | n11317 ;
  assign n36705 = ~n11315 ;
  assign n11319 = n36705 & n11318 ;
  assign n36706 = ~n11319 ;
  assign n11320 = n170 & n36706 ;
  assign n10826 = n10668 & n36404 ;
  assign n36707 = ~n10832 ;
  assign n10863 = n10826 & n36707 ;
  assign n11084 = n10863 & n11067 ;
  assign n10864 = n10832 | n10843 ;
  assign n36708 = ~n10864 ;
  assign n11163 = n36708 & n155 ;
  assign n11164 = n10668 | n11163 ;
  assign n36709 = ~n11084 ;
  assign n11165 = n36709 & n11164 ;
  assign n11316 = n170 | n11315 ;
  assign n36710 = ~n11316 ;
  assign n11321 = n36710 & n11318 ;
  assign n11322 = n11165 | n11321 ;
  assign n36711 = ~n11320 ;
  assign n11323 = n36711 & n11322 ;
  assign n36712 = ~n11323 ;
  assign n11324 = n3940 & n36712 ;
  assign n11325 = n3631 | n11324 ;
  assign n36713 = ~n10836 ;
  assign n10860 = n10664 & n36713 ;
  assign n10861 = n36431 & n10860 ;
  assign n11100 = n10861 & n11067 ;
  assign n10862 = n10836 | n10845 ;
  assign n36714 = ~n10862 ;
  assign n11299 = n36714 & n155 ;
  assign n11300 = n10664 | n11299 ;
  assign n36715 = ~n11100 ;
  assign n11301 = n36715 & n11300 ;
  assign n36716 = ~n11297 ;
  assign n11332 = n36716 & n11313 ;
  assign n36717 = ~n11332 ;
  assign n11333 = n169 & n36717 ;
  assign n36718 = ~n11333 ;
  assign n11334 = n11318 & n36718 ;
  assign n36719 = ~n11334 ;
  assign n11335 = n170 & n36719 ;
  assign n11336 = n3940 | n11335 ;
  assign n36720 = ~n11336 ;
  assign n11337 = n11322 & n36720 ;
  assign n11338 = n11301 | n11337 ;
  assign n36721 = ~n11325 ;
  assign n11341 = n36721 & n11338 ;
  assign n11342 = n11162 | n11341 ;
  assign n36722 = ~n11335 ;
  assign n11352 = n11322 & n36722 ;
  assign n36723 = ~n11352 ;
  assign n11353 = n171 & n36723 ;
  assign n36724 = ~n11353 ;
  assign n11354 = n11338 & n36724 ;
  assign n36725 = ~n11354 ;
  assign n11355 = n3631 & n36725 ;
  assign n36726 = ~n11355 ;
  assign n11361 = n11342 & n36726 ;
  assign n36727 = ~n11361 ;
  assign n11362 = n173 & n36727 ;
  assign n11356 = n173 | n11355 ;
  assign n36728 = ~n11356 ;
  assign n11357 = n11342 & n36728 ;
  assign n36729 = ~n10851 ;
  assign n10929 = n36729 & n10913 ;
  assign n10930 = n36447 & n10929 ;
  assign n11068 = n10930 & n11067 ;
  assign n10857 = n10851 | n10855 ;
  assign n36730 = ~n10857 ;
  assign n11309 = n36730 & n155 ;
  assign n11468 = n10913 | n11309 ;
  assign n36731 = ~n11068 ;
  assign n11469 = n36731 & n11468 ;
  assign n11470 = n11357 | n11469 ;
  assign n36732 = ~n11362 ;
  assign n11471 = n36732 & n11470 ;
  assign n36733 = ~n11471 ;
  assign n11472 = n174 & n36733 ;
  assign n10918 = n10682 & n36436 ;
  assign n36734 = ~n10919 ;
  assign n11462 = n10918 & n36734 ;
  assign n11463 = n11067 & n11462 ;
  assign n11464 = n10916 | n10919 ;
  assign n36735 = ~n11464 ;
  assign n11465 = n155 & n36735 ;
  assign n11466 = n10682 | n11465 ;
  assign n36736 = ~n11463 ;
  assign n11467 = n36736 & n11466 ;
  assign n36737 = ~n11324 ;
  assign n11339 = n36737 & n11338 ;
  assign n36738 = ~n11339 ;
  assign n11340 = n172 & n36738 ;
  assign n36739 = ~n11340 ;
  assign n11343 = n36739 & n11342 ;
  assign n36740 = ~n11343 ;
  assign n11344 = n173 & n36740 ;
  assign n11345 = n174 | n11344 ;
  assign n36741 = ~n11345 ;
  assign n11475 = n36741 & n11470 ;
  assign n11476 = n11467 | n11475 ;
  assign n36742 = ~n11472 ;
  assign n11477 = n36742 & n11476 ;
  assign n36743 = ~n11477 ;
  assign n11478 = n175 & n36743 ;
  assign n36744 = ~n10923 ;
  assign n11455 = n10659 & n36744 ;
  assign n11456 = n36463 & n11455 ;
  assign n11457 = n11067 & n11456 ;
  assign n11458 = n10923 | n10934 ;
  assign n36745 = ~n11458 ;
  assign n11459 = n155 & n36745 ;
  assign n11460 = n10659 | n11459 ;
  assign n36746 = ~n11457 ;
  assign n11461 = n36746 & n11460 ;
  assign n11473 = n2753 | n11472 ;
  assign n36747 = ~n11473 ;
  assign n11479 = n36747 & n11476 ;
  assign n11480 = n11461 | n11479 ;
  assign n36748 = ~n11478 ;
  assign n11481 = n36748 & n11480 ;
  assign n36749 = ~n11481 ;
  assign n11482 = n2431 & n36749 ;
  assign n10928 = n10714 & n36452 ;
  assign n36750 = ~n10936 ;
  assign n11449 = n10928 & n36750 ;
  assign n11450 = n11067 & n11449 ;
  assign n11451 = n10926 | n10936 ;
  assign n36751 = ~n11451 ;
  assign n11452 = n155 & n36751 ;
  assign n11453 = n10714 | n11452 ;
  assign n36752 = ~n11450 ;
  assign n11454 = n36752 & n11453 ;
  assign n36753 = ~n11344 ;
  assign n11487 = n36753 & n11470 ;
  assign n36754 = ~n11487 ;
  assign n11488 = n174 & n36754 ;
  assign n36755 = ~n11488 ;
  assign n11489 = n11476 & n36755 ;
  assign n36756 = ~n11489 ;
  assign n11490 = n2753 & n36756 ;
  assign n11491 = n2431 | n11490 ;
  assign n36757 = ~n11491 ;
  assign n11492 = n11480 & n36757 ;
  assign n11493 = n11454 | n11492 ;
  assign n36758 = ~n11482 ;
  assign n11494 = n36758 & n11493 ;
  assign n36759 = ~n11494 ;
  assign n11495 = n177 & n36759 ;
  assign n36760 = ~n10940 ;
  assign n11442 = n10729 & n36760 ;
  assign n11443 = n36479 & n11442 ;
  assign n11444 = n11067 & n11443 ;
  assign n11445 = n10940 | n10949 ;
  assign n36761 = ~n11445 ;
  assign n11446 = n155 & n36761 ;
  assign n11447 = n10729 | n11446 ;
  assign n36762 = ~n11444 ;
  assign n11448 = n36762 & n11447 ;
  assign n11483 = n177 | n11482 ;
  assign n36763 = ~n11483 ;
  assign n11496 = n36763 & n11493 ;
  assign n11497 = n11448 | n11496 ;
  assign n36764 = ~n11495 ;
  assign n11498 = n36764 & n11497 ;
  assign n36765 = ~n11498 ;
  assign n11499 = n178 & n36765 ;
  assign n10945 = n10731 & n36468 ;
  assign n36766 = ~n10951 ;
  assign n10963 = n10945 & n36766 ;
  assign n11107 = n10963 & n11067 ;
  assign n10964 = n10943 | n10951 ;
  assign n36767 = ~n10964 ;
  assign n11153 = n36767 & n155 ;
  assign n11154 = n10731 | n11153 ;
  assign n36768 = ~n11107 ;
  assign n11155 = n36768 & n11154 ;
  assign n36769 = ~n11490 ;
  assign n11502 = n11480 & n36769 ;
  assign n36770 = ~n11502 ;
  assign n11503 = n176 & n36770 ;
  assign n36771 = ~n11503 ;
  assign n11504 = n11493 & n36771 ;
  assign n36772 = ~n11504 ;
  assign n11505 = n177 & n36772 ;
  assign n11506 = n178 | n11505 ;
  assign n36773 = ~n11506 ;
  assign n11507 = n11497 & n36773 ;
  assign n11508 = n11155 | n11507 ;
  assign n36774 = ~n11499 ;
  assign n11509 = n36774 & n11508 ;
  assign n36775 = ~n11509 ;
  assign n11510 = n179 & n36775 ;
  assign n36776 = ~n10955 ;
  assign n11435 = n10733 & n36776 ;
  assign n11436 = n36495 & n11435 ;
  assign n11437 = n11067 & n11436 ;
  assign n11438 = n10955 | n10966 ;
  assign n36777 = ~n11438 ;
  assign n11439 = n155 & n36777 ;
  assign n11440 = n10733 | n11439 ;
  assign n36778 = ~n11437 ;
  assign n11441 = n36778 & n11440 ;
  assign n11500 = n1707 | n11499 ;
  assign n36779 = ~n11500 ;
  assign n11511 = n36779 & n11508 ;
  assign n11512 = n11441 | n11511 ;
  assign n36780 = ~n11510 ;
  assign n11513 = n36780 & n11512 ;
  assign n36781 = ~n11513 ;
  assign n11514 = n1487 & n36781 ;
  assign n10960 = n10712 & n36484 ;
  assign n36782 = ~n10968 ;
  assign n11429 = n10960 & n36782 ;
  assign n11430 = n11067 & n11429 ;
  assign n11431 = n10958 | n10968 ;
  assign n36783 = ~n11431 ;
  assign n11432 = n155 & n36783 ;
  assign n11433 = n10712 | n11432 ;
  assign n36784 = ~n11430 ;
  assign n11434 = n36784 & n11433 ;
  assign n36785 = ~n11505 ;
  assign n11517 = n11497 & n36785 ;
  assign n36786 = ~n11517 ;
  assign n11518 = n178 & n36786 ;
  assign n36787 = ~n11518 ;
  assign n11519 = n11508 & n36787 ;
  assign n36788 = ~n11519 ;
  assign n11520 = n1707 & n36788 ;
  assign n11521 = n1487 | n11520 ;
  assign n36789 = ~n11521 ;
  assign n11522 = n11512 & n36789 ;
  assign n11523 = n11434 | n11522 ;
  assign n36790 = ~n11514 ;
  assign n11524 = n36790 & n11523 ;
  assign n36791 = ~n11524 ;
  assign n11525 = n181 & n36791 ;
  assign n36792 = ~n10972 ;
  assign n11422 = n10735 & n36792 ;
  assign n11423 = n36511 & n11422 ;
  assign n11424 = n11067 & n11423 ;
  assign n11425 = n10972 | n10981 ;
  assign n36793 = ~n11425 ;
  assign n11426 = n155 & n36793 ;
  assign n11427 = n10735 | n11426 ;
  assign n36794 = ~n11424 ;
  assign n11428 = n36794 & n11427 ;
  assign n11515 = n181 | n11514 ;
  assign n36795 = ~n11515 ;
  assign n11526 = n36795 & n11523 ;
  assign n11527 = n11428 | n11526 ;
  assign n36796 = ~n11525 ;
  assign n11528 = n36796 & n11527 ;
  assign n36797 = ~n11528 ;
  assign n11529 = n182 & n36797 ;
  assign n10977 = n10737 & n36500 ;
  assign n36798 = ~n10983 ;
  assign n11416 = n10977 & n36798 ;
  assign n11417 = n11067 & n11416 ;
  assign n11418 = n10983 | n10994 ;
  assign n36799 = ~n11418 ;
  assign n11419 = n11067 & n36799 ;
  assign n11420 = n10737 | n11419 ;
  assign n36800 = ~n11417 ;
  assign n11421 = n36800 & n11420 ;
  assign n36801 = ~n11520 ;
  assign n11532 = n11512 & n36801 ;
  assign n36802 = ~n11532 ;
  assign n11533 = n180 & n36802 ;
  assign n36803 = ~n11533 ;
  assign n11536 = n11523 & n36803 ;
  assign n36804 = ~n11536 ;
  assign n11537 = n181 & n36804 ;
  assign n11538 = n182 | n11537 ;
  assign n36805 = ~n11538 ;
  assign n11539 = n11527 & n36805 ;
  assign n11540 = n11421 | n11539 ;
  assign n36806 = ~n11529 ;
  assign n11541 = n36806 & n11540 ;
  assign n36807 = ~n11541 ;
  assign n11542 = n183 & n36807 ;
  assign n36808 = ~n10987 ;
  assign n11409 = n10739 & n36808 ;
  assign n11410 = n36527 & n11409 ;
  assign n11411 = n11067 & n11410 ;
  assign n11412 = n10987 | n10996 ;
  assign n36809 = ~n11412 ;
  assign n11413 = n155 & n36809 ;
  assign n11414 = n10739 | n11413 ;
  assign n36810 = ~n11411 ;
  assign n11415 = n36810 & n11414 ;
  assign n11530 = n183 | n11529 ;
  assign n36811 = ~n11530 ;
  assign n11543 = n36811 & n11540 ;
  assign n11544 = n11415 | n11543 ;
  assign n36812 = ~n11542 ;
  assign n11545 = n36812 & n11544 ;
  assign n36813 = ~n11545 ;
  assign n11546 = n838 & n36813 ;
  assign n10992 = n10741 & n36516 ;
  assign n36814 = ~n10998 ;
  assign n11403 = n10992 & n36814 ;
  assign n11404 = n11067 & n11403 ;
  assign n11405 = n10998 | n11009 ;
  assign n36815 = ~n11405 ;
  assign n11406 = n155 & n36815 ;
  assign n11407 = n10741 | n11406 ;
  assign n36816 = ~n11404 ;
  assign n11408 = n36816 & n11407 ;
  assign n36817 = ~n11537 ;
  assign n11549 = n11527 & n36817 ;
  assign n36818 = ~n11549 ;
  assign n11550 = n182 & n36818 ;
  assign n36819 = ~n11550 ;
  assign n11551 = n11540 & n36819 ;
  assign n36820 = ~n11551 ;
  assign n11552 = n996 & n36820 ;
  assign n11553 = n838 | n11552 ;
  assign n36821 = ~n11553 ;
  assign n11554 = n11544 & n36821 ;
  assign n11555 = n11408 | n11554 ;
  assign n36822 = ~n11546 ;
  assign n11556 = n36822 & n11555 ;
  assign n36823 = ~n11556 ;
  assign n11557 = n185 & n36823 ;
  assign n36824 = ~n11002 ;
  assign n11396 = n10699 & n36824 ;
  assign n11397 = n36543 & n11396 ;
  assign n11398 = n11067 & n11397 ;
  assign n11399 = n11002 | n11011 ;
  assign n36825 = ~n11399 ;
  assign n11400 = n155 & n36825 ;
  assign n11401 = n10699 | n11400 ;
  assign n36826 = ~n11398 ;
  assign n11402 = n36826 & n11401 ;
  assign n11547 = n185 | n11546 ;
  assign n36827 = ~n11547 ;
  assign n11558 = n36827 & n11555 ;
  assign n11559 = n11402 | n11558 ;
  assign n36828 = ~n11557 ;
  assign n11560 = n36828 & n11559 ;
  assign n36829 = ~n11560 ;
  assign n11561 = n186 & n36829 ;
  assign n11007 = n10727 & n36532 ;
  assign n36830 = ~n11013 ;
  assign n11390 = n11007 & n36830 ;
  assign n11391 = n11067 & n11390 ;
  assign n11392 = n11013 | n11024 ;
  assign n36831 = ~n11392 ;
  assign n11393 = n155 & n36831 ;
  assign n11394 = n10727 | n11393 ;
  assign n36832 = ~n11391 ;
  assign n11395 = n36832 & n11394 ;
  assign n36833 = ~n11552 ;
  assign n11564 = n11544 & n36833 ;
  assign n36834 = ~n11564 ;
  assign n11565 = n184 & n36834 ;
  assign n36835 = ~n11565 ;
  assign n11566 = n11555 & n36835 ;
  assign n36836 = ~n11566 ;
  assign n11567 = n185 & n36836 ;
  assign n11568 = n186 | n11567 ;
  assign n36837 = ~n11568 ;
  assign n11569 = n11559 & n36837 ;
  assign n11570 = n11395 | n11569 ;
  assign n36838 = ~n11561 ;
  assign n11571 = n36838 & n11570 ;
  assign n36839 = ~n11571 ;
  assign n11572 = n187 & n36839 ;
  assign n36840 = ~n11017 ;
  assign n11383 = n10678 & n36840 ;
  assign n11384 = n36559 & n11383 ;
  assign n11385 = n11067 & n11384 ;
  assign n11386 = n11017 | n11026 ;
  assign n36841 = ~n11386 ;
  assign n11387 = n155 & n36841 ;
  assign n11388 = n10678 | n11387 ;
  assign n36842 = ~n11385 ;
  assign n11389 = n36842 & n11388 ;
  assign n11562 = n528 | n11561 ;
  assign n36843 = ~n11562 ;
  assign n11573 = n36843 & n11570 ;
  assign n11574 = n11389 | n11573 ;
  assign n36844 = ~n11572 ;
  assign n11575 = n36844 & n11574 ;
  assign n36845 = ~n11575 ;
  assign n11576 = n413 & n36845 ;
  assign n11577 = n189 | n11576 ;
  assign n11022 = n10725 & n36548 ;
  assign n36846 = ~n11028 ;
  assign n11040 = n11022 & n36846 ;
  assign n11108 = n11040 & n11067 ;
  assign n11041 = n11028 | n11039 ;
  assign n36847 = ~n11041 ;
  assign n11156 = n36847 & n155 ;
  assign n11157 = n10725 | n11156 ;
  assign n36848 = ~n11108 ;
  assign n11158 = n36848 & n11157 ;
  assign n36849 = ~n11567 ;
  assign n11579 = n11559 & n36849 ;
  assign n36850 = ~n11579 ;
  assign n11580 = n186 & n36850 ;
  assign n36851 = ~n11580 ;
  assign n11581 = n11570 & n36851 ;
  assign n36852 = ~n11581 ;
  assign n11582 = n528 & n36852 ;
  assign n11583 = n413 | n11582 ;
  assign n36853 = ~n11583 ;
  assign n11584 = n11574 & n36853 ;
  assign n11585 = n11158 | n11584 ;
  assign n36854 = ~n11577 ;
  assign n11588 = n36854 & n11585 ;
  assign n11589 = n11382 | n11588 ;
  assign n36855 = ~n11582 ;
  assign n11594 = n11574 & n36855 ;
  assign n36856 = ~n11594 ;
  assign n11595 = n188 & n36856 ;
  assign n36857 = ~n11595 ;
  assign n11596 = n11585 & n36857 ;
  assign n36858 = ~n11596 ;
  assign n11597 = n189 & n36858 ;
  assign n36859 = ~n11597 ;
  assign n11599 = n11589 & n36859 ;
  assign n36860 = ~n11599 ;
  assign n11600 = n190 & n36860 ;
  assign n11037 = n10723 & n36564 ;
  assign n36861 = ~n11045 ;
  assign n11370 = n11037 & n36861 ;
  assign n11371 = n155 & n11370 ;
  assign n11372 = n11035 | n11045 ;
  assign n36862 = ~n11372 ;
  assign n11373 = n155 & n36862 ;
  assign n11374 = n10723 | n11373 ;
  assign n36863 = ~n11371 ;
  assign n11375 = n36863 & n11374 ;
  assign n11598 = n190 | n11597 ;
  assign n36864 = ~n11598 ;
  assign n11601 = n11589 & n36864 ;
  assign n11602 = n11375 | n11601 ;
  assign n36865 = ~n11600 ;
  assign n11605 = n36865 & n11602 ;
  assign n36866 = ~n11605 ;
  assign n11606 = n287 & n36866 ;
  assign n36867 = ~n11049 ;
  assign n11363 = n10911 & n36867 ;
  assign n11364 = n36588 & n11363 ;
  assign n11365 = n155 & n11364 ;
  assign n11366 = n11049 | n11058 ;
  assign n36868 = ~n11366 ;
  assign n11367 = n155 & n36868 ;
  assign n11368 = n10911 | n11367 ;
  assign n36869 = ~n11365 ;
  assign n11369 = n36869 & n11368 ;
  assign n36870 = ~n11576 ;
  assign n11586 = n36870 & n11585 ;
  assign n36871 = ~n11586 ;
  assign n11587 = n189 & n36871 ;
  assign n36872 = ~n11587 ;
  assign n11590 = n36872 & n11589 ;
  assign n36873 = ~n11590 ;
  assign n11591 = n190 & n36873 ;
  assign n11592 = n287 | n11591 ;
  assign n36874 = ~n11592 ;
  assign n11603 = n36874 & n11602 ;
  assign n11610 = n11369 | n11603 ;
  assign n36875 = ~n11606 ;
  assign n11611 = n36875 & n11610 ;
  assign n11612 = n11151 | n11611 ;
  assign n11613 = n31336 & n11612 ;
  assign n10896 = n10886 | n10895 ;
  assign n36876 = ~n10896 ;
  assign n10902 = n36876 & n10899 ;
  assign n10903 = n36608 & n10902 ;
  assign n11120 = n10903 & n36609 ;
  assign n11121 = n36610 & n11120 ;
  assign n11129 = n192 & n11126 ;
  assign n36877 = ~n10900 ;
  assign n11302 = n36877 & n155 ;
  assign n36878 = ~n11302 ;
  assign n11303 = n11062 & n36878 ;
  assign n36879 = ~n11303 ;
  assign n11304 = n11129 & n36879 ;
  assign n11305 = n11121 | n11304 ;
  assign n11607 = n11150 & n36875 ;
  assign n11616 = n11607 & n11610 ;
  assign n11617 = n11305 | n11616 ;
  assign n154 = n11613 | n11617 ;
  assign n11609 = n11603 | n11606 ;
  assign n36880 = ~n11609 ;
  assign n11686 = n36880 & n154 ;
  assign n11687 = n11369 | n11686 ;
  assign n36881 = ~n11603 ;
  assign n11604 = n11369 & n36881 ;
  assign n11608 = n11604 & n36875 ;
  assign n11705 = n11608 & n154 ;
  assign n36882 = ~n11705 ;
  assign n11706 = n11687 & n36882 ;
  assign n11614 = n11150 | n11611 ;
  assign n36883 = ~n11614 ;
  assign n11688 = n36883 & n154 ;
  assign n11947 = n11616 | n11688 ;
  assign n11948 = n11706 | n11947 ;
  assign n197 = x48 | x49 ;
  assign n198 = x50 | n197 ;
  assign n11656 = x50 & n154 ;
  assign n36884 = ~n11656 ;
  assign n11657 = n198 & n36884 ;
  assign n36885 = ~n11657 ;
  assign n11658 = n155 & n36885 ;
  assign n10890 = n198 & n36607 ;
  assign n10891 = n36608 & n10890 ;
  assign n11124 = n10891 & n36609 ;
  assign n11125 = n36610 & n11124 ;
  assign n11700 = n11125 & n36884 ;
  assign n36886 = ~n194 ;
  assign n11655 = n36886 & n154 ;
  assign n36887 = ~x50 ;
  assign n11712 = n36887 & n154 ;
  assign n36888 = ~n11712 ;
  assign n11713 = x51 & n36888 ;
  assign n11714 = n11655 | n11713 ;
  assign n11715 = n11700 | n11714 ;
  assign n36889 = ~n11658 ;
  assign n11718 = n36889 & n11715 ;
  assign n36890 = ~n11718 ;
  assign n11719 = n10657 & n36890 ;
  assign n199 = n36887 & n197 ;
  assign n36891 = ~n154 ;
  assign n11707 = x50 & n36891 ;
  assign n11708 = n199 | n11707 ;
  assign n36892 = ~n11708 ;
  assign n11709 = n11067 & n36892 ;
  assign n11710 = n10657 | n11709 ;
  assign n36893 = ~n11710 ;
  assign n11716 = n36893 & n11715 ;
  assign n36894 = ~n11121 ;
  assign n11122 = n11067 & n36894 ;
  assign n36895 = ~n11304 ;
  assign n11306 = n11122 & n36895 ;
  assign n36896 = ~n11616 ;
  assign n11724 = n11306 & n36896 ;
  assign n36897 = ~n11613 ;
  assign n11725 = n36897 & n11724 ;
  assign n11726 = n11655 | n11725 ;
  assign n11727 = x52 & n11726 ;
  assign n11728 = x52 | n11725 ;
  assign n11729 = n11655 | n11728 ;
  assign n36898 = ~n11727 ;
  assign n11730 = n36898 & n11729 ;
  assign n11731 = n11716 | n11730 ;
  assign n36899 = ~n11719 ;
  assign n11732 = n36899 & n11731 ;
  assign n36900 = ~n11732 ;
  assign n11733 = n157 & n36900 ;
  assign n11087 = n11071 | n11086 ;
  assign n36901 = ~n11087 ;
  assign n11695 = n36901 & n154 ;
  assign n11696 = n11092 | n11695 ;
  assign n11093 = n36901 & n11092 ;
  assign n11701 = n11093 & n154 ;
  assign n36902 = ~n11701 ;
  assign n11702 = n11696 & n36902 ;
  assign n11721 = n157 | n11719 ;
  assign n36903 = ~n11721 ;
  assign n11736 = n36903 & n11731 ;
  assign n11737 = n11702 | n11736 ;
  assign n36904 = ~n11733 ;
  assign n11738 = n36904 & n11737 ;
  assign n36905 = ~n11738 ;
  assign n11739 = n158 & n36905 ;
  assign n11099 = n11096 | n11098 ;
  assign n36906 = ~n11099 ;
  assign n11693 = n36906 & n154 ;
  assign n11694 = n11115 | n11693 ;
  assign n36907 = ~n11098 ;
  assign n11116 = n36907 & n11115 ;
  assign n11117 = n36615 & n11116 ;
  assign n11703 = n11117 & n154 ;
  assign n36908 = ~n11703 ;
  assign n11704 = n11694 & n36908 ;
  assign n11734 = n158 | n11733 ;
  assign n36909 = ~n11734 ;
  assign n11740 = n36909 & n11737 ;
  assign n11741 = n11704 | n11740 ;
  assign n36910 = ~n11739 ;
  assign n11742 = n36910 & n11741 ;
  assign n36911 = ~n11742 ;
  assign n11743 = n8857 & n36911 ;
  assign n11217 = n36621 & n11199 ;
  assign n36912 = ~n11119 ;
  assign n11218 = n36912 & n11217 ;
  assign n11689 = n11218 & n154 ;
  assign n11192 = n11119 | n11191 ;
  assign n36913 = ~n11192 ;
  assign n11690 = n36913 & n154 ;
  assign n11691 = n11199 | n11690 ;
  assign n36914 = ~n11689 ;
  assign n11692 = n36914 & n11691 ;
  assign n11722 = n156 & n36890 ;
  assign n11659 = n156 | n11658 ;
  assign n36915 = ~n11659 ;
  assign n11723 = n36915 & n11715 ;
  assign n11752 = n11723 | n11730 ;
  assign n36916 = ~n11722 ;
  assign n11753 = n36916 & n11752 ;
  assign n36917 = ~n11753 ;
  assign n11754 = n157 & n36917 ;
  assign n11755 = n36903 & n11752 ;
  assign n11756 = n11702 | n11755 ;
  assign n36918 = ~n11754 ;
  assign n11757 = n36918 & n11756 ;
  assign n36919 = ~n11757 ;
  assign n11758 = n158 & n36919 ;
  assign n11759 = n8857 | n11758 ;
  assign n36920 = ~n11759 ;
  assign n11760 = n11741 & n36920 ;
  assign n11761 = n11692 | n11760 ;
  assign n36921 = ~n11743 ;
  assign n11762 = n36921 & n11761 ;
  assign n36922 = ~n11762 ;
  assign n11763 = n160 & n36922 ;
  assign n36923 = ~n11204 ;
  assign n11214 = n11196 & n36923 ;
  assign n11215 = n36627 & n11214 ;
  assign n11647 = n11215 & n154 ;
  assign n11216 = n11202 | n11204 ;
  assign n36924 = ~n11216 ;
  assign n11669 = n36924 & n154 ;
  assign n11670 = n11196 | n11669 ;
  assign n36925 = ~n11647 ;
  assign n11671 = n36925 & n11670 ;
  assign n11744 = n160 | n11743 ;
  assign n36926 = ~n11744 ;
  assign n11764 = n36926 & n11761 ;
  assign n11765 = n11671 | n11764 ;
  assign n36927 = ~n11763 ;
  assign n11766 = n36927 & n11765 ;
  assign n36928 = ~n11766 ;
  assign n11767 = n161 & n36928 ;
  assign n11213 = n11207 | n11208 ;
  assign n36929 = ~n11213 ;
  assign n11619 = n36929 & n154 ;
  assign n11620 = n11177 | n11619 ;
  assign n11236 = n11177 & n36652 ;
  assign n36930 = ~n11208 ;
  assign n11237 = n36930 & n11236 ;
  assign n11648 = n11237 & n154 ;
  assign n36931 = ~n11648 ;
  assign n11649 = n11620 & n36931 ;
  assign n11775 = n36909 & n11756 ;
  assign n11776 = n11704 | n11775 ;
  assign n36932 = ~n11758 ;
  assign n11777 = n36932 & n11776 ;
  assign n36933 = ~n11777 ;
  assign n11778 = n159 & n36933 ;
  assign n11779 = n36920 & n11776 ;
  assign n11780 = n11692 | n11779 ;
  assign n36934 = ~n11778 ;
  assign n11781 = n36934 & n11780 ;
  assign n36935 = ~n11781 ;
  assign n11782 = n8534 & n36935 ;
  assign n11783 = n161 | n11782 ;
  assign n36936 = ~n11783 ;
  assign n11784 = n11765 & n36936 ;
  assign n11785 = n11649 | n11784 ;
  assign n36937 = ~n11767 ;
  assign n11786 = n36937 & n11785 ;
  assign n36938 = ~n11786 ;
  assign n11787 = n162 & n36938 ;
  assign n11235 = n11211 | n11223 ;
  assign n36939 = ~n11235 ;
  assign n11641 = n36939 & n154 ;
  assign n11642 = n11171 | n11641 ;
  assign n36940 = ~n11223 ;
  assign n11233 = n11171 & n36940 ;
  assign n11234 = n36641 & n11233 ;
  assign n11643 = n11234 & n154 ;
  assign n36941 = ~n11643 ;
  assign n11644 = n11642 & n36941 ;
  assign n11768 = n162 | n11767 ;
  assign n36942 = ~n11768 ;
  assign n11788 = n36942 & n11785 ;
  assign n11789 = n11644 | n11788 ;
  assign n36943 = ~n11787 ;
  assign n11790 = n36943 & n11789 ;
  assign n36944 = ~n11790 ;
  assign n11791 = n6889 & n36944 ;
  assign n11256 = n11105 & n36668 ;
  assign n36945 = ~n11227 ;
  assign n11257 = n36945 & n11256 ;
  assign n11636 = n11257 & n154 ;
  assign n11232 = n11226 | n11227 ;
  assign n36946 = ~n11232 ;
  assign n11637 = n36946 & n154 ;
  assign n11638 = n11105 | n11637 ;
  assign n36947 = ~n11636 ;
  assign n11639 = n36947 & n11638 ;
  assign n11799 = n36926 & n11780 ;
  assign n11800 = n11671 | n11799 ;
  assign n36948 = ~n11782 ;
  assign n11801 = n36948 & n11800 ;
  assign n36949 = ~n11801 ;
  assign n11802 = n161 & n36949 ;
  assign n11803 = n36936 & n11800 ;
  assign n11804 = n11649 | n11803 ;
  assign n36950 = ~n11802 ;
  assign n11805 = n36950 & n11804 ;
  assign n36951 = ~n11805 ;
  assign n11806 = n162 & n36951 ;
  assign n11807 = n6889 | n11806 ;
  assign n36952 = ~n11807 ;
  assign n11808 = n11789 & n36952 ;
  assign n11809 = n11639 | n11808 ;
  assign n36953 = ~n11791 ;
  assign n11810 = n36953 & n11809 ;
  assign n36954 = ~n11810 ;
  assign n11811 = n164 & n36954 ;
  assign n11253 = n11230 | n11243 ;
  assign n36955 = ~n11253 ;
  assign n11634 = n36955 & n154 ;
  assign n11635 = n11174 | n11634 ;
  assign n36956 = ~n11243 ;
  assign n11254 = n11174 & n36956 ;
  assign n11255 = n36657 & n11254 ;
  assign n11660 = n11255 & n154 ;
  assign n36957 = ~n11660 ;
  assign n11661 = n11635 & n36957 ;
  assign n11792 = n6600 | n11791 ;
  assign n36958 = ~n11792 ;
  assign n11812 = n36958 & n11809 ;
  assign n11815 = n11661 | n11812 ;
  assign n36959 = ~n11811 ;
  assign n11816 = n36959 & n11815 ;
  assign n36960 = ~n11816 ;
  assign n11817 = n165 & n36960 ;
  assign n11252 = n11246 | n11247 ;
  assign n36961 = ~n11252 ;
  assign n11645 = n36961 & n154 ;
  assign n11646 = n11102 | n11645 ;
  assign n11276 = n11102 & n36684 ;
  assign n36962 = ~n11247 ;
  assign n11277 = n36962 & n11276 ;
  assign n11662 = n11277 & n154 ;
  assign n36963 = ~n11662 ;
  assign n11663 = n11646 & n36963 ;
  assign n11823 = n36942 & n11804 ;
  assign n11824 = n11644 | n11823 ;
  assign n36964 = ~n11806 ;
  assign n11825 = n36964 & n11824 ;
  assign n36965 = ~n11825 ;
  assign n11826 = n163 & n36965 ;
  assign n11827 = n36952 & n11824 ;
  assign n11828 = n11639 | n11827 ;
  assign n36966 = ~n11826 ;
  assign n11829 = n36966 & n11828 ;
  assign n36967 = ~n11829 ;
  assign n11830 = n6600 & n36967 ;
  assign n11831 = n165 | n11830 ;
  assign n36968 = ~n11831 ;
  assign n11832 = n11815 & n36968 ;
  assign n11833 = n11663 | n11832 ;
  assign n36969 = ~n11817 ;
  assign n11834 = n36969 & n11833 ;
  assign n36970 = ~n11834 ;
  assign n11835 = n166 & n36970 ;
  assign n11275 = n11250 | n11263 ;
  assign n36971 = ~n11275 ;
  assign n11624 = n36971 & n154 ;
  assign n11625 = n11168 | n11624 ;
  assign n36972 = ~n11263 ;
  assign n11273 = n11168 & n36972 ;
  assign n11274 = n36673 & n11273 ;
  assign n11664 = n11274 & n154 ;
  assign n36973 = ~n11664 ;
  assign n11665 = n11625 & n36973 ;
  assign n11818 = n166 | n11817 ;
  assign n36974 = ~n11818 ;
  assign n11836 = n36974 & n11833 ;
  assign n11837 = n11665 | n11836 ;
  assign n36975 = ~n11835 ;
  assign n11838 = n36975 & n11837 ;
  assign n36976 = ~n11838 ;
  assign n11839 = n5352 & n36976 ;
  assign n11272 = n11266 | n11267 ;
  assign n36977 = ~n11272 ;
  assign n11631 = n36977 & n154 ;
  assign n11632 = n11183 | n11631 ;
  assign n11292 = n11183 & n36700 ;
  assign n36978 = ~n11267 ;
  assign n11293 = n36978 & n11292 ;
  assign n11650 = n11293 & n154 ;
  assign n36979 = ~n11650 ;
  assign n11651 = n11632 & n36979 ;
  assign n11847 = n36958 & n11828 ;
  assign n11848 = n11661 | n11847 ;
  assign n36980 = ~n11830 ;
  assign n11849 = n36980 & n11848 ;
  assign n36981 = ~n11849 ;
  assign n11850 = n165 & n36981 ;
  assign n11851 = n36968 & n11848 ;
  assign n11852 = n11663 | n11851 ;
  assign n36982 = ~n11850 ;
  assign n11853 = n36982 & n11852 ;
  assign n36983 = ~n11853 ;
  assign n11854 = n166 & n36983 ;
  assign n11855 = n5352 | n11854 ;
  assign n36984 = ~n11855 ;
  assign n11856 = n11837 & n36984 ;
  assign n11857 = n11651 | n11856 ;
  assign n36985 = ~n11839 ;
  assign n11858 = n36985 & n11857 ;
  assign n36986 = ~n11858 ;
  assign n11859 = n168 & n36986 ;
  assign n11291 = n11270 | n11283 ;
  assign n36987 = ~n11291 ;
  assign n11667 = n36987 & n154 ;
  assign n11668 = n11180 | n11667 ;
  assign n36988 = ~n11283 ;
  assign n11289 = n11180 & n36988 ;
  assign n11290 = n36689 & n11289 ;
  assign n11678 = n11290 & n154 ;
  assign n36989 = ~n11678 ;
  assign n11679 = n11668 & n36989 ;
  assign n11840 = n4934 | n11839 ;
  assign n36990 = ~n11840 ;
  assign n11860 = n36990 & n11857 ;
  assign n11861 = n11679 | n11860 ;
  assign n36991 = ~n11859 ;
  assign n11862 = n36991 & n11861 ;
  assign n36992 = ~n11862 ;
  assign n11863 = n169 & n36992 ;
  assign n11288 = n11286 | n11287 ;
  assign n36993 = ~n11288 ;
  assign n11621 = n36993 & n154 ;
  assign n11622 = n11312 | n11621 ;
  assign n11330 = n36716 & n11312 ;
  assign n36994 = ~n11287 ;
  assign n11331 = n36994 & n11330 ;
  assign n11674 = n11331 & n154 ;
  assign n36995 = ~n11674 ;
  assign n11675 = n11622 & n36995 ;
  assign n11871 = n36974 & n11852 ;
  assign n11872 = n11665 | n11871 ;
  assign n36996 = ~n11854 ;
  assign n11873 = n36996 & n11872 ;
  assign n36997 = ~n11873 ;
  assign n11874 = n167 & n36997 ;
  assign n11875 = n36984 & n11872 ;
  assign n11876 = n11651 | n11875 ;
  assign n36998 = ~n11874 ;
  assign n11877 = n36998 & n11876 ;
  assign n36999 = ~n11877 ;
  assign n11878 = n4934 & n36999 ;
  assign n11879 = n169 | n11878 ;
  assign n37000 = ~n11879 ;
  assign n11880 = n11861 & n37000 ;
  assign n11881 = n11675 | n11880 ;
  assign n37001 = ~n11863 ;
  assign n11882 = n37001 & n11881 ;
  assign n37002 = ~n11882 ;
  assign n11883 = n170 & n37002 ;
  assign n11329 = n11315 | n11317 ;
  assign n37003 = ~n11329 ;
  assign n11672 = n37003 & n154 ;
  assign n11673 = n11147 | n11672 ;
  assign n37004 = ~n11317 ;
  assign n11327 = n11147 & n37004 ;
  assign n11328 = n36705 & n11327 ;
  assign n11676 = n11328 & n154 ;
  assign n37005 = ~n11676 ;
  assign n11677 = n11673 & n37005 ;
  assign n11864 = n170 | n11863 ;
  assign n37006 = ~n11864 ;
  assign n11884 = n37006 & n11881 ;
  assign n11885 = n11677 | n11884 ;
  assign n37007 = ~n11883 ;
  assign n11886 = n37007 & n11885 ;
  assign n37008 = ~n11886 ;
  assign n11887 = n3940 & n37008 ;
  assign n11350 = n11165 & n36722 ;
  assign n37009 = ~n11321 ;
  assign n11351 = n37009 & n11350 ;
  assign n11666 = n11351 & n154 ;
  assign n11326 = n11320 | n11321 ;
  assign n37010 = ~n11326 ;
  assign n11680 = n37010 & n154 ;
  assign n11681 = n11165 | n11680 ;
  assign n37011 = ~n11666 ;
  assign n11682 = n37011 & n11681 ;
  assign n11895 = n36990 & n11876 ;
  assign n11896 = n11679 | n11895 ;
  assign n37012 = ~n11878 ;
  assign n11897 = n37012 & n11896 ;
  assign n37013 = ~n11897 ;
  assign n11898 = n169 & n37013 ;
  assign n11899 = n37000 & n11896 ;
  assign n11900 = n11675 | n11899 ;
  assign n37014 = ~n11898 ;
  assign n11901 = n37014 & n11900 ;
  assign n37015 = ~n11901 ;
  assign n11902 = n170 & n37015 ;
  assign n11903 = n3940 | n11902 ;
  assign n37016 = ~n11903 ;
  assign n11904 = n11885 & n37016 ;
  assign n11905 = n11682 | n11904 ;
  assign n37017 = ~n11887 ;
  assign n11906 = n37017 & n11905 ;
  assign n37018 = ~n11906 ;
  assign n11907 = n172 & n37018 ;
  assign n37019 = ~n11337 ;
  assign n11347 = n11301 & n37019 ;
  assign n11348 = n36737 & n11347 ;
  assign n11633 = n11348 & n154 ;
  assign n11349 = n11324 | n11337 ;
  assign n37020 = ~n11349 ;
  assign n11683 = n37020 & n154 ;
  assign n11684 = n11301 | n11683 ;
  assign n37021 = ~n11633 ;
  assign n11685 = n37021 & n11684 ;
  assign n11888 = n3631 | n11887 ;
  assign n37022 = ~n11888 ;
  assign n11908 = n37022 & n11905 ;
  assign n11909 = n11685 | n11908 ;
  assign n37023 = ~n11907 ;
  assign n11910 = n37023 & n11909 ;
  assign n37024 = ~n11910 ;
  assign n11911 = n173 & n37024 ;
  assign n11359 = n11162 & n36726 ;
  assign n37025 = ~n11341 ;
  assign n11360 = n37025 & n11359 ;
  assign n11627 = n11360 & n154 ;
  assign n11346 = n11340 | n11341 ;
  assign n37026 = ~n11346 ;
  assign n11628 = n37026 & n154 ;
  assign n11629 = n11162 | n11628 ;
  assign n37027 = ~n11627 ;
  assign n11630 = n37027 & n11629 ;
  assign n11919 = n37006 & n11900 ;
  assign n11920 = n11677 | n11919 ;
  assign n37028 = ~n11902 ;
  assign n11921 = n37028 & n11920 ;
  assign n37029 = ~n11921 ;
  assign n11922 = n171 & n37029 ;
  assign n11923 = n37016 & n11920 ;
  assign n11924 = n11682 | n11923 ;
  assign n37030 = ~n11922 ;
  assign n11925 = n37030 & n11924 ;
  assign n37031 = ~n11925 ;
  assign n11926 = n3631 & n37031 ;
  assign n11927 = n173 | n11926 ;
  assign n37032 = ~n11927 ;
  assign n11928 = n11909 & n37032 ;
  assign n11929 = n11630 | n11928 ;
  assign n37033 = ~n11911 ;
  assign n11930 = n37033 & n11929 ;
  assign n37034 = ~n11930 ;
  assign n11931 = n174 & n37034 ;
  assign n11913 = n174 | n11911 ;
  assign n37035 = ~n11913 ;
  assign n11932 = n37035 & n11929 ;
  assign n37036 = ~n11357 ;
  assign n11485 = n37036 & n11469 ;
  assign n11486 = n36753 & n11485 ;
  assign n11640 = n11486 & n154 ;
  assign n11358 = n11344 | n11357 ;
  assign n37037 = ~n11358 ;
  assign n11626 = n37037 & n154 ;
  assign n12065 = n11469 | n11626 ;
  assign n37038 = ~n11640 ;
  assign n12066 = n37038 & n12065 ;
  assign n12067 = n11932 | n12066 ;
  assign n37039 = ~n11931 ;
  assign n12068 = n37039 & n12067 ;
  assign n37040 = ~n12068 ;
  assign n12069 = n2753 & n37040 ;
  assign n11474 = n11467 & n36742 ;
  assign n37041 = ~n11475 ;
  assign n12059 = n11474 & n37041 ;
  assign n12060 = n154 & n12059 ;
  assign n12061 = n11475 | n11488 ;
  assign n37042 = ~n12061 ;
  assign n12062 = n154 & n37042 ;
  assign n12063 = n11467 | n12062 ;
  assign n37043 = ~n12060 ;
  assign n12064 = n37043 & n12063 ;
  assign n11936 = n37022 & n11924 ;
  assign n11937 = n11685 | n11936 ;
  assign n37044 = ~n11926 ;
  assign n11938 = n37044 & n11937 ;
  assign n37045 = ~n11938 ;
  assign n11939 = n173 & n37045 ;
  assign n11940 = n37032 & n11937 ;
  assign n11941 = n11630 | n11940 ;
  assign n37046 = ~n11939 ;
  assign n11942 = n37046 & n11941 ;
  assign n37047 = ~n11942 ;
  assign n11943 = n174 & n37047 ;
  assign n11944 = n2753 | n11943 ;
  assign n37048 = ~n11944 ;
  assign n12072 = n37048 & n12067 ;
  assign n12073 = n12064 | n12072 ;
  assign n37049 = ~n12069 ;
  assign n12074 = n37049 & n12073 ;
  assign n37050 = ~n12074 ;
  assign n12075 = n176 & n37050 ;
  assign n37051 = ~n11479 ;
  assign n12052 = n11461 & n37051 ;
  assign n12053 = n36769 & n12052 ;
  assign n12054 = n154 & n12053 ;
  assign n12055 = n11479 | n11490 ;
  assign n37052 = ~n12055 ;
  assign n12056 = n154 & n37052 ;
  assign n12057 = n11461 | n12056 ;
  assign n37053 = ~n12054 ;
  assign n12058 = n37053 & n12057 ;
  assign n12070 = n2431 | n12069 ;
  assign n37054 = ~n12070 ;
  assign n12076 = n37054 & n12073 ;
  assign n12077 = n12058 | n12076 ;
  assign n37055 = ~n12075 ;
  assign n12078 = n37055 & n12077 ;
  assign n37056 = ~n12078 ;
  assign n12079 = n177 & n37056 ;
  assign n11484 = n11454 & n36758 ;
  assign n37057 = ~n11492 ;
  assign n12046 = n11484 & n37057 ;
  assign n12047 = n154 & n12046 ;
  assign n12048 = n11492 | n11503 ;
  assign n37058 = ~n12048 ;
  assign n12049 = n154 & n37058 ;
  assign n12050 = n11454 | n12049 ;
  assign n37059 = ~n12047 ;
  assign n12051 = n37059 & n12050 ;
  assign n11946 = n37035 & n11941 ;
  assign n12088 = n11946 | n12066 ;
  assign n37060 = ~n11943 ;
  assign n12089 = n37060 & n12088 ;
  assign n37061 = ~n12089 ;
  assign n12090 = n175 & n37061 ;
  assign n12091 = n37048 & n12088 ;
  assign n12092 = n12064 | n12091 ;
  assign n37062 = ~n12090 ;
  assign n12093 = n37062 & n12092 ;
  assign n37063 = ~n12093 ;
  assign n12094 = n2431 & n37063 ;
  assign n12095 = n177 | n12094 ;
  assign n37064 = ~n12095 ;
  assign n12096 = n12077 & n37064 ;
  assign n12097 = n12051 | n12096 ;
  assign n37065 = ~n12079 ;
  assign n12098 = n37065 & n12097 ;
  assign n37066 = ~n12098 ;
  assign n12099 = n178 & n37066 ;
  assign n12039 = n11496 | n11505 ;
  assign n37067 = ~n12039 ;
  assign n12040 = n154 & n37067 ;
  assign n12041 = n11448 | n12040 ;
  assign n37068 = ~n11496 ;
  assign n12042 = n11448 & n37068 ;
  assign n12043 = n36785 & n12042 ;
  assign n12044 = n154 & n12043 ;
  assign n37069 = ~n12044 ;
  assign n12045 = n12041 & n37069 ;
  assign n12080 = n178 | n12079 ;
  assign n37070 = ~n12080 ;
  assign n12100 = n37070 & n12097 ;
  assign n12101 = n12045 | n12100 ;
  assign n37071 = ~n12099 ;
  assign n12102 = n37071 & n12101 ;
  assign n37072 = ~n12102 ;
  assign n12103 = n1707 & n37072 ;
  assign n11501 = n11155 & n36774 ;
  assign n37073 = ~n11507 ;
  assign n12033 = n11501 & n37073 ;
  assign n12034 = n154 & n12033 ;
  assign n12035 = n11507 | n11518 ;
  assign n37074 = ~n12035 ;
  assign n12036 = n154 & n37074 ;
  assign n12037 = n11155 | n12036 ;
  assign n37075 = ~n12034 ;
  assign n12038 = n37075 & n12037 ;
  assign n12111 = n37054 & n12092 ;
  assign n12112 = n12058 | n12111 ;
  assign n37076 = ~n12094 ;
  assign n12113 = n37076 & n12112 ;
  assign n37077 = ~n12113 ;
  assign n12114 = n177 & n37077 ;
  assign n12115 = n37064 & n12112 ;
  assign n12116 = n12051 | n12115 ;
  assign n37078 = ~n12114 ;
  assign n12117 = n37078 & n12116 ;
  assign n37079 = ~n12117 ;
  assign n12118 = n178 & n37079 ;
  assign n12119 = n1707 | n12118 ;
  assign n37080 = ~n12119 ;
  assign n12120 = n12101 & n37080 ;
  assign n12121 = n12038 | n12120 ;
  assign n37081 = ~n12103 ;
  assign n12122 = n37081 & n12121 ;
  assign n37082 = ~n12122 ;
  assign n12123 = n180 & n37082 ;
  assign n37083 = ~n11511 ;
  assign n12026 = n11441 & n37083 ;
  assign n12027 = n36801 & n12026 ;
  assign n12028 = n154 & n12027 ;
  assign n12029 = n11511 | n11520 ;
  assign n37084 = ~n12029 ;
  assign n12030 = n154 & n37084 ;
  assign n12031 = n11441 | n12030 ;
  assign n37085 = ~n12028 ;
  assign n12032 = n37085 & n12031 ;
  assign n12104 = n1487 | n12103 ;
  assign n37086 = ~n12104 ;
  assign n12124 = n37086 & n12121 ;
  assign n12125 = n12032 | n12124 ;
  assign n37087 = ~n12123 ;
  assign n12126 = n37087 & n12125 ;
  assign n37088 = ~n12126 ;
  assign n12127 = n181 & n37088 ;
  assign n11516 = n11434 & n36790 ;
  assign n37089 = ~n11522 ;
  assign n11534 = n11516 & n37089 ;
  assign n11623 = n11534 & n154 ;
  assign n11535 = n11522 | n11533 ;
  assign n37090 = ~n11535 ;
  assign n11652 = n37090 & n154 ;
  assign n11653 = n11434 | n11652 ;
  assign n37091 = ~n11623 ;
  assign n11654 = n37091 & n11653 ;
  assign n12135 = n37070 & n12116 ;
  assign n12136 = n12045 | n12135 ;
  assign n37092 = ~n12118 ;
  assign n12137 = n37092 & n12136 ;
  assign n37093 = ~n12137 ;
  assign n12138 = n179 & n37093 ;
  assign n12139 = n37080 & n12136 ;
  assign n12140 = n12038 | n12139 ;
  assign n37094 = ~n12138 ;
  assign n12141 = n37094 & n12140 ;
  assign n37095 = ~n12141 ;
  assign n12142 = n1487 & n37095 ;
  assign n12143 = n181 | n12142 ;
  assign n37096 = ~n12143 ;
  assign n12144 = n12125 & n37096 ;
  assign n12145 = n11654 | n12144 ;
  assign n37097 = ~n12127 ;
  assign n12146 = n37097 & n12145 ;
  assign n37098 = ~n12146 ;
  assign n12147 = n182 & n37098 ;
  assign n37099 = ~n11526 ;
  assign n12019 = n11428 & n37099 ;
  assign n12020 = n36817 & n12019 ;
  assign n12021 = n154 & n12020 ;
  assign n12022 = n11526 | n11537 ;
  assign n37100 = ~n12022 ;
  assign n12023 = n154 & n37100 ;
  assign n12024 = n11428 | n12023 ;
  assign n37101 = ~n12021 ;
  assign n12025 = n37101 & n12024 ;
  assign n12128 = n182 | n12127 ;
  assign n37102 = ~n12128 ;
  assign n12148 = n37102 & n12145 ;
  assign n12149 = n12025 | n12148 ;
  assign n37103 = ~n12147 ;
  assign n12150 = n37103 & n12149 ;
  assign n37104 = ~n12150 ;
  assign n12151 = n996 & n37104 ;
  assign n11531 = n11421 & n36806 ;
  assign n37105 = ~n11539 ;
  assign n12013 = n11531 & n37105 ;
  assign n12014 = n154 & n12013 ;
  assign n12015 = n11539 | n11550 ;
  assign n37106 = ~n12015 ;
  assign n12016 = n154 & n37106 ;
  assign n12017 = n11421 | n12016 ;
  assign n37107 = ~n12014 ;
  assign n12018 = n37107 & n12017 ;
  assign n12159 = n37086 & n12140 ;
  assign n12160 = n12032 | n12159 ;
  assign n37108 = ~n12142 ;
  assign n12161 = n37108 & n12160 ;
  assign n37109 = ~n12161 ;
  assign n12162 = n181 & n37109 ;
  assign n12163 = n37096 & n12160 ;
  assign n12164 = n11654 | n12163 ;
  assign n37110 = ~n12162 ;
  assign n12165 = n37110 & n12164 ;
  assign n37111 = ~n12165 ;
  assign n12166 = n182 & n37111 ;
  assign n12167 = n183 | n12166 ;
  assign n37112 = ~n12167 ;
  assign n12168 = n12149 & n37112 ;
  assign n12169 = n12018 | n12168 ;
  assign n37113 = ~n12151 ;
  assign n12170 = n37113 & n12169 ;
  assign n37114 = ~n12170 ;
  assign n12171 = n184 & n37114 ;
  assign n37115 = ~n11543 ;
  assign n12006 = n11415 & n37115 ;
  assign n12007 = n36833 & n12006 ;
  assign n12008 = n154 & n12007 ;
  assign n12009 = n11543 | n11552 ;
  assign n37116 = ~n12009 ;
  assign n12010 = n154 & n37116 ;
  assign n12011 = n11415 | n12010 ;
  assign n37117 = ~n12008 ;
  assign n12012 = n37117 & n12011 ;
  assign n12152 = n838 | n12151 ;
  assign n37118 = ~n12152 ;
  assign n12172 = n37118 & n12169 ;
  assign n12173 = n12012 | n12172 ;
  assign n37119 = ~n12171 ;
  assign n12174 = n37119 & n12173 ;
  assign n37120 = ~n12174 ;
  assign n12175 = n185 & n37120 ;
  assign n11548 = n11408 & n36822 ;
  assign n37121 = ~n11554 ;
  assign n12000 = n11548 & n37121 ;
  assign n12001 = n154 & n12000 ;
  assign n12002 = n11554 | n11565 ;
  assign n37122 = ~n12002 ;
  assign n12003 = n154 & n37122 ;
  assign n12004 = n11408 | n12003 ;
  assign n37123 = ~n12001 ;
  assign n12005 = n37123 & n12004 ;
  assign n12183 = n37102 & n12164 ;
  assign n12184 = n12025 | n12183 ;
  assign n37124 = ~n12166 ;
  assign n12185 = n37124 & n12184 ;
  assign n37125 = ~n12185 ;
  assign n12186 = n183 & n37125 ;
  assign n12187 = n37112 & n12184 ;
  assign n12188 = n12018 | n12187 ;
  assign n37126 = ~n12186 ;
  assign n12189 = n37126 & n12188 ;
  assign n37127 = ~n12189 ;
  assign n12190 = n838 & n37127 ;
  assign n12191 = n185 | n12190 ;
  assign n37128 = ~n12191 ;
  assign n12192 = n12173 & n37128 ;
  assign n12193 = n12005 | n12192 ;
  assign n37129 = ~n12175 ;
  assign n12194 = n37129 & n12193 ;
  assign n37130 = ~n12194 ;
  assign n12195 = n186 & n37130 ;
  assign n37131 = ~n11558 ;
  assign n11993 = n11402 & n37131 ;
  assign n11994 = n36849 & n11993 ;
  assign n11995 = n154 & n11994 ;
  assign n11996 = n11558 | n11567 ;
  assign n37132 = ~n11996 ;
  assign n11997 = n154 & n37132 ;
  assign n11998 = n11402 | n11997 ;
  assign n37133 = ~n11995 ;
  assign n11999 = n37133 & n11998 ;
  assign n12176 = n186 | n12175 ;
  assign n37134 = ~n12176 ;
  assign n12196 = n37134 & n12193 ;
  assign n12197 = n11999 | n12196 ;
  assign n37135 = ~n12195 ;
  assign n12198 = n37135 & n12197 ;
  assign n37136 = ~n12198 ;
  assign n12199 = n528 & n37136 ;
  assign n11563 = n11395 & n36838 ;
  assign n37137 = ~n11569 ;
  assign n11987 = n11563 & n37137 ;
  assign n11988 = n154 & n11987 ;
  assign n11989 = n11569 | n11580 ;
  assign n37138 = ~n11989 ;
  assign n11990 = n154 & n37138 ;
  assign n11991 = n11395 | n11990 ;
  assign n37139 = ~n11988 ;
  assign n11992 = n37139 & n11991 ;
  assign n12207 = n37118 & n12188 ;
  assign n12208 = n12012 | n12207 ;
  assign n37140 = ~n12190 ;
  assign n12209 = n37140 & n12208 ;
  assign n37141 = ~n12209 ;
  assign n12210 = n185 & n37141 ;
  assign n12211 = n37128 & n12208 ;
  assign n12212 = n12005 | n12211 ;
  assign n37142 = ~n12210 ;
  assign n12213 = n37142 & n12212 ;
  assign n37143 = ~n12213 ;
  assign n12214 = n186 & n37143 ;
  assign n12215 = n528 | n12214 ;
  assign n37144 = ~n12215 ;
  assign n12216 = n12197 & n37144 ;
  assign n12217 = n11992 | n12216 ;
  assign n37145 = ~n12199 ;
  assign n12218 = n37145 & n12217 ;
  assign n37146 = ~n12218 ;
  assign n12219 = n188 & n37146 ;
  assign n11980 = n11573 | n11582 ;
  assign n37147 = ~n11980 ;
  assign n11981 = n154 & n37147 ;
  assign n11982 = n11389 | n11981 ;
  assign n37148 = ~n11573 ;
  assign n11983 = n11389 & n37148 ;
  assign n11984 = n36855 & n11983 ;
  assign n11985 = n154 & n11984 ;
  assign n37149 = ~n11985 ;
  assign n11986 = n11982 & n37149 ;
  assign n12200 = n413 | n12199 ;
  assign n37150 = ~n12200 ;
  assign n12220 = n37150 & n12217 ;
  assign n12221 = n11986 | n12220 ;
  assign n37151 = ~n12219 ;
  assign n12222 = n37151 & n12221 ;
  assign n37152 = ~n12222 ;
  assign n12223 = n189 & n37152 ;
  assign n11578 = n11158 & n36870 ;
  assign n37153 = ~n11584 ;
  assign n11974 = n11578 & n37153 ;
  assign n11975 = n154 & n11974 ;
  assign n11976 = n11584 | n11595 ;
  assign n37154 = ~n11976 ;
  assign n11977 = n154 & n37154 ;
  assign n11978 = n11158 | n11977 ;
  assign n37155 = ~n11975 ;
  assign n11979 = n37155 & n11978 ;
  assign n12231 = n37134 & n12212 ;
  assign n12232 = n11999 | n12231 ;
  assign n37156 = ~n12214 ;
  assign n12233 = n37156 & n12232 ;
  assign n37157 = ~n12233 ;
  assign n12234 = n187 & n37157 ;
  assign n12235 = n37144 & n12232 ;
  assign n12236 = n11992 | n12235 ;
  assign n37158 = ~n12234 ;
  assign n12237 = n37158 & n12236 ;
  assign n37159 = ~n12237 ;
  assign n12238 = n413 & n37159 ;
  assign n12239 = n189 | n12238 ;
  assign n37160 = ~n12239 ;
  assign n12240 = n12221 & n37160 ;
  assign n12241 = n11979 | n12240 ;
  assign n37161 = ~n12223 ;
  assign n12242 = n37161 & n12241 ;
  assign n37162 = ~n12242 ;
  assign n12243 = n190 & n37162 ;
  assign n37163 = ~n11588 ;
  assign n11967 = n11382 & n37163 ;
  assign n11968 = n36859 & n11967 ;
  assign n11969 = n154 & n11968 ;
  assign n11970 = n11588 | n11597 ;
  assign n37164 = ~n11970 ;
  assign n11971 = n154 & n37164 ;
  assign n11972 = n11382 | n11971 ;
  assign n37165 = ~n11969 ;
  assign n11973 = n37165 & n11972 ;
  assign n12224 = n190 | n12223 ;
  assign n37166 = ~n12224 ;
  assign n12244 = n37166 & n12241 ;
  assign n12245 = n11973 | n12244 ;
  assign n37167 = ~n12243 ;
  assign n12246 = n37167 & n12245 ;
  assign n37168 = ~n12246 ;
  assign n12247 = n287 & n37168 ;
  assign n37169 = ~n11591 ;
  assign n11593 = n11375 & n37169 ;
  assign n37170 = ~n11601 ;
  assign n11961 = n11593 & n37170 ;
  assign n11962 = n154 & n11961 ;
  assign n11963 = n11600 | n11601 ;
  assign n37171 = ~n11963 ;
  assign n11964 = n154 & n37171 ;
  assign n11965 = n11375 | n11964 ;
  assign n37172 = ~n11962 ;
  assign n11966 = n37172 & n11965 ;
  assign n12255 = n37150 & n12236 ;
  assign n12256 = n11986 | n12255 ;
  assign n37173 = ~n12238 ;
  assign n12257 = n37173 & n12256 ;
  assign n37174 = ~n12257 ;
  assign n12258 = n189 & n37174 ;
  assign n12259 = n37160 & n12256 ;
  assign n12260 = n11979 | n12259 ;
  assign n37175 = ~n12258 ;
  assign n12261 = n37175 & n12260 ;
  assign n37176 = ~n12261 ;
  assign n12262 = n190 & n37176 ;
  assign n12263 = n287 | n12262 ;
  assign n37177 = ~n12263 ;
  assign n12264 = n12245 & n37177 ;
  assign n12267 = n11966 | n12264 ;
  assign n37178 = ~n12247 ;
  assign n12268 = n37178 & n12267 ;
  assign n12271 = n11948 | n12268 ;
  assign n12272 = n31336 & n12271 ;
  assign n11615 = n192 & n11614 ;
  assign n37179 = ~n11150 ;
  assign n11697 = n37179 & n154 ;
  assign n37180 = ~n11697 ;
  assign n11698 = n11611 & n37180 ;
  assign n37181 = ~n11698 ;
  assign n11699 = n11615 & n37181 ;
  assign n11134 = n11121 | n11133 ;
  assign n37182 = ~n11134 ;
  assign n11152 = n37182 & n11149 ;
  assign n11307 = n11152 & n36895 ;
  assign n11949 = n11307 & n36896 ;
  assign n11950 = n36897 & n11949 ;
  assign n11951 = n11699 | n11950 ;
  assign n12248 = n11706 & n37178 ;
  assign n12273 = n12248 & n12267 ;
  assign n12274 = n11951 | n12273 ;
  assign n153 = n12272 | n12274 ;
  assign n12249 = n11966 & n37178 ;
  assign n37183 = ~n12264 ;
  assign n12265 = n12249 & n37183 ;
  assign n12420 = n12265 & n153 ;
  assign n12266 = n12247 | n12264 ;
  assign n37184 = ~n12266 ;
  assign n12421 = n37184 & n153 ;
  assign n12422 = n11966 | n12421 ;
  assign n37185 = ~n12420 ;
  assign n12423 = n37185 & n12422 ;
  assign n12269 = n11706 | n12268 ;
  assign n37186 = ~n12269 ;
  assign n12433 = n37186 & n153 ;
  assign n12693 = n12273 | n12433 ;
  assign n12694 = n12423 | n12693 ;
  assign n200 = x46 | x47 ;
  assign n201 = x48 | n200 ;
  assign n12361 = x48 & n153 ;
  assign n37187 = ~n12361 ;
  assign n12386 = n201 & n37187 ;
  assign n37188 = ~n12386 ;
  assign n12387 = n154 & n37188 ;
  assign n11123 = n201 & n36894 ;
  assign n11308 = n11123 & n36895 ;
  assign n11959 = n11308 & n36896 ;
  assign n11960 = n36897 & n11959 ;
  assign n12362 = n11960 & n37187 ;
  assign n37189 = ~n197 ;
  assign n12309 = n37189 & n153 ;
  assign n37190 = ~x48 ;
  assign n12434 = n37190 & n153 ;
  assign n37191 = ~n12434 ;
  assign n12435 = x49 & n37191 ;
  assign n12436 = n12309 | n12435 ;
  assign n12438 = n12362 | n12436 ;
  assign n37192 = ~n12387 ;
  assign n12439 = n37192 & n12438 ;
  assign n37193 = ~n12439 ;
  assign n12440 = n11067 & n37193 ;
  assign n202 = n37190 & n200 ;
  assign n37194 = ~n153 ;
  assign n12429 = x48 & n37194 ;
  assign n12430 = n202 | n12429 ;
  assign n37195 = ~n12430 ;
  assign n12431 = n154 & n37195 ;
  assign n12432 = n11067 | n12431 ;
  assign n37196 = ~n12432 ;
  assign n12443 = n37196 & n12438 ;
  assign n37197 = ~n11950 ;
  assign n11952 = n154 & n37197 ;
  assign n37198 = ~n11699 ;
  assign n11953 = n37198 & n11952 ;
  assign n37199 = ~n12273 ;
  assign n12446 = n11953 & n37199 ;
  assign n37200 = ~n12272 ;
  assign n12447 = n37200 & n12446 ;
  assign n12448 = n12309 | n12447 ;
  assign n12449 = x50 & n12448 ;
  assign n12450 = x50 | n12447 ;
  assign n12451 = n12309 | n12450 ;
  assign n37201 = ~n12449 ;
  assign n12452 = n37201 & n12451 ;
  assign n12453 = n12443 | n12452 ;
  assign n37202 = ~n12440 ;
  assign n12454 = n37202 & n12453 ;
  assign n37203 = ~n12454 ;
  assign n12455 = n10657 & n37203 ;
  assign n11711 = n11700 | n11709 ;
  assign n37204 = ~n11711 ;
  assign n12350 = n37204 & n153 ;
  assign n12351 = n11714 | n12350 ;
  assign n11717 = n37204 & n11714 ;
  assign n12357 = n11717 & n153 ;
  assign n37205 = ~n12357 ;
  assign n12358 = n12351 & n37205 ;
  assign n12441 = n10657 | n12440 ;
  assign n37206 = ~n12441 ;
  assign n12458 = n37206 & n12453 ;
  assign n12459 = n12358 | n12458 ;
  assign n37207 = ~n12455 ;
  assign n12460 = n37207 & n12459 ;
  assign n37208 = ~n12460 ;
  assign n12461 = n157 & n37208 ;
  assign n37209 = ~n11716 ;
  assign n11750 = n37209 & n11730 ;
  assign n11751 = n36899 & n11750 ;
  assign n12345 = n11751 & n153 ;
  assign n11720 = n11716 | n11719 ;
  assign n37210 = ~n11720 ;
  assign n12347 = n37210 & n153 ;
  assign n12348 = n11730 | n12347 ;
  assign n37211 = ~n12345 ;
  assign n12349 = n37211 & n12348 ;
  assign n12456 = n157 | n12455 ;
  assign n37212 = ~n12456 ;
  assign n12462 = n37212 & n12459 ;
  assign n12463 = n12349 | n12462 ;
  assign n37213 = ~n12461 ;
  assign n12464 = n37213 & n12463 ;
  assign n37214 = ~n12464 ;
  assign n12465 = n158 & n37214 ;
  assign n11749 = n11733 | n11736 ;
  assign n37215 = ~n11749 ;
  assign n12320 = n37215 & n153 ;
  assign n12321 = n11702 | n12320 ;
  assign n11735 = n11702 & n36904 ;
  assign n37216 = ~n11736 ;
  assign n11748 = n11735 & n37216 ;
  assign n12427 = n11748 & n153 ;
  assign n37217 = ~n12427 ;
  assign n12428 = n12321 & n37217 ;
  assign n12442 = n155 & n37193 ;
  assign n12388 = n155 | n12387 ;
  assign n37218 = ~n12388 ;
  assign n12445 = n37218 & n12438 ;
  assign n12475 = n12445 | n12452 ;
  assign n37219 = ~n12442 ;
  assign n12476 = n37219 & n12475 ;
  assign n37220 = ~n12476 ;
  assign n12477 = n156 & n37220 ;
  assign n12478 = n37206 & n12475 ;
  assign n12479 = n12358 | n12478 ;
  assign n37221 = ~n12477 ;
  assign n12480 = n37221 & n12479 ;
  assign n37222 = ~n12480 ;
  assign n12481 = n157 & n37222 ;
  assign n12482 = n158 | n12481 ;
  assign n37223 = ~n12482 ;
  assign n12483 = n12463 & n37223 ;
  assign n12484 = n12428 | n12483 ;
  assign n37224 = ~n12465 ;
  assign n12485 = n37224 & n12484 ;
  assign n37225 = ~n12485 ;
  assign n12486 = n159 & n37225 ;
  assign n37226 = ~n11740 ;
  assign n11746 = n11704 & n37226 ;
  assign n11747 = n36910 & n11746 ;
  assign n12314 = n11747 & n153 ;
  assign n11774 = n11740 | n11758 ;
  assign n37227 = ~n11774 ;
  assign n12322 = n37227 & n153 ;
  assign n12323 = n11704 | n12322 ;
  assign n37228 = ~n12314 ;
  assign n12324 = n37228 & n12323 ;
  assign n12467 = n8857 | n12465 ;
  assign n37229 = ~n12467 ;
  assign n12487 = n37229 & n12484 ;
  assign n12488 = n12324 | n12487 ;
  assign n37230 = ~n12486 ;
  assign n12489 = n37230 & n12488 ;
  assign n37231 = ~n12489 ;
  assign n12490 = n8534 & n37231 ;
  assign n11773 = n11743 | n11760 ;
  assign n37232 = ~n11773 ;
  assign n12298 = n37232 & n153 ;
  assign n12299 = n11692 | n12298 ;
  assign n11745 = n11692 & n36921 ;
  assign n37233 = ~n11760 ;
  assign n11772 = n11745 & n37233 ;
  assign n12353 = n11772 & n153 ;
  assign n37234 = ~n12353 ;
  assign n12354 = n12299 & n37234 ;
  assign n12498 = n37212 & n12479 ;
  assign n12499 = n12349 | n12498 ;
  assign n37235 = ~n12481 ;
  assign n12500 = n37235 & n12499 ;
  assign n37236 = ~n12500 ;
  assign n12501 = n158 & n37236 ;
  assign n12502 = n37223 & n12499 ;
  assign n12503 = n12428 | n12502 ;
  assign n37237 = ~n12501 ;
  assign n12504 = n37237 & n12503 ;
  assign n37238 = ~n12504 ;
  assign n12505 = n8857 & n37238 ;
  assign n12506 = n160 | n12505 ;
  assign n37239 = ~n12506 ;
  assign n12507 = n12488 & n37239 ;
  assign n12508 = n12354 | n12507 ;
  assign n37240 = ~n12490 ;
  assign n12509 = n37240 & n12508 ;
  assign n37241 = ~n12509 ;
  assign n12510 = n161 & n37241 ;
  assign n11798 = n11764 | n11782 ;
  assign n37242 = ~n11798 ;
  assign n12366 = n37242 & n153 ;
  assign n12367 = n11671 | n12366 ;
  assign n37243 = ~n11764 ;
  assign n11770 = n11671 & n37243 ;
  assign n11771 = n36927 & n11770 ;
  assign n12376 = n11771 & n153 ;
  assign n37244 = ~n12376 ;
  assign n12377 = n12367 & n37244 ;
  assign n12491 = n161 | n12490 ;
  assign n37245 = ~n12491 ;
  assign n12511 = n37245 & n12508 ;
  assign n12512 = n12377 | n12511 ;
  assign n37246 = ~n12510 ;
  assign n12513 = n37246 & n12512 ;
  assign n37247 = ~n12513 ;
  assign n12514 = n162 & n37247 ;
  assign n11769 = n11649 & n36937 ;
  assign n37248 = ~n11784 ;
  assign n11796 = n11769 & n37248 ;
  assign n12352 = n11796 & n153 ;
  assign n11797 = n11767 | n11784 ;
  assign n37249 = ~n11797 ;
  assign n12368 = n37249 & n153 ;
  assign n12369 = n11649 | n12368 ;
  assign n37250 = ~n12352 ;
  assign n12370 = n37250 & n12369 ;
  assign n12522 = n37229 & n12503 ;
  assign n12523 = n12324 | n12522 ;
  assign n37251 = ~n12505 ;
  assign n12524 = n37251 & n12523 ;
  assign n37252 = ~n12524 ;
  assign n12525 = n160 & n37252 ;
  assign n12526 = n37239 & n12523 ;
  assign n12527 = n12354 | n12526 ;
  assign n37253 = ~n12525 ;
  assign n12528 = n37253 & n12527 ;
  assign n37254 = ~n12528 ;
  assign n12529 = n161 & n37254 ;
  assign n12530 = n162 | n12529 ;
  assign n37255 = ~n12530 ;
  assign n12531 = n12512 & n37255 ;
  assign n12532 = n12370 | n12531 ;
  assign n37256 = ~n12514 ;
  assign n12533 = n37256 & n12532 ;
  assign n37257 = ~n12533 ;
  assign n12534 = n163 & n37257 ;
  assign n11822 = n11788 | n11806 ;
  assign n37258 = ~n11822 ;
  assign n12325 = n37258 & n153 ;
  assign n12326 = n11644 | n12325 ;
  assign n37259 = ~n11788 ;
  assign n11794 = n11644 & n37259 ;
  assign n11795 = n36943 & n11794 ;
  assign n12374 = n11795 & n153 ;
  assign n37260 = ~n12374 ;
  assign n12375 = n12326 & n37260 ;
  assign n12515 = n6889 | n12514 ;
  assign n37261 = ~n12515 ;
  assign n12535 = n37261 & n12532 ;
  assign n12536 = n12375 | n12535 ;
  assign n37262 = ~n12534 ;
  assign n12537 = n37262 & n12536 ;
  assign n37263 = ~n12537 ;
  assign n12538 = n6600 & n37263 ;
  assign n11793 = n11639 & n36953 ;
  assign n37264 = ~n11808 ;
  assign n11820 = n11793 & n37264 ;
  assign n12340 = n11820 & n153 ;
  assign n11821 = n11791 | n11808 ;
  assign n37265 = ~n11821 ;
  assign n12379 = n37265 & n153 ;
  assign n12380 = n11639 | n12379 ;
  assign n37266 = ~n12340 ;
  assign n12381 = n37266 & n12380 ;
  assign n12546 = n37245 & n12527 ;
  assign n12547 = n12377 | n12546 ;
  assign n37267 = ~n12529 ;
  assign n12548 = n37267 & n12547 ;
  assign n37268 = ~n12548 ;
  assign n12549 = n162 & n37268 ;
  assign n12550 = n37255 & n12547 ;
  assign n12551 = n12370 | n12550 ;
  assign n37269 = ~n12549 ;
  assign n12552 = n37269 & n12551 ;
  assign n37270 = ~n12552 ;
  assign n12553 = n6889 & n37270 ;
  assign n12554 = n6600 | n12553 ;
  assign n37271 = ~n12554 ;
  assign n12555 = n12536 & n37271 ;
  assign n12556 = n12381 | n12555 ;
  assign n37272 = ~n12538 ;
  assign n12557 = n37272 & n12556 ;
  assign n37273 = ~n12557 ;
  assign n12558 = n165 & n37273 ;
  assign n11846 = n11812 | n11830 ;
  assign n37274 = ~n11846 ;
  assign n12341 = n37274 & n153 ;
  assign n12342 = n11661 | n12341 ;
  assign n37275 = ~n11812 ;
  assign n11813 = n11661 & n37275 ;
  assign n11814 = n36959 & n11813 ;
  assign n12343 = n11814 & n153 ;
  assign n37276 = ~n12343 ;
  assign n12344 = n12342 & n37276 ;
  assign n12539 = n165 | n12538 ;
  assign n37277 = ~n12539 ;
  assign n12559 = n37277 & n12556 ;
  assign n12560 = n12344 | n12559 ;
  assign n37278 = ~n12558 ;
  assign n12561 = n37278 & n12560 ;
  assign n37279 = ~n12561 ;
  assign n12562 = n166 & n37279 ;
  assign n11819 = n11663 & n36969 ;
  assign n37280 = ~n11832 ;
  assign n11844 = n11819 & n37280 ;
  assign n12312 = n11844 & n153 ;
  assign n11845 = n11817 | n11832 ;
  assign n37281 = ~n11845 ;
  assign n12327 = n37281 & n153 ;
  assign n12328 = n11663 | n12327 ;
  assign n37282 = ~n12312 ;
  assign n12329 = n37282 & n12328 ;
  assign n12570 = n37261 & n12551 ;
  assign n12571 = n12375 | n12570 ;
  assign n37283 = ~n12553 ;
  assign n12572 = n37283 & n12571 ;
  assign n37284 = ~n12572 ;
  assign n12573 = n164 & n37284 ;
  assign n12574 = n37271 & n12571 ;
  assign n12575 = n12381 | n12574 ;
  assign n37285 = ~n12573 ;
  assign n12576 = n37285 & n12575 ;
  assign n37286 = ~n12576 ;
  assign n12577 = n165 & n37286 ;
  assign n12578 = n166 | n12577 ;
  assign n37287 = ~n12578 ;
  assign n12579 = n12560 & n37287 ;
  assign n12580 = n12329 | n12579 ;
  assign n37288 = ~n12562 ;
  assign n12581 = n37288 & n12580 ;
  assign n37289 = ~n12581 ;
  assign n12582 = n167 & n37289 ;
  assign n11870 = n11836 | n11854 ;
  assign n37290 = ~n11870 ;
  assign n12401 = n37290 & n153 ;
  assign n12402 = n11665 | n12401 ;
  assign n37291 = ~n11836 ;
  assign n11842 = n11665 & n37291 ;
  assign n11843 = n36975 & n11842 ;
  assign n12405 = n11843 & n153 ;
  assign n37292 = ~n12405 ;
  assign n12406 = n12402 & n37292 ;
  assign n12563 = n5352 | n12562 ;
  assign n37293 = ~n12563 ;
  assign n12583 = n37293 & n12580 ;
  assign n12584 = n12406 | n12583 ;
  assign n37294 = ~n12582 ;
  assign n12585 = n37294 & n12584 ;
  assign n37295 = ~n12585 ;
  assign n12586 = n4934 & n37295 ;
  assign n11841 = n11651 & n36985 ;
  assign n37296 = ~n11856 ;
  assign n11869 = n11841 & n37296 ;
  assign n12356 = n11869 & n153 ;
  assign n11868 = n11839 | n11856 ;
  assign n37297 = ~n11868 ;
  assign n12395 = n37297 & n153 ;
  assign n12396 = n11651 | n12395 ;
  assign n37298 = ~n12356 ;
  assign n12397 = n37298 & n12396 ;
  assign n12594 = n37277 & n12575 ;
  assign n12595 = n12344 | n12594 ;
  assign n37299 = ~n12577 ;
  assign n12596 = n37299 & n12595 ;
  assign n37300 = ~n12596 ;
  assign n12597 = n166 & n37300 ;
  assign n12598 = n37287 & n12595 ;
  assign n12599 = n12329 | n12598 ;
  assign n37301 = ~n12597 ;
  assign n12600 = n37301 & n12599 ;
  assign n37302 = ~n12600 ;
  assign n12601 = n5352 & n37302 ;
  assign n12602 = n4934 | n12601 ;
  assign n37303 = ~n12602 ;
  assign n12603 = n12584 & n37303 ;
  assign n12604 = n12397 | n12603 ;
  assign n37304 = ~n12586 ;
  assign n12605 = n37304 & n12604 ;
  assign n37305 = ~n12605 ;
  assign n12606 = n169 & n37305 ;
  assign n37306 = ~n11860 ;
  assign n11866 = n11679 & n37306 ;
  assign n11867 = n36991 & n11866 ;
  assign n12332 = n11867 & n153 ;
  assign n11894 = n11860 | n11878 ;
  assign n37307 = ~n11894 ;
  assign n12398 = n37307 & n153 ;
  assign n12399 = n11679 | n12398 ;
  assign n37308 = ~n12332 ;
  assign n12400 = n37308 & n12399 ;
  assign n12587 = n169 | n12586 ;
  assign n37309 = ~n12587 ;
  assign n12607 = n37309 & n12604 ;
  assign n12608 = n12400 | n12607 ;
  assign n37310 = ~n12606 ;
  assign n12609 = n37310 & n12608 ;
  assign n37311 = ~n12609 ;
  assign n12610 = n170 & n37311 ;
  assign n11865 = n11675 & n37001 ;
  assign n37312 = ~n11880 ;
  assign n11892 = n11865 & n37312 ;
  assign n12355 = n11892 & n153 ;
  assign n11893 = n11863 | n11880 ;
  assign n37313 = ~n11893 ;
  assign n12371 = n37313 & n153 ;
  assign n12372 = n11675 | n12371 ;
  assign n37314 = ~n12355 ;
  assign n12373 = n37314 & n12372 ;
  assign n12618 = n37293 & n12599 ;
  assign n12619 = n12406 | n12618 ;
  assign n37315 = ~n12601 ;
  assign n12620 = n37315 & n12619 ;
  assign n37316 = ~n12620 ;
  assign n12621 = n168 & n37316 ;
  assign n12622 = n37303 & n12619 ;
  assign n12623 = n12397 | n12622 ;
  assign n37317 = ~n12621 ;
  assign n12624 = n37317 & n12623 ;
  assign n37318 = ~n12624 ;
  assign n12625 = n169 & n37318 ;
  assign n12626 = n170 | n12625 ;
  assign n37319 = ~n12626 ;
  assign n12627 = n12608 & n37319 ;
  assign n12628 = n12373 | n12627 ;
  assign n37320 = ~n12610 ;
  assign n12629 = n37320 & n12628 ;
  assign n37321 = ~n12629 ;
  assign n12630 = n171 & n37321 ;
  assign n11918 = n11884 | n11902 ;
  assign n37322 = ~n11918 ;
  assign n12293 = n37322 & n153 ;
  assign n12294 = n11677 | n12293 ;
  assign n37323 = ~n11884 ;
  assign n11890 = n11677 & n37323 ;
  assign n11891 = n37007 & n11890 ;
  assign n12330 = n11891 & n153 ;
  assign n37324 = ~n12330 ;
  assign n12331 = n12294 & n37324 ;
  assign n12611 = n3940 | n12610 ;
  assign n37325 = ~n12611 ;
  assign n12631 = n37325 & n12628 ;
  assign n12632 = n12331 | n12631 ;
  assign n37326 = ~n12630 ;
  assign n12633 = n37326 & n12632 ;
  assign n37327 = ~n12633 ;
  assign n12634 = n3631 & n37327 ;
  assign n11917 = n11887 | n11904 ;
  assign n37328 = ~n11917 ;
  assign n12310 = n37328 & n153 ;
  assign n12311 = n11682 | n12310 ;
  assign n11889 = n11682 & n37017 ;
  assign n37329 = ~n11904 ;
  assign n11916 = n11889 & n37329 ;
  assign n12359 = n11916 & n153 ;
  assign n37330 = ~n12359 ;
  assign n12360 = n12311 & n37330 ;
  assign n12642 = n37309 & n12623 ;
  assign n12643 = n12400 | n12642 ;
  assign n37331 = ~n12625 ;
  assign n12644 = n37331 & n12643 ;
  assign n37332 = ~n12644 ;
  assign n12645 = n170 & n37332 ;
  assign n12646 = n37319 & n12643 ;
  assign n12647 = n12373 | n12646 ;
  assign n37333 = ~n12645 ;
  assign n12648 = n37333 & n12647 ;
  assign n37334 = ~n12648 ;
  assign n12649 = n3940 & n37334 ;
  assign n12650 = n3631 | n12649 ;
  assign n37335 = ~n12650 ;
  assign n12651 = n12632 & n37335 ;
  assign n12652 = n12360 | n12651 ;
  assign n37336 = ~n12634 ;
  assign n12653 = n37336 & n12652 ;
  assign n37337 = ~n12653 ;
  assign n12654 = n173 & n37337 ;
  assign n37338 = ~n11908 ;
  assign n11914 = n11685 & n37338 ;
  assign n11915 = n37023 & n11914 ;
  assign n12290 = n11915 & n153 ;
  assign n11935 = n11908 | n11926 ;
  assign n37339 = ~n11935 ;
  assign n12306 = n37339 & n153 ;
  assign n12307 = n11685 | n12306 ;
  assign n37340 = ~n12290 ;
  assign n12308 = n37340 & n12307 ;
  assign n12635 = n173 | n12634 ;
  assign n37341 = ~n12635 ;
  assign n12655 = n37341 & n12652 ;
  assign n12656 = n12308 | n12655 ;
  assign n37342 = ~n12654 ;
  assign n12657 = n37342 & n12656 ;
  assign n37343 = ~n12657 ;
  assign n12658 = n174 & n37343 ;
  assign n11934 = n11911 | n11928 ;
  assign n37344 = ~n11934 ;
  assign n12288 = n37344 & n153 ;
  assign n12289 = n11630 | n12288 ;
  assign n11912 = n11630 & n37033 ;
  assign n37345 = ~n11928 ;
  assign n11933 = n11912 & n37345 ;
  assign n12338 = n11933 & n153 ;
  assign n37346 = ~n12338 ;
  assign n12339 = n12289 & n37346 ;
  assign n12666 = n37325 & n12647 ;
  assign n12667 = n12331 | n12666 ;
  assign n37347 = ~n12649 ;
  assign n12668 = n37347 & n12667 ;
  assign n37348 = ~n12668 ;
  assign n12669 = n172 & n37348 ;
  assign n12670 = n37335 & n12667 ;
  assign n12671 = n12360 | n12670 ;
  assign n37349 = ~n12669 ;
  assign n12672 = n37349 & n12671 ;
  assign n37350 = ~n12672 ;
  assign n12673 = n173 & n37350 ;
  assign n12674 = n174 | n12673 ;
  assign n37351 = ~n12674 ;
  assign n12675 = n12656 & n37351 ;
  assign n12676 = n12339 | n12675 ;
  assign n37352 = ~n12658 ;
  assign n12677 = n37352 & n12676 ;
  assign n37353 = ~n12677 ;
  assign n12678 = n175 & n37353 ;
  assign n12659 = n2753 | n12658 ;
  assign n37354 = ~n12659 ;
  assign n12679 = n37354 & n12676 ;
  assign n37355 = ~n11932 ;
  assign n12086 = n37355 & n12066 ;
  assign n12087 = n37039 & n12086 ;
  assign n12313 = n12087 & n153 ;
  assign n11945 = n11932 | n11943 ;
  assign n37356 = ~n11945 ;
  assign n12346 = n37356 & n153 ;
  assign n12711 = n12066 | n12346 ;
  assign n37357 = ~n12313 ;
  assign n12712 = n37357 & n12711 ;
  assign n12713 = n12679 | n12712 ;
  assign n37358 = ~n12678 ;
  assign n12714 = n37358 & n12713 ;
  assign n37359 = ~n12714 ;
  assign n12715 = n2431 & n37359 ;
  assign n12085 = n12069 | n12072 ;
  assign n37360 = ~n12085 ;
  assign n12286 = n37360 & n153 ;
  assign n12287 = n12064 | n12286 ;
  assign n12071 = n12064 & n37049 ;
  assign n37361 = ~n12072 ;
  assign n12084 = n12071 & n37361 ;
  assign n12302 = n12084 & n153 ;
  assign n37362 = ~n12302 ;
  assign n12303 = n12287 & n37362 ;
  assign n12683 = n37341 & n12671 ;
  assign n12684 = n12308 | n12683 ;
  assign n37363 = ~n12673 ;
  assign n12685 = n37363 & n12684 ;
  assign n37364 = ~n12685 ;
  assign n12686 = n174 & n37364 ;
  assign n12687 = n37351 & n12684 ;
  assign n12688 = n12339 | n12687 ;
  assign n37365 = ~n12686 ;
  assign n12689 = n37365 & n12688 ;
  assign n37366 = ~n12689 ;
  assign n12690 = n2753 & n37366 ;
  assign n12691 = n2431 | n12690 ;
  assign n37367 = ~n12691 ;
  assign n12718 = n37367 & n12713 ;
  assign n12719 = n12303 | n12718 ;
  assign n37368 = ~n12715 ;
  assign n12720 = n37368 & n12719 ;
  assign n37369 = ~n12720 ;
  assign n12721 = n177 & n37369 ;
  assign n12110 = n12076 | n12094 ;
  assign n37370 = ~n12110 ;
  assign n12284 = n37370 & n153 ;
  assign n12285 = n12058 | n12284 ;
  assign n37371 = ~n12076 ;
  assign n12082 = n12058 & n37371 ;
  assign n12083 = n37055 & n12082 ;
  assign n12296 = n12083 & n153 ;
  assign n37372 = ~n12296 ;
  assign n12297 = n12285 & n37372 ;
  assign n12716 = n177 | n12715 ;
  assign n37373 = ~n12716 ;
  assign n12722 = n37373 & n12719 ;
  assign n12723 = n12297 | n12722 ;
  assign n37374 = ~n12721 ;
  assign n12724 = n37374 & n12723 ;
  assign n37375 = ~n12724 ;
  assign n12725 = n178 & n37375 ;
  assign n12109 = n12079 | n12096 ;
  assign n37376 = ~n12109 ;
  assign n12300 = n37376 & n153 ;
  assign n12301 = n12051 | n12300 ;
  assign n12081 = n12051 & n37065 ;
  assign n37377 = ~n12096 ;
  assign n12108 = n12081 & n37377 ;
  assign n12304 = n12108 & n153 ;
  assign n37378 = ~n12304 ;
  assign n12305 = n12301 & n37378 ;
  assign n12692 = n37354 & n12688 ;
  assign n12735 = n12692 | n12712 ;
  assign n37379 = ~n12690 ;
  assign n12736 = n37379 & n12735 ;
  assign n37380 = ~n12736 ;
  assign n12737 = n176 & n37380 ;
  assign n12738 = n37367 & n12735 ;
  assign n12739 = n12303 | n12738 ;
  assign n37381 = ~n12737 ;
  assign n12740 = n37381 & n12739 ;
  assign n37382 = ~n12740 ;
  assign n12741 = n177 & n37382 ;
  assign n12742 = n178 | n12741 ;
  assign n37383 = ~n12742 ;
  assign n12743 = n12723 & n37383 ;
  assign n12744 = n12305 | n12743 ;
  assign n37384 = ~n12725 ;
  assign n12745 = n37384 & n12744 ;
  assign n37385 = ~n12745 ;
  assign n12746 = n179 & n37385 ;
  assign n12134 = n12100 | n12118 ;
  assign n37386 = ~n12134 ;
  assign n12281 = n37386 & n153 ;
  assign n12282 = n12045 | n12281 ;
  assign n37387 = ~n12100 ;
  assign n12106 = n12045 & n37387 ;
  assign n12107 = n37071 & n12106 ;
  assign n12336 = n12107 & n153 ;
  assign n37388 = ~n12336 ;
  assign n12337 = n12282 & n37388 ;
  assign n12726 = n1707 | n12725 ;
  assign n37389 = ~n12726 ;
  assign n12747 = n37389 & n12744 ;
  assign n12748 = n12337 | n12747 ;
  assign n37390 = ~n12746 ;
  assign n12749 = n37390 & n12748 ;
  assign n37391 = ~n12749 ;
  assign n12750 = n1487 & n37391 ;
  assign n12105 = n12038 & n37081 ;
  assign n37392 = ~n12120 ;
  assign n12132 = n12105 & n37392 ;
  assign n12280 = n12132 & n153 ;
  assign n12133 = n12103 | n12120 ;
  assign n37393 = ~n12133 ;
  assign n12383 = n37393 & n153 ;
  assign n12384 = n12038 | n12383 ;
  assign n37394 = ~n12280 ;
  assign n12385 = n37394 & n12384 ;
  assign n12758 = n37373 & n12739 ;
  assign n12759 = n12297 | n12758 ;
  assign n37395 = ~n12741 ;
  assign n12760 = n37395 & n12759 ;
  assign n37396 = ~n12760 ;
  assign n12761 = n178 & n37396 ;
  assign n12762 = n37383 & n12759 ;
  assign n12763 = n12305 | n12762 ;
  assign n37397 = ~n12761 ;
  assign n12764 = n37397 & n12763 ;
  assign n37398 = ~n12764 ;
  assign n12765 = n1707 & n37398 ;
  assign n12766 = n1487 | n12765 ;
  assign n37399 = ~n12766 ;
  assign n12767 = n12748 & n37399 ;
  assign n12768 = n12385 | n12767 ;
  assign n37400 = ~n12750 ;
  assign n12769 = n37400 & n12768 ;
  assign n37401 = ~n12769 ;
  assign n12770 = n181 & n37401 ;
  assign n37402 = ~n12124 ;
  assign n12130 = n12032 & n37402 ;
  assign n12131 = n37087 & n12130 ;
  assign n12295 = n12131 & n153 ;
  assign n12158 = n12124 | n12142 ;
  assign n37403 = ~n12158 ;
  assign n12317 = n37403 & n153 ;
  assign n12318 = n12032 | n12317 ;
  assign n37404 = ~n12295 ;
  assign n12319 = n37404 & n12318 ;
  assign n12751 = n181 | n12750 ;
  assign n37405 = ~n12751 ;
  assign n12771 = n37405 & n12768 ;
  assign n12772 = n12319 | n12771 ;
  assign n37406 = ~n12770 ;
  assign n12773 = n37406 & n12772 ;
  assign n37407 = ~n12773 ;
  assign n12774 = n182 & n37407 ;
  assign n12129 = n11654 & n37097 ;
  assign n37408 = ~n12144 ;
  assign n12156 = n12129 & n37408 ;
  assign n12279 = n12156 & n153 ;
  assign n12157 = n12127 | n12144 ;
  assign n37409 = ~n12157 ;
  assign n12333 = n37409 & n153 ;
  assign n12334 = n11654 | n12333 ;
  assign n37410 = ~n12279 ;
  assign n12335 = n37410 & n12334 ;
  assign n12782 = n37389 & n12763 ;
  assign n12783 = n12337 | n12782 ;
  assign n37411 = ~n12765 ;
  assign n12784 = n37411 & n12783 ;
  assign n37412 = ~n12784 ;
  assign n12785 = n180 & n37412 ;
  assign n12786 = n37399 & n12783 ;
  assign n12787 = n12385 | n12786 ;
  assign n37413 = ~n12785 ;
  assign n12788 = n37413 & n12787 ;
  assign n37414 = ~n12788 ;
  assign n12789 = n181 & n37414 ;
  assign n12790 = n182 | n12789 ;
  assign n37415 = ~n12790 ;
  assign n12791 = n12772 & n37415 ;
  assign n12792 = n12335 | n12791 ;
  assign n37416 = ~n12774 ;
  assign n12793 = n37416 & n12792 ;
  assign n37417 = ~n12793 ;
  assign n12794 = n183 & n37417 ;
  assign n37418 = ~n12148 ;
  assign n12154 = n12025 & n37418 ;
  assign n12155 = n37103 & n12154 ;
  assign n12276 = n12155 & n153 ;
  assign n12182 = n12148 | n12166 ;
  assign n37419 = ~n12182 ;
  assign n12392 = n37419 & n153 ;
  assign n12393 = n12025 | n12392 ;
  assign n37420 = ~n12276 ;
  assign n12394 = n37420 & n12393 ;
  assign n12775 = n183 | n12774 ;
  assign n37421 = ~n12775 ;
  assign n12795 = n37421 & n12792 ;
  assign n12796 = n12394 | n12795 ;
  assign n37422 = ~n12794 ;
  assign n12797 = n37422 & n12796 ;
  assign n37423 = ~n12797 ;
  assign n12798 = n838 & n37423 ;
  assign n12181 = n12151 | n12168 ;
  assign n37424 = ~n12181 ;
  assign n12407 = n37424 & n153 ;
  assign n12408 = n12018 | n12407 ;
  assign n12153 = n12018 & n37113 ;
  assign n37425 = ~n12168 ;
  assign n12180 = n12153 & n37425 ;
  assign n12409 = n12180 & n153 ;
  assign n37426 = ~n12409 ;
  assign n12410 = n12408 & n37426 ;
  assign n12806 = n37405 & n12787 ;
  assign n12807 = n12319 | n12806 ;
  assign n37427 = ~n12789 ;
  assign n12808 = n37427 & n12807 ;
  assign n37428 = ~n12808 ;
  assign n12809 = n182 & n37428 ;
  assign n12810 = n37415 & n12807 ;
  assign n12811 = n12335 | n12810 ;
  assign n37429 = ~n12809 ;
  assign n12812 = n37429 & n12811 ;
  assign n37430 = ~n12812 ;
  assign n12813 = n996 & n37430 ;
  assign n12814 = n838 | n12813 ;
  assign n37431 = ~n12814 ;
  assign n12815 = n12796 & n37431 ;
  assign n12816 = n12410 | n12815 ;
  assign n37432 = ~n12798 ;
  assign n12817 = n37432 & n12816 ;
  assign n37433 = ~n12817 ;
  assign n12818 = n185 & n37433 ;
  assign n12206 = n12172 | n12190 ;
  assign n37434 = ~n12206 ;
  assign n12291 = n37434 & n153 ;
  assign n12292 = n12012 | n12291 ;
  assign n37435 = ~n12172 ;
  assign n12178 = n12012 & n37435 ;
  assign n12179 = n37119 & n12178 ;
  assign n12315 = n12179 & n153 ;
  assign n37436 = ~n12315 ;
  assign n12316 = n12292 & n37436 ;
  assign n12799 = n185 | n12798 ;
  assign n37437 = ~n12799 ;
  assign n12819 = n37437 & n12816 ;
  assign n12820 = n12316 | n12819 ;
  assign n37438 = ~n12818 ;
  assign n12821 = n37438 & n12820 ;
  assign n37439 = ~n12821 ;
  assign n12822 = n186 & n37439 ;
  assign n12205 = n12175 | n12192 ;
  assign n37440 = ~n12205 ;
  assign n12277 = n37440 & n153 ;
  assign n12278 = n12005 | n12277 ;
  assign n12177 = n12005 & n37129 ;
  assign n37441 = ~n12192 ;
  assign n12204 = n12177 & n37441 ;
  assign n12390 = n12204 & n153 ;
  assign n37442 = ~n12390 ;
  assign n12391 = n12278 & n37442 ;
  assign n12830 = n37421 & n12811 ;
  assign n12831 = n12394 | n12830 ;
  assign n37443 = ~n12813 ;
  assign n12832 = n37443 & n12831 ;
  assign n37444 = ~n12832 ;
  assign n12833 = n184 & n37444 ;
  assign n12834 = n37431 & n12831 ;
  assign n12835 = n12410 | n12834 ;
  assign n37445 = ~n12833 ;
  assign n12836 = n37445 & n12835 ;
  assign n37446 = ~n12836 ;
  assign n12837 = n185 & n37446 ;
  assign n12838 = n186 | n12837 ;
  assign n37447 = ~n12838 ;
  assign n12839 = n12820 & n37447 ;
  assign n12840 = n12391 | n12839 ;
  assign n37448 = ~n12822 ;
  assign n12841 = n37448 & n12840 ;
  assign n37449 = ~n12841 ;
  assign n12842 = n187 & n37449 ;
  assign n12230 = n12196 | n12214 ;
  assign n37450 = ~n12230 ;
  assign n12411 = n37450 & n153 ;
  assign n12412 = n11999 | n12411 ;
  assign n37451 = ~n12196 ;
  assign n12202 = n11999 & n37451 ;
  assign n12203 = n37135 & n12202 ;
  assign n12413 = n12203 & n153 ;
  assign n37452 = ~n12413 ;
  assign n12414 = n12412 & n37452 ;
  assign n12823 = n528 | n12822 ;
  assign n37453 = ~n12823 ;
  assign n12843 = n37453 & n12840 ;
  assign n12844 = n12414 | n12843 ;
  assign n37454 = ~n12842 ;
  assign n12845 = n37454 & n12844 ;
  assign n37455 = ~n12845 ;
  assign n12846 = n413 & n37455 ;
  assign n12201 = n11992 & n37145 ;
  assign n37456 = ~n12216 ;
  assign n12228 = n12201 & n37456 ;
  assign n12382 = n12228 & n153 ;
  assign n12229 = n12199 | n12216 ;
  assign n37457 = ~n12229 ;
  assign n12415 = n37457 & n153 ;
  assign n12416 = n11992 | n12415 ;
  assign n37458 = ~n12382 ;
  assign n12417 = n37458 & n12416 ;
  assign n12854 = n37437 & n12835 ;
  assign n12855 = n12316 | n12854 ;
  assign n37459 = ~n12837 ;
  assign n12856 = n37459 & n12855 ;
  assign n37460 = ~n12856 ;
  assign n12857 = n186 & n37460 ;
  assign n12858 = n37447 & n12855 ;
  assign n12859 = n12391 | n12858 ;
  assign n37461 = ~n12857 ;
  assign n12860 = n37461 & n12859 ;
  assign n37462 = ~n12860 ;
  assign n12861 = n528 & n37462 ;
  assign n12862 = n413 | n12861 ;
  assign n37463 = ~n12862 ;
  assign n12863 = n12844 & n37463 ;
  assign n12864 = n12417 | n12863 ;
  assign n37464 = ~n12846 ;
  assign n12865 = n37464 & n12864 ;
  assign n37465 = ~n12865 ;
  assign n12866 = n189 & n37465 ;
  assign n12254 = n12220 | n12238 ;
  assign n37466 = ~n12254 ;
  assign n12403 = n37466 & n153 ;
  assign n12404 = n11986 | n12403 ;
  assign n37467 = ~n12220 ;
  assign n12226 = n11986 & n37467 ;
  assign n12227 = n37151 & n12226 ;
  assign n12418 = n12227 & n153 ;
  assign n37468 = ~n12418 ;
  assign n12419 = n12404 & n37468 ;
  assign n12847 = n189 | n12846 ;
  assign n37469 = ~n12847 ;
  assign n12867 = n37469 & n12864 ;
  assign n12868 = n12419 | n12867 ;
  assign n37470 = ~n12866 ;
  assign n12869 = n37470 & n12868 ;
  assign n37471 = ~n12869 ;
  assign n12870 = n190 & n37471 ;
  assign n12225 = n11979 & n37161 ;
  assign n37472 = ~n12240 ;
  assign n12252 = n12225 & n37472 ;
  assign n12283 = n12252 & n153 ;
  assign n12253 = n12223 | n12240 ;
  assign n37473 = ~n12253 ;
  assign n12363 = n37473 & n153 ;
  assign n12364 = n11979 | n12363 ;
  assign n37474 = ~n12283 ;
  assign n12365 = n37474 & n12364 ;
  assign n12876 = n37453 & n12859 ;
  assign n12877 = n12414 | n12876 ;
  assign n37475 = ~n12861 ;
  assign n12878 = n37475 & n12877 ;
  assign n37476 = ~n12878 ;
  assign n12879 = n188 & n37476 ;
  assign n12880 = n37463 & n12877 ;
  assign n12881 = n12417 | n12880 ;
  assign n37477 = ~n12879 ;
  assign n12882 = n37477 & n12881 ;
  assign n37478 = ~n12882 ;
  assign n12883 = n189 & n37478 ;
  assign n12884 = n190 | n12883 ;
  assign n37479 = ~n12884 ;
  assign n12885 = n12868 & n37479 ;
  assign n12886 = n12365 | n12885 ;
  assign n37480 = ~n12870 ;
  assign n12891 = n37480 & n12886 ;
  assign n37481 = ~n12891 ;
  assign n12892 = n191 & n37481 ;
  assign n37482 = ~n12244 ;
  assign n12250 = n11973 & n37482 ;
  assign n12251 = n37167 & n12250 ;
  assign n12378 = n12251 & n153 ;
  assign n12707 = n12244 | n12262 ;
  assign n37483 = ~n12707 ;
  assign n12708 = n153 & n37483 ;
  assign n12709 = n11973 | n12708 ;
  assign n37484 = ~n12378 ;
  assign n12710 = n37484 & n12709 ;
  assign n12871 = n191 | n12870 ;
  assign n37485 = ~n12871 ;
  assign n12902 = n37485 & n12886 ;
  assign n12903 = n12710 | n12902 ;
  assign n37486 = ~n12892 ;
  assign n12904 = n37486 & n12903 ;
  assign n12905 = n12694 | n12904 ;
  assign n12906 = n31336 & n12905 ;
  assign n12270 = n192 & n12269 ;
  assign n37487 = ~n11706 ;
  assign n12424 = n37487 & n153 ;
  assign n37488 = ~n12424 ;
  assign n12425 = n12268 & n37488 ;
  assign n37489 = ~n12425 ;
  assign n12426 = n12270 & n37489 ;
  assign n11954 = n11705 | n11950 ;
  assign n37490 = ~n11954 ;
  assign n11955 = n11687 & n37490 ;
  assign n11956 = n37198 & n11955 ;
  assign n12695 = n11956 & n37199 ;
  assign n12696 = n37200 & n12695 ;
  assign n12697 = n12426 | n12696 ;
  assign n12893 = n12423 & n37486 ;
  assign n12912 = n12893 & n12903 ;
  assign n12913 = n12697 | n12912 ;
  assign n152 = n12906 | n12913 ;
  assign n12700 = n12420 | n12696 ;
  assign n37491 = ~n12700 ;
  assign n12701 = n12422 & n37491 ;
  assign n37492 = ~n12426 ;
  assign n12702 = n37492 & n12701 ;
  assign n12872 = n287 | n12870 ;
  assign n37493 = ~n12872 ;
  assign n12887 = n37493 & n12886 ;
  assign n12888 = n12710 | n12887 ;
  assign n12894 = n12888 & n12893 ;
  assign n37494 = ~n12894 ;
  assign n12898 = n12702 & n37494 ;
  assign n37495 = ~n12906 ;
  assign n12909 = n12898 & n37495 ;
  assign n12899 = n12888 & n37486 ;
  assign n12900 = n12423 | n12899 ;
  assign n12901 = n192 & n12900 ;
  assign n37496 = ~n12423 ;
  assign n12923 = n37496 & n152 ;
  assign n37497 = ~n12923 ;
  assign n12924 = n12899 & n37497 ;
  assign n37498 = ~n12924 ;
  assign n12925 = n12901 & n37498 ;
  assign n12926 = n12909 | n12925 ;
  assign n12873 = n12365 & n37480 ;
  assign n37499 = ~n12885 ;
  assign n12889 = n12873 & n37499 ;
  assign n12943 = n12889 & n152 ;
  assign n12890 = n12870 | n12885 ;
  assign n37500 = ~n12890 ;
  assign n12967 = n37500 & n152 ;
  assign n12968 = n12365 | n12967 ;
  assign n37501 = ~n12943 ;
  assign n12969 = n37501 & n12968 ;
  assign n13372 = n37469 & n12881 ;
  assign n37502 = ~n13372 ;
  assign n13373 = n12419 & n37502 ;
  assign n13374 = n37470 & n13373 ;
  assign n13375 = n152 & n13374 ;
  assign n13376 = n12866 | n13372 ;
  assign n37503 = ~n13376 ;
  assign n13377 = n152 & n37503 ;
  assign n13378 = n12419 | n13377 ;
  assign n37504 = ~n13375 ;
  assign n13379 = n37504 & n13378 ;
  assign n37505 = ~n12696 ;
  assign n12698 = n153 & n37505 ;
  assign n12699 = n37492 & n12698 ;
  assign n12896 = n12699 & n37494 ;
  assign n12907 = n12896 & n37495 ;
  assign n12908 = x48 | n12907 ;
  assign n37506 = ~n200 ;
  assign n12988 = n37506 & n152 ;
  assign n12990 = n12908 | n12988 ;
  assign n12991 = n12907 | n12988 ;
  assign n12992 = x48 & n12991 ;
  assign n37507 = ~n12992 ;
  assign n12993 = n12990 & n37507 ;
  assign n37508 = ~x46 ;
  assign n12933 = n37508 & n152 ;
  assign n37509 = ~n12933 ;
  assign n12934 = x47 & n37509 ;
  assign n12989 = n12934 | n12988 ;
  assign n203 = x44 | x45 ;
  assign n204 = x46 | n203 ;
  assign n11957 = n204 & n37197 ;
  assign n11958 = n37198 & n11957 ;
  assign n12705 = n11958 & n37199 ;
  assign n12706 = n37200 & n12705 ;
  assign n12998 = x46 & n152 ;
  assign n37510 = ~n12998 ;
  assign n12999 = n12706 & n37510 ;
  assign n13000 = n12989 | n12999 ;
  assign n13013 = n204 & n37510 ;
  assign n37511 = ~n13013 ;
  assign n13014 = n153 & n37511 ;
  assign n13015 = n154 | n13014 ;
  assign n37512 = ~n13015 ;
  assign n13016 = n13000 & n37512 ;
  assign n13017 = n12993 | n13016 ;
  assign n205 = n37508 & n203 ;
  assign n12895 = n12697 | n12894 ;
  assign n13077 = n12694 | n12899 ;
  assign n13078 = n31336 & n13077 ;
  assign n13079 = n12895 | n13078 ;
  assign n37513 = ~n13079 ;
  assign n13082 = x46 & n37513 ;
  assign n13083 = n205 | n13082 ;
  assign n37514 = ~n13083 ;
  assign n13084 = n153 & n37514 ;
  assign n37515 = ~n13084 ;
  assign n13085 = n13000 & n37515 ;
  assign n37516 = ~n13085 ;
  assign n13086 = n154 & n37516 ;
  assign n37517 = ~n13086 ;
  assign n13087 = n13017 & n37517 ;
  assign n37518 = ~n13087 ;
  assign n13090 = n155 & n37518 ;
  assign n12389 = n12362 | n12387 ;
  assign n37519 = ~n12389 ;
  assign n12921 = n37519 & n152 ;
  assign n12922 = n12436 | n12921 ;
  assign n12437 = n37519 & n12436 ;
  assign n13005 = n12437 & n152 ;
  assign n37520 = ~n13005 ;
  assign n13006 = n12922 & n37520 ;
  assign n13092 = n155 | n13086 ;
  assign n13095 = n154 | n13084 ;
  assign n37521 = ~n13095 ;
  assign n13096 = n13000 & n37521 ;
  assign n13097 = n12993 | n13096 ;
  assign n37522 = ~n13092 ;
  assign n13116 = n37522 & n13097 ;
  assign n13117 = n13006 | n13116 ;
  assign n37523 = ~n13090 ;
  assign n13118 = n37523 & n13117 ;
  assign n37524 = ~n13118 ;
  assign n13119 = n156 & n37524 ;
  assign n12444 = n12442 | n12443 ;
  assign n37525 = ~n12444 ;
  assign n12941 = n37525 & n152 ;
  assign n12942 = n12452 | n12941 ;
  assign n37526 = ~n12443 ;
  assign n12473 = n37526 & n12452 ;
  assign n12474 = n37219 & n12473 ;
  assign n12983 = n12474 & n152 ;
  assign n37527 = ~n12983 ;
  assign n12984 = n12942 & n37527 ;
  assign n13088 = n11067 & n37518 ;
  assign n13089 = n10657 | n13088 ;
  assign n37528 = ~n13089 ;
  assign n13120 = n37528 & n13117 ;
  assign n13121 = n12984 | n13120 ;
  assign n37529 = ~n13119 ;
  assign n13122 = n37529 & n13121 ;
  assign n37530 = ~n13122 ;
  assign n13123 = n157 & n37530 ;
  assign n12472 = n12455 | n12458 ;
  assign n37531 = ~n12472 ;
  assign n13009 = n37531 & n152 ;
  assign n13010 = n12358 | n13009 ;
  assign n12457 = n12358 & n37207 ;
  assign n37532 = ~n12458 ;
  assign n12471 = n12457 & n37532 ;
  assign n13055 = n12471 & n152 ;
  assign n37533 = ~n13055 ;
  assign n13056 = n13010 & n37533 ;
  assign n37534 = ~n13014 ;
  assign n13018 = n13000 & n37534 ;
  assign n37535 = ~n13018 ;
  assign n13019 = n154 & n37535 ;
  assign n13020 = n11067 | n13019 ;
  assign n37536 = ~n13020 ;
  assign n13098 = n37536 & n13097 ;
  assign n13099 = n13006 | n13098 ;
  assign n37537 = ~n13088 ;
  assign n13100 = n37537 & n13099 ;
  assign n37538 = ~n13100 ;
  assign n13101 = n10657 & n37538 ;
  assign n13102 = n157 | n13101 ;
  assign n37539 = ~n13102 ;
  assign n13129 = n37539 & n13121 ;
  assign n13130 = n13056 | n13129 ;
  assign n37540 = ~n13123 ;
  assign n13131 = n37540 & n13130 ;
  assign n37541 = ~n13131 ;
  assign n13132 = n158 & n37541 ;
  assign n13124 = n158 | n13123 ;
  assign n37542 = ~n13124 ;
  assign n13133 = n37542 & n13130 ;
  assign n12470 = n12461 | n12462 ;
  assign n37543 = ~n12470 ;
  assign n12929 = n37543 & n152 ;
  assign n12930 = n12349 | n12929 ;
  assign n37544 = ~n12462 ;
  assign n12468 = n12349 & n37544 ;
  assign n12469 = n37213 & n12468 ;
  assign n13141 = n12469 & n13079 ;
  assign n37545 = ~n13141 ;
  assign n13142 = n12930 & n37545 ;
  assign n13154 = n13133 | n13142 ;
  assign n37546 = ~n13132 ;
  assign n13155 = n37546 & n13154 ;
  assign n37547 = ~n13155 ;
  assign n13156 = n8857 & n37547 ;
  assign n12466 = n12428 & n37224 ;
  assign n37548 = ~n12483 ;
  assign n12496 = n12466 & n37548 ;
  assign n12970 = n12496 & n152 ;
  assign n12497 = n12465 | n12483 ;
  assign n37549 = ~n12497 ;
  assign n13001 = n37549 & n152 ;
  assign n13002 = n12428 | n13001 ;
  assign n37550 = ~n12970 ;
  assign n13003 = n37550 & n13002 ;
  assign n13103 = n37528 & n13099 ;
  assign n13104 = n12984 | n13103 ;
  assign n37551 = ~n13101 ;
  assign n13105 = n37551 & n13104 ;
  assign n37552 = ~n13105 ;
  assign n13106 = n157 & n37552 ;
  assign n13107 = n37539 & n13104 ;
  assign n13108 = n13056 | n13107 ;
  assign n37553 = ~n13106 ;
  assign n13109 = n37553 & n13108 ;
  assign n37554 = ~n13109 ;
  assign n13110 = n158 & n37554 ;
  assign n13111 = n8857 | n13110 ;
  assign n37555 = ~n13111 ;
  assign n13172 = n37555 & n13154 ;
  assign n13173 = n13003 | n13172 ;
  assign n37556 = ~n13156 ;
  assign n13174 = n37556 & n13173 ;
  assign n37557 = ~n13174 ;
  assign n13175 = n160 & n37557 ;
  assign n12495 = n12486 | n12487 ;
  assign n37558 = ~n12495 ;
  assign n12918 = n37558 & n152 ;
  assign n12919 = n12324 | n12918 ;
  assign n37559 = ~n12487 ;
  assign n12493 = n12324 & n37559 ;
  assign n12494 = n37230 & n12493 ;
  assign n12939 = n12494 & n152 ;
  assign n37560 = ~n12939 ;
  assign n12940 = n12919 & n37560 ;
  assign n13157 = n160 | n13156 ;
  assign n37561 = ~n13157 ;
  assign n13176 = n37561 & n13173 ;
  assign n13177 = n12940 | n13176 ;
  assign n37562 = ~n13175 ;
  assign n13178 = n37562 & n13177 ;
  assign n37563 = ~n13178 ;
  assign n13179 = n161 & n37563 ;
  assign n12492 = n12354 & n37240 ;
  assign n37564 = ~n12507 ;
  assign n12520 = n12492 & n37564 ;
  assign n13011 = n12520 & n152 ;
  assign n12521 = n12490 | n12507 ;
  assign n37565 = ~n12521 ;
  assign n13033 = n37565 & n152 ;
  assign n13034 = n12354 | n13033 ;
  assign n37566 = ~n13011 ;
  assign n13035 = n37566 & n13034 ;
  assign n13125 = n13108 & n37542 ;
  assign n13145 = n13125 | n13142 ;
  assign n37567 = ~n13110 ;
  assign n13146 = n37567 & n13145 ;
  assign n37568 = ~n13146 ;
  assign n13147 = n159 & n37568 ;
  assign n13148 = n37555 & n13145 ;
  assign n13149 = n13003 | n13148 ;
  assign n37569 = ~n13147 ;
  assign n13150 = n37569 & n13149 ;
  assign n37570 = ~n13150 ;
  assign n13151 = n8534 & n37570 ;
  assign n13152 = n161 | n13151 ;
  assign n37571 = ~n13152 ;
  assign n13196 = n37571 & n13177 ;
  assign n13197 = n13035 | n13196 ;
  assign n37572 = ~n13179 ;
  assign n13198 = n37572 & n13197 ;
  assign n37573 = ~n13198 ;
  assign n13199 = n162 & n37573 ;
  assign n37574 = ~n12511 ;
  assign n12517 = n12377 & n37574 ;
  assign n12518 = n37246 & n12517 ;
  assign n13027 = n12518 & n152 ;
  assign n12519 = n12510 | n12511 ;
  assign n37575 = ~n12519 ;
  assign n13060 = n37575 & n152 ;
  assign n13061 = n12377 | n13060 ;
  assign n37576 = ~n13027 ;
  assign n13062 = n37576 & n13061 ;
  assign n13180 = n162 | n13179 ;
  assign n37577 = ~n13180 ;
  assign n13200 = n37577 & n13197 ;
  assign n13201 = n13062 | n13200 ;
  assign n37578 = ~n13199 ;
  assign n13202 = n37578 & n13201 ;
  assign n37579 = ~n13202 ;
  assign n13203 = n6889 & n37579 ;
  assign n12545 = n12514 | n12531 ;
  assign n37580 = ~n12545 ;
  assign n12915 = n37580 & n152 ;
  assign n12916 = n12370 | n12915 ;
  assign n12516 = n12370 & n37256 ;
  assign n37581 = ~n12531 ;
  assign n12544 = n12516 & n37581 ;
  assign n12981 = n12544 & n152 ;
  assign n37582 = ~n12981 ;
  assign n12982 = n12916 & n37582 ;
  assign n13158 = n13149 & n37561 ;
  assign n13159 = n12940 | n13158 ;
  assign n37583 = ~n13151 ;
  assign n13160 = n37583 & n13159 ;
  assign n37584 = ~n13160 ;
  assign n13161 = n161 & n37584 ;
  assign n13162 = n37571 & n13159 ;
  assign n13163 = n13035 | n13162 ;
  assign n37585 = ~n13161 ;
  assign n13164 = n37585 & n13163 ;
  assign n37586 = ~n13164 ;
  assign n13165 = n162 & n37586 ;
  assign n13166 = n6889 | n13165 ;
  assign n37587 = ~n13166 ;
  assign n13221 = n37587 & n13201 ;
  assign n13222 = n12982 | n13221 ;
  assign n37588 = ~n13203 ;
  assign n13223 = n37588 & n13222 ;
  assign n37589 = ~n13223 ;
  assign n13224 = n164 & n37589 ;
  assign n12543 = n12534 | n12535 ;
  assign n37590 = ~n12543 ;
  assign n12975 = n37590 & n152 ;
  assign n12976 = n12375 | n12975 ;
  assign n37591 = ~n12535 ;
  assign n12541 = n12375 & n37591 ;
  assign n12542 = n37262 & n12541 ;
  assign n12977 = n12542 & n152 ;
  assign n37592 = ~n12977 ;
  assign n12978 = n12976 & n37592 ;
  assign n13204 = n6600 | n13203 ;
  assign n37593 = ~n13204 ;
  assign n13225 = n37593 & n13222 ;
  assign n13226 = n12978 | n13225 ;
  assign n37594 = ~n13224 ;
  assign n13227 = n37594 & n13226 ;
  assign n37595 = ~n13227 ;
  assign n13228 = n165 & n37595 ;
  assign n12540 = n12381 & n37272 ;
  assign n37596 = ~n12555 ;
  assign n12568 = n12540 & n37596 ;
  assign n12987 = n12568 & n152 ;
  assign n12569 = n12538 | n12555 ;
  assign n37597 = ~n12569 ;
  assign n13065 = n37597 & n152 ;
  assign n13066 = n12381 | n13065 ;
  assign n37598 = ~n12987 ;
  assign n13067 = n37598 & n13066 ;
  assign n13181 = n13163 & n37577 ;
  assign n13182 = n13062 | n13181 ;
  assign n37599 = ~n13165 ;
  assign n13183 = n37599 & n13182 ;
  assign n37600 = ~n13183 ;
  assign n13184 = n163 & n37600 ;
  assign n13185 = n37587 & n13182 ;
  assign n13186 = n12982 | n13185 ;
  assign n37601 = ~n13184 ;
  assign n13187 = n37601 & n13186 ;
  assign n37602 = ~n13187 ;
  assign n13188 = n6600 & n37602 ;
  assign n13189 = n165 | n13188 ;
  assign n37603 = ~n13189 ;
  assign n13244 = n37603 & n13226 ;
  assign n13245 = n13067 | n13244 ;
  assign n37604 = ~n13228 ;
  assign n13246 = n37604 & n13245 ;
  assign n37605 = ~n13246 ;
  assign n13247 = n166 & n37605 ;
  assign n37606 = ~n12559 ;
  assign n12565 = n12344 & n37606 ;
  assign n12566 = n37278 & n12565 ;
  assign n12971 = n12566 & n152 ;
  assign n12567 = n12558 | n12559 ;
  assign n37607 = ~n12567 ;
  assign n13021 = n37607 & n152 ;
  assign n13022 = n12344 | n13021 ;
  assign n37608 = ~n12971 ;
  assign n13023 = n37608 & n13022 ;
  assign n13229 = n166 | n13228 ;
  assign n37609 = ~n13229 ;
  assign n13248 = n37609 & n13245 ;
  assign n13249 = n13023 | n13248 ;
  assign n37610 = ~n13247 ;
  assign n13250 = n37610 & n13249 ;
  assign n37611 = ~n13250 ;
  assign n13251 = n5352 & n37611 ;
  assign n12564 = n12329 & n37288 ;
  assign n37612 = ~n12579 ;
  assign n12592 = n12564 & n37612 ;
  assign n12966 = n12592 & n152 ;
  assign n12593 = n12562 | n12579 ;
  assign n37613 = ~n12593 ;
  assign n13039 = n37613 & n152 ;
  assign n13040 = n12329 | n13039 ;
  assign n37614 = ~n12966 ;
  assign n13041 = n37614 & n13040 ;
  assign n13205 = n13186 & n37593 ;
  assign n13206 = n12978 | n13205 ;
  assign n37615 = ~n13188 ;
  assign n13207 = n37615 & n13206 ;
  assign n37616 = ~n13207 ;
  assign n13208 = n165 & n37616 ;
  assign n13209 = n37603 & n13206 ;
  assign n13210 = n13067 | n13209 ;
  assign n37617 = ~n13208 ;
  assign n13211 = n37617 & n13210 ;
  assign n37618 = ~n13211 ;
  assign n13212 = n166 & n37618 ;
  assign n13213 = n5352 | n13212 ;
  assign n37619 = ~n13213 ;
  assign n13258 = n37619 & n13249 ;
  assign n13259 = n13041 | n13258 ;
  assign n37620 = ~n13251 ;
  assign n13260 = n37620 & n13259 ;
  assign n37621 = ~n13260 ;
  assign n13261 = n168 & n37621 ;
  assign n13252 = n4934 | n13251 ;
  assign n37622 = ~n13252 ;
  assign n13262 = n37622 & n13259 ;
  assign n12591 = n12582 | n12583 ;
  assign n37623 = ~n12591 ;
  assign n13028 = n37623 & n152 ;
  assign n13029 = n12406 | n13028 ;
  assign n37624 = ~n12583 ;
  assign n12589 = n12406 & n37624 ;
  assign n12590 = n37294 & n12589 ;
  assign n13263 = n12590 & n13079 ;
  assign n37625 = ~n13263 ;
  assign n13264 = n13029 & n37625 ;
  assign n13276 = n13262 | n13264 ;
  assign n37626 = ~n13261 ;
  assign n13277 = n37626 & n13276 ;
  assign n37627 = ~n13277 ;
  assign n13278 = n169 & n37627 ;
  assign n12588 = n12397 & n37304 ;
  assign n37628 = ~n12603 ;
  assign n12616 = n12588 & n37628 ;
  assign n13026 = n12616 & n152 ;
  assign n12617 = n12586 | n12603 ;
  assign n37629 = ~n12617 ;
  assign n13071 = n37629 & n152 ;
  assign n13072 = n12397 | n13071 ;
  assign n37630 = ~n13026 ;
  assign n13073 = n37630 & n13072 ;
  assign n13230 = n13210 & n37609 ;
  assign n13231 = n13023 | n13230 ;
  assign n37631 = ~n13212 ;
  assign n13232 = n37631 & n13231 ;
  assign n37632 = ~n13232 ;
  assign n13233 = n167 & n37632 ;
  assign n13234 = n37619 & n13231 ;
  assign n13235 = n13041 | n13234 ;
  assign n37633 = ~n13233 ;
  assign n13236 = n37633 & n13235 ;
  assign n37634 = ~n13236 ;
  assign n13237 = n4934 & n37634 ;
  assign n13238 = n169 | n13237 ;
  assign n37635 = ~n13238 ;
  assign n13295 = n37635 & n13276 ;
  assign n13296 = n13073 | n13295 ;
  assign n37636 = ~n13278 ;
  assign n13297 = n37636 & n13296 ;
  assign n37637 = ~n13297 ;
  assign n13298 = n170 & n37637 ;
  assign n12615 = n12606 | n12607 ;
  assign n37638 = ~n12615 ;
  assign n13007 = n37638 & n152 ;
  assign n13008 = n12400 | n13007 ;
  assign n37639 = ~n12607 ;
  assign n12613 = n12400 & n37639 ;
  assign n12614 = n37310 & n12613 ;
  assign n13042 = n12614 & n152 ;
  assign n37640 = ~n13042 ;
  assign n13043 = n13008 & n37640 ;
  assign n13279 = n170 | n13278 ;
  assign n37641 = ~n13279 ;
  assign n13299 = n37641 & n13296 ;
  assign n13300 = n13043 | n13299 ;
  assign n37642 = ~n13298 ;
  assign n13301 = n37642 & n13300 ;
  assign n37643 = ~n13301 ;
  assign n13302 = n3940 & n37643 ;
  assign n12641 = n12610 | n12627 ;
  assign n37644 = ~n12641 ;
  assign n12996 = n37644 & n152 ;
  assign n12997 = n12373 | n12996 ;
  assign n12612 = n12373 & n37320 ;
  assign n37645 = ~n12627 ;
  assign n12640 = n12612 & n37645 ;
  assign n13024 = n12640 & n152 ;
  assign n37646 = ~n13024 ;
  assign n13025 = n12997 & n37646 ;
  assign n13253 = n13235 & n37622 ;
  assign n13267 = n13253 | n13264 ;
  assign n37647 = ~n13237 ;
  assign n13268 = n37647 & n13267 ;
  assign n37648 = ~n13268 ;
  assign n13269 = n169 & n37648 ;
  assign n13270 = n37635 & n13267 ;
  assign n13271 = n13073 | n13270 ;
  assign n37649 = ~n13269 ;
  assign n13272 = n37649 & n13271 ;
  assign n37650 = ~n13272 ;
  assign n13273 = n170 & n37650 ;
  assign n13274 = n3940 | n13273 ;
  assign n37651 = ~n13274 ;
  assign n13319 = n37651 & n13300 ;
  assign n13320 = n13025 | n13319 ;
  assign n37652 = ~n13302 ;
  assign n13321 = n37652 & n13320 ;
  assign n37653 = ~n13321 ;
  assign n13322 = n172 & n37653 ;
  assign n37654 = ~n12631 ;
  assign n12637 = n12331 & n37654 ;
  assign n12638 = n37326 & n12637 ;
  assign n13051 = n12638 & n152 ;
  assign n12639 = n12630 | n12631 ;
  assign n37655 = ~n12639 ;
  assign n13052 = n37655 & n152 ;
  assign n13053 = n12331 | n13052 ;
  assign n37656 = ~n13051 ;
  assign n13054 = n37656 & n13053 ;
  assign n13303 = n3631 | n13302 ;
  assign n37657 = ~n13303 ;
  assign n13323 = n37657 & n13320 ;
  assign n13324 = n13054 | n13323 ;
  assign n37658 = ~n13322 ;
  assign n13325 = n37658 & n13324 ;
  assign n37659 = ~n13325 ;
  assign n13326 = n173 & n37659 ;
  assign n12636 = n12360 & n37336 ;
  assign n37660 = ~n12651 ;
  assign n12664 = n12636 & n37660 ;
  assign n12937 = n12664 & n152 ;
  assign n12665 = n12634 | n12651 ;
  assign n37661 = ~n12665 ;
  assign n13057 = n37661 & n152 ;
  assign n13058 = n12360 | n13057 ;
  assign n37662 = ~n12937 ;
  assign n13059 = n37662 & n13058 ;
  assign n13280 = n13271 & n37641 ;
  assign n13281 = n13043 | n13280 ;
  assign n37663 = ~n13273 ;
  assign n13282 = n37663 & n13281 ;
  assign n37664 = ~n13282 ;
  assign n13283 = n171 & n37664 ;
  assign n13284 = n37651 & n13281 ;
  assign n13285 = n13025 | n13284 ;
  assign n37665 = ~n13283 ;
  assign n13286 = n37665 & n13285 ;
  assign n37666 = ~n13286 ;
  assign n13287 = n3631 & n37666 ;
  assign n13288 = n173 | n13287 ;
  assign n37667 = ~n13288 ;
  assign n13343 = n37667 & n13324 ;
  assign n13344 = n13059 | n13343 ;
  assign n37668 = ~n13326 ;
  assign n13345 = n37668 & n13344 ;
  assign n37669 = ~n13345 ;
  assign n13346 = n174 & n37669 ;
  assign n37670 = ~n12655 ;
  assign n12661 = n12308 & n37670 ;
  assign n12662 = n37342 & n12661 ;
  assign n12949 = n12662 & n152 ;
  assign n12663 = n12654 | n12655 ;
  assign n37671 = ~n12663 ;
  assign n12972 = n37671 & n152 ;
  assign n12973 = n12308 | n12972 ;
  assign n37672 = ~n12949 ;
  assign n12974 = n37672 & n12973 ;
  assign n13327 = n174 | n13326 ;
  assign n37673 = ~n13327 ;
  assign n13347 = n37673 & n13344 ;
  assign n13348 = n12974 | n13347 ;
  assign n37674 = ~n13346 ;
  assign n13349 = n37674 & n13348 ;
  assign n37675 = ~n13349 ;
  assign n13350 = n2753 & n37675 ;
  assign n12682 = n12658 | n12675 ;
  assign n37676 = ~n12682 ;
  assign n12985 = n37676 & n152 ;
  assign n12986 = n12339 | n12985 ;
  assign n12660 = n12339 & n37352 ;
  assign n37677 = ~n12675 ;
  assign n12681 = n12660 & n37677 ;
  assign n13063 = n12681 & n152 ;
  assign n37678 = ~n13063 ;
  assign n13064 = n12986 & n37678 ;
  assign n13304 = n13285 & n37657 ;
  assign n13305 = n13054 | n13304 ;
  assign n37679 = ~n13287 ;
  assign n13306 = n37679 & n13305 ;
  assign n37680 = ~n13306 ;
  assign n13307 = n173 & n37680 ;
  assign n13308 = n37667 & n13305 ;
  assign n13309 = n13059 | n13308 ;
  assign n37681 = ~n13307 ;
  assign n13310 = n37681 & n13309 ;
  assign n37682 = ~n13310 ;
  assign n13311 = n174 & n37682 ;
  assign n13312 = n2753 | n13311 ;
  assign n37683 = ~n13312 ;
  assign n13356 = n37683 & n13348 ;
  assign n13357 = n13064 | n13356 ;
  assign n37684 = ~n13350 ;
  assign n13358 = n37684 & n13357 ;
  assign n37685 = ~n13358 ;
  assign n13359 = n176 & n37685 ;
  assign n13351 = n2431 | n13350 ;
  assign n37686 = ~n13351 ;
  assign n13360 = n37686 & n13357 ;
  assign n37687 = ~n12679 ;
  assign n12733 = n37687 & n12712 ;
  assign n12734 = n37358 & n12733 ;
  assign n12917 = n12734 & n152 ;
  assign n12680 = n12678 | n12679 ;
  assign n37688 = ~n12680 ;
  assign n13012 = n37688 & n152 ;
  assign n13380 = n12712 | n13012 ;
  assign n37689 = ~n12917 ;
  assign n13381 = n37689 & n13380 ;
  assign n13382 = n13360 | n13381 ;
  assign n37690 = ~n13359 ;
  assign n13383 = n37690 & n13382 ;
  assign n37691 = ~n13383 ;
  assign n13384 = n177 & n37691 ;
  assign n12717 = n12303 & n37368 ;
  assign n37692 = ~n12718 ;
  assign n12731 = n12717 & n37692 ;
  assign n13004 = n12731 & n152 ;
  assign n12732 = n12715 | n12718 ;
  assign n37693 = ~n12732 ;
  assign n13048 = n37693 & n152 ;
  assign n13049 = n12303 | n13048 ;
  assign n37694 = ~n13004 ;
  assign n13050 = n37694 & n13049 ;
  assign n13328 = n13309 & n37673 ;
  assign n13329 = n12974 | n13328 ;
  assign n37695 = ~n13311 ;
  assign n13330 = n37695 & n13329 ;
  assign n37696 = ~n13330 ;
  assign n13331 = n175 & n37696 ;
  assign n13332 = n37683 & n13329 ;
  assign n13333 = n13064 | n13332 ;
  assign n37697 = ~n13331 ;
  assign n13334 = n37697 & n13333 ;
  assign n37698 = ~n13334 ;
  assign n13335 = n2431 & n37698 ;
  assign n13336 = n177 | n13335 ;
  assign n37699 = ~n13336 ;
  assign n13387 = n37699 & n13382 ;
  assign n13388 = n13050 | n13387 ;
  assign n37700 = ~n13384 ;
  assign n13389 = n37700 & n13388 ;
  assign n37701 = ~n13389 ;
  assign n13390 = n178 & n37701 ;
  assign n12730 = n12721 | n12722 ;
  assign n37702 = ~n12730 ;
  assign n13044 = n37702 & n152 ;
  assign n13045 = n12297 | n13044 ;
  assign n37703 = ~n12722 ;
  assign n12728 = n12297 & n37703 ;
  assign n12729 = n37374 & n12728 ;
  assign n13069 = n12729 & n152 ;
  assign n37704 = ~n13069 ;
  assign n13070 = n13045 & n37704 ;
  assign n13385 = n178 | n13384 ;
  assign n37705 = ~n13385 ;
  assign n13391 = n37705 & n13388 ;
  assign n13392 = n13070 | n13391 ;
  assign n37706 = ~n13390 ;
  assign n13393 = n37706 & n13392 ;
  assign n37707 = ~n13393 ;
  assign n13394 = n1707 & n37707 ;
  assign n12727 = n12305 & n37384 ;
  assign n37708 = ~n12743 ;
  assign n12756 = n12727 & n37708 ;
  assign n12928 = n12756 & n152 ;
  assign n12757 = n12725 | n12743 ;
  assign n37709 = ~n12757 ;
  assign n13030 = n37709 & n152 ;
  assign n13031 = n12305 | n13030 ;
  assign n37710 = ~n12928 ;
  assign n13032 = n37710 & n13031 ;
  assign n13352 = n13333 & n37686 ;
  assign n13399 = n13352 | n13381 ;
  assign n37711 = ~n13335 ;
  assign n13400 = n37711 & n13399 ;
  assign n37712 = ~n13400 ;
  assign n13401 = n177 & n37712 ;
  assign n13402 = n37699 & n13399 ;
  assign n13403 = n13050 | n13402 ;
  assign n37713 = ~n13401 ;
  assign n13404 = n37713 & n13403 ;
  assign n37714 = ~n13404 ;
  assign n13405 = n178 & n37714 ;
  assign n13406 = n1707 | n13405 ;
  assign n37715 = ~n13406 ;
  assign n13407 = n13392 & n37715 ;
  assign n13408 = n13032 | n13407 ;
  assign n37716 = ~n13394 ;
  assign n13409 = n37716 & n13408 ;
  assign n37717 = ~n13409 ;
  assign n13410 = n180 & n37717 ;
  assign n37718 = ~n12747 ;
  assign n12753 = n12337 & n37718 ;
  assign n12754 = n37390 & n12753 ;
  assign n12920 = n12754 & n152 ;
  assign n12755 = n12746 | n12747 ;
  assign n37719 = ~n12755 ;
  assign n13036 = n37719 & n152 ;
  assign n13037 = n12337 | n13036 ;
  assign n37720 = ~n12920 ;
  assign n13038 = n37720 & n13037 ;
  assign n13395 = n1487 | n13394 ;
  assign n37721 = ~n13395 ;
  assign n13411 = n37721 & n13408 ;
  assign n13412 = n13038 | n13411 ;
  assign n37722 = ~n13410 ;
  assign n13413 = n37722 & n13412 ;
  assign n37723 = ~n13413 ;
  assign n13414 = n181 & n37723 ;
  assign n12780 = n12750 | n12767 ;
  assign n37724 = ~n12780 ;
  assign n12979 = n37724 & n152 ;
  assign n12980 = n12385 | n12979 ;
  assign n12752 = n12385 & n37400 ;
  assign n37725 = ~n12767 ;
  assign n12781 = n12752 & n37725 ;
  assign n12994 = n12781 & n152 ;
  assign n37726 = ~n12994 ;
  assign n12995 = n12980 & n37726 ;
  assign n13417 = n37705 & n13403 ;
  assign n13418 = n13070 | n13417 ;
  assign n37727 = ~n13405 ;
  assign n13419 = n37727 & n13418 ;
  assign n37728 = ~n13419 ;
  assign n13420 = n179 & n37728 ;
  assign n13421 = n37715 & n13418 ;
  assign n13422 = n13032 | n13421 ;
  assign n37729 = ~n13420 ;
  assign n13423 = n37729 & n13422 ;
  assign n37730 = ~n13423 ;
  assign n13424 = n1487 & n37730 ;
  assign n13425 = n181 | n13424 ;
  assign n37731 = ~n13425 ;
  assign n13426 = n13412 & n37731 ;
  assign n13427 = n12995 | n13426 ;
  assign n37732 = ~n13414 ;
  assign n13428 = n37732 & n13427 ;
  assign n37733 = ~n13428 ;
  assign n13429 = n182 & n37733 ;
  assign n37734 = ~n12771 ;
  assign n12777 = n12319 & n37734 ;
  assign n12778 = n37406 & n12777 ;
  assign n13068 = n12778 & n152 ;
  assign n12779 = n12770 | n12771 ;
  assign n37735 = ~n12779 ;
  assign n13074 = n37735 & n152 ;
  assign n13075 = n12319 | n13074 ;
  assign n37736 = ~n13068 ;
  assign n13076 = n37736 & n13075 ;
  assign n13415 = n182 | n13414 ;
  assign n37737 = ~n13415 ;
  assign n13430 = n37737 & n13427 ;
  assign n13431 = n13076 | n13430 ;
  assign n37738 = ~n13429 ;
  assign n13432 = n37738 & n13431 ;
  assign n37739 = ~n13432 ;
  assign n13433 = n996 & n37739 ;
  assign n12805 = n12774 | n12791 ;
  assign n37740 = ~n12805 ;
  assign n12962 = n37740 & n152 ;
  assign n12963 = n12335 | n12962 ;
  assign n12776 = n12335 & n37416 ;
  assign n37741 = ~n12791 ;
  assign n12804 = n12776 & n37741 ;
  assign n12964 = n12804 & n152 ;
  assign n37742 = ~n12964 ;
  assign n12965 = n12963 & n37742 ;
  assign n13436 = n37721 & n13422 ;
  assign n13437 = n13038 | n13436 ;
  assign n37743 = ~n13424 ;
  assign n13438 = n37743 & n13437 ;
  assign n37744 = ~n13438 ;
  assign n13439 = n181 & n37744 ;
  assign n13440 = n37731 & n13437 ;
  assign n13441 = n12995 | n13440 ;
  assign n37745 = ~n13439 ;
  assign n13442 = n37745 & n13441 ;
  assign n37746 = ~n13442 ;
  assign n13443 = n182 & n37746 ;
  assign n13444 = n183 | n13443 ;
  assign n37747 = ~n13444 ;
  assign n13445 = n13431 & n37747 ;
  assign n13446 = n12965 | n13445 ;
  assign n37748 = ~n13433 ;
  assign n13447 = n37748 & n13446 ;
  assign n37749 = ~n13447 ;
  assign n13448 = n184 & n37749 ;
  assign n12803 = n12794 | n12795 ;
  assign n37750 = ~n12803 ;
  assign n12954 = n37750 & n152 ;
  assign n12955 = n12394 | n12954 ;
  assign n37751 = ~n12795 ;
  assign n12801 = n12394 & n37751 ;
  assign n12802 = n37422 & n12801 ;
  assign n12960 = n12802 & n152 ;
  assign n37752 = ~n12960 ;
  assign n12961 = n12955 & n37752 ;
  assign n13434 = n838 | n13433 ;
  assign n37753 = ~n13434 ;
  assign n13449 = n37753 & n13446 ;
  assign n13450 = n12961 | n13449 ;
  assign n37754 = ~n13448 ;
  assign n13451 = n37754 & n13450 ;
  assign n37755 = ~n13451 ;
  assign n13452 = n185 & n37755 ;
  assign n12829 = n12798 | n12815 ;
  assign n37756 = ~n12829 ;
  assign n12952 = n37756 & n152 ;
  assign n12953 = n12410 | n12952 ;
  assign n12800 = n12410 & n37432 ;
  assign n37757 = ~n12815 ;
  assign n12828 = n12800 & n37757 ;
  assign n13139 = n12828 & n13079 ;
  assign n37758 = ~n13139 ;
  assign n13140 = n12953 & n37758 ;
  assign n13455 = n37737 & n13441 ;
  assign n13456 = n13076 | n13455 ;
  assign n37759 = ~n13443 ;
  assign n13457 = n37759 & n13456 ;
  assign n37760 = ~n13457 ;
  assign n13458 = n183 & n37760 ;
  assign n13459 = n37747 & n13456 ;
  assign n13462 = n12965 | n13459 ;
  assign n37761 = ~n13458 ;
  assign n13463 = n37761 & n13462 ;
  assign n37762 = ~n13463 ;
  assign n13464 = n838 & n37762 ;
  assign n13465 = n185 | n13464 ;
  assign n37763 = ~n13465 ;
  assign n13466 = n13450 & n37763 ;
  assign n13467 = n13140 | n13466 ;
  assign n37764 = ~n13452 ;
  assign n13468 = n37764 & n13467 ;
  assign n37765 = ~n13468 ;
  assign n13469 = n186 & n37765 ;
  assign n12827 = n12818 | n12819 ;
  assign n37766 = ~n12827 ;
  assign n13046 = n37766 & n152 ;
  assign n13047 = n12316 | n13046 ;
  assign n37767 = ~n12819 ;
  assign n12825 = n12316 & n37767 ;
  assign n12826 = n37438 & n12825 ;
  assign n13080 = n12826 & n13079 ;
  assign n37768 = ~n13080 ;
  assign n13081 = n13047 & n37768 ;
  assign n13453 = n186 | n13452 ;
  assign n37769 = ~n13453 ;
  assign n13470 = n37769 & n13467 ;
  assign n13471 = n13081 | n13470 ;
  assign n37770 = ~n13469 ;
  assign n13472 = n37770 & n13471 ;
  assign n37771 = ~n13472 ;
  assign n13473 = n528 & n37771 ;
  assign n12853 = n12822 | n12839 ;
  assign n37772 = ~n12853 ;
  assign n12956 = n37772 & n152 ;
  assign n12957 = n12391 | n12956 ;
  assign n12824 = n12391 & n37448 ;
  assign n37773 = ~n12839 ;
  assign n12852 = n12824 & n37773 ;
  assign n12958 = n12852 & n152 ;
  assign n37774 = ~n12958 ;
  assign n12959 = n12957 & n37774 ;
  assign n13476 = n37753 & n13462 ;
  assign n13477 = n12961 | n13476 ;
  assign n37775 = ~n13464 ;
  assign n13478 = n37775 & n13477 ;
  assign n37776 = ~n13478 ;
  assign n13479 = n185 & n37776 ;
  assign n13480 = n37763 & n13477 ;
  assign n13481 = n13140 | n13480 ;
  assign n37777 = ~n13479 ;
  assign n13482 = n37777 & n13481 ;
  assign n37778 = ~n13482 ;
  assign n13483 = n186 & n37778 ;
  assign n13484 = n528 | n13483 ;
  assign n37779 = ~n13484 ;
  assign n13485 = n13471 & n37779 ;
  assign n13486 = n12959 | n13485 ;
  assign n37780 = ~n13473 ;
  assign n13487 = n37780 & n13486 ;
  assign n37781 = ~n13487 ;
  assign n13488 = n188 & n37781 ;
  assign n12851 = n12842 | n12843 ;
  assign n37782 = ~n12851 ;
  assign n12947 = n37782 & n152 ;
  assign n12948 = n12414 | n12947 ;
  assign n37783 = ~n12843 ;
  assign n12849 = n12414 & n37783 ;
  assign n12850 = n37454 & n12849 ;
  assign n12950 = n12850 & n152 ;
  assign n37784 = ~n12950 ;
  assign n12951 = n12948 & n37784 ;
  assign n13474 = n413 | n13473 ;
  assign n37785 = ~n13474 ;
  assign n13489 = n37785 & n13486 ;
  assign n13490 = n12951 | n13489 ;
  assign n37786 = ~n13488 ;
  assign n13491 = n37786 & n13490 ;
  assign n37787 = ~n13491 ;
  assign n13492 = n189 & n37787 ;
  assign n13493 = n190 | n13492 ;
  assign n12848 = n12417 & n37464 ;
  assign n37788 = ~n12863 ;
  assign n12874 = n12848 & n37788 ;
  assign n12938 = n12874 & n152 ;
  assign n12875 = n12846 | n12863 ;
  assign n37789 = ~n12875 ;
  assign n12944 = n37789 & n152 ;
  assign n12945 = n12417 | n12944 ;
  assign n37790 = ~n12938 ;
  assign n12946 = n37790 & n12945 ;
  assign n13495 = n37769 & n13481 ;
  assign n13496 = n13081 | n13495 ;
  assign n37791 = ~n13483 ;
  assign n13497 = n37791 & n13496 ;
  assign n37792 = ~n13497 ;
  assign n13498 = n187 & n37792 ;
  assign n13499 = n37779 & n13496 ;
  assign n13500 = n12959 | n13499 ;
  assign n37793 = ~n13498 ;
  assign n13501 = n37793 & n13500 ;
  assign n37794 = ~n13501 ;
  assign n13502 = n413 & n37794 ;
  assign n13503 = n189 | n13502 ;
  assign n13504 = n37785 & n13500 ;
  assign n13505 = n12951 | n13504 ;
  assign n37795 = ~n13503 ;
  assign n13508 = n37795 & n13505 ;
  assign n13509 = n12946 | n13508 ;
  assign n37796 = ~n13493 ;
  assign n13510 = n37796 & n13509 ;
  assign n13511 = n13379 | n13510 ;
  assign n37797 = ~n13502 ;
  assign n13506 = n37797 & n13505 ;
  assign n37798 = ~n13506 ;
  assign n13507 = n189 & n37798 ;
  assign n37799 = ~n13507 ;
  assign n13513 = n37799 & n13509 ;
  assign n37800 = ~n13513 ;
  assign n13514 = n190 & n37800 ;
  assign n13516 = n287 | n13514 ;
  assign n37801 = ~n13516 ;
  assign n13517 = n13511 & n37801 ;
  assign n13518 = n12969 | n13517 ;
  assign n37802 = ~n12902 ;
  assign n13361 = n12710 & n37802 ;
  assign n13362 = n37486 & n13361 ;
  assign n13363 = n152 & n13362 ;
  assign n13365 = n12892 | n12902 ;
  assign n37803 = ~n13365 ;
  assign n13366 = n152 & n37803 ;
  assign n13367 = n12710 | n13366 ;
  assign n37804 = ~n13363 ;
  assign n13368 = n37804 & n13367 ;
  assign n37805 = ~n13514 ;
  assign n13521 = n13511 & n37805 ;
  assign n37806 = ~n13521 ;
  assign n13522 = n191 & n37806 ;
  assign n37807 = ~n13522 ;
  assign n13523 = n13368 & n37807 ;
  assign n13524 = n13518 & n13523 ;
  assign n13525 = n12926 | n13524 ;
  assign n37808 = ~n12900 ;
  assign n12935 = n37808 & n152 ;
  assign n12936 = n12894 | n12935 ;
  assign n13369 = n12936 | n13368 ;
  assign n13530 = n13518 & n37807 ;
  assign n13660 = n13369 | n13530 ;
  assign n13661 = n31336 & n13660 ;
  assign n13662 = n13525 | n13661 ;
  assign n13531 = n13368 | n13530 ;
  assign n13515 = n191 | n13514 ;
  assign n37809 = ~n13515 ;
  assign n13533 = n13511 & n37809 ;
  assign n13534 = n12969 | n13533 ;
  assign n13535 = n37807 & n13534 ;
  assign n13536 = n13369 | n13535 ;
  assign n13537 = n31336 & n13536 ;
  assign n13538 = n13523 & n13534 ;
  assign n13539 = n12926 | n13538 ;
  assign n151 = n13537 | n13539 ;
  assign n37810 = ~n13531 ;
  assign n13610 = n37810 & n151 ;
  assign n13611 = n13524 | n13610 ;
  assign n13529 = n12969 & n37807 ;
  assign n37811 = ~n13533 ;
  assign n13653 = n13529 & n37811 ;
  assign n13654 = n151 & n13653 ;
  assign n13655 = n13522 | n13533 ;
  assign n37812 = ~n13655 ;
  assign n13656 = n151 & n37812 ;
  assign n13657 = n12969 | n13656 ;
  assign n37813 = ~n13654 ;
  assign n13658 = n37813 & n13657 ;
  assign n13659 = n13611 | n13658 ;
  assign n13520 = n13510 | n13514 ;
  assign n37814 = ~n13520 ;
  assign n13649 = n37814 & n151 ;
  assign n13650 = n13379 | n13649 ;
  assign n37815 = ~n13510 ;
  assign n13512 = n13379 & n37815 ;
  assign n13519 = n13512 & n37805 ;
  assign n13651 = n13519 & n151 ;
  assign n37816 = ~n13651 ;
  assign n13652 = n13650 & n37816 ;
  assign n37817 = ~x44 ;
  assign n13556 = n37817 & n151 ;
  assign n37818 = ~n13556 ;
  assign n13557 = x45 & n37818 ;
  assign n37819 = ~n203 ;
  assign n13616 = n37819 & n151 ;
  assign n13631 = n13557 | n13616 ;
  assign n206 = x42 | x43 ;
  assign n207 = x44 | n206 ;
  assign n12703 = n207 & n37505 ;
  assign n12704 = n37492 & n12703 ;
  assign n12897 = n12704 & n37494 ;
  assign n12911 = n12897 & n37495 ;
  assign n13600 = x44 & n151 ;
  assign n37820 = ~n13600 ;
  assign n13634 = n12911 & n37820 ;
  assign n13635 = n13631 | n13634 ;
  assign n208 = n37817 & n206 ;
  assign n37821 = ~n13662 ;
  assign n13663 = x44 & n37821 ;
  assign n13664 = n208 | n13663 ;
  assign n37822 = ~n13664 ;
  assign n13665 = n13079 & n37822 ;
  assign n37823 = ~n13665 ;
  assign n13666 = n13635 & n37823 ;
  assign n37824 = ~n13666 ;
  assign n13667 = n153 & n37824 ;
  assign n13601 = n207 & n37820 ;
  assign n37825 = ~n13601 ;
  assign n13602 = n152 & n37825 ;
  assign n13603 = n153 | n13602 ;
  assign n37826 = ~n13603 ;
  assign n13636 = n37826 & n13635 ;
  assign n37827 = ~n12909 ;
  assign n12931 = n37827 & n152 ;
  assign n37828 = ~n12925 ;
  assign n12932 = n37828 & n12931 ;
  assign n37829 = ~n13524 ;
  assign n13526 = n12932 & n37829 ;
  assign n37830 = ~n13661 ;
  assign n13684 = n13526 & n37830 ;
  assign n13685 = n13616 | n13684 ;
  assign n13686 = x46 & n13685 ;
  assign n13687 = x46 | n13684 ;
  assign n13688 = n13616 | n13687 ;
  assign n37831 = ~n13686 ;
  assign n13689 = n37831 & n13688 ;
  assign n13690 = n13636 | n13689 ;
  assign n37832 = ~n13667 ;
  assign n13691 = n37832 & n13690 ;
  assign n37833 = ~n13691 ;
  assign n13692 = n154 & n37833 ;
  assign n13093 = n12999 | n13084 ;
  assign n37834 = ~n13093 ;
  assign n13094 = n12989 & n37834 ;
  assign n13541 = n13094 & n151 ;
  assign n13597 = n37834 & n151 ;
  assign n13598 = n12989 | n13597 ;
  assign n37835 = ~n13541 ;
  assign n13599 = n37835 & n13598 ;
  assign n13668 = n154 | n13667 ;
  assign n13669 = n153 | n13665 ;
  assign n37836 = ~n13669 ;
  assign n13670 = n13635 & n37836 ;
  assign n13697 = n13670 | n13689 ;
  assign n37837 = ~n13668 ;
  assign n13716 = n37837 & n13697 ;
  assign n13717 = n13599 | n13716 ;
  assign n37838 = ~n13692 ;
  assign n13718 = n37838 & n13717 ;
  assign n37839 = ~n13718 ;
  assign n13719 = n155 & n37839 ;
  assign n37840 = ~n13096 ;
  assign n13137 = n12993 & n37840 ;
  assign n37841 = ~n13019 ;
  assign n13138 = n37841 & n13137 ;
  assign n13547 = n13138 & n151 ;
  assign n13136 = n13019 | n13096 ;
  assign n37842 = ~n13136 ;
  assign n13588 = n37842 & n151 ;
  assign n13589 = n12993 | n13588 ;
  assign n37843 = ~n13547 ;
  assign n13590 = n37843 & n13589 ;
  assign n13694 = n11067 | n13692 ;
  assign n37844 = ~n13694 ;
  assign n13720 = n37844 & n13717 ;
  assign n13721 = n13590 | n13720 ;
  assign n37845 = ~n13719 ;
  assign n13722 = n37845 & n13721 ;
  assign n37846 = ~n13722 ;
  assign n13723 = n10657 & n37846 ;
  assign n13135 = n13090 | n13098 ;
  assign n37847 = ~n13135 ;
  assign n13573 = n37847 & n151 ;
  assign n13574 = n13006 | n13573 ;
  assign n13091 = n13006 & n37523 ;
  assign n37848 = ~n13098 ;
  assign n13134 = n13091 & n37848 ;
  assign n13608 = n13134 & n151 ;
  assign n37849 = ~n13608 ;
  assign n13609 = n13574 & n37849 ;
  assign n13671 = n152 & n37822 ;
  assign n37850 = ~n13671 ;
  assign n13672 = n13635 & n37850 ;
  assign n37851 = ~n13672 ;
  assign n13673 = n153 & n37851 ;
  assign n13674 = n154 | n13673 ;
  assign n37852 = ~n13674 ;
  assign n13698 = n37852 & n13697 ;
  assign n13699 = n13599 | n13698 ;
  assign n13700 = n37838 & n13699 ;
  assign n37853 = ~n13700 ;
  assign n13701 = n11067 & n37853 ;
  assign n13702 = n10657 | n13701 ;
  assign n37854 = ~n13702 ;
  assign n13740 = n37854 & n13721 ;
  assign n13741 = n13609 | n13740 ;
  assign n37855 = ~n13723 ;
  assign n13742 = n37855 & n13741 ;
  assign n37856 = ~n13742 ;
  assign n13743 = n157 & n37856 ;
  assign n13115 = n13101 | n13103 ;
  assign n37857 = ~n13115 ;
  assign n13586 = n37857 & n151 ;
  assign n13587 = n12984 | n13586 ;
  assign n37858 = ~n13103 ;
  assign n13113 = n12984 & n37858 ;
  assign n13114 = n37551 & n13113 ;
  assign n13678 = n13114 & n13662 ;
  assign n37859 = ~n13678 ;
  assign n13679 = n13587 & n37859 ;
  assign n13724 = n157 | n13723 ;
  assign n37860 = ~n13724 ;
  assign n13744 = n37860 & n13741 ;
  assign n13745 = n13679 | n13744 ;
  assign n37861 = ~n13743 ;
  assign n13746 = n37861 & n13745 ;
  assign n37862 = ~n13746 ;
  assign n13747 = n158 & n37862 ;
  assign n13127 = n13056 & n37540 ;
  assign n37863 = ~n13107 ;
  assign n13128 = n37863 & n13127 ;
  assign n13572 = n13128 & n151 ;
  assign n13112 = n13106 | n13107 ;
  assign n37864 = ~n13112 ;
  assign n13605 = n37864 & n151 ;
  assign n13606 = n13056 | n13605 ;
  assign n37865 = ~n13572 ;
  assign n13607 = n37865 & n13606 ;
  assign n13703 = n37844 & n13699 ;
  assign n13704 = n13590 | n13703 ;
  assign n37866 = ~n13701 ;
  assign n13705 = n37866 & n13704 ;
  assign n37867 = ~n13705 ;
  assign n13706 = n156 & n37867 ;
  assign n13707 = n37854 & n13704 ;
  assign n13708 = n13609 | n13707 ;
  assign n37868 = ~n13706 ;
  assign n13709 = n37868 & n13708 ;
  assign n37869 = ~n13709 ;
  assign n13710 = n157 & n37869 ;
  assign n13711 = n158 | n13710 ;
  assign n37870 = ~n13711 ;
  assign n13764 = n37870 & n13745 ;
  assign n13765 = n13607 | n13764 ;
  assign n37871 = ~n13747 ;
  assign n13766 = n37871 & n13765 ;
  assign n37872 = ~n13766 ;
  assign n13767 = n159 & n37872 ;
  assign n37873 = ~n13125 ;
  assign n13143 = n37873 & n13142 ;
  assign n13144 = n37567 & n13143 ;
  assign n13612 = n13144 & n151 ;
  assign n13126 = n13110 | n13125 ;
  assign n37874 = ~n13126 ;
  assign n13623 = n37874 & n151 ;
  assign n13624 = n13142 | n13623 ;
  assign n37875 = ~n13612 ;
  assign n13625 = n37875 & n13624 ;
  assign n13748 = n8857 | n13747 ;
  assign n37876 = ~n13748 ;
  assign n13768 = n37876 & n13765 ;
  assign n13769 = n13625 | n13768 ;
  assign n37877 = ~n13767 ;
  assign n13770 = n37877 & n13769 ;
  assign n37878 = ~n13770 ;
  assign n13771 = n8534 & n37878 ;
  assign n13153 = n13147 | n13148 ;
  assign n37879 = ~n13153 ;
  assign n13570 = n37879 & n151 ;
  assign n13571 = n13003 | n13570 ;
  assign n13170 = n13003 & n37556 ;
  assign n37880 = ~n13148 ;
  assign n13171 = n37880 & n13170 ;
  assign n13628 = n13171 & n151 ;
  assign n37881 = ~n13628 ;
  assign n13629 = n13571 & n37881 ;
  assign n13725 = n13708 & n37860 ;
  assign n13726 = n13679 | n13725 ;
  assign n37882 = ~n13710 ;
  assign n13727 = n37882 & n13726 ;
  assign n37883 = ~n13727 ;
  assign n13728 = n158 & n37883 ;
  assign n13729 = n37870 & n13726 ;
  assign n13731 = n13607 | n13729 ;
  assign n37884 = ~n13728 ;
  assign n13732 = n37884 & n13731 ;
  assign n37885 = ~n13732 ;
  assign n13733 = n8857 & n37885 ;
  assign n13734 = n160 | n13733 ;
  assign n37886 = ~n13734 ;
  assign n13788 = n37886 & n13769 ;
  assign n13789 = n13629 | n13788 ;
  assign n37887 = ~n13771 ;
  assign n13790 = n37887 & n13789 ;
  assign n37888 = ~n13790 ;
  assign n13791 = n161 & n37888 ;
  assign n13169 = n13151 | n13158 ;
  assign n37889 = ~n13169 ;
  assign n13578 = n37889 & n151 ;
  assign n13579 = n12940 | n13578 ;
  assign n37890 = ~n13158 ;
  assign n13167 = n12940 & n37890 ;
  assign n13168 = n37583 & n13167 ;
  assign n13632 = n13168 & n151 ;
  assign n37891 = ~n13632 ;
  assign n13633 = n13579 & n37891 ;
  assign n13772 = n161 | n13771 ;
  assign n37892 = ~n13772 ;
  assign n13792 = n37892 & n13789 ;
  assign n13793 = n13633 | n13792 ;
  assign n37893 = ~n13791 ;
  assign n13794 = n37893 & n13793 ;
  assign n37894 = ~n13794 ;
  assign n13795 = n162 & n37894 ;
  assign n13195 = n13162 | n13179 ;
  assign n37895 = ~n13195 ;
  assign n13584 = n37895 & n151 ;
  assign n13585 = n13035 | n13584 ;
  assign n13193 = n13035 & n37572 ;
  assign n37896 = ~n13162 ;
  assign n13194 = n37896 & n13193 ;
  assign n13637 = n13194 & n151 ;
  assign n37897 = ~n13637 ;
  assign n13638 = n13585 & n37897 ;
  assign n13749 = n13731 & n37876 ;
  assign n13750 = n13625 | n13749 ;
  assign n37898 = ~n13733 ;
  assign n13751 = n37898 & n13750 ;
  assign n37899 = ~n13751 ;
  assign n13752 = n160 & n37899 ;
  assign n13753 = n37886 & n13750 ;
  assign n13754 = n13629 | n13753 ;
  assign n37900 = ~n13752 ;
  assign n13755 = n37900 & n13754 ;
  assign n37901 = ~n13755 ;
  assign n13756 = n161 & n37901 ;
  assign n13757 = n162 | n13756 ;
  assign n37902 = ~n13757 ;
  assign n13812 = n37902 & n13793 ;
  assign n13813 = n13638 | n13812 ;
  assign n37903 = ~n13795 ;
  assign n13814 = n37903 & n13813 ;
  assign n37904 = ~n13814 ;
  assign n13815 = n163 & n37904 ;
  assign n37905 = ~n13181 ;
  assign n13190 = n13062 & n37905 ;
  assign n13191 = n37599 & n13190 ;
  assign n13604 = n13191 & n151 ;
  assign n13192 = n13165 | n13181 ;
  assign n37906 = ~n13192 ;
  assign n13639 = n37906 & n151 ;
  assign n13640 = n13062 | n13639 ;
  assign n37907 = ~n13604 ;
  assign n13641 = n37907 & n13640 ;
  assign n13796 = n6889 | n13795 ;
  assign n37908 = ~n13796 ;
  assign n13816 = n37908 & n13813 ;
  assign n13817 = n13641 | n13816 ;
  assign n37909 = ~n13815 ;
  assign n13818 = n37909 & n13817 ;
  assign n37910 = ~n13818 ;
  assign n13819 = n6600 & n37910 ;
  assign n13218 = n12982 & n37588 ;
  assign n37911 = ~n13185 ;
  assign n13219 = n37911 & n13218 ;
  assign n13630 = n13219 & n151 ;
  assign n13220 = n13185 | n13203 ;
  assign n37912 = ~n13220 ;
  assign n13642 = n37912 & n151 ;
  assign n13643 = n12982 | n13642 ;
  assign n37913 = ~n13630 ;
  assign n13644 = n37913 & n13643 ;
  assign n13773 = n13754 & n37892 ;
  assign n13774 = n13633 | n13773 ;
  assign n37914 = ~n13756 ;
  assign n13775 = n37914 & n13774 ;
  assign n37915 = ~n13775 ;
  assign n13776 = n162 & n37915 ;
  assign n13777 = n37902 & n13774 ;
  assign n13778 = n13638 | n13777 ;
  assign n37916 = ~n13776 ;
  assign n13779 = n37916 & n13778 ;
  assign n37917 = ~n13779 ;
  assign n13780 = n6889 & n37917 ;
  assign n13781 = n6600 | n13780 ;
  assign n37918 = ~n13781 ;
  assign n13836 = n37918 & n13817 ;
  assign n13837 = n13644 | n13836 ;
  assign n37919 = ~n13819 ;
  assign n13838 = n37919 & n13837 ;
  assign n37920 = ~n13838 ;
  assign n13839 = n165 & n37920 ;
  assign n13217 = n13188 | n13205 ;
  assign n37921 = ~n13217 ;
  assign n13617 = n37921 & n151 ;
  assign n13618 = n12978 | n13617 ;
  assign n37922 = ~n13205 ;
  assign n13215 = n12978 & n37922 ;
  assign n13216 = n37615 & n13215 ;
  assign n13645 = n13216 & n151 ;
  assign n37923 = ~n13645 ;
  assign n13646 = n13618 & n37923 ;
  assign n13820 = n165 | n13819 ;
  assign n37924 = ~n13820 ;
  assign n13840 = n37924 & n13837 ;
  assign n13841 = n13646 | n13840 ;
  assign n37925 = ~n13839 ;
  assign n13842 = n37925 & n13841 ;
  assign n37926 = ~n13842 ;
  assign n13843 = n166 & n37926 ;
  assign n13214 = n13208 | n13209 ;
  assign n37927 = ~n13214 ;
  assign n13568 = n37927 & n151 ;
  assign n13569 = n13067 | n13568 ;
  assign n13242 = n13067 & n37604 ;
  assign n37928 = ~n13209 ;
  assign n13243 = n37928 & n13242 ;
  assign n13593 = n13243 & n151 ;
  assign n37929 = ~n13593 ;
  assign n13594 = n13569 & n37929 ;
  assign n13797 = n13778 & n37908 ;
  assign n13798 = n13641 | n13797 ;
  assign n37930 = ~n13780 ;
  assign n13799 = n37930 & n13798 ;
  assign n37931 = ~n13799 ;
  assign n13800 = n164 & n37931 ;
  assign n13801 = n37918 & n13798 ;
  assign n13802 = n13644 | n13801 ;
  assign n37932 = ~n13800 ;
  assign n13803 = n37932 & n13802 ;
  assign n37933 = ~n13803 ;
  assign n13804 = n165 & n37933 ;
  assign n13805 = n166 | n13804 ;
  assign n37934 = ~n13805 ;
  assign n13860 = n37934 & n13841 ;
  assign n13861 = n13594 | n13860 ;
  assign n37935 = ~n13843 ;
  assign n13862 = n37935 & n13861 ;
  assign n37936 = ~n13862 ;
  assign n13863 = n167 & n37936 ;
  assign n13241 = n13212 | n13230 ;
  assign n37937 = ~n13241 ;
  assign n13564 = n37937 & n151 ;
  assign n13565 = n13023 | n13564 ;
  assign n37938 = ~n13230 ;
  assign n13239 = n13023 & n37938 ;
  assign n13240 = n37631 & n13239 ;
  assign n13566 = n13240 & n151 ;
  assign n37939 = ~n13566 ;
  assign n13567 = n13565 & n37939 ;
  assign n13844 = n5352 | n13843 ;
  assign n37940 = ~n13844 ;
  assign n13864 = n37940 & n13861 ;
  assign n13865 = n13567 | n13864 ;
  assign n37941 = ~n13863 ;
  assign n13866 = n37941 & n13865 ;
  assign n37942 = ~n13866 ;
  assign n13867 = n4934 & n37942 ;
  assign n13257 = n13234 | n13251 ;
  assign n37943 = ~n13257 ;
  assign n13591 = n37943 & n151 ;
  assign n13592 = n13041 | n13591 ;
  assign n13255 = n13041 & n37620 ;
  assign n37944 = ~n13234 ;
  assign n13256 = n37944 & n13255 ;
  assign n13595 = n13256 & n151 ;
  assign n37945 = ~n13595 ;
  assign n13596 = n13592 & n37945 ;
  assign n13821 = n13802 & n37924 ;
  assign n13822 = n13646 | n13821 ;
  assign n37946 = ~n13804 ;
  assign n13823 = n37946 & n13822 ;
  assign n37947 = ~n13823 ;
  assign n13824 = n166 & n37947 ;
  assign n13825 = n37934 & n13822 ;
  assign n13826 = n13594 | n13825 ;
  assign n37948 = ~n13824 ;
  assign n13827 = n37948 & n13826 ;
  assign n37949 = ~n13827 ;
  assign n13828 = n5352 & n37949 ;
  assign n13829 = n4934 | n13828 ;
  assign n37950 = ~n13829 ;
  assign n13884 = n37950 & n13865 ;
  assign n13885 = n13596 | n13884 ;
  assign n37951 = ~n13867 ;
  assign n13886 = n37951 & n13885 ;
  assign n37952 = ~n13886 ;
  assign n13887 = n169 & n37952 ;
  assign n13254 = n13237 | n13253 ;
  assign n37953 = ~n13254 ;
  assign n13561 = n37953 & n151 ;
  assign n13562 = n13264 | n13561 ;
  assign n37954 = ~n13253 ;
  assign n13265 = n37954 & n13264 ;
  assign n13266 = n37647 & n13265 ;
  assign n13680 = n13266 & n13662 ;
  assign n37955 = ~n13680 ;
  assign n13681 = n13562 & n37955 ;
  assign n13868 = n169 | n13867 ;
  assign n37956 = ~n13868 ;
  assign n13888 = n37956 & n13885 ;
  assign n13889 = n13681 | n13888 ;
  assign n37957 = ~n13887 ;
  assign n13890 = n37957 & n13889 ;
  assign n37958 = ~n13890 ;
  assign n13891 = n170 & n37958 ;
  assign n13275 = n13269 | n13270 ;
  assign n37959 = ~n13275 ;
  assign n13559 = n37959 & n151 ;
  assign n13560 = n13073 | n13559 ;
  assign n13293 = n13073 & n37636 ;
  assign n37960 = ~n13270 ;
  assign n13294 = n37960 & n13293 ;
  assign n13682 = n13294 & n13662 ;
  assign n37961 = ~n13682 ;
  assign n13683 = n13560 & n37961 ;
  assign n13845 = n13826 & n37940 ;
  assign n13846 = n13567 | n13845 ;
  assign n37962 = ~n13828 ;
  assign n13847 = n37962 & n13846 ;
  assign n37963 = ~n13847 ;
  assign n13848 = n168 & n37963 ;
  assign n13849 = n37950 & n13846 ;
  assign n13850 = n13596 | n13849 ;
  assign n37964 = ~n13848 ;
  assign n13851 = n37964 & n13850 ;
  assign n37965 = ~n13851 ;
  assign n13852 = n169 & n37965 ;
  assign n13853 = n170 | n13852 ;
  assign n37966 = ~n13853 ;
  assign n13908 = n37966 & n13889 ;
  assign n13909 = n13683 | n13908 ;
  assign n37967 = ~n13891 ;
  assign n13910 = n37967 & n13909 ;
  assign n37968 = ~n13910 ;
  assign n13911 = n171 & n37968 ;
  assign n37969 = ~n13280 ;
  assign n13290 = n13043 & n37969 ;
  assign n13291 = n37663 & n13290 ;
  assign n13558 = n13291 & n151 ;
  assign n13292 = n13273 | n13280 ;
  assign n37970 = ~n13292 ;
  assign n13580 = n37970 & n151 ;
  assign n13581 = n13043 | n13580 ;
  assign n37971 = ~n13558 ;
  assign n13582 = n37971 & n13581 ;
  assign n13892 = n3940 | n13891 ;
  assign n37972 = ~n13892 ;
  assign n13912 = n37972 & n13909 ;
  assign n13913 = n13582 | n13912 ;
  assign n37973 = ~n13911 ;
  assign n13914 = n37973 & n13913 ;
  assign n37974 = ~n13914 ;
  assign n13915 = n3631 & n37974 ;
  assign n13317 = n13025 & n37652 ;
  assign n37975 = ~n13284 ;
  assign n13318 = n37975 & n13317 ;
  assign n13550 = n13318 & n151 ;
  assign n13289 = n13283 | n13284 ;
  assign n37976 = ~n13289 ;
  assign n13553 = n37976 & n151 ;
  assign n13554 = n13025 | n13553 ;
  assign n37977 = ~n13550 ;
  assign n13555 = n37977 & n13554 ;
  assign n13869 = n13850 & n37956 ;
  assign n13870 = n13681 | n13869 ;
  assign n37978 = ~n13852 ;
  assign n13871 = n37978 & n13870 ;
  assign n37979 = ~n13871 ;
  assign n13872 = n170 & n37979 ;
  assign n13873 = n37966 & n13870 ;
  assign n13874 = n13683 | n13873 ;
  assign n37980 = ~n13872 ;
  assign n13875 = n37980 & n13874 ;
  assign n37981 = ~n13875 ;
  assign n13876 = n3940 & n37981 ;
  assign n13877 = n3631 | n13876 ;
  assign n37982 = ~n13877 ;
  assign n13932 = n37982 & n13913 ;
  assign n13933 = n13555 | n13932 ;
  assign n37983 = ~n13915 ;
  assign n13934 = n37983 & n13933 ;
  assign n37984 = ~n13934 ;
  assign n13935 = n173 & n37984 ;
  assign n37985 = ~n13304 ;
  assign n13314 = n13054 & n37985 ;
  assign n13315 = n37679 & n13314 ;
  assign n13563 = n13315 & n151 ;
  assign n13316 = n13287 | n13304 ;
  assign n37986 = ~n13316 ;
  assign n13575 = n37986 & n151 ;
  assign n13576 = n13054 | n13575 ;
  assign n37987 = ~n13563 ;
  assign n13577 = n37987 & n13576 ;
  assign n13916 = n173 | n13915 ;
  assign n37988 = ~n13916 ;
  assign n13936 = n37988 & n13933 ;
  assign n13937 = n13577 | n13936 ;
  assign n37989 = ~n13935 ;
  assign n13938 = n37989 & n13937 ;
  assign n37990 = ~n13938 ;
  assign n13939 = n174 & n37990 ;
  assign n13313 = n13307 | n13308 ;
  assign n37991 = ~n13313 ;
  assign n13619 = n37991 & n151 ;
  assign n13620 = n13059 | n13619 ;
  assign n13341 = n13059 & n37668 ;
  assign n37992 = ~n13308 ;
  assign n13342 = n37992 & n13341 ;
  assign n13626 = n13342 & n151 ;
  assign n37993 = ~n13626 ;
  assign n13627 = n13620 & n37993 ;
  assign n13893 = n13874 & n37972 ;
  assign n13894 = n13582 | n13893 ;
  assign n37994 = ~n13876 ;
  assign n13895 = n37994 & n13894 ;
  assign n37995 = ~n13895 ;
  assign n13896 = n172 & n37995 ;
  assign n13897 = n37982 & n13894 ;
  assign n13898 = n13555 | n13897 ;
  assign n37996 = ~n13896 ;
  assign n13899 = n37996 & n13898 ;
  assign n37997 = ~n13899 ;
  assign n13900 = n173 & n37997 ;
  assign n13901 = n174 | n13900 ;
  assign n37998 = ~n13901 ;
  assign n13956 = n37998 & n13937 ;
  assign n13957 = n13627 | n13956 ;
  assign n37999 = ~n13939 ;
  assign n13958 = n37999 & n13957 ;
  assign n38000 = ~n13958 ;
  assign n13959 = n175 & n38000 ;
  assign n13340 = n13311 | n13328 ;
  assign n38001 = ~n13340 ;
  assign n13548 = n38001 & n151 ;
  assign n13549 = n12974 | n13548 ;
  assign n38002 = ~n13328 ;
  assign n13338 = n12974 & n38002 ;
  assign n13339 = n37695 & n13338 ;
  assign n13551 = n13339 & n151 ;
  assign n38003 = ~n13551 ;
  assign n13552 = n13549 & n38003 ;
  assign n13940 = n2753 | n13939 ;
  assign n38004 = ~n13940 ;
  assign n13960 = n38004 & n13957 ;
  assign n13961 = n13552 | n13960 ;
  assign n38005 = ~n13959 ;
  assign n13962 = n38005 & n13961 ;
  assign n38006 = ~n13962 ;
  assign n13963 = n2431 & n38006 ;
  assign n13354 = n13064 & n37684 ;
  assign n38007 = ~n13332 ;
  assign n13355 = n38007 & n13354 ;
  assign n13543 = n13355 & n151 ;
  assign n13337 = n13331 | n13332 ;
  assign n38008 = ~n13337 ;
  assign n13544 = n38008 & n151 ;
  assign n13545 = n13064 | n13544 ;
  assign n38009 = ~n13543 ;
  assign n13546 = n38009 & n13545 ;
  assign n13917 = n13898 & n37988 ;
  assign n13918 = n13577 | n13917 ;
  assign n38010 = ~n13900 ;
  assign n13919 = n38010 & n13918 ;
  assign n38011 = ~n13919 ;
  assign n13920 = n174 & n38011 ;
  assign n13921 = n37998 & n13918 ;
  assign n13922 = n13627 | n13921 ;
  assign n38012 = ~n13920 ;
  assign n13923 = n38012 & n13922 ;
  assign n38013 = ~n13923 ;
  assign n13924 = n2753 & n38013 ;
  assign n13925 = n2431 | n13924 ;
  assign n38014 = ~n13925 ;
  assign n13969 = n38014 & n13961 ;
  assign n13970 = n13546 | n13969 ;
  assign n38015 = ~n13963 ;
  assign n13971 = n38015 & n13970 ;
  assign n38016 = ~n13971 ;
  assign n13972 = n177 & n38016 ;
  assign n13964 = n177 | n13963 ;
  assign n38017 = ~n13964 ;
  assign n13973 = n38017 & n13970 ;
  assign n38018 = ~n13352 ;
  assign n13397 = n38018 & n13381 ;
  assign n13398 = n37711 & n13397 ;
  assign n13583 = n13398 & n151 ;
  assign n13353 = n13335 | n13352 ;
  assign n38019 = ~n13353 ;
  assign n13542 = n38019 & n151 ;
  assign n14064 = n13381 | n13542 ;
  assign n38020 = ~n13583 ;
  assign n14065 = n38020 & n14064 ;
  assign n14066 = n13973 | n14065 ;
  assign n38021 = ~n13972 ;
  assign n14067 = n38021 & n14066 ;
  assign n38022 = ~n14067 ;
  assign n14068 = n178 & n38022 ;
  assign n13386 = n13050 & n37700 ;
  assign n38023 = ~n13402 ;
  assign n14058 = n13386 & n38023 ;
  assign n14059 = n151 & n14058 ;
  assign n14060 = n13401 | n13402 ;
  assign n38024 = ~n14060 ;
  assign n14061 = n151 & n38024 ;
  assign n14062 = n13050 | n14061 ;
  assign n38025 = ~n14059 ;
  assign n14063 = n38025 & n14062 ;
  assign n13941 = n13922 & n38004 ;
  assign n13942 = n13552 | n13941 ;
  assign n38026 = ~n13924 ;
  assign n13943 = n38026 & n13942 ;
  assign n38027 = ~n13943 ;
  assign n13944 = n176 & n38027 ;
  assign n13945 = n38014 & n13942 ;
  assign n13946 = n13546 | n13945 ;
  assign n38028 = ~n13944 ;
  assign n13947 = n38028 & n13946 ;
  assign n38029 = ~n13947 ;
  assign n13948 = n177 & n38029 ;
  assign n13949 = n178 | n13948 ;
  assign n38030 = ~n13949 ;
  assign n14071 = n38030 & n14066 ;
  assign n14072 = n14063 | n14071 ;
  assign n38031 = ~n14068 ;
  assign n14073 = n38031 & n14072 ;
  assign n38032 = ~n14073 ;
  assign n14074 = n179 & n38032 ;
  assign n38033 = ~n13417 ;
  assign n14051 = n13070 & n38033 ;
  assign n14052 = n37727 & n14051 ;
  assign n14053 = n151 & n14052 ;
  assign n14054 = n13405 | n13417 ;
  assign n38034 = ~n14054 ;
  assign n14055 = n151 & n38034 ;
  assign n14056 = n13070 | n14055 ;
  assign n38035 = ~n14053 ;
  assign n14057 = n38035 & n14056 ;
  assign n14069 = n1707 | n14068 ;
  assign n38036 = ~n14069 ;
  assign n14075 = n38036 & n14072 ;
  assign n14076 = n14057 | n14075 ;
  assign n38037 = ~n14074 ;
  assign n14077 = n38037 & n14076 ;
  assign n38038 = ~n14077 ;
  assign n14078 = n1487 & n38038 ;
  assign n13396 = n13032 & n37716 ;
  assign n38039 = ~n13421 ;
  assign n14045 = n13396 & n38039 ;
  assign n14046 = n151 & n14045 ;
  assign n14047 = n13394 | n13421 ;
  assign n38040 = ~n14047 ;
  assign n14048 = n151 & n38040 ;
  assign n14049 = n13032 | n14048 ;
  assign n38041 = ~n14046 ;
  assign n14050 = n38041 & n14049 ;
  assign n13965 = n13946 & n38017 ;
  assign n14083 = n13965 | n14065 ;
  assign n38042 = ~n13948 ;
  assign n14084 = n38042 & n14083 ;
  assign n38043 = ~n14084 ;
  assign n14085 = n178 & n38043 ;
  assign n14086 = n38030 & n14083 ;
  assign n14087 = n14063 | n14086 ;
  assign n38044 = ~n14085 ;
  assign n14088 = n38044 & n14087 ;
  assign n38045 = ~n14088 ;
  assign n14089 = n1707 & n38045 ;
  assign n14090 = n1487 | n14089 ;
  assign n38046 = ~n14090 ;
  assign n14091 = n14076 & n38046 ;
  assign n14092 = n14050 | n14091 ;
  assign n38047 = ~n14078 ;
  assign n14093 = n38047 & n14092 ;
  assign n38048 = ~n14093 ;
  assign n14094 = n181 & n38048 ;
  assign n38049 = ~n13436 ;
  assign n14038 = n13038 & n38049 ;
  assign n14039 = n37743 & n14038 ;
  assign n14040 = n151 & n14039 ;
  assign n14041 = n13424 | n13436 ;
  assign n38050 = ~n14041 ;
  assign n14042 = n151 & n38050 ;
  assign n14043 = n13038 | n14042 ;
  assign n38051 = ~n14040 ;
  assign n14044 = n38051 & n14043 ;
  assign n14079 = n181 | n14078 ;
  assign n38052 = ~n14079 ;
  assign n14095 = n38052 & n14092 ;
  assign n14096 = n14044 | n14095 ;
  assign n38053 = ~n14094 ;
  assign n14097 = n38053 & n14096 ;
  assign n38054 = ~n14097 ;
  assign n14098 = n182 & n38054 ;
  assign n13416 = n12995 & n37732 ;
  assign n38055 = ~n13440 ;
  assign n14032 = n13416 & n38055 ;
  assign n14033 = n13662 & n14032 ;
  assign n14034 = n13439 | n13440 ;
  assign n38056 = ~n14034 ;
  assign n14035 = n151 & n38056 ;
  assign n14036 = n12995 | n14035 ;
  assign n38057 = ~n14033 ;
  assign n14037 = n38057 & n14036 ;
  assign n14101 = n38036 & n14087 ;
  assign n14102 = n14057 | n14101 ;
  assign n38058 = ~n14089 ;
  assign n14103 = n38058 & n14102 ;
  assign n38059 = ~n14103 ;
  assign n14104 = n180 & n38059 ;
  assign n14105 = n38046 & n14102 ;
  assign n14106 = n14050 | n14105 ;
  assign n38060 = ~n14104 ;
  assign n14107 = n38060 & n14106 ;
  assign n38061 = ~n14107 ;
  assign n14108 = n181 & n38061 ;
  assign n14109 = n182 | n14108 ;
  assign n38062 = ~n14109 ;
  assign n14110 = n14096 & n38062 ;
  assign n14111 = n14037 | n14110 ;
  assign n38063 = ~n14098 ;
  assign n14112 = n38063 & n14111 ;
  assign n38064 = ~n14112 ;
  assign n14113 = n183 & n38064 ;
  assign n38065 = ~n13455 ;
  assign n14025 = n13076 & n38065 ;
  assign n14026 = n37759 & n14025 ;
  assign n14027 = n151 & n14026 ;
  assign n14028 = n13443 | n13455 ;
  assign n38066 = ~n14028 ;
  assign n14029 = n151 & n38066 ;
  assign n14030 = n13076 | n14029 ;
  assign n38067 = ~n14027 ;
  assign n14031 = n38067 & n14030 ;
  assign n14099 = n183 | n14098 ;
  assign n38068 = ~n14099 ;
  assign n14114 = n38068 & n14111 ;
  assign n14115 = n14031 | n14114 ;
  assign n38069 = ~n14113 ;
  assign n14116 = n38069 & n14115 ;
  assign n38070 = ~n14116 ;
  assign n14117 = n838 & n38070 ;
  assign n13461 = n13458 | n13459 ;
  assign n38071 = ~n13461 ;
  assign n13621 = n38071 & n151 ;
  assign n13622 = n12965 | n13621 ;
  assign n13435 = n12965 & n37748 ;
  assign n38072 = ~n13459 ;
  assign n13460 = n13435 & n38072 ;
  assign n13647 = n13460 & n151 ;
  assign n38073 = ~n13647 ;
  assign n13648 = n13622 & n38073 ;
  assign n14120 = n38052 & n14106 ;
  assign n14121 = n14044 | n14120 ;
  assign n38074 = ~n14108 ;
  assign n14122 = n38074 & n14121 ;
  assign n38075 = ~n14122 ;
  assign n14123 = n182 & n38075 ;
  assign n14124 = n38062 & n14121 ;
  assign n14125 = n14037 | n14124 ;
  assign n38076 = ~n14123 ;
  assign n14126 = n38076 & n14125 ;
  assign n38077 = ~n14126 ;
  assign n14127 = n996 & n38077 ;
  assign n14128 = n838 | n14127 ;
  assign n38078 = ~n14128 ;
  assign n14129 = n14115 & n38078 ;
  assign n14130 = n13648 | n14129 ;
  assign n38079 = ~n14117 ;
  assign n14131 = n38079 & n14130 ;
  assign n38080 = ~n14131 ;
  assign n14132 = n185 & n38080 ;
  assign n38081 = ~n13476 ;
  assign n14018 = n12961 & n38081 ;
  assign n14019 = n37775 & n14018 ;
  assign n14020 = n151 & n14019 ;
  assign n14021 = n13464 | n13476 ;
  assign n38082 = ~n14021 ;
  assign n14022 = n151 & n38082 ;
  assign n14023 = n12961 | n14022 ;
  assign n38083 = ~n14020 ;
  assign n14024 = n38083 & n14023 ;
  assign n14118 = n185 | n14117 ;
  assign n38084 = ~n14118 ;
  assign n14133 = n38084 & n14130 ;
  assign n14134 = n14024 | n14133 ;
  assign n38085 = ~n14132 ;
  assign n14135 = n38085 & n14134 ;
  assign n38086 = ~n14135 ;
  assign n14136 = n186 & n38086 ;
  assign n13454 = n13140 & n37764 ;
  assign n38087 = ~n13480 ;
  assign n14012 = n13454 & n38087 ;
  assign n14013 = n151 & n14012 ;
  assign n14014 = n13479 | n13480 ;
  assign n38088 = ~n14014 ;
  assign n14015 = n151 & n38088 ;
  assign n14016 = n13140 | n14015 ;
  assign n38089 = ~n14013 ;
  assign n14017 = n38089 & n14016 ;
  assign n14139 = n38068 & n14125 ;
  assign n14140 = n14031 | n14139 ;
  assign n38090 = ~n14127 ;
  assign n14141 = n38090 & n14140 ;
  assign n38091 = ~n14141 ;
  assign n14142 = n184 & n38091 ;
  assign n14143 = n38078 & n14140 ;
  assign n14144 = n13648 | n14143 ;
  assign n38092 = ~n14142 ;
  assign n14145 = n38092 & n14144 ;
  assign n38093 = ~n14145 ;
  assign n14146 = n185 & n38093 ;
  assign n14147 = n186 | n14146 ;
  assign n38094 = ~n14147 ;
  assign n14148 = n14134 & n38094 ;
  assign n14149 = n14017 | n14148 ;
  assign n38095 = ~n14136 ;
  assign n14150 = n38095 & n14149 ;
  assign n38096 = ~n14150 ;
  assign n14151 = n187 & n38096 ;
  assign n38097 = ~n13495 ;
  assign n14005 = n13081 & n38097 ;
  assign n14006 = n37791 & n14005 ;
  assign n14007 = n13662 & n14006 ;
  assign n14008 = n13483 | n13495 ;
  assign n38098 = ~n14008 ;
  assign n14009 = n151 & n38098 ;
  assign n14010 = n13081 | n14009 ;
  assign n38099 = ~n14007 ;
  assign n14011 = n38099 & n14010 ;
  assign n14137 = n528 | n14136 ;
  assign n38100 = ~n14137 ;
  assign n14152 = n38100 & n14149 ;
  assign n14153 = n14011 | n14152 ;
  assign n38101 = ~n14151 ;
  assign n14154 = n38101 & n14153 ;
  assign n38102 = ~n14154 ;
  assign n14155 = n413 & n38102 ;
  assign n13475 = n12959 & n37780 ;
  assign n38103 = ~n13499 ;
  assign n13999 = n13475 & n38103 ;
  assign n14000 = n151 & n13999 ;
  assign n14001 = n13498 | n13499 ;
  assign n38104 = ~n14001 ;
  assign n14002 = n151 & n38104 ;
  assign n14003 = n12959 | n14002 ;
  assign n38105 = ~n14000 ;
  assign n14004 = n38105 & n14003 ;
  assign n14158 = n38084 & n14144 ;
  assign n14159 = n14024 | n14158 ;
  assign n38106 = ~n14146 ;
  assign n14160 = n38106 & n14159 ;
  assign n38107 = ~n14160 ;
  assign n14161 = n186 & n38107 ;
  assign n14162 = n38094 & n14159 ;
  assign n14165 = n14017 | n14162 ;
  assign n38108 = ~n14161 ;
  assign n14166 = n38108 & n14165 ;
  assign n38109 = ~n14166 ;
  assign n14167 = n528 & n38109 ;
  assign n14168 = n413 | n14167 ;
  assign n38110 = ~n14168 ;
  assign n14169 = n14153 & n38110 ;
  assign n14170 = n14004 | n14169 ;
  assign n38111 = ~n14155 ;
  assign n14171 = n38111 & n14170 ;
  assign n38112 = ~n14171 ;
  assign n14172 = n189 & n38112 ;
  assign n38113 = ~n13504 ;
  assign n13992 = n12951 & n38113 ;
  assign n13993 = n37797 & n13992 ;
  assign n13994 = n151 & n13993 ;
  assign n13995 = n13502 | n13504 ;
  assign n38114 = ~n13995 ;
  assign n13996 = n151 & n38114 ;
  assign n13997 = n12951 | n13996 ;
  assign n38115 = ~n13994 ;
  assign n13998 = n38115 & n13997 ;
  assign n14156 = n189 | n14155 ;
  assign n38116 = ~n14156 ;
  assign n14173 = n38116 & n14170 ;
  assign n14174 = n13998 | n14173 ;
  assign n38117 = ~n14172 ;
  assign n14175 = n38117 & n14174 ;
  assign n38118 = ~n14175 ;
  assign n14176 = n190 & n38118 ;
  assign n14177 = n287 | n14176 ;
  assign n38119 = ~n13492 ;
  assign n13494 = n12946 & n38119 ;
  assign n38120 = ~n13508 ;
  assign n13986 = n13494 & n38120 ;
  assign n13987 = n13662 & n13986 ;
  assign n13988 = n13507 | n13508 ;
  assign n38121 = ~n13988 ;
  assign n13989 = n151 & n38121 ;
  assign n13990 = n12946 | n13989 ;
  assign n38122 = ~n13987 ;
  assign n13991 = n38122 & n13990 ;
  assign n14179 = n38100 & n14165 ;
  assign n14180 = n14011 | n14179 ;
  assign n38123 = ~n14167 ;
  assign n14181 = n38123 & n14180 ;
  assign n38124 = ~n14181 ;
  assign n14182 = n188 & n38124 ;
  assign n14183 = n38110 & n14180 ;
  assign n14184 = n14004 | n14183 ;
  assign n38125 = ~n14182 ;
  assign n14185 = n38125 & n14184 ;
  assign n38126 = ~n14185 ;
  assign n14186 = n189 & n38126 ;
  assign n14187 = n190 | n14186 ;
  assign n14188 = n38116 & n14184 ;
  assign n14189 = n13998 | n14188 ;
  assign n38127 = ~n14187 ;
  assign n14192 = n38127 & n14189 ;
  assign n14193 = n13991 | n14192 ;
  assign n38128 = ~n14177 ;
  assign n14194 = n38128 & n14193 ;
  assign n14196 = n13652 | n14194 ;
  assign n38129 = ~n14186 ;
  assign n14190 = n38129 & n14189 ;
  assign n38130 = ~n14190 ;
  assign n14191 = n190 & n38130 ;
  assign n38131 = ~n14191 ;
  assign n14197 = n38131 & n14193 ;
  assign n38132 = ~n14197 ;
  assign n14198 = n287 & n38132 ;
  assign n38133 = ~n14198 ;
  assign n14199 = n14196 & n38133 ;
  assign n14200 = n13659 | n14199 ;
  assign n14201 = n31336 & n14200 ;
  assign n13532 = n192 & n13531 ;
  assign n38134 = ~n13368 ;
  assign n13613 = n38134 & n151 ;
  assign n38135 = ~n13613 ;
  assign n13614 = n13530 & n38135 ;
  assign n38136 = ~n13614 ;
  assign n13615 = n13532 & n38136 ;
  assign n13364 = n12909 | n13363 ;
  assign n38137 = ~n13364 ;
  assign n13370 = n38137 & n13367 ;
  assign n13371 = n37828 & n13370 ;
  assign n13527 = n13371 & n37829 ;
  assign n13976 = n13527 & n37830 ;
  assign n13977 = n13615 | n13976 ;
  assign n14204 = n13658 & n38133 ;
  assign n14205 = n14196 & n14204 ;
  assign n14206 = n13977 | n14205 ;
  assign n150 = n14201 | n14206 ;
  assign n14202 = n13658 | n14199 ;
  assign n38138 = ~n14202 ;
  assign n14307 = n38138 & n150 ;
  assign n14660 = n14205 | n14307 ;
  assign n38139 = ~n14194 ;
  assign n14195 = n13652 & n38139 ;
  assign n14670 = n14195 & n38133 ;
  assign n14671 = n150 & n14670 ;
  assign n14673 = n14194 | n14198 ;
  assign n38140 = ~n14673 ;
  assign n14674 = n150 & n38140 ;
  assign n14675 = n13652 | n14674 ;
  assign n38141 = ~n14671 ;
  assign n14676 = n38141 & n14675 ;
  assign n14677 = n14660 | n14676 ;
  assign n209 = x40 | x41 ;
  assign n210 = x42 | n209 ;
  assign n14263 = x42 & n150 ;
  assign n38142 = ~n14263 ;
  assign n14264 = n210 & n38142 ;
  assign n38143 = ~n14264 ;
  assign n14265 = n151 & n38143 ;
  assign n12910 = n210 & n37827 ;
  assign n12927 = n12910 & n37828 ;
  assign n13528 = n12927 & n37829 ;
  assign n13985 = n13528 & n37830 ;
  assign n14308 = n13985 & n38142 ;
  assign n38144 = ~n206 ;
  assign n14259 = n38144 & n150 ;
  assign n38145 = ~x42 ;
  assign n14329 = n38145 & n150 ;
  assign n38146 = ~n14329 ;
  assign n14330 = x43 & n38146 ;
  assign n14331 = n14259 | n14330 ;
  assign n14332 = n14308 | n14331 ;
  assign n38147 = ~n14265 ;
  assign n14335 = n38147 & n14332 ;
  assign n38148 = ~n14335 ;
  assign n14336 = n13079 & n38148 ;
  assign n211 = n38145 & n209 ;
  assign n38149 = ~n150 ;
  assign n14309 = x42 & n38149 ;
  assign n14310 = n211 | n14309 ;
  assign n38150 = ~n14310 ;
  assign n14311 = n13662 & n38150 ;
  assign n14312 = n13079 | n14311 ;
  assign n38151 = ~n14312 ;
  assign n14333 = n38151 & n14332 ;
  assign n38152 = ~n13976 ;
  assign n13978 = n13662 & n38152 ;
  assign n38153 = ~n13615 ;
  assign n13979 = n38153 & n13978 ;
  assign n38154 = ~n14205 ;
  assign n14341 = n13979 & n38154 ;
  assign n38155 = ~n14201 ;
  assign n14342 = n38155 & n14341 ;
  assign n14343 = n14259 | n14342 ;
  assign n14344 = x44 & n14343 ;
  assign n14345 = x44 | n14342 ;
  assign n14346 = n14259 | n14345 ;
  assign n38156 = ~n14344 ;
  assign n14347 = n38156 & n14346 ;
  assign n14348 = n14333 | n14347 ;
  assign n38157 = ~n14336 ;
  assign n14349 = n38157 & n14348 ;
  assign n38158 = ~n14349 ;
  assign n14350 = n153 & n38158 ;
  assign n13676 = n13634 | n13671 ;
  assign n38159 = ~n13676 ;
  assign n13677 = n13631 & n38159 ;
  assign n14316 = n13677 & n150 ;
  assign n14317 = n38159 & n150 ;
  assign n14318 = n13631 | n14317 ;
  assign n38160 = ~n14316 ;
  assign n14319 = n38160 & n14318 ;
  assign n14337 = n153 | n14336 ;
  assign n38161 = ~n14337 ;
  assign n14353 = n38161 & n14348 ;
  assign n14354 = n14319 | n14353 ;
  assign n38162 = ~n14350 ;
  assign n14355 = n38162 & n14354 ;
  assign n38163 = ~n14355 ;
  assign n14356 = n154 & n38163 ;
  assign n13675 = n13670 | n13673 ;
  assign n38164 = ~n13675 ;
  assign n14314 = n38164 & n150 ;
  assign n14315 = n13689 | n14314 ;
  assign n38165 = ~n13670 ;
  assign n13695 = n38165 & n13689 ;
  assign n38166 = ~n13673 ;
  assign n13696 = n38166 & n13695 ;
  assign n14320 = n13696 & n150 ;
  assign n38167 = ~n14320 ;
  assign n14321 = n14315 & n38167 ;
  assign n14351 = n154 | n14350 ;
  assign n38168 = ~n14351 ;
  assign n14357 = n38168 & n14354 ;
  assign n14358 = n14321 | n14357 ;
  assign n38169 = ~n14356 ;
  assign n14359 = n38169 & n14358 ;
  assign n38170 = ~n14359 ;
  assign n14360 = n11067 & n38170 ;
  assign n13975 = n13692 | n13698 ;
  assign n38171 = ~n13975 ;
  assign n14322 = n38171 & n150 ;
  assign n14323 = n13599 | n14322 ;
  assign n13693 = n13599 & n37838 ;
  assign n38172 = ~n13698 ;
  assign n13974 = n13693 & n38172 ;
  assign n14324 = n13974 & n150 ;
  assign n38173 = ~n14324 ;
  assign n14325 = n14323 & n38173 ;
  assign n14338 = n152 & n38148 ;
  assign n14266 = n152 | n14265 ;
  assign n38174 = ~n14266 ;
  assign n14340 = n38174 & n14332 ;
  assign n14369 = n14340 | n14347 ;
  assign n38175 = ~n14338 ;
  assign n14370 = n38175 & n14369 ;
  assign n38176 = ~n14370 ;
  assign n14371 = n153 & n38176 ;
  assign n14372 = n38161 & n14369 ;
  assign n14373 = n14319 | n14372 ;
  assign n38177 = ~n14371 ;
  assign n14374 = n38177 & n14373 ;
  assign n38178 = ~n14374 ;
  assign n14375 = n154 & n38178 ;
  assign n14376 = n11067 | n14375 ;
  assign n38179 = ~n14376 ;
  assign n14377 = n14358 & n38179 ;
  assign n14378 = n14325 | n14377 ;
  assign n38180 = ~n14360 ;
  assign n14379 = n38180 & n14378 ;
  assign n38181 = ~n14379 ;
  assign n14380 = n156 & n38181 ;
  assign n13715 = n13701 | n13703 ;
  assign n38182 = ~n13715 ;
  assign n14237 = n38182 & n150 ;
  assign n14238 = n13590 | n14237 ;
  assign n38183 = ~n13703 ;
  assign n13713 = n13590 & n38183 ;
  assign n13714 = n37866 & n13713 ;
  assign n14254 = n13714 & n150 ;
  assign n38184 = ~n14254 ;
  assign n14255 = n14238 & n38184 ;
  assign n14361 = n10657 | n14360 ;
  assign n38185 = ~n14361 ;
  assign n14381 = n38185 & n14378 ;
  assign n14382 = n14255 | n14381 ;
  assign n38186 = ~n14380 ;
  assign n14383 = n38186 & n14382 ;
  assign n38187 = ~n14383 ;
  assign n14384 = n157 & n38187 ;
  assign n13738 = n13609 & n37855 ;
  assign n38188 = ~n13707 ;
  assign n13739 = n38188 & n13738 ;
  assign n14236 = n13739 & n150 ;
  assign n13712 = n13706 | n13707 ;
  assign n38189 = ~n13712 ;
  assign n14270 = n38189 & n150 ;
  assign n14271 = n13609 | n14270 ;
  assign n38190 = ~n14236 ;
  assign n14272 = n38190 & n14271 ;
  assign n14392 = n38168 & n14373 ;
  assign n14393 = n14321 | n14392 ;
  assign n38191 = ~n14375 ;
  assign n14394 = n38191 & n14393 ;
  assign n38192 = ~n14394 ;
  assign n14395 = n155 & n38192 ;
  assign n14396 = n38179 & n14393 ;
  assign n14397 = n14325 | n14396 ;
  assign n38193 = ~n14395 ;
  assign n14398 = n38193 & n14397 ;
  assign n38194 = ~n14398 ;
  assign n14399 = n10657 & n38194 ;
  assign n14400 = n157 | n14399 ;
  assign n38195 = ~n14400 ;
  assign n14401 = n14382 & n38195 ;
  assign n14402 = n14272 | n14401 ;
  assign n38196 = ~n14384 ;
  assign n14403 = n38196 & n14402 ;
  assign n38197 = ~n14403 ;
  assign n14404 = n158 & n38197 ;
  assign n38198 = ~n13725 ;
  assign n13735 = n13679 & n38198 ;
  assign n13736 = n37882 & n13735 ;
  assign n14239 = n13736 & n150 ;
  assign n13737 = n13710 | n13725 ;
  assign n38199 = ~n13737 ;
  assign n14240 = n38199 & n150 ;
  assign n14241 = n13679 | n14240 ;
  assign n38200 = ~n14239 ;
  assign n14242 = n38200 & n14241 ;
  assign n14385 = n158 | n14384 ;
  assign n38201 = ~n14385 ;
  assign n14405 = n38201 & n14402 ;
  assign n14406 = n14242 | n14405 ;
  assign n38202 = ~n14404 ;
  assign n14407 = n38202 & n14406 ;
  assign n38203 = ~n14407 ;
  assign n14408 = n8857 & n38203 ;
  assign n13762 = n13607 & n37871 ;
  assign n38204 = ~n13729 ;
  assign n13763 = n38204 & n13762 ;
  assign n14227 = n13763 & n150 ;
  assign n13730 = n13728 | n13729 ;
  assign n38205 = ~n13730 ;
  assign n14230 = n38205 & n150 ;
  assign n14231 = n13607 | n14230 ;
  assign n38206 = ~n14227 ;
  assign n14232 = n38206 & n14231 ;
  assign n14416 = n38185 & n14397 ;
  assign n14417 = n14255 | n14416 ;
  assign n38207 = ~n14399 ;
  assign n14418 = n38207 & n14417 ;
  assign n38208 = ~n14418 ;
  assign n14419 = n157 & n38208 ;
  assign n14420 = n38195 & n14417 ;
  assign n14421 = n14272 | n14420 ;
  assign n38209 = ~n14419 ;
  assign n14422 = n38209 & n14421 ;
  assign n38210 = ~n14422 ;
  assign n14423 = n158 & n38210 ;
  assign n14424 = n8857 | n14423 ;
  assign n38211 = ~n14424 ;
  assign n14425 = n14406 & n38211 ;
  assign n14426 = n14232 | n14425 ;
  assign n38212 = ~n14408 ;
  assign n14427 = n38212 & n14426 ;
  assign n38213 = ~n14427 ;
  assign n14428 = n160 & n38213 ;
  assign n13761 = n13733 | n13749 ;
  assign n38214 = ~n13761 ;
  assign n14228 = n38214 & n150 ;
  assign n14229 = n13625 | n14228 ;
  assign n38215 = ~n13749 ;
  assign n13759 = n13625 & n38215 ;
  assign n13760 = n37898 & n13759 ;
  assign n14276 = n13760 & n150 ;
  assign n38216 = ~n14276 ;
  assign n14277 = n14229 & n38216 ;
  assign n14409 = n160 | n14408 ;
  assign n38217 = ~n14409 ;
  assign n14429 = n38217 & n14426 ;
  assign n14430 = n14277 | n14429 ;
  assign n38218 = ~n14428 ;
  assign n14431 = n38218 & n14430 ;
  assign n38219 = ~n14431 ;
  assign n14432 = n161 & n38219 ;
  assign n13786 = n13629 & n37887 ;
  assign n38220 = ~n13753 ;
  assign n13787 = n38220 & n13786 ;
  assign n14275 = n13787 & n150 ;
  assign n13758 = n13752 | n13753 ;
  assign n38221 = ~n13758 ;
  assign n14289 = n38221 & n150 ;
  assign n14290 = n13629 | n14289 ;
  assign n38222 = ~n14275 ;
  assign n14291 = n38222 & n14290 ;
  assign n14440 = n38201 & n14421 ;
  assign n14441 = n14242 | n14440 ;
  assign n38223 = ~n14423 ;
  assign n14442 = n38223 & n14441 ;
  assign n38224 = ~n14442 ;
  assign n14443 = n159 & n38224 ;
  assign n14444 = n38211 & n14441 ;
  assign n14445 = n14232 | n14444 ;
  assign n38225 = ~n14443 ;
  assign n14446 = n38225 & n14445 ;
  assign n38226 = ~n14446 ;
  assign n14447 = n8534 & n38226 ;
  assign n14448 = n161 | n14447 ;
  assign n38227 = ~n14448 ;
  assign n14449 = n14430 & n38227 ;
  assign n14450 = n14291 | n14449 ;
  assign n38228 = ~n14432 ;
  assign n14451 = n38228 & n14450 ;
  assign n38229 = ~n14451 ;
  assign n14452 = n162 & n38229 ;
  assign n13785 = n13756 | n13773 ;
  assign n38230 = ~n13785 ;
  assign n14243 = n38230 & n150 ;
  assign n14244 = n13633 | n14243 ;
  assign n38231 = ~n13773 ;
  assign n13783 = n13633 & n38231 ;
  assign n13784 = n37914 & n13783 ;
  assign n14278 = n13784 & n150 ;
  assign n38232 = ~n14278 ;
  assign n14279 = n14244 & n38232 ;
  assign n14433 = n162 | n14432 ;
  assign n38233 = ~n14433 ;
  assign n14453 = n38233 & n14450 ;
  assign n14454 = n14279 | n14453 ;
  assign n38234 = ~n14452 ;
  assign n14455 = n38234 & n14454 ;
  assign n38235 = ~n14455 ;
  assign n14456 = n6889 & n38235 ;
  assign n13810 = n13638 & n37903 ;
  assign n38236 = ~n13777 ;
  assign n13811 = n38236 & n13810 ;
  assign n14284 = n13811 & n150 ;
  assign n13782 = n13776 | n13777 ;
  assign n38237 = ~n13782 ;
  assign n14292 = n38237 & n150 ;
  assign n14293 = n13638 | n14292 ;
  assign n38238 = ~n14284 ;
  assign n14294 = n38238 & n14293 ;
  assign n14464 = n38217 & n14445 ;
  assign n14465 = n14277 | n14464 ;
  assign n38239 = ~n14447 ;
  assign n14466 = n38239 & n14465 ;
  assign n38240 = ~n14466 ;
  assign n14467 = n161 & n38240 ;
  assign n14468 = n38227 & n14465 ;
  assign n14469 = n14291 | n14468 ;
  assign n38241 = ~n14467 ;
  assign n14470 = n38241 & n14469 ;
  assign n38242 = ~n14470 ;
  assign n14471 = n162 & n38242 ;
  assign n14472 = n6889 | n14471 ;
  assign n38243 = ~n14472 ;
  assign n14473 = n14454 & n38243 ;
  assign n14474 = n14294 | n14473 ;
  assign n38244 = ~n14456 ;
  assign n14475 = n38244 & n14474 ;
  assign n38245 = ~n14475 ;
  assign n14476 = n164 & n38245 ;
  assign n13809 = n13780 | n13797 ;
  assign n38246 = ~n13809 ;
  assign n14285 = n38246 & n150 ;
  assign n14286 = n13641 | n14285 ;
  assign n38247 = ~n13797 ;
  assign n13807 = n13641 & n38247 ;
  assign n13808 = n37930 & n13807 ;
  assign n14287 = n13808 & n150 ;
  assign n38248 = ~n14287 ;
  assign n14288 = n14286 & n38248 ;
  assign n14457 = n6600 | n14456 ;
  assign n38249 = ~n14457 ;
  assign n14477 = n38249 & n14474 ;
  assign n14478 = n14288 | n14477 ;
  assign n38250 = ~n14476 ;
  assign n14479 = n38250 & n14478 ;
  assign n38251 = ~n14479 ;
  assign n14480 = n165 & n38251 ;
  assign n13834 = n13644 & n37919 ;
  assign n38252 = ~n13801 ;
  assign n13835 = n38252 & n13834 ;
  assign n14297 = n13835 & n150 ;
  assign n13806 = n13800 | n13801 ;
  assign n38253 = ~n13806 ;
  assign n14298 = n38253 & n150 ;
  assign n14299 = n13644 | n14298 ;
  assign n38254 = ~n14297 ;
  assign n14300 = n38254 & n14299 ;
  assign n14488 = n38233 & n14469 ;
  assign n14489 = n14279 | n14488 ;
  assign n38255 = ~n14471 ;
  assign n14490 = n38255 & n14489 ;
  assign n38256 = ~n14490 ;
  assign n14491 = n163 & n38256 ;
  assign n14492 = n38243 & n14489 ;
  assign n14493 = n14294 | n14492 ;
  assign n38257 = ~n14491 ;
  assign n14494 = n38257 & n14493 ;
  assign n38258 = ~n14494 ;
  assign n14495 = n6600 & n38258 ;
  assign n14496 = n165 | n14495 ;
  assign n38259 = ~n14496 ;
  assign n14497 = n14478 & n38259 ;
  assign n14498 = n14300 | n14497 ;
  assign n38260 = ~n14480 ;
  assign n14499 = n38260 & n14498 ;
  assign n38261 = ~n14499 ;
  assign n14500 = n166 & n38261 ;
  assign n38262 = ~n13821 ;
  assign n13831 = n13646 & n38262 ;
  assign n13832 = n37946 & n13831 ;
  assign n14211 = n13832 & n150 ;
  assign n13833 = n13804 | n13821 ;
  assign n38263 = ~n13833 ;
  assign n14301 = n38263 & n150 ;
  assign n14302 = n13646 | n14301 ;
  assign n38264 = ~n14211 ;
  assign n14303 = n38264 & n14302 ;
  assign n14481 = n166 | n14480 ;
  assign n38265 = ~n14481 ;
  assign n14501 = n38265 & n14498 ;
  assign n14502 = n14303 | n14501 ;
  assign n38266 = ~n14500 ;
  assign n14503 = n38266 & n14502 ;
  assign n38267 = ~n14503 ;
  assign n14504 = n5352 & n38267 ;
  assign n13830 = n13824 | n13825 ;
  assign n38268 = ~n13830 ;
  assign n14249 = n38268 & n150 ;
  assign n14250 = n13594 | n14249 ;
  assign n13858 = n13594 & n37935 ;
  assign n38269 = ~n13825 ;
  assign n13859 = n38269 & n13858 ;
  assign n14295 = n13859 & n150 ;
  assign n38270 = ~n14295 ;
  assign n14296 = n14250 & n38270 ;
  assign n14512 = n38249 & n14493 ;
  assign n14513 = n14288 | n14512 ;
  assign n38271 = ~n14495 ;
  assign n14514 = n38271 & n14513 ;
  assign n38272 = ~n14514 ;
  assign n14515 = n165 & n38272 ;
  assign n14516 = n38259 & n14513 ;
  assign n14517 = n14300 | n14516 ;
  assign n38273 = ~n14515 ;
  assign n14518 = n38273 & n14517 ;
  assign n38274 = ~n14518 ;
  assign n14519 = n166 & n38274 ;
  assign n14520 = n5352 | n14519 ;
  assign n38275 = ~n14520 ;
  assign n14521 = n14502 & n38275 ;
  assign n14522 = n14296 | n14521 ;
  assign n38276 = ~n14504 ;
  assign n14523 = n38276 & n14522 ;
  assign n38277 = ~n14523 ;
  assign n14524 = n168 & n38277 ;
  assign n38278 = ~n13845 ;
  assign n13855 = n13567 & n38278 ;
  assign n13856 = n37962 & n13855 ;
  assign n14226 = n13856 & n150 ;
  assign n13857 = n13828 | n13845 ;
  assign n38279 = ~n13857 ;
  assign n14260 = n38279 & n150 ;
  assign n14261 = n13567 | n14260 ;
  assign n38280 = ~n14226 ;
  assign n14262 = n38280 & n14261 ;
  assign n14505 = n4934 | n14504 ;
  assign n38281 = ~n14505 ;
  assign n14525 = n38281 & n14522 ;
  assign n14526 = n14262 | n14525 ;
  assign n38282 = ~n14524 ;
  assign n14527 = n38282 & n14526 ;
  assign n38283 = ~n14527 ;
  assign n14528 = n169 & n38283 ;
  assign n13854 = n13848 | n13849 ;
  assign n38284 = ~n13854 ;
  assign n14224 = n38284 & n150 ;
  assign n14225 = n13596 | n14224 ;
  assign n13882 = n13596 & n37951 ;
  assign n38285 = ~n13849 ;
  assign n13883 = n38285 & n13882 ;
  assign n14273 = n13883 & n150 ;
  assign n38286 = ~n14273 ;
  assign n14274 = n14225 & n38286 ;
  assign n14536 = n38265 & n14517 ;
  assign n14537 = n14303 | n14536 ;
  assign n38287 = ~n14519 ;
  assign n14538 = n38287 & n14537 ;
  assign n38288 = ~n14538 ;
  assign n14539 = n167 & n38288 ;
  assign n14540 = n38275 & n14537 ;
  assign n14541 = n14296 | n14540 ;
  assign n38289 = ~n14539 ;
  assign n14542 = n38289 & n14541 ;
  assign n38290 = ~n14542 ;
  assign n14543 = n4934 & n38290 ;
  assign n14544 = n169 | n14543 ;
  assign n38291 = ~n14544 ;
  assign n14545 = n14526 & n38291 ;
  assign n14546 = n14274 | n14545 ;
  assign n38292 = ~n14528 ;
  assign n14547 = n38292 & n14546 ;
  assign n38293 = ~n14547 ;
  assign n14548 = n170 & n38293 ;
  assign n13881 = n13852 | n13869 ;
  assign n38294 = ~n13881 ;
  assign n14222 = n38294 & n150 ;
  assign n14223 = n13681 | n14222 ;
  assign n38295 = ~n13869 ;
  assign n13879 = n13681 & n38295 ;
  assign n13880 = n37978 & n13879 ;
  assign n14282 = n13880 & n150 ;
  assign n38296 = ~n14282 ;
  assign n14283 = n14223 & n38296 ;
  assign n14529 = n170 | n14528 ;
  assign n38297 = ~n14529 ;
  assign n14549 = n38297 & n14546 ;
  assign n14550 = n14283 | n14549 ;
  assign n38298 = ~n14548 ;
  assign n14551 = n38298 & n14550 ;
  assign n38299 = ~n14551 ;
  assign n14552 = n3940 & n38299 ;
  assign n13878 = n13872 | n13873 ;
  assign n38300 = ~n13878 ;
  assign n14217 = n38300 & n150 ;
  assign n14218 = n13683 | n14217 ;
  assign n13906 = n13683 & n37967 ;
  assign n38301 = ~n13873 ;
  assign n13907 = n38301 & n13906 ;
  assign n14247 = n13907 & n150 ;
  assign n38302 = ~n14247 ;
  assign n14248 = n14218 & n38302 ;
  assign n14560 = n38281 & n14541 ;
  assign n14561 = n14262 | n14560 ;
  assign n38303 = ~n14543 ;
  assign n14562 = n38303 & n14561 ;
  assign n38304 = ~n14562 ;
  assign n14563 = n169 & n38304 ;
  assign n14564 = n38291 & n14561 ;
  assign n14565 = n14274 | n14564 ;
  assign n38305 = ~n14563 ;
  assign n14566 = n38305 & n14565 ;
  assign n38306 = ~n14566 ;
  assign n14567 = n170 & n38306 ;
  assign n14568 = n3940 | n14567 ;
  assign n38307 = ~n14568 ;
  assign n14569 = n14550 & n38307 ;
  assign n14570 = n14248 | n14569 ;
  assign n38308 = ~n14552 ;
  assign n14571 = n38308 & n14570 ;
  assign n38309 = ~n14571 ;
  assign n14572 = n172 & n38309 ;
  assign n13905 = n13876 | n13893 ;
  assign n38310 = ~n13905 ;
  assign n14233 = n38310 & n150 ;
  assign n14234 = n13582 | n14233 ;
  assign n38311 = ~n13893 ;
  assign n13903 = n13582 & n38311 ;
  assign n13904 = n37994 & n13903 ;
  assign n14280 = n13904 & n150 ;
  assign n38312 = ~n14280 ;
  assign n14281 = n14234 & n38312 ;
  assign n14553 = n3631 | n14552 ;
  assign n38313 = ~n14553 ;
  assign n14573 = n38313 & n14570 ;
  assign n14574 = n14281 | n14573 ;
  assign n38314 = ~n14572 ;
  assign n14575 = n38314 & n14574 ;
  assign n38315 = ~n14575 ;
  assign n14576 = n173 & n38315 ;
  assign n13930 = n13555 & n37983 ;
  assign n38316 = ~n13897 ;
  assign n13931 = n38316 & n13930 ;
  assign n14220 = n13931 & n150 ;
  assign n13902 = n13896 | n13897 ;
  assign n38317 = ~n13902 ;
  assign n14267 = n38317 & n150 ;
  assign n14268 = n13555 | n14267 ;
  assign n38318 = ~n14220 ;
  assign n14269 = n38318 & n14268 ;
  assign n14584 = n38297 & n14565 ;
  assign n14585 = n14283 | n14584 ;
  assign n38319 = ~n14567 ;
  assign n14586 = n38319 & n14585 ;
  assign n38320 = ~n14586 ;
  assign n14587 = n171 & n38320 ;
  assign n14588 = n38307 & n14585 ;
  assign n14589 = n14248 | n14588 ;
  assign n38321 = ~n14587 ;
  assign n14590 = n38321 & n14589 ;
  assign n38322 = ~n14590 ;
  assign n14591 = n3631 & n38322 ;
  assign n14592 = n173 | n14591 ;
  assign n38323 = ~n14592 ;
  assign n14593 = n14574 & n38323 ;
  assign n14594 = n14269 | n14593 ;
  assign n38324 = ~n14576 ;
  assign n14595 = n38324 & n14594 ;
  assign n38325 = ~n14595 ;
  assign n14596 = n174 & n38325 ;
  assign n38326 = ~n13917 ;
  assign n13927 = n13577 & n38326 ;
  assign n13928 = n38010 & n13927 ;
  assign n14219 = n13928 & n150 ;
  assign n13929 = n13900 | n13917 ;
  assign n38327 = ~n13929 ;
  assign n14251 = n38327 & n150 ;
  assign n14252 = n13577 | n14251 ;
  assign n38328 = ~n14219 ;
  assign n14253 = n38328 & n14252 ;
  assign n14577 = n174 | n14576 ;
  assign n38329 = ~n14577 ;
  assign n14597 = n38329 & n14594 ;
  assign n14598 = n14253 | n14597 ;
  assign n38330 = ~n14596 ;
  assign n14599 = n38330 & n14598 ;
  assign n38331 = ~n14599 ;
  assign n14600 = n2753 & n38331 ;
  assign n13926 = n13920 | n13921 ;
  assign n38332 = ~n13926 ;
  assign n14213 = n38332 & n150 ;
  assign n14214 = n13627 | n14213 ;
  assign n13954 = n13627 & n37999 ;
  assign n38333 = ~n13921 ;
  assign n13955 = n38333 & n13954 ;
  assign n14215 = n13955 & n150 ;
  assign n38334 = ~n14215 ;
  assign n14216 = n14214 & n38334 ;
  assign n14608 = n38313 & n14589 ;
  assign n14609 = n14281 | n14608 ;
  assign n38335 = ~n14591 ;
  assign n14610 = n38335 & n14609 ;
  assign n38336 = ~n14610 ;
  assign n14611 = n173 & n38336 ;
  assign n14612 = n38323 & n14609 ;
  assign n14613 = n14269 | n14612 ;
  assign n38337 = ~n14611 ;
  assign n14614 = n38337 & n14613 ;
  assign n38338 = ~n14614 ;
  assign n14615 = n174 & n38338 ;
  assign n14616 = n2753 | n14615 ;
  assign n38339 = ~n14616 ;
  assign n14617 = n14598 & n38339 ;
  assign n14618 = n14216 | n14617 ;
  assign n38340 = ~n14600 ;
  assign n14619 = n38340 & n14618 ;
  assign n38341 = ~n14619 ;
  assign n14620 = n176 & n38341 ;
  assign n13953 = n13924 | n13941 ;
  assign n38342 = ~n13953 ;
  assign n14208 = n38342 & n150 ;
  assign n14209 = n13552 | n14208 ;
  assign n38343 = ~n13941 ;
  assign n13951 = n13552 & n38343 ;
  assign n13952 = n38026 & n13951 ;
  assign n14245 = n13952 & n150 ;
  assign n38344 = ~n14245 ;
  assign n14246 = n14209 & n38344 ;
  assign n14601 = n2431 | n14600 ;
  assign n38345 = ~n14601 ;
  assign n14621 = n38345 & n14618 ;
  assign n14622 = n14246 | n14621 ;
  assign n38346 = ~n14620 ;
  assign n14623 = n38346 & n14622 ;
  assign n38347 = ~n14623 ;
  assign n14624 = n177 & n38347 ;
  assign n13967 = n13546 & n38015 ;
  assign n38348 = ~n13945 ;
  assign n13968 = n38348 & n13967 ;
  assign n14212 = n13968 & n150 ;
  assign n13950 = n13944 | n13945 ;
  assign n38349 = ~n13950 ;
  assign n14256 = n38349 & n150 ;
  assign n14257 = n13546 | n14256 ;
  assign n38350 = ~n14212 ;
  assign n14258 = n38350 & n14257 ;
  assign n14632 = n38329 & n14613 ;
  assign n14633 = n14253 | n14632 ;
  assign n38351 = ~n14615 ;
  assign n14634 = n38351 & n14633 ;
  assign n38352 = ~n14634 ;
  assign n14635 = n175 & n38352 ;
  assign n14636 = n38339 & n14633 ;
  assign n14637 = n14216 | n14636 ;
  assign n38353 = ~n14635 ;
  assign n14638 = n38353 & n14637 ;
  assign n38354 = ~n14638 ;
  assign n14639 = n2431 & n38354 ;
  assign n14640 = n177 | n14639 ;
  assign n38355 = ~n14640 ;
  assign n14641 = n14622 & n38355 ;
  assign n14642 = n14258 | n14641 ;
  assign n38356 = ~n14624 ;
  assign n14643 = n38356 & n14642 ;
  assign n38357 = ~n14643 ;
  assign n14644 = n178 & n38357 ;
  assign n14625 = n178 | n14624 ;
  assign n38358 = ~n14625 ;
  assign n14645 = n38358 & n14642 ;
  assign n38359 = ~n13965 ;
  assign n14081 = n38359 & n14065 ;
  assign n14082 = n38042 & n14081 ;
  assign n14210 = n14082 & n150 ;
  assign n13966 = n13948 | n13965 ;
  assign n38360 = ~n13966 ;
  assign n14235 = n38360 & n150 ;
  assign n14758 = n14065 | n14235 ;
  assign n38361 = ~n14210 ;
  assign n14759 = n38361 & n14758 ;
  assign n14760 = n14645 | n14759 ;
  assign n38362 = ~n14644 ;
  assign n14761 = n38362 & n14760 ;
  assign n38363 = ~n14761 ;
  assign n14762 = n1707 & n38363 ;
  assign n14070 = n14063 & n38031 ;
  assign n38364 = ~n14086 ;
  assign n14752 = n14070 & n38364 ;
  assign n14753 = n150 & n14752 ;
  assign n14754 = n14085 | n14086 ;
  assign n38365 = ~n14754 ;
  assign n14755 = n150 & n38365 ;
  assign n14756 = n14063 | n14755 ;
  assign n38366 = ~n14753 ;
  assign n14757 = n38366 & n14756 ;
  assign n14649 = n38345 & n14637 ;
  assign n14650 = n14246 | n14649 ;
  assign n38367 = ~n14639 ;
  assign n14651 = n38367 & n14650 ;
  assign n38368 = ~n14651 ;
  assign n14652 = n177 & n38368 ;
  assign n14653 = n38355 & n14650 ;
  assign n14654 = n14258 | n14653 ;
  assign n38369 = ~n14652 ;
  assign n14655 = n38369 & n14654 ;
  assign n38370 = ~n14655 ;
  assign n14656 = n178 & n38370 ;
  assign n14657 = n1707 | n14656 ;
  assign n38371 = ~n14657 ;
  assign n14765 = n38371 & n14760 ;
  assign n14766 = n14757 | n14765 ;
  assign n38372 = ~n14762 ;
  assign n14767 = n38372 & n14766 ;
  assign n38373 = ~n14767 ;
  assign n14768 = n180 & n38373 ;
  assign n38374 = ~n14101 ;
  assign n14745 = n14057 & n38374 ;
  assign n14746 = n38058 & n14745 ;
  assign n14747 = n150 & n14746 ;
  assign n14748 = n14089 | n14101 ;
  assign n38375 = ~n14748 ;
  assign n14749 = n150 & n38375 ;
  assign n14750 = n14057 | n14749 ;
  assign n38376 = ~n14747 ;
  assign n14751 = n38376 & n14750 ;
  assign n14763 = n1487 | n14762 ;
  assign n38377 = ~n14763 ;
  assign n14769 = n38377 & n14766 ;
  assign n14770 = n14751 | n14769 ;
  assign n38378 = ~n14768 ;
  assign n14771 = n38378 & n14770 ;
  assign n38379 = ~n14771 ;
  assign n14772 = n181 & n38379 ;
  assign n14080 = n14050 & n38047 ;
  assign n38380 = ~n14105 ;
  assign n14739 = n14080 & n38380 ;
  assign n14740 = n150 & n14739 ;
  assign n14741 = n14104 | n14105 ;
  assign n38381 = ~n14741 ;
  assign n14742 = n150 & n38381 ;
  assign n14743 = n14050 | n14742 ;
  assign n38382 = ~n14740 ;
  assign n14744 = n38382 & n14743 ;
  assign n14659 = n38358 & n14654 ;
  assign n14779 = n14659 | n14759 ;
  assign n38383 = ~n14656 ;
  assign n14780 = n38383 & n14779 ;
  assign n38384 = ~n14780 ;
  assign n14781 = n179 & n38384 ;
  assign n14782 = n38371 & n14779 ;
  assign n14783 = n14757 | n14782 ;
  assign n38385 = ~n14781 ;
  assign n14784 = n38385 & n14783 ;
  assign n38386 = ~n14784 ;
  assign n14785 = n1487 & n38386 ;
  assign n14786 = n181 | n14785 ;
  assign n38387 = ~n14786 ;
  assign n14787 = n14770 & n38387 ;
  assign n14788 = n14744 | n14787 ;
  assign n38388 = ~n14772 ;
  assign n14789 = n38388 & n14788 ;
  assign n38389 = ~n14789 ;
  assign n14790 = n182 & n38389 ;
  assign n14732 = n14108 | n14120 ;
  assign n38390 = ~n14732 ;
  assign n14733 = n150 & n38390 ;
  assign n14734 = n14044 | n14733 ;
  assign n38391 = ~n14120 ;
  assign n14735 = n14044 & n38391 ;
  assign n14736 = n38074 & n14735 ;
  assign n14737 = n150 & n14736 ;
  assign n38392 = ~n14737 ;
  assign n14738 = n14734 & n38392 ;
  assign n14773 = n182 | n14772 ;
  assign n38393 = ~n14773 ;
  assign n14791 = n38393 & n14788 ;
  assign n14792 = n14738 | n14791 ;
  assign n38394 = ~n14790 ;
  assign n14793 = n38394 & n14792 ;
  assign n38395 = ~n14793 ;
  assign n14794 = n996 & n38395 ;
  assign n14100 = n14037 & n38063 ;
  assign n38396 = ~n14124 ;
  assign n14726 = n14100 & n38396 ;
  assign n14727 = n150 & n14726 ;
  assign n14728 = n14123 | n14124 ;
  assign n38397 = ~n14728 ;
  assign n14729 = n150 & n38397 ;
  assign n14730 = n14037 | n14729 ;
  assign n38398 = ~n14727 ;
  assign n14731 = n38398 & n14730 ;
  assign n14802 = n38377 & n14783 ;
  assign n14803 = n14751 | n14802 ;
  assign n38399 = ~n14785 ;
  assign n14804 = n38399 & n14803 ;
  assign n38400 = ~n14804 ;
  assign n14805 = n181 & n38400 ;
  assign n14806 = n38387 & n14803 ;
  assign n14807 = n14744 | n14806 ;
  assign n38401 = ~n14805 ;
  assign n14808 = n38401 & n14807 ;
  assign n38402 = ~n14808 ;
  assign n14809 = n182 & n38402 ;
  assign n14810 = n183 | n14809 ;
  assign n38403 = ~n14810 ;
  assign n14811 = n14792 & n38403 ;
  assign n14812 = n14731 | n14811 ;
  assign n38404 = ~n14794 ;
  assign n14813 = n38404 & n14812 ;
  assign n38405 = ~n14813 ;
  assign n14814 = n184 & n38405 ;
  assign n38406 = ~n14139 ;
  assign n14719 = n14031 & n38406 ;
  assign n14720 = n38090 & n14719 ;
  assign n14721 = n150 & n14720 ;
  assign n14722 = n14127 | n14139 ;
  assign n38407 = ~n14722 ;
  assign n14723 = n150 & n38407 ;
  assign n14724 = n14031 | n14723 ;
  assign n38408 = ~n14721 ;
  assign n14725 = n38408 & n14724 ;
  assign n14795 = n838 | n14794 ;
  assign n38409 = ~n14795 ;
  assign n14815 = n38409 & n14812 ;
  assign n14816 = n14725 | n14815 ;
  assign n38410 = ~n14814 ;
  assign n14817 = n38410 & n14816 ;
  assign n38411 = ~n14817 ;
  assign n14818 = n185 & n38411 ;
  assign n14119 = n13648 & n38079 ;
  assign n38412 = ~n14143 ;
  assign n14713 = n14119 & n38412 ;
  assign n14714 = n150 & n14713 ;
  assign n14715 = n14142 | n14143 ;
  assign n38413 = ~n14715 ;
  assign n14716 = n150 & n38413 ;
  assign n14717 = n13648 | n14716 ;
  assign n38414 = ~n14714 ;
  assign n14718 = n38414 & n14717 ;
  assign n14826 = n38393 & n14807 ;
  assign n14827 = n14738 | n14826 ;
  assign n38415 = ~n14809 ;
  assign n14828 = n38415 & n14827 ;
  assign n38416 = ~n14828 ;
  assign n14829 = n183 & n38416 ;
  assign n14830 = n38403 & n14827 ;
  assign n14831 = n14731 | n14830 ;
  assign n38417 = ~n14829 ;
  assign n14832 = n38417 & n14831 ;
  assign n38418 = ~n14832 ;
  assign n14833 = n838 & n38418 ;
  assign n14834 = n185 | n14833 ;
  assign n38419 = ~n14834 ;
  assign n14835 = n14816 & n38419 ;
  assign n14836 = n14718 | n14835 ;
  assign n38420 = ~n14818 ;
  assign n14837 = n38420 & n14836 ;
  assign n38421 = ~n14837 ;
  assign n14838 = n186 & n38421 ;
  assign n14706 = n14146 | n14158 ;
  assign n38422 = ~n14706 ;
  assign n14707 = n150 & n38422 ;
  assign n14708 = n14024 | n14707 ;
  assign n38423 = ~n14158 ;
  assign n14709 = n14024 & n38423 ;
  assign n14710 = n38106 & n14709 ;
  assign n14711 = n150 & n14710 ;
  assign n38424 = ~n14711 ;
  assign n14712 = n14708 & n38424 ;
  assign n14819 = n186 | n14818 ;
  assign n38425 = ~n14819 ;
  assign n14839 = n38425 & n14836 ;
  assign n14840 = n14712 | n14839 ;
  assign n38426 = ~n14838 ;
  assign n14841 = n38426 & n14840 ;
  assign n38427 = ~n14841 ;
  assign n14842 = n528 & n38427 ;
  assign n14138 = n14017 & n38095 ;
  assign n38428 = ~n14162 ;
  assign n14163 = n14138 & n38428 ;
  assign n14221 = n14163 & n150 ;
  assign n14164 = n14161 | n14162 ;
  assign n38429 = ~n14164 ;
  assign n14304 = n38429 & n150 ;
  assign n14305 = n14017 | n14304 ;
  assign n38430 = ~n14221 ;
  assign n14306 = n38430 & n14305 ;
  assign n14850 = n38409 & n14831 ;
  assign n14851 = n14725 | n14850 ;
  assign n38431 = ~n14833 ;
  assign n14852 = n38431 & n14851 ;
  assign n38432 = ~n14852 ;
  assign n14853 = n185 & n38432 ;
  assign n14854 = n38419 & n14851 ;
  assign n14855 = n14718 | n14854 ;
  assign n38433 = ~n14853 ;
  assign n14856 = n38433 & n14855 ;
  assign n38434 = ~n14856 ;
  assign n14857 = n186 & n38434 ;
  assign n14858 = n528 | n14857 ;
  assign n38435 = ~n14858 ;
  assign n14859 = n14840 & n38435 ;
  assign n14860 = n14306 | n14859 ;
  assign n38436 = ~n14842 ;
  assign n14861 = n38436 & n14860 ;
  assign n38437 = ~n14861 ;
  assign n14862 = n188 & n38437 ;
  assign n38438 = ~n14179 ;
  assign n14699 = n14011 & n38438 ;
  assign n14700 = n38123 & n14699 ;
  assign n14701 = n150 & n14700 ;
  assign n14702 = n14167 | n14179 ;
  assign n38439 = ~n14702 ;
  assign n14703 = n150 & n38439 ;
  assign n14704 = n14011 | n14703 ;
  assign n38440 = ~n14701 ;
  assign n14705 = n38440 & n14704 ;
  assign n14843 = n413 | n14842 ;
  assign n38441 = ~n14843 ;
  assign n14863 = n38441 & n14860 ;
  assign n14864 = n14705 | n14863 ;
  assign n38442 = ~n14862 ;
  assign n14865 = n38442 & n14864 ;
  assign n38443 = ~n14865 ;
  assign n14866 = n189 & n38443 ;
  assign n14157 = n14004 & n38111 ;
  assign n38444 = ~n14183 ;
  assign n14693 = n14157 & n38444 ;
  assign n14694 = n150 & n14693 ;
  assign n14695 = n14182 | n14183 ;
  assign n38445 = ~n14695 ;
  assign n14696 = n150 & n38445 ;
  assign n14697 = n14004 | n14696 ;
  assign n38446 = ~n14694 ;
  assign n14698 = n38446 & n14697 ;
  assign n14874 = n38425 & n14855 ;
  assign n14875 = n14712 | n14874 ;
  assign n38447 = ~n14857 ;
  assign n14876 = n38447 & n14875 ;
  assign n38448 = ~n14876 ;
  assign n14877 = n187 & n38448 ;
  assign n14878 = n38435 & n14875 ;
  assign n14879 = n14306 | n14878 ;
  assign n38449 = ~n14877 ;
  assign n14880 = n38449 & n14879 ;
  assign n38450 = ~n14880 ;
  assign n14881 = n413 & n38450 ;
  assign n14882 = n189 | n14881 ;
  assign n38451 = ~n14882 ;
  assign n14883 = n14864 & n38451 ;
  assign n14884 = n14698 | n14883 ;
  assign n38452 = ~n14866 ;
  assign n14885 = n38452 & n14884 ;
  assign n38453 = ~n14885 ;
  assign n14886 = n190 & n38453 ;
  assign n38454 = ~n14188 ;
  assign n14686 = n13998 & n38454 ;
  assign n14687 = n38129 & n14686 ;
  assign n14688 = n150 & n14687 ;
  assign n14689 = n14186 | n14188 ;
  assign n38455 = ~n14689 ;
  assign n14690 = n150 & n38455 ;
  assign n14691 = n13998 | n14690 ;
  assign n38456 = ~n14688 ;
  assign n14692 = n38456 & n14691 ;
  assign n14867 = n190 | n14866 ;
  assign n38457 = ~n14867 ;
  assign n14887 = n38457 & n14884 ;
  assign n14888 = n14692 | n14887 ;
  assign n38458 = ~n14886 ;
  assign n14889 = n38458 & n14888 ;
  assign n38459 = ~n14889 ;
  assign n14890 = n287 & n38459 ;
  assign n38460 = ~n14176 ;
  assign n14178 = n13991 & n38460 ;
  assign n38461 = ~n14192 ;
  assign n14680 = n14178 & n38461 ;
  assign n14681 = n150 & n14680 ;
  assign n14682 = n14191 | n14192 ;
  assign n38462 = ~n14682 ;
  assign n14683 = n150 & n38462 ;
  assign n14684 = n13991 | n14683 ;
  assign n38463 = ~n14681 ;
  assign n14685 = n38463 & n14684 ;
  assign n14898 = n38441 & n14879 ;
  assign n14899 = n14705 | n14898 ;
  assign n38464 = ~n14881 ;
  assign n14900 = n38464 & n14899 ;
  assign n38465 = ~n14900 ;
  assign n14901 = n189 & n38465 ;
  assign n14902 = n38451 & n14899 ;
  assign n14903 = n14698 | n14902 ;
  assign n38466 = ~n14901 ;
  assign n14904 = n38466 & n14903 ;
  assign n38467 = ~n14904 ;
  assign n14905 = n190 & n38467 ;
  assign n14906 = n287 | n14905 ;
  assign n38468 = ~n14906 ;
  assign n14907 = n14888 & n38468 ;
  assign n14910 = n14685 | n14907 ;
  assign n38469 = ~n14890 ;
  assign n14911 = n38469 & n14910 ;
  assign n14914 = n14677 | n14911 ;
  assign n14915 = n31336 & n14914 ;
  assign n14203 = n192 & n14202 ;
  assign n38470 = ~n13658 ;
  assign n14326 = n38470 & n150 ;
  assign n38471 = ~n14326 ;
  assign n14327 = n14199 & n38471 ;
  assign n38472 = ~n14327 ;
  assign n14328 = n14203 & n38472 ;
  assign n13982 = n13654 | n13976 ;
  assign n38473 = ~n13982 ;
  assign n13983 = n13657 & n38473 ;
  assign n13984 = n38153 & n13983 ;
  assign n14661 = n13984 & n38154 ;
  assign n14662 = n38155 & n14661 ;
  assign n14663 = n14328 | n14662 ;
  assign n14891 = n14676 & n38469 ;
  assign n14916 = n14891 & n14910 ;
  assign n14917 = n14663 | n14916 ;
  assign n149 = n14915 | n14917 ;
  assign n14909 = n14890 | n14907 ;
  assign n38474 = ~n14909 ;
  assign n14924 = n38474 & n149 ;
  assign n14925 = n14685 | n14924 ;
  assign n14892 = n14685 & n38469 ;
  assign n38475 = ~n14907 ;
  assign n14908 = n14892 & n38475 ;
  assign n15078 = n14908 & n149 ;
  assign n38476 = ~n15078 ;
  assign n15079 = n14925 & n38476 ;
  assign n14912 = n14676 | n14911 ;
  assign n38477 = ~n14912 ;
  assign n15082 = n38477 & n149 ;
  assign n15447 = n14916 | n15082 ;
  assign n15448 = n15079 | n15447 ;
  assign n212 = x38 | x39 ;
  assign n213 = x40 | n212 ;
  assign n15003 = x40 & n149 ;
  assign n38478 = ~n15003 ;
  assign n15022 = n213 & n38478 ;
  assign n38479 = ~n15022 ;
  assign n15023 = n150 & n38479 ;
  assign n13980 = n213 & n38152 ;
  assign n13981 = n38153 & n13980 ;
  assign n14668 = n13981 & n38154 ;
  assign n14669 = n38155 & n14668 ;
  assign n15004 = n14669 & n38478 ;
  assign n38480 = ~n209 ;
  assign n14997 = n38480 & n149 ;
  assign n38481 = ~x40 ;
  assign n15092 = n38481 & n149 ;
  assign n38482 = ~n15092 ;
  assign n15093 = x41 & n38482 ;
  assign n15094 = n14997 | n15093 ;
  assign n15096 = n15004 | n15094 ;
  assign n38483 = ~n15023 ;
  assign n15097 = n38483 & n15096 ;
  assign n38484 = ~n15097 ;
  assign n15098 = n13662 & n38484 ;
  assign n214 = n38481 & n212 ;
  assign n38485 = ~n149 ;
  assign n15085 = x40 & n38485 ;
  assign n15086 = n214 | n15085 ;
  assign n38486 = ~n15086 ;
  assign n15087 = n150 & n38486 ;
  assign n15088 = n13662 | n15087 ;
  assign n38487 = ~n15088 ;
  assign n15101 = n38487 & n15096 ;
  assign n38488 = ~n14662 ;
  assign n14664 = n150 & n38488 ;
  assign n38489 = ~n14328 ;
  assign n14665 = n38489 & n14664 ;
  assign n38490 = ~n14916 ;
  assign n15104 = n14665 & n38490 ;
  assign n38491 = ~n14915 ;
  assign n15105 = n38491 & n15104 ;
  assign n15106 = n14997 | n15105 ;
  assign n15107 = x42 & n15106 ;
  assign n15108 = x42 | n15105 ;
  assign n15109 = n14997 | n15108 ;
  assign n38492 = ~n15107 ;
  assign n15110 = n38492 & n15109 ;
  assign n15111 = n15101 | n15110 ;
  assign n38493 = ~n15098 ;
  assign n15112 = n38493 & n15111 ;
  assign n38494 = ~n15112 ;
  assign n15113 = n13079 & n38494 ;
  assign n14313 = n14308 | n14311 ;
  assign n38495 = ~n14313 ;
  assign n14334 = n38495 & n14331 ;
  assign n14996 = n14334 & n149 ;
  assign n15036 = n38495 & n149 ;
  assign n15037 = n14331 | n15036 ;
  assign n38496 = ~n14996 ;
  assign n15038 = n38496 & n15037 ;
  assign n15099 = n13079 | n15098 ;
  assign n38497 = ~n15099 ;
  assign n15116 = n38497 & n15111 ;
  assign n15117 = n15038 | n15116 ;
  assign n38498 = ~n15113 ;
  assign n15118 = n38498 & n15117 ;
  assign n38499 = ~n15118 ;
  assign n15119 = n153 & n38499 ;
  assign n14339 = n14333 | n14338 ;
  assign n38500 = ~n14339 ;
  assign n15029 = n38500 & n149 ;
  assign n15030 = n14347 | n15029 ;
  assign n38501 = ~n14333 ;
  assign n14367 = n38501 & n14347 ;
  assign n14368 = n38157 & n14367 ;
  assign n15080 = n14368 & n149 ;
  assign n38502 = ~n15080 ;
  assign n15081 = n15030 & n38502 ;
  assign n15114 = n153 | n15113 ;
  assign n38503 = ~n15114 ;
  assign n15120 = n38503 & n15117 ;
  assign n15121 = n15081 | n15120 ;
  assign n38504 = ~n15119 ;
  assign n15122 = n38504 & n15121 ;
  assign n38505 = ~n15122 ;
  assign n15123 = n154 & n38505 ;
  assign n14365 = n14350 | n14353 ;
  assign n38506 = ~n14365 ;
  assign n14976 = n38506 & n149 ;
  assign n14977 = n14319 | n14976 ;
  assign n14352 = n14319 & n38162 ;
  assign n38507 = ~n14353 ;
  assign n14366 = n14352 & n38507 ;
  assign n15083 = n14366 & n149 ;
  assign n38508 = ~n15083 ;
  assign n15084 = n14977 & n38508 ;
  assign n15100 = n151 & n38484 ;
  assign n15024 = n151 | n15023 ;
  assign n38509 = ~n15024 ;
  assign n15103 = n38509 & n15096 ;
  assign n15133 = n15103 | n15110 ;
  assign n38510 = ~n15100 ;
  assign n15134 = n38510 & n15133 ;
  assign n38511 = ~n15134 ;
  assign n15135 = n152 & n38511 ;
  assign n15136 = n38497 & n15133 ;
  assign n15137 = n15038 | n15136 ;
  assign n38512 = ~n15135 ;
  assign n15138 = n38512 & n15137 ;
  assign n38513 = ~n15138 ;
  assign n15139 = n153 & n38513 ;
  assign n15140 = n154 | n15139 ;
  assign n38514 = ~n15140 ;
  assign n15141 = n15121 & n38514 ;
  assign n15142 = n15084 | n15141 ;
  assign n38515 = ~n15123 ;
  assign n15143 = n38515 & n15142 ;
  assign n38516 = ~n15143 ;
  assign n15144 = n155 & n38516 ;
  assign n38517 = ~n14357 ;
  assign n14363 = n14321 & n38517 ;
  assign n14364 = n38169 & n14363 ;
  assign n14965 = n14364 & n149 ;
  assign n14391 = n14357 | n14375 ;
  assign n38518 = ~n14391 ;
  assign n14978 = n38518 & n149 ;
  assign n14979 = n14321 | n14978 ;
  assign n38519 = ~n14965 ;
  assign n14980 = n38519 & n14979 ;
  assign n15124 = n11067 | n15123 ;
  assign n38520 = ~n15124 ;
  assign n15145 = n38520 & n15142 ;
  assign n15146 = n14980 | n15145 ;
  assign n38521 = ~n15144 ;
  assign n15147 = n38521 & n15146 ;
  assign n38522 = ~n15147 ;
  assign n15148 = n10657 & n38522 ;
  assign n14362 = n14325 & n38180 ;
  assign n38523 = ~n14377 ;
  assign n14390 = n14362 & n38523 ;
  assign n14953 = n14390 & n149 ;
  assign n14389 = n14360 | n14377 ;
  assign n38524 = ~n14389 ;
  assign n14973 = n38524 & n149 ;
  assign n14974 = n14325 | n14973 ;
  assign n38525 = ~n14953 ;
  assign n14975 = n38525 & n14974 ;
  assign n15156 = n38503 & n15137 ;
  assign n15157 = n15081 | n15156 ;
  assign n38526 = ~n15139 ;
  assign n15158 = n38526 & n15157 ;
  assign n38527 = ~n15158 ;
  assign n15159 = n154 & n38527 ;
  assign n15160 = n38514 & n15157 ;
  assign n15161 = n15084 | n15160 ;
  assign n38528 = ~n15159 ;
  assign n15162 = n38528 & n15161 ;
  assign n38529 = ~n15162 ;
  assign n15163 = n11067 & n38529 ;
  assign n15164 = n10657 | n15163 ;
  assign n38530 = ~n15164 ;
  assign n15165 = n15146 & n38530 ;
  assign n15166 = n14975 | n15165 ;
  assign n38531 = ~n15148 ;
  assign n15167 = n38531 & n15166 ;
  assign n38532 = ~n15167 ;
  assign n15168 = n157 & n38532 ;
  assign n14415 = n14381 | n14399 ;
  assign n38533 = ~n14415 ;
  assign n14981 = n38533 & n149 ;
  assign n14982 = n14255 | n14981 ;
  assign n38534 = ~n14381 ;
  assign n14387 = n14255 & n38534 ;
  assign n14388 = n38186 & n14387 ;
  assign n14983 = n14388 & n149 ;
  assign n38535 = ~n14983 ;
  assign n14984 = n14982 & n38535 ;
  assign n15149 = n157 | n15148 ;
  assign n38536 = ~n15149 ;
  assign n15169 = n38536 & n15166 ;
  assign n15170 = n14984 | n15169 ;
  assign n38537 = ~n15168 ;
  assign n15171 = n38537 & n15170 ;
  assign n38538 = ~n15171 ;
  assign n15172 = n158 & n38538 ;
  assign n14413 = n14384 | n14401 ;
  assign n38539 = ~n14413 ;
  assign n14945 = n38539 & n149 ;
  assign n14946 = n14272 | n14945 ;
  assign n14386 = n14272 & n38196 ;
  assign n38540 = ~n14401 ;
  assign n14414 = n14386 & n38540 ;
  assign n15015 = n14414 & n149 ;
  assign n38541 = ~n15015 ;
  assign n15016 = n14946 & n38541 ;
  assign n15180 = n38520 & n15161 ;
  assign n15181 = n14980 | n15180 ;
  assign n38542 = ~n15163 ;
  assign n15182 = n38542 & n15181 ;
  assign n38543 = ~n15182 ;
  assign n15183 = n156 & n38543 ;
  assign n15184 = n38530 & n15181 ;
  assign n15185 = n14975 | n15184 ;
  assign n38544 = ~n15183 ;
  assign n15186 = n38544 & n15185 ;
  assign n38545 = ~n15186 ;
  assign n15187 = n157 & n38545 ;
  assign n15188 = n158 | n15187 ;
  assign n38546 = ~n15188 ;
  assign n15189 = n15170 & n38546 ;
  assign n15190 = n15016 | n15189 ;
  assign n38547 = ~n15172 ;
  assign n15191 = n38547 & n15190 ;
  assign n38548 = ~n15191 ;
  assign n15192 = n159 & n38548 ;
  assign n38549 = ~n14405 ;
  assign n14411 = n14242 & n38549 ;
  assign n14412 = n38202 & n14411 ;
  assign n14969 = n14412 & n149 ;
  assign n14439 = n14405 | n14423 ;
  assign n38550 = ~n14439 ;
  assign n15026 = n38550 & n149 ;
  assign n15027 = n14242 | n15026 ;
  assign n38551 = ~n14969 ;
  assign n15028 = n38551 & n15027 ;
  assign n15173 = n8857 | n15172 ;
  assign n38552 = ~n15173 ;
  assign n15193 = n38552 & n15190 ;
  assign n15194 = n15028 | n15193 ;
  assign n38553 = ~n15192 ;
  assign n15195 = n38553 & n15194 ;
  assign n38554 = ~n15195 ;
  assign n15196 = n8534 & n38554 ;
  assign n14410 = n14232 & n38212 ;
  assign n38555 = ~n14425 ;
  assign n14437 = n14410 & n38555 ;
  assign n14929 = n14437 & n149 ;
  assign n14438 = n14408 | n14425 ;
  assign n38556 = ~n14438 ;
  assign n14970 = n38556 & n149 ;
  assign n14971 = n14232 | n14970 ;
  assign n38557 = ~n14929 ;
  assign n14972 = n38557 & n14971 ;
  assign n15204 = n38536 & n15185 ;
  assign n15205 = n14984 | n15204 ;
  assign n38558 = ~n15187 ;
  assign n15206 = n38558 & n15205 ;
  assign n38559 = ~n15206 ;
  assign n15207 = n158 & n38559 ;
  assign n15208 = n38546 & n15205 ;
  assign n15209 = n15016 | n15208 ;
  assign n38560 = ~n15207 ;
  assign n15210 = n38560 & n15209 ;
  assign n38561 = ~n15210 ;
  assign n15211 = n8857 & n38561 ;
  assign n15212 = n160 | n15211 ;
  assign n38562 = ~n15212 ;
  assign n15213 = n15194 & n38562 ;
  assign n15214 = n14972 | n15213 ;
  assign n38563 = ~n15196 ;
  assign n15215 = n38563 & n15214 ;
  assign n38564 = ~n15215 ;
  assign n15216 = n161 & n38564 ;
  assign n38565 = ~n14429 ;
  assign n14435 = n14277 & n38565 ;
  assign n14436 = n38218 & n14435 ;
  assign n14992 = n14436 & n149 ;
  assign n14463 = n14429 | n14447 ;
  assign n38566 = ~n14463 ;
  assign n15033 = n38566 & n149 ;
  assign n15034 = n14277 | n15033 ;
  assign n38567 = ~n14992 ;
  assign n15035 = n38567 & n15034 ;
  assign n15197 = n161 | n15196 ;
  assign n38568 = ~n15197 ;
  assign n15217 = n38568 & n15214 ;
  assign n15221 = n15035 | n15217 ;
  assign n38569 = ~n15216 ;
  assign n15222 = n38569 & n15221 ;
  assign n38570 = ~n15222 ;
  assign n15223 = n162 & n38570 ;
  assign n14462 = n14432 | n14449 ;
  assign n38571 = ~n14462 ;
  assign n14987 = n38571 & n149 ;
  assign n14988 = n14291 | n14987 ;
  assign n14434 = n14291 & n38228 ;
  assign n38572 = ~n14449 ;
  assign n14461 = n14434 & n38572 ;
  assign n15039 = n14461 & n149 ;
  assign n38573 = ~n15039 ;
  assign n15040 = n14988 & n38573 ;
  assign n15228 = n38552 & n15209 ;
  assign n15229 = n15028 | n15228 ;
  assign n38574 = ~n15211 ;
  assign n15230 = n38574 & n15229 ;
  assign n38575 = ~n15230 ;
  assign n15231 = n160 & n38575 ;
  assign n15232 = n38562 & n15229 ;
  assign n15233 = n14972 | n15232 ;
  assign n38576 = ~n15231 ;
  assign n15234 = n38576 & n15233 ;
  assign n38577 = ~n15234 ;
  assign n15235 = n161 & n38577 ;
  assign n15236 = n162 | n15235 ;
  assign n38578 = ~n15236 ;
  assign n15237 = n15221 & n38578 ;
  assign n15238 = n15040 | n15237 ;
  assign n38579 = ~n15223 ;
  assign n15239 = n38579 & n15238 ;
  assign n38580 = ~n15239 ;
  assign n15240 = n163 & n38580 ;
  assign n14487 = n14453 | n14471 ;
  assign n38581 = ~n14487 ;
  assign n15010 = n38581 & n149 ;
  assign n15011 = n14279 | n15010 ;
  assign n38582 = ~n14453 ;
  assign n14459 = n14279 & n38582 ;
  assign n14460 = n38234 & n14459 ;
  assign n15017 = n14460 & n149 ;
  assign n38583 = ~n15017 ;
  assign n15018 = n15011 & n38583 ;
  assign n15224 = n6889 | n15223 ;
  assign n38584 = ~n15224 ;
  assign n15241 = n38584 & n15238 ;
  assign n15242 = n15018 | n15241 ;
  assign n38585 = ~n15240 ;
  assign n15243 = n38585 & n15242 ;
  assign n38586 = ~n15243 ;
  assign n15244 = n6600 & n38586 ;
  assign n14458 = n14294 & n38244 ;
  assign n38587 = ~n14473 ;
  assign n14485 = n14458 & n38587 ;
  assign n14950 = n14485 & n149 ;
  assign n14486 = n14456 | n14473 ;
  assign n38588 = ~n14486 ;
  assign n15012 = n38588 & n149 ;
  assign n15013 = n14294 | n15012 ;
  assign n38589 = ~n14950 ;
  assign n15014 = n38589 & n15013 ;
  assign n15252 = n38568 & n15233 ;
  assign n15253 = n15035 | n15252 ;
  assign n38590 = ~n15235 ;
  assign n15254 = n38590 & n15253 ;
  assign n38591 = ~n15254 ;
  assign n15255 = n162 & n38591 ;
  assign n15256 = n38578 & n15253 ;
  assign n15257 = n15040 | n15256 ;
  assign n38592 = ~n15255 ;
  assign n15258 = n38592 & n15257 ;
  assign n38593 = ~n15258 ;
  assign n15259 = n6889 & n38593 ;
  assign n15260 = n6600 | n15259 ;
  assign n38594 = ~n15260 ;
  assign n15261 = n15242 & n38594 ;
  assign n15262 = n15014 | n15261 ;
  assign n38595 = ~n15244 ;
  assign n15263 = n38595 & n15262 ;
  assign n38596 = ~n15263 ;
  assign n15264 = n165 & n38596 ;
  assign n38597 = ~n14477 ;
  assign n14483 = n14288 & n38597 ;
  assign n14484 = n38250 & n14483 ;
  assign n14928 = n14484 & n149 ;
  assign n14511 = n14477 | n14495 ;
  assign n38598 = ~n14511 ;
  assign n14962 = n38598 & n149 ;
  assign n14963 = n14288 | n14962 ;
  assign n38599 = ~n14928 ;
  assign n14964 = n38599 & n14963 ;
  assign n15245 = n165 | n15244 ;
  assign n38600 = ~n15245 ;
  assign n15265 = n38600 & n15262 ;
  assign n15266 = n14964 | n15265 ;
  assign n38601 = ~n15264 ;
  assign n15267 = n38601 & n15266 ;
  assign n38602 = ~n15267 ;
  assign n15268 = n166 & n38602 ;
  assign n14510 = n14480 | n14497 ;
  assign n38603 = ~n14510 ;
  assign n14958 = n38603 & n149 ;
  assign n14959 = n14300 | n14958 ;
  assign n14482 = n14300 & n38260 ;
  assign n38604 = ~n14497 ;
  assign n14509 = n14482 & n38604 ;
  assign n14993 = n14509 & n149 ;
  assign n38605 = ~n14993 ;
  assign n14994 = n14959 & n38605 ;
  assign n15276 = n38584 & n15257 ;
  assign n15277 = n15018 | n15276 ;
  assign n38606 = ~n15259 ;
  assign n15278 = n38606 & n15277 ;
  assign n38607 = ~n15278 ;
  assign n15279 = n164 & n38607 ;
  assign n15280 = n38594 & n15277 ;
  assign n15281 = n15014 | n15280 ;
  assign n38608 = ~n15279 ;
  assign n15282 = n38608 & n15281 ;
  assign n38609 = ~n15282 ;
  assign n15283 = n165 & n38609 ;
  assign n15284 = n166 | n15283 ;
  assign n38610 = ~n15284 ;
  assign n15285 = n15266 & n38610 ;
  assign n15286 = n14994 | n15285 ;
  assign n38611 = ~n15268 ;
  assign n15287 = n38611 & n15286 ;
  assign n38612 = ~n15287 ;
  assign n15288 = n167 & n38612 ;
  assign n38613 = ~n14501 ;
  assign n14507 = n14303 & n38613 ;
  assign n14508 = n38266 & n14507 ;
  assign n14954 = n14508 & n149 ;
  assign n14535 = n14501 | n14519 ;
  assign n38614 = ~n14535 ;
  assign n14955 = n38614 & n149 ;
  assign n14956 = n14303 | n14955 ;
  assign n38615 = ~n14954 ;
  assign n14957 = n38615 & n14956 ;
  assign n15269 = n5352 | n15268 ;
  assign n38616 = ~n15269 ;
  assign n15289 = n38616 & n15286 ;
  assign n15290 = n14957 | n15289 ;
  assign n38617 = ~n15288 ;
  assign n15291 = n38617 & n15290 ;
  assign n38618 = ~n15291 ;
  assign n15292 = n4934 & n38618 ;
  assign n14506 = n14296 & n38276 ;
  assign n38619 = ~n14521 ;
  assign n14533 = n14506 & n38619 ;
  assign n14944 = n14533 & n149 ;
  assign n14534 = n14504 | n14521 ;
  assign n38620 = ~n14534 ;
  assign n14947 = n38620 & n149 ;
  assign n14948 = n14296 | n14947 ;
  assign n38621 = ~n14944 ;
  assign n14949 = n38621 & n14948 ;
  assign n15300 = n38600 & n15281 ;
  assign n15301 = n14964 | n15300 ;
  assign n38622 = ~n15283 ;
  assign n15302 = n38622 & n15301 ;
  assign n38623 = ~n15302 ;
  assign n15303 = n166 & n38623 ;
  assign n15304 = n38610 & n15301 ;
  assign n15305 = n14994 | n15304 ;
  assign n38624 = ~n15303 ;
  assign n15306 = n38624 & n15305 ;
  assign n38625 = ~n15306 ;
  assign n15307 = n5352 & n38625 ;
  assign n15308 = n4934 | n15307 ;
  assign n38626 = ~n15308 ;
  assign n15309 = n15290 & n38626 ;
  assign n15310 = n14949 | n15309 ;
  assign n38627 = ~n15292 ;
  assign n15311 = n38627 & n15310 ;
  assign n38628 = ~n15311 ;
  assign n15312 = n169 & n38628 ;
  assign n14559 = n14525 | n14543 ;
  assign n38629 = ~n14559 ;
  assign n14922 = n38629 & n149 ;
  assign n14923 = n14262 | n14922 ;
  assign n38630 = ~n14525 ;
  assign n14531 = n14262 & n38630 ;
  assign n14532 = n38282 & n14531 ;
  assign n14951 = n14532 & n149 ;
  assign n38631 = ~n14951 ;
  assign n14952 = n14923 & n38631 ;
  assign n15293 = n169 | n15292 ;
  assign n38632 = ~n15293 ;
  assign n15313 = n38632 & n15310 ;
  assign n15314 = n14952 | n15313 ;
  assign n38633 = ~n15312 ;
  assign n15315 = n38633 & n15314 ;
  assign n38634 = ~n15315 ;
  assign n15316 = n170 & n38634 ;
  assign n14530 = n14274 & n38292 ;
  assign n38635 = ~n14545 ;
  assign n14557 = n14530 & n38635 ;
  assign n14943 = n14557 & n149 ;
  assign n14558 = n14528 | n14545 ;
  assign n38636 = ~n14558 ;
  assign n14966 = n38636 & n149 ;
  assign n14967 = n14274 | n14966 ;
  assign n38637 = ~n14943 ;
  assign n14968 = n38637 & n14967 ;
  assign n15324 = n38616 & n15305 ;
  assign n15325 = n14957 | n15324 ;
  assign n38638 = ~n15307 ;
  assign n15326 = n38638 & n15325 ;
  assign n38639 = ~n15326 ;
  assign n15327 = n168 & n38639 ;
  assign n15328 = n38626 & n15325 ;
  assign n15329 = n14949 | n15328 ;
  assign n38640 = ~n15327 ;
  assign n15330 = n38640 & n15329 ;
  assign n38641 = ~n15330 ;
  assign n15331 = n169 & n38641 ;
  assign n15332 = n170 | n15331 ;
  assign n38642 = ~n15332 ;
  assign n15333 = n15314 & n38642 ;
  assign n15334 = n14968 | n15333 ;
  assign n38643 = ~n15316 ;
  assign n15335 = n38643 & n15334 ;
  assign n38644 = ~n15335 ;
  assign n15336 = n171 & n38644 ;
  assign n14583 = n14549 | n14567 ;
  assign n38645 = ~n14583 ;
  assign n14941 = n38645 & n149 ;
  assign n14942 = n14283 | n14941 ;
  assign n38646 = ~n14549 ;
  assign n14555 = n14283 & n38646 ;
  assign n14556 = n38298 & n14555 ;
  assign n14960 = n14556 & n149 ;
  assign n38647 = ~n14960 ;
  assign n14961 = n14942 & n38647 ;
  assign n15317 = n3940 | n15316 ;
  assign n38648 = ~n15317 ;
  assign n15337 = n38648 & n15334 ;
  assign n15338 = n14961 | n15337 ;
  assign n38649 = ~n15336 ;
  assign n15339 = n38649 & n15338 ;
  assign n38650 = ~n15339 ;
  assign n15340 = n3631 & n38650 ;
  assign n14554 = n14248 & n38308 ;
  assign n38651 = ~n14569 ;
  assign n14581 = n14554 & n38651 ;
  assign n14937 = n14581 & n149 ;
  assign n14582 = n14552 | n14569 ;
  assign n38652 = ~n14582 ;
  assign n14938 = n38652 & n149 ;
  assign n14939 = n14248 | n14938 ;
  assign n38653 = ~n14937 ;
  assign n14940 = n38653 & n14939 ;
  assign n15348 = n38632 & n15329 ;
  assign n15349 = n14952 | n15348 ;
  assign n38654 = ~n15331 ;
  assign n15350 = n38654 & n15349 ;
  assign n38655 = ~n15350 ;
  assign n15351 = n170 & n38655 ;
  assign n15352 = n38642 & n15349 ;
  assign n15353 = n14968 | n15352 ;
  assign n38656 = ~n15351 ;
  assign n15354 = n38656 & n15353 ;
  assign n38657 = ~n15354 ;
  assign n15355 = n3940 & n38657 ;
  assign n15356 = n3631 | n15355 ;
  assign n38658 = ~n15356 ;
  assign n15357 = n15338 & n38658 ;
  assign n15358 = n14940 | n15357 ;
  assign n38659 = ~n15340 ;
  assign n15359 = n38659 & n15358 ;
  assign n38660 = ~n15359 ;
  assign n15360 = n173 & n38660 ;
  assign n38661 = ~n14573 ;
  assign n14579 = n14281 & n38661 ;
  assign n14580 = n38314 & n14579 ;
  assign n14936 = n14580 & n149 ;
  assign n14607 = n14573 | n14591 ;
  assign n38662 = ~n14607 ;
  assign n15019 = n38662 & n149 ;
  assign n15020 = n14281 | n15019 ;
  assign n38663 = ~n14936 ;
  assign n15021 = n38663 & n15020 ;
  assign n15341 = n173 | n15340 ;
  assign n38664 = ~n15341 ;
  assign n15361 = n38664 & n15358 ;
  assign n15362 = n15021 | n15361 ;
  assign n38665 = ~n15360 ;
  assign n15363 = n38665 & n15362 ;
  assign n38666 = ~n15363 ;
  assign n15364 = n174 & n38666 ;
  assign n14606 = n14576 | n14593 ;
  assign n38667 = ~n14606 ;
  assign n14934 = n38667 & n149 ;
  assign n14935 = n14269 | n14934 ;
  assign n14578 = n14269 & n38324 ;
  assign n38668 = ~n14593 ;
  assign n14605 = n14578 & n38668 ;
  assign n15005 = n14605 & n149 ;
  assign n38669 = ~n15005 ;
  assign n15006 = n14935 & n38669 ;
  assign n15372 = n38648 & n15353 ;
  assign n15373 = n14961 | n15372 ;
  assign n38670 = ~n15355 ;
  assign n15374 = n38670 & n15373 ;
  assign n38671 = ~n15374 ;
  assign n15375 = n172 & n38671 ;
  assign n15376 = n38658 & n15373 ;
  assign n15377 = n14940 | n15376 ;
  assign n38672 = ~n15375 ;
  assign n15378 = n38672 & n15377 ;
  assign n38673 = ~n15378 ;
  assign n15379 = n173 & n38673 ;
  assign n15380 = n174 | n15379 ;
  assign n38674 = ~n15380 ;
  assign n15381 = n15362 & n38674 ;
  assign n15382 = n15006 | n15381 ;
  assign n38675 = ~n15364 ;
  assign n15383 = n38675 & n15382 ;
  assign n38676 = ~n15383 ;
  assign n15384 = n175 & n38676 ;
  assign n38677 = ~n14597 ;
  assign n14603 = n14253 & n38677 ;
  assign n14604 = n38330 & n14603 ;
  assign n14991 = n14604 & n149 ;
  assign n14631 = n14597 | n14615 ;
  assign n38678 = ~n14631 ;
  assign n15007 = n38678 & n149 ;
  assign n15008 = n14253 | n15007 ;
  assign n38679 = ~n14991 ;
  assign n15009 = n38679 & n15008 ;
  assign n15365 = n2753 | n15364 ;
  assign n38680 = ~n15365 ;
  assign n15385 = n38680 & n15382 ;
  assign n15386 = n15009 | n15385 ;
  assign n38681 = ~n15384 ;
  assign n15387 = n38681 & n15386 ;
  assign n38682 = ~n15387 ;
  assign n15388 = n2431 & n38682 ;
  assign n14630 = n14600 | n14617 ;
  assign n38683 = ~n14630 ;
  assign n14919 = n38683 & n149 ;
  assign n14920 = n14216 | n14919 ;
  assign n14602 = n14216 & n38340 ;
  assign n38684 = ~n14617 ;
  assign n14629 = n14602 & n38684 ;
  assign n14926 = n14629 & n149 ;
  assign n38685 = ~n14926 ;
  assign n14927 = n14920 & n38685 ;
  assign n15396 = n38664 & n15377 ;
  assign n15397 = n15021 | n15396 ;
  assign n38686 = ~n15379 ;
  assign n15398 = n38686 & n15397 ;
  assign n38687 = ~n15398 ;
  assign n15399 = n174 & n38687 ;
  assign n15400 = n38674 & n15397 ;
  assign n15401 = n15006 | n15400 ;
  assign n38688 = ~n15399 ;
  assign n15402 = n38688 & n15401 ;
  assign n38689 = ~n15402 ;
  assign n15403 = n2753 & n38689 ;
  assign n15404 = n2431 | n15403 ;
  assign n38690 = ~n15404 ;
  assign n15405 = n15386 & n38690 ;
  assign n15406 = n14927 | n15405 ;
  assign n38691 = ~n15388 ;
  assign n15407 = n38691 & n15406 ;
  assign n38692 = ~n15407 ;
  assign n15408 = n177 & n38692 ;
  assign n14648 = n14621 | n14639 ;
  assign n38693 = ~n14648 ;
  assign n14932 = n38693 & n149 ;
  assign n14933 = n14246 | n14932 ;
  assign n38694 = ~n14621 ;
  assign n14627 = n14246 & n38694 ;
  assign n14628 = n38346 & n14627 ;
  assign n14989 = n14628 & n149 ;
  assign n38695 = ~n14989 ;
  assign n14990 = n14933 & n38695 ;
  assign n15390 = n177 | n15388 ;
  assign n38696 = ~n15390 ;
  assign n15409 = n38696 & n15406 ;
  assign n15410 = n14990 | n15409 ;
  assign n38697 = ~n15408 ;
  assign n15411 = n38697 & n15410 ;
  assign n38698 = ~n15411 ;
  assign n15412 = n178 & n38698 ;
  assign n14647 = n14624 | n14641 ;
  assign n38699 = ~n14647 ;
  assign n14930 = n38699 & n149 ;
  assign n14931 = n14258 | n14930 ;
  assign n14626 = n14258 & n38356 ;
  assign n38700 = ~n14641 ;
  assign n14646 = n14626 & n38700 ;
  assign n14998 = n14646 & n149 ;
  assign n38701 = ~n14998 ;
  assign n14999 = n14931 & n38701 ;
  assign n15420 = n38680 & n15401 ;
  assign n15421 = n15009 | n15420 ;
  assign n38702 = ~n15403 ;
  assign n15422 = n38702 & n15421 ;
  assign n38703 = ~n15422 ;
  assign n15423 = n176 & n38703 ;
  assign n15424 = n38690 & n15421 ;
  assign n15425 = n14927 | n15424 ;
  assign n38704 = ~n15423 ;
  assign n15426 = n38704 & n15425 ;
  assign n38705 = ~n15426 ;
  assign n15427 = n177 & n38705 ;
  assign n15428 = n178 | n15427 ;
  assign n38706 = ~n15428 ;
  assign n15429 = n15410 & n38706 ;
  assign n15430 = n14999 | n15429 ;
  assign n38707 = ~n15412 ;
  assign n15431 = n38707 & n15430 ;
  assign n38708 = ~n15431 ;
  assign n15432 = n179 & n38708 ;
  assign n15413 = n1707 | n15412 ;
  assign n38709 = ~n15413 ;
  assign n15433 = n38709 & n15430 ;
  assign n38710 = ~n14645 ;
  assign n15465 = n38710 & n14759 ;
  assign n15466 = n38362 & n15465 ;
  assign n15467 = n149 & n15466 ;
  assign n14658 = n14645 | n14656 ;
  assign n38711 = ~n14658 ;
  assign n14921 = n38711 & n149 ;
  assign n15468 = n14759 | n14921 ;
  assign n38712 = ~n15467 ;
  assign n15469 = n38712 & n15468 ;
  assign n15470 = n15433 | n15469 ;
  assign n38713 = ~n15432 ;
  assign n15471 = n38713 & n15470 ;
  assign n38714 = ~n15471 ;
  assign n15472 = n1487 & n38714 ;
  assign n14778 = n14762 | n14765 ;
  assign n38715 = ~n14778 ;
  assign n14985 = n38715 & n149 ;
  assign n14986 = n14757 | n14985 ;
  assign n14764 = n14757 & n38372 ;
  assign n38716 = ~n14765 ;
  assign n14777 = n14764 & n38716 ;
  assign n15041 = n14777 & n149 ;
  assign n38717 = ~n15041 ;
  assign n15042 = n14986 & n38717 ;
  assign n15436 = n38696 & n15425 ;
  assign n15437 = n14990 | n15436 ;
  assign n38718 = ~n15427 ;
  assign n15438 = n38718 & n15437 ;
  assign n38719 = ~n15438 ;
  assign n15439 = n178 & n38719 ;
  assign n15440 = n38706 & n15437 ;
  assign n15441 = n14999 | n15440 ;
  assign n38720 = ~n15439 ;
  assign n15442 = n38720 & n15441 ;
  assign n38721 = ~n15442 ;
  assign n15443 = n1707 & n38721 ;
  assign n15444 = n1487 | n15443 ;
  assign n38722 = ~n15444 ;
  assign n15475 = n38722 & n15470 ;
  assign n15476 = n15042 | n15475 ;
  assign n38723 = ~n15472 ;
  assign n15477 = n38723 & n15476 ;
  assign n38724 = ~n15477 ;
  assign n15478 = n181 & n38724 ;
  assign n14801 = n14769 | n14785 ;
  assign n38725 = ~n14801 ;
  assign n15043 = n38725 & n149 ;
  assign n15044 = n14751 | n15043 ;
  assign n38726 = ~n14769 ;
  assign n14775 = n14751 & n38726 ;
  assign n14776 = n38378 & n14775 ;
  assign n15047 = n14776 & n149 ;
  assign n38727 = ~n15047 ;
  assign n15048 = n15044 & n38727 ;
  assign n15473 = n181 | n15472 ;
  assign n38728 = ~n15473 ;
  assign n15479 = n38728 & n15476 ;
  assign n15480 = n15048 | n15479 ;
  assign n38729 = ~n15478 ;
  assign n15481 = n38729 & n15480 ;
  assign n38730 = ~n15481 ;
  assign n15482 = n182 & n38730 ;
  assign n14800 = n14772 | n14787 ;
  assign n38731 = ~n14800 ;
  assign n15045 = n38731 & n149 ;
  assign n15046 = n14744 | n15045 ;
  assign n14774 = n14744 & n38388 ;
  assign n38732 = ~n14787 ;
  assign n14799 = n14774 & n38732 ;
  assign n15049 = n14799 & n149 ;
  assign n38733 = ~n15049 ;
  assign n15050 = n15046 & n38733 ;
  assign n15446 = n38709 & n15441 ;
  assign n15492 = n15446 | n15469 ;
  assign n38734 = ~n15443 ;
  assign n15493 = n38734 & n15492 ;
  assign n38735 = ~n15493 ;
  assign n15494 = n180 & n38735 ;
  assign n15495 = n38722 & n15492 ;
  assign n15496 = n15042 | n15495 ;
  assign n38736 = ~n15494 ;
  assign n15497 = n38736 & n15496 ;
  assign n38737 = ~n15497 ;
  assign n15498 = n181 & n38737 ;
  assign n15499 = n182 | n15498 ;
  assign n38738 = ~n15499 ;
  assign n15500 = n15480 & n38738 ;
  assign n15501 = n15050 | n15500 ;
  assign n38739 = ~n15482 ;
  assign n15502 = n38739 & n15501 ;
  assign n38740 = ~n15502 ;
  assign n15503 = n183 & n38740 ;
  assign n14825 = n14791 | n14809 ;
  assign n38741 = ~n14825 ;
  assign n15051 = n38741 & n149 ;
  assign n15052 = n14738 | n15051 ;
  assign n38742 = ~n14791 ;
  assign n14797 = n14738 & n38742 ;
  assign n14798 = n38394 & n14797 ;
  assign n15053 = n14798 & n149 ;
  assign n38743 = ~n15053 ;
  assign n15054 = n15052 & n38743 ;
  assign n15483 = n183 | n15482 ;
  assign n38744 = ~n15483 ;
  assign n15504 = n38744 & n15501 ;
  assign n15508 = n15054 | n15504 ;
  assign n38745 = ~n15503 ;
  assign n15509 = n38745 & n15508 ;
  assign n38746 = ~n15509 ;
  assign n15510 = n838 & n38746 ;
  assign n14796 = n14731 & n38404 ;
  assign n38747 = ~n14811 ;
  assign n14824 = n14796 & n38747 ;
  assign n15000 = n14824 & n149 ;
  assign n14823 = n14794 | n14811 ;
  assign n38748 = ~n14823 ;
  assign n15055 = n38748 & n149 ;
  assign n15056 = n14731 | n15055 ;
  assign n38749 = ~n15000 ;
  assign n15057 = n38749 & n15056 ;
  assign n15515 = n38728 & n15496 ;
  assign n15516 = n15048 | n15515 ;
  assign n38750 = ~n15498 ;
  assign n15517 = n38750 & n15516 ;
  assign n38751 = ~n15517 ;
  assign n15518 = n182 & n38751 ;
  assign n15519 = n38738 & n15516 ;
  assign n15520 = n15050 | n15519 ;
  assign n38752 = ~n15518 ;
  assign n15521 = n38752 & n15520 ;
  assign n38753 = ~n15521 ;
  assign n15522 = n996 & n38753 ;
  assign n15523 = n838 | n15522 ;
  assign n38754 = ~n15523 ;
  assign n15524 = n15508 & n38754 ;
  assign n15525 = n15057 | n15524 ;
  assign n38755 = ~n15510 ;
  assign n15526 = n38755 & n15525 ;
  assign n38756 = ~n15526 ;
  assign n15527 = n185 & n38756 ;
  assign n14849 = n14815 | n14833 ;
  assign n38757 = ~n14849 ;
  assign n15058 = n38757 & n149 ;
  assign n15059 = n14725 | n15058 ;
  assign n38758 = ~n14815 ;
  assign n14821 = n14725 & n38758 ;
  assign n14822 = n38410 & n14821 ;
  assign n15060 = n14822 & n149 ;
  assign n38759 = ~n15060 ;
  assign n15061 = n15059 & n38759 ;
  assign n15511 = n185 | n15510 ;
  assign n38760 = ~n15511 ;
  assign n15528 = n38760 & n15525 ;
  assign n15529 = n15061 | n15528 ;
  assign n38761 = ~n15527 ;
  assign n15530 = n38761 & n15529 ;
  assign n38762 = ~n15530 ;
  assign n15531 = n186 & n38762 ;
  assign n14848 = n14818 | n14835 ;
  assign n38763 = ~n14848 ;
  assign n15062 = n38763 & n149 ;
  assign n15063 = n14718 | n15062 ;
  assign n14820 = n14718 & n38420 ;
  assign n38764 = ~n14835 ;
  assign n14847 = n14820 & n38764 ;
  assign n15064 = n14847 & n149 ;
  assign n38765 = ~n15064 ;
  assign n15065 = n15063 & n38765 ;
  assign n15539 = n38744 & n15520 ;
  assign n15540 = n15054 | n15539 ;
  assign n38766 = ~n15522 ;
  assign n15541 = n38766 & n15540 ;
  assign n38767 = ~n15541 ;
  assign n15542 = n184 & n38767 ;
  assign n15543 = n38754 & n15540 ;
  assign n15544 = n15057 | n15543 ;
  assign n38768 = ~n15542 ;
  assign n15545 = n38768 & n15544 ;
  assign n38769 = ~n15545 ;
  assign n15546 = n185 & n38769 ;
  assign n15547 = n186 | n15546 ;
  assign n38770 = ~n15547 ;
  assign n15548 = n15529 & n38770 ;
  assign n15549 = n15065 | n15548 ;
  assign n38771 = ~n15531 ;
  assign n15550 = n38771 & n15549 ;
  assign n38772 = ~n15550 ;
  assign n15551 = n187 & n38772 ;
  assign n14873 = n14839 | n14857 ;
  assign n38773 = ~n14873 ;
  assign n15001 = n38773 & n149 ;
  assign n15002 = n14712 | n15001 ;
  assign n38774 = ~n14839 ;
  assign n14845 = n14712 & n38774 ;
  assign n14846 = n38426 & n14845 ;
  assign n15066 = n14846 & n149 ;
  assign n38775 = ~n15066 ;
  assign n15067 = n15002 & n38775 ;
  assign n15532 = n528 | n15531 ;
  assign n38776 = ~n15532 ;
  assign n15552 = n38776 & n15549 ;
  assign n15553 = n15067 | n15552 ;
  assign n38777 = ~n15551 ;
  assign n15554 = n38777 & n15553 ;
  assign n38778 = ~n15554 ;
  assign n15555 = n413 & n38778 ;
  assign n14872 = n14842 | n14859 ;
  assign n38779 = ~n14872 ;
  assign n15068 = n38779 & n149 ;
  assign n15069 = n14306 | n15068 ;
  assign n14844 = n14306 & n38436 ;
  assign n38780 = ~n14859 ;
  assign n14871 = n14844 & n38780 ;
  assign n15070 = n14871 & n149 ;
  assign n38781 = ~n15070 ;
  assign n15071 = n15069 & n38781 ;
  assign n15563 = n38760 & n15544 ;
  assign n15564 = n15061 | n15563 ;
  assign n38782 = ~n15546 ;
  assign n15565 = n38782 & n15564 ;
  assign n38783 = ~n15565 ;
  assign n15566 = n186 & n38783 ;
  assign n15567 = n38770 & n15564 ;
  assign n15568 = n15065 | n15567 ;
  assign n38784 = ~n15566 ;
  assign n15569 = n38784 & n15568 ;
  assign n38785 = ~n15569 ;
  assign n15570 = n528 & n38785 ;
  assign n15571 = n413 | n15570 ;
  assign n38786 = ~n15571 ;
  assign n15572 = n15553 & n38786 ;
  assign n15573 = n15071 | n15572 ;
  assign n38787 = ~n15555 ;
  assign n15574 = n38787 & n15573 ;
  assign n38788 = ~n15574 ;
  assign n15575 = n189 & n38788 ;
  assign n14897 = n14863 | n14881 ;
  assign n38789 = ~n14897 ;
  assign n15031 = n38789 & n149 ;
  assign n15032 = n14705 | n15031 ;
  assign n38790 = ~n14863 ;
  assign n14869 = n14705 & n38790 ;
  assign n14870 = n38442 & n14869 ;
  assign n15072 = n14870 & n149 ;
  assign n38791 = ~n15072 ;
  assign n15073 = n15032 & n38791 ;
  assign n15556 = n189 | n15555 ;
  assign n38792 = ~n15556 ;
  assign n15576 = n38792 & n15573 ;
  assign n15577 = n15073 | n15576 ;
  assign n38793 = ~n15575 ;
  assign n15578 = n38793 & n15577 ;
  assign n38794 = ~n15578 ;
  assign n15579 = n190 & n38794 ;
  assign n14896 = n14866 | n14883 ;
  assign n38795 = ~n14896 ;
  assign n15074 = n38795 & n149 ;
  assign n15075 = n14698 | n15074 ;
  assign n14868 = n14698 & n38452 ;
  assign n38796 = ~n14883 ;
  assign n14895 = n14868 & n38796 ;
  assign n15076 = n14895 & n149 ;
  assign n38797 = ~n15076 ;
  assign n15077 = n15075 & n38797 ;
  assign n15585 = n38776 & n15568 ;
  assign n15586 = n15067 | n15585 ;
  assign n38798 = ~n15570 ;
  assign n15587 = n38798 & n15586 ;
  assign n38799 = ~n15587 ;
  assign n15588 = n188 & n38799 ;
  assign n15589 = n38786 & n15586 ;
  assign n15590 = n15071 | n15589 ;
  assign n38800 = ~n15588 ;
  assign n15591 = n38800 & n15590 ;
  assign n38801 = ~n15591 ;
  assign n15592 = n189 & n38801 ;
  assign n15593 = n190 | n15592 ;
  assign n38802 = ~n15593 ;
  assign n15594 = n15577 & n38802 ;
  assign n15595 = n15077 | n15594 ;
  assign n38803 = ~n15579 ;
  assign n15600 = n38803 & n15595 ;
  assign n38804 = ~n15600 ;
  assign n15601 = n191 & n38804 ;
  assign n38805 = ~n14887 ;
  assign n14893 = n14692 & n38805 ;
  assign n14894 = n38458 & n14893 ;
  assign n14995 = n14894 & n149 ;
  assign n15461 = n14887 | n14905 ;
  assign n38806 = ~n15461 ;
  assign n15462 = n149 & n38806 ;
  assign n15463 = n14692 | n15462 ;
  assign n38807 = ~n14995 ;
  assign n15464 = n38807 & n15463 ;
  assign n15580 = n191 | n15579 ;
  assign n38808 = ~n15580 ;
  assign n15611 = n38808 & n15595 ;
  assign n15612 = n15464 | n15611 ;
  assign n38809 = ~n15601 ;
  assign n15613 = n38809 & n15612 ;
  assign n15614 = n15448 | n15613 ;
  assign n15615 = n31336 & n15614 ;
  assign n14913 = n192 & n14912 ;
  assign n38810 = ~n14676 ;
  assign n15089 = n38810 & n149 ;
  assign n38811 = ~n15089 ;
  assign n15090 = n14911 & n38811 ;
  assign n38812 = ~n15090 ;
  assign n15091 = n14913 & n38812 ;
  assign n14672 = n14662 | n14671 ;
  assign n38813 = ~n14672 ;
  assign n14678 = n38813 & n14675 ;
  assign n14679 = n38489 & n14678 ;
  assign n15449 = n14679 & n38490 ;
  assign n15450 = n38491 & n15449 ;
  assign n15451 = n15091 | n15450 ;
  assign n15602 = n15079 & n38809 ;
  assign n15621 = n15602 & n15612 ;
  assign n15622 = n15451 | n15621 ;
  assign n148 = n15615 | n15622 ;
  assign n15581 = n287 | n15579 ;
  assign n38814 = ~n15581 ;
  assign n15596 = n38814 & n15595 ;
  assign n15597 = n15464 | n15596 ;
  assign n15603 = n15597 & n15602 ;
  assign n15608 = n15597 & n38809 ;
  assign n15609 = n15079 | n15608 ;
  assign n38815 = ~n15609 ;
  assign n15643 = n38815 & n148 ;
  assign n15644 = n15603 | n15643 ;
  assign n38816 = ~n15611 ;
  assign n16179 = n15464 & n38816 ;
  assign n16180 = n38809 & n16179 ;
  assign n16181 = n148 & n16180 ;
  assign n16183 = n15601 | n15611 ;
  assign n38817 = ~n16183 ;
  assign n16184 = n148 & n38817 ;
  assign n16185 = n15464 | n16184 ;
  assign n38818 = ~n16181 ;
  assign n16186 = n38818 & n16185 ;
  assign n16187 = n15644 | n16186 ;
  assign n215 = x36 | x37 ;
  assign n216 = x38 | n215 ;
  assign n15681 = x38 & n148 ;
  assign n38819 = ~n15681 ;
  assign n15688 = n216 & n38819 ;
  assign n38820 = ~n15688 ;
  assign n15689 = n149 & n38820 ;
  assign n15690 = n150 | n15689 ;
  assign n14666 = n216 & n38488 ;
  assign n14667 = n38489 & n14666 ;
  assign n15459 = n14667 & n38490 ;
  assign n15460 = n38491 & n15459 ;
  assign n15682 = n15460 & n38819 ;
  assign n38821 = ~n212 ;
  assign n15692 = n38821 & n148 ;
  assign n38822 = ~x38 ;
  assign n15705 = n38822 & n148 ;
  assign n38823 = ~n15705 ;
  assign n15706 = x39 & n38823 ;
  assign n15720 = n15692 | n15706 ;
  assign n15721 = n15682 | n15720 ;
  assign n38824 = ~n15690 ;
  assign n15722 = n38824 & n15721 ;
  assign n38825 = ~n15450 ;
  assign n15455 = n149 & n38825 ;
  assign n38826 = ~n15091 ;
  assign n15456 = n38826 & n15455 ;
  assign n38827 = ~n15603 ;
  assign n15605 = n15456 & n38827 ;
  assign n38828 = ~n15615 ;
  assign n15616 = n15605 & n38828 ;
  assign n15617 = x40 | n15616 ;
  assign n15693 = n15617 | n15692 ;
  assign n15723 = n15616 | n15692 ;
  assign n15724 = x40 & n15723 ;
  assign n38829 = ~n15724 ;
  assign n15725 = n15693 & n38829 ;
  assign n15726 = n15722 | n15725 ;
  assign n217 = n38822 & n215 ;
  assign n15604 = n15451 | n15603 ;
  assign n15805 = n15448 | n15608 ;
  assign n15806 = n31336 & n15805 ;
  assign n15807 = n15604 | n15806 ;
  assign n38830 = ~n15807 ;
  assign n15818 = x38 & n38830 ;
  assign n15819 = n217 | n15818 ;
  assign n38831 = ~n15819 ;
  assign n15820 = n149 & n38831 ;
  assign n38832 = ~n15820 ;
  assign n15821 = n15721 & n38832 ;
  assign n38833 = ~n15821 ;
  assign n15822 = n150 & n38833 ;
  assign n38834 = ~n15822 ;
  assign n15823 = n15726 & n38834 ;
  assign n38835 = ~n15823 ;
  assign n15828 = n151 & n38835 ;
  assign n15025 = n15004 | n15023 ;
  assign n38836 = ~n15025 ;
  assign n15647 = n38836 & n148 ;
  assign n15648 = n15094 | n15647 ;
  assign n15095 = n38836 & n15094 ;
  assign n15715 = n15095 & n148 ;
  assign n38837 = ~n15715 ;
  assign n15716 = n15648 & n38837 ;
  assign n15845 = n151 | n15822 ;
  assign n38838 = ~n15845 ;
  assign n15846 = n15726 & n38838 ;
  assign n15847 = n15716 | n15846 ;
  assign n38839 = ~n15828 ;
  assign n15848 = n38839 & n15847 ;
  assign n38840 = ~n15848 ;
  assign n15849 = n152 & n38840 ;
  assign n38841 = ~n15101 ;
  assign n15131 = n38841 & n15110 ;
  assign n15132 = n38493 & n15131 ;
  assign n15701 = n15132 & n148 ;
  assign n15102 = n15100 | n15101 ;
  assign n38842 = ~n15102 ;
  assign n15738 = n38842 & n148 ;
  assign n15739 = n15110 | n15738 ;
  assign n38843 = ~n15701 ;
  assign n15740 = n38843 & n15739 ;
  assign n15824 = n13662 & n38835 ;
  assign n15832 = n13079 | n15824 ;
  assign n38844 = ~n15832 ;
  assign n15850 = n38844 & n15847 ;
  assign n15851 = n15740 | n15850 ;
  assign n38845 = ~n15849 ;
  assign n15852 = n38845 & n15851 ;
  assign n38846 = ~n15852 ;
  assign n15853 = n153 & n38846 ;
  assign n15130 = n15113 | n15116 ;
  assign n38847 = ~n15130 ;
  assign n15653 = n38847 & n148 ;
  assign n15654 = n15038 | n15653 ;
  assign n15115 = n15038 & n38498 ;
  assign n38848 = ~n15116 ;
  assign n15129 = n15115 & n38848 ;
  assign n15694 = n15129 & n148 ;
  assign n38849 = ~n15694 ;
  assign n15695 = n15654 & n38849 ;
  assign n38850 = ~n15689 ;
  assign n15728 = n38850 & n15721 ;
  assign n38851 = ~n15728 ;
  assign n15729 = n150 & n38851 ;
  assign n15730 = n13662 | n15729 ;
  assign n38852 = ~n15730 ;
  assign n15731 = n15726 & n38852 ;
  assign n15732 = n15716 | n15731 ;
  assign n38853 = ~n15824 ;
  assign n15825 = n15732 & n38853 ;
  assign n38854 = ~n15825 ;
  assign n15826 = n13079 & n38854 ;
  assign n15827 = n153 | n15826 ;
  assign n38855 = ~n15827 ;
  assign n15871 = n38855 & n15851 ;
  assign n15872 = n15695 | n15871 ;
  assign n38856 = ~n15853 ;
  assign n15873 = n38856 & n15872 ;
  assign n38857 = ~n15873 ;
  assign n15874 = n154 & n38857 ;
  assign n38858 = ~n15120 ;
  assign n15126 = n15081 & n38858 ;
  assign n15127 = n38504 & n15126 ;
  assign n15656 = n15127 & n148 ;
  assign n15128 = n15119 | n15120 ;
  assign n38859 = ~n15128 ;
  assign n15696 = n38859 & n148 ;
  assign n15697 = n15081 | n15696 ;
  assign n38860 = ~n15656 ;
  assign n15698 = n38860 & n15697 ;
  assign n15854 = n154 | n15853 ;
  assign n38861 = ~n15854 ;
  assign n15875 = n38861 & n15872 ;
  assign n15876 = n15698 | n15875 ;
  assign n38862 = ~n15874 ;
  assign n15877 = n38862 & n15876 ;
  assign n38863 = ~n15877 ;
  assign n15878 = n11067 & n38863 ;
  assign n15125 = n15084 & n38515 ;
  assign n38864 = ~n15141 ;
  assign n15154 = n15125 & n38864 ;
  assign n15691 = n15154 & n148 ;
  assign n15155 = n15123 | n15141 ;
  assign n38865 = ~n15155 ;
  assign n15735 = n38865 & n148 ;
  assign n15736 = n15084 | n15735 ;
  assign n38866 = ~n15691 ;
  assign n15737 = n38866 & n15736 ;
  assign n15833 = n15732 & n38844 ;
  assign n15834 = n15740 | n15833 ;
  assign n38867 = ~n15826 ;
  assign n15835 = n38867 & n15834 ;
  assign n38868 = ~n15835 ;
  assign n15836 = n153 & n38868 ;
  assign n15837 = n38855 & n15834 ;
  assign n15838 = n15695 | n15837 ;
  assign n38869 = ~n15836 ;
  assign n15839 = n38869 & n15838 ;
  assign n38870 = ~n15839 ;
  assign n15840 = n154 & n38870 ;
  assign n15841 = n11067 | n15840 ;
  assign n38871 = ~n15841 ;
  assign n15895 = n38871 & n15876 ;
  assign n15896 = n15737 | n15895 ;
  assign n38872 = ~n15878 ;
  assign n15897 = n38872 & n15896 ;
  assign n38873 = ~n15897 ;
  assign n15898 = n156 & n38873 ;
  assign n15153 = n15144 | n15145 ;
  assign n38874 = ~n15153 ;
  assign n15628 = n38874 & n148 ;
  assign n15629 = n14980 | n15628 ;
  assign n38875 = ~n15145 ;
  assign n15151 = n14980 & n38875 ;
  assign n15152 = n38521 & n15151 ;
  assign n15816 = n15152 & n15807 ;
  assign n38876 = ~n15816 ;
  assign n15817 = n15629 & n38876 ;
  assign n15879 = n10657 | n15878 ;
  assign n38877 = ~n15879 ;
  assign n15899 = n38877 & n15896 ;
  assign n15900 = n15817 | n15899 ;
  assign n38878 = ~n15898 ;
  assign n15901 = n38878 & n15900 ;
  assign n38879 = ~n15901 ;
  assign n15902 = n157 & n38879 ;
  assign n15179 = n15148 | n15165 ;
  assign n38880 = ~n15179 ;
  assign n15747 = n38880 & n148 ;
  assign n15748 = n14975 | n15747 ;
  assign n15150 = n14975 & n38531 ;
  assign n38881 = ~n15165 ;
  assign n15178 = n15150 & n38881 ;
  assign n15757 = n15178 & n148 ;
  assign n38882 = ~n15757 ;
  assign n15758 = n15748 & n38882 ;
  assign n15855 = n15838 & n38861 ;
  assign n15856 = n15698 | n15855 ;
  assign n38883 = ~n15840 ;
  assign n15857 = n38883 & n15856 ;
  assign n38884 = ~n15857 ;
  assign n15858 = n155 & n38884 ;
  assign n15859 = n38871 & n15856 ;
  assign n15860 = n15737 | n15859 ;
  assign n38885 = ~n15858 ;
  assign n15861 = n38885 & n15860 ;
  assign n38886 = ~n15861 ;
  assign n15862 = n10657 & n38886 ;
  assign n15863 = n157 | n15862 ;
  assign n38887 = ~n15863 ;
  assign n15919 = n38887 & n15900 ;
  assign n15920 = n15758 | n15919 ;
  assign n38888 = ~n15902 ;
  assign n15921 = n38888 & n15920 ;
  assign n38889 = ~n15921 ;
  assign n15922 = n158 & n38889 ;
  assign n15177 = n15168 | n15169 ;
  assign n38890 = ~n15177 ;
  assign n15637 = n38890 & n148 ;
  assign n15638 = n14984 | n15637 ;
  assign n38891 = ~n15169 ;
  assign n15175 = n14984 & n38891 ;
  assign n15176 = n38537 & n15175 ;
  assign n15676 = n15176 & n148 ;
  assign n38892 = ~n15676 ;
  assign n15677 = n15638 & n38892 ;
  assign n15903 = n158 | n15902 ;
  assign n38893 = ~n15903 ;
  assign n15923 = n38893 & n15920 ;
  assign n15924 = n15677 | n15923 ;
  assign n38894 = ~n15922 ;
  assign n15925 = n38894 & n15924 ;
  assign n38895 = ~n15925 ;
  assign n15926 = n8857 & n38895 ;
  assign n15203 = n15172 | n15189 ;
  assign n38896 = ~n15203 ;
  assign n15745 = n38896 & n148 ;
  assign n15746 = n15016 | n15745 ;
  assign n15174 = n15016 & n38547 ;
  assign n38897 = ~n15189 ;
  assign n15202 = n15174 & n38897 ;
  assign n15755 = n15202 & n148 ;
  assign n38898 = ~n15755 ;
  assign n15756 = n15746 & n38898 ;
  assign n15880 = n15860 & n38877 ;
  assign n15881 = n15817 | n15880 ;
  assign n38899 = ~n15862 ;
  assign n15882 = n38899 & n15881 ;
  assign n38900 = ~n15882 ;
  assign n15883 = n157 & n38900 ;
  assign n15884 = n38887 & n15881 ;
  assign n15885 = n15758 | n15884 ;
  assign n38901 = ~n15883 ;
  assign n15886 = n38901 & n15885 ;
  assign n38902 = ~n15886 ;
  assign n15887 = n158 & n38902 ;
  assign n15888 = n8857 | n15887 ;
  assign n38903 = ~n15888 ;
  assign n15943 = n38903 & n15924 ;
  assign n15944 = n15756 | n15943 ;
  assign n38904 = ~n15926 ;
  assign n15945 = n38904 & n15944 ;
  assign n38905 = ~n15945 ;
  assign n15946 = n160 & n38905 ;
  assign n15201 = n15192 | n15193 ;
  assign n38906 = ~n15201 ;
  assign n15759 = n38906 & n148 ;
  assign n15760 = n15028 | n15759 ;
  assign n38907 = ~n15193 ;
  assign n15199 = n15028 & n38907 ;
  assign n15200 = n38553 & n15199 ;
  assign n15814 = n15200 & n15807 ;
  assign n38908 = ~n15814 ;
  assign n15815 = n15760 & n38908 ;
  assign n15927 = n160 | n15926 ;
  assign n38909 = ~n15927 ;
  assign n15947 = n38909 & n15944 ;
  assign n15948 = n15815 | n15947 ;
  assign n38910 = ~n15946 ;
  assign n15949 = n38910 & n15948 ;
  assign n38911 = ~n15949 ;
  assign n15950 = n161 & n38911 ;
  assign n15198 = n14972 & n38563 ;
  assign n38912 = ~n15213 ;
  assign n15227 = n15198 & n38912 ;
  assign n15651 = n15227 & n148 ;
  assign n15226 = n15196 | n15213 ;
  assign n38913 = ~n15226 ;
  assign n15752 = n38913 & n148 ;
  assign n15753 = n14972 | n15752 ;
  assign n38914 = ~n15651 ;
  assign n15754 = n38914 & n15753 ;
  assign n15904 = n15885 & n38893 ;
  assign n15905 = n15677 | n15904 ;
  assign n38915 = ~n15887 ;
  assign n15906 = n38915 & n15905 ;
  assign n38916 = ~n15906 ;
  assign n15907 = n159 & n38916 ;
  assign n15908 = n38903 & n15905 ;
  assign n15909 = n15756 | n15908 ;
  assign n38917 = ~n15907 ;
  assign n15910 = n38917 & n15909 ;
  assign n38918 = ~n15910 ;
  assign n15911 = n8534 & n38918 ;
  assign n15912 = n161 | n15911 ;
  assign n38919 = ~n15912 ;
  assign n15966 = n38919 & n15948 ;
  assign n15967 = n15754 | n15966 ;
  assign n38920 = ~n15950 ;
  assign n15968 = n38920 & n15967 ;
  assign n38921 = ~n15968 ;
  assign n15969 = n162 & n38921 ;
  assign n15220 = n15216 | n15217 ;
  assign n38922 = ~n15220 ;
  assign n15699 = n38922 & n148 ;
  assign n15700 = n15035 | n15699 ;
  assign n38923 = ~n15217 ;
  assign n15218 = n15035 & n38923 ;
  assign n15219 = n38569 & n15218 ;
  assign n15763 = n15219 & n148 ;
  assign n38924 = ~n15763 ;
  assign n15764 = n15700 & n38924 ;
  assign n15951 = n162 | n15950 ;
  assign n38925 = ~n15951 ;
  assign n15970 = n38925 & n15967 ;
  assign n15971 = n15764 | n15970 ;
  assign n38926 = ~n15969 ;
  assign n15972 = n38926 & n15971 ;
  assign n38927 = ~n15972 ;
  assign n15973 = n6889 & n38927 ;
  assign n15251 = n15223 | n15237 ;
  assign n38928 = ~n15251 ;
  assign n15632 = n38928 & n148 ;
  assign n15633 = n15040 | n15632 ;
  assign n15225 = n15040 & n38579 ;
  assign n38929 = ~n15237 ;
  assign n15250 = n15225 & n38929 ;
  assign n15761 = n15250 & n148 ;
  assign n38930 = ~n15761 ;
  assign n15762 = n15633 & n38930 ;
  assign n15928 = n15909 & n38909 ;
  assign n15929 = n15815 | n15928 ;
  assign n38931 = ~n15911 ;
  assign n15930 = n38931 & n15929 ;
  assign n38932 = ~n15930 ;
  assign n15931 = n161 & n38932 ;
  assign n15932 = n38919 & n15929 ;
  assign n15933 = n15754 | n15932 ;
  assign n38933 = ~n15931 ;
  assign n15934 = n38933 & n15933 ;
  assign n38934 = ~n15934 ;
  assign n15935 = n162 & n38934 ;
  assign n15936 = n6889 | n15935 ;
  assign n38935 = ~n15936 ;
  assign n15990 = n38935 & n15971 ;
  assign n15991 = n15762 | n15990 ;
  assign n38936 = ~n15973 ;
  assign n15992 = n38936 & n15991 ;
  assign n38937 = ~n15992 ;
  assign n15993 = n164 & n38937 ;
  assign n15249 = n15240 | n15241 ;
  assign n38938 = ~n15249 ;
  assign n15679 = n38938 & n148 ;
  assign n15680 = n15018 | n15679 ;
  assign n38939 = ~n15241 ;
  assign n15247 = n15018 & n38939 ;
  assign n15248 = n38585 & n15247 ;
  assign n15685 = n15248 & n148 ;
  assign n38940 = ~n15685 ;
  assign n15686 = n15680 & n38940 ;
  assign n15974 = n6600 | n15973 ;
  assign n38941 = ~n15974 ;
  assign n15994 = n38941 & n15991 ;
  assign n15995 = n15686 | n15994 ;
  assign n38942 = ~n15993 ;
  assign n15996 = n38942 & n15995 ;
  assign n38943 = ~n15996 ;
  assign n15997 = n165 & n38943 ;
  assign n15246 = n15014 & n38595 ;
  assign n38944 = ~n15261 ;
  assign n15274 = n15246 & n38944 ;
  assign n15678 = n15274 & n148 ;
  assign n15275 = n15244 | n15261 ;
  assign n38945 = ~n15275 ;
  assign n15712 = n38945 & n148 ;
  assign n15713 = n15014 | n15712 ;
  assign n38946 = ~n15678 ;
  assign n15714 = n38946 & n15713 ;
  assign n15952 = n15933 & n38925 ;
  assign n15953 = n15764 | n15952 ;
  assign n38947 = ~n15935 ;
  assign n15954 = n38947 & n15953 ;
  assign n38948 = ~n15954 ;
  assign n15955 = n163 & n38948 ;
  assign n15956 = n38935 & n15953 ;
  assign n15957 = n15762 | n15956 ;
  assign n38949 = ~n15955 ;
  assign n15958 = n38949 & n15957 ;
  assign n38950 = ~n15958 ;
  assign n15959 = n6600 & n38950 ;
  assign n15960 = n165 | n15959 ;
  assign n38951 = ~n15960 ;
  assign n16014 = n38951 & n15995 ;
  assign n16015 = n15714 | n16014 ;
  assign n38952 = ~n15997 ;
  assign n16016 = n38952 & n16015 ;
  assign n38953 = ~n16016 ;
  assign n16017 = n166 & n38953 ;
  assign n15273 = n15264 | n15265 ;
  assign n38954 = ~n15273 ;
  assign n15670 = n38954 & n148 ;
  assign n15671 = n14964 | n15670 ;
  assign n38955 = ~n15265 ;
  assign n15271 = n14964 & n38955 ;
  assign n15272 = n38601 & n15271 ;
  assign n15674 = n15272 & n148 ;
  assign n38956 = ~n15674 ;
  assign n15675 = n15671 & n38956 ;
  assign n15998 = n166 | n15997 ;
  assign n38957 = ~n15998 ;
  assign n16018 = n38957 & n16015 ;
  assign n16019 = n15675 | n16018 ;
  assign n38958 = ~n16017 ;
  assign n16020 = n38958 & n16019 ;
  assign n38959 = ~n16020 ;
  assign n16021 = n5352 & n38959 ;
  assign n15299 = n15268 | n15285 ;
  assign n38960 = ~n15299 ;
  assign n15662 = n38960 & n148 ;
  assign n15663 = n14994 | n15662 ;
  assign n15270 = n14994 & n38611 ;
  assign n38961 = ~n15285 ;
  assign n15298 = n15270 & n38961 ;
  assign n15664 = n15298 & n148 ;
  assign n38962 = ~n15664 ;
  assign n15665 = n15663 & n38962 ;
  assign n15975 = n15957 & n38941 ;
  assign n15976 = n15686 | n15975 ;
  assign n38963 = ~n15959 ;
  assign n15977 = n38963 & n15976 ;
  assign n38964 = ~n15977 ;
  assign n15978 = n165 & n38964 ;
  assign n15979 = n38951 & n15976 ;
  assign n15980 = n15714 | n15979 ;
  assign n38965 = ~n15978 ;
  assign n15981 = n38965 & n15980 ;
  assign n38966 = ~n15981 ;
  assign n15982 = n166 & n38966 ;
  assign n15983 = n5352 | n15982 ;
  assign n38967 = ~n15983 ;
  assign n16039 = n38967 & n16019 ;
  assign n16040 = n15665 | n16039 ;
  assign n38968 = ~n16021 ;
  assign n16041 = n38968 & n16040 ;
  assign n38969 = ~n16041 ;
  assign n16042 = n168 & n38969 ;
  assign n15297 = n15288 | n15289 ;
  assign n38970 = ~n15297 ;
  assign n15660 = n38970 & n148 ;
  assign n15661 = n14957 | n15660 ;
  assign n38971 = ~n15289 ;
  assign n15295 = n14957 & n38971 ;
  assign n15296 = n38617 & n15295 ;
  assign n15743 = n15296 & n148 ;
  assign n38972 = ~n15743 ;
  assign n15744 = n15661 & n38972 ;
  assign n16022 = n4934 | n16021 ;
  assign n38973 = ~n16022 ;
  assign n16043 = n38973 & n16040 ;
  assign n16044 = n15744 | n16043 ;
  assign n38974 = ~n16042 ;
  assign n16045 = n38974 & n16044 ;
  assign n38975 = ~n16045 ;
  assign n16046 = n169 & n38975 ;
  assign n15294 = n14949 & n38627 ;
  assign n38976 = ~n15309 ;
  assign n15322 = n15294 & n38976 ;
  assign n15655 = n15322 & n148 ;
  assign n15323 = n15292 | n15309 ;
  assign n38977 = ~n15323 ;
  assign n15657 = n38977 & n148 ;
  assign n15658 = n14949 | n15657 ;
  assign n38978 = ~n15655 ;
  assign n15659 = n38978 & n15658 ;
  assign n15999 = n15980 & n38957 ;
  assign n16000 = n15675 | n15999 ;
  assign n38979 = ~n15982 ;
  assign n16001 = n38979 & n16000 ;
  assign n38980 = ~n16001 ;
  assign n16002 = n167 & n38980 ;
  assign n16003 = n38967 & n16000 ;
  assign n16004 = n15665 | n16003 ;
  assign n38981 = ~n16002 ;
  assign n16005 = n38981 & n16004 ;
  assign n38982 = ~n16005 ;
  assign n16006 = n4934 & n38982 ;
  assign n16007 = n169 | n16006 ;
  assign n38983 = ~n16007 ;
  assign n16063 = n38983 & n16044 ;
  assign n16064 = n15659 | n16063 ;
  assign n38984 = ~n16046 ;
  assign n16065 = n38984 & n16064 ;
  assign n38985 = ~n16065 ;
  assign n16066 = n170 & n38985 ;
  assign n38986 = ~n15313 ;
  assign n15319 = n14952 & n38986 ;
  assign n15320 = n38633 & n15319 ;
  assign n15652 = n15320 & n148 ;
  assign n15321 = n15312 | n15313 ;
  assign n38987 = ~n15321 ;
  assign n15667 = n38987 & n148 ;
  assign n15668 = n14952 | n15667 ;
  assign n38988 = ~n15652 ;
  assign n15669 = n38988 & n15668 ;
  assign n16047 = n170 | n16046 ;
  assign n38989 = ~n16047 ;
  assign n16067 = n38989 & n16064 ;
  assign n16068 = n15669 | n16067 ;
  assign n38990 = ~n16066 ;
  assign n16069 = n38990 & n16068 ;
  assign n38991 = ~n16069 ;
  assign n16070 = n3940 & n38991 ;
  assign n15347 = n15316 | n15333 ;
  assign n38992 = ~n15347 ;
  assign n15703 = n38992 & n148 ;
  assign n15704 = n14968 | n15703 ;
  assign n15318 = n14968 & n38643 ;
  assign n38993 = ~n15333 ;
  assign n15346 = n15318 & n38993 ;
  assign n15709 = n15346 & n148 ;
  assign n38994 = ~n15709 ;
  assign n15710 = n15704 & n38994 ;
  assign n16023 = n16004 & n38973 ;
  assign n16024 = n15744 | n16023 ;
  assign n38995 = ~n16006 ;
  assign n16025 = n38995 & n16024 ;
  assign n38996 = ~n16025 ;
  assign n16026 = n169 & n38996 ;
  assign n16027 = n38983 & n16024 ;
  assign n16028 = n15659 | n16027 ;
  assign n38997 = ~n16026 ;
  assign n16029 = n38997 & n16028 ;
  assign n38998 = ~n16029 ;
  assign n16030 = n170 & n38998 ;
  assign n16031 = n3940 | n16030 ;
  assign n38999 = ~n16031 ;
  assign n16087 = n38999 & n16068 ;
  assign n16088 = n15710 | n16087 ;
  assign n39000 = ~n16070 ;
  assign n16089 = n39000 & n16088 ;
  assign n39001 = ~n16089 ;
  assign n16090 = n172 & n39001 ;
  assign n39002 = ~n15337 ;
  assign n15343 = n14961 & n39002 ;
  assign n15344 = n38649 & n15343 ;
  assign n15666 = n15344 & n148 ;
  assign n15345 = n15336 | n15337 ;
  assign n39003 = ~n15345 ;
  assign n15749 = n39003 & n148 ;
  assign n15750 = n14961 | n15749 ;
  assign n39004 = ~n15666 ;
  assign n15751 = n39004 & n15750 ;
  assign n16071 = n3631 | n16070 ;
  assign n39005 = ~n16071 ;
  assign n16091 = n39005 & n16088 ;
  assign n16092 = n15751 | n16091 ;
  assign n39006 = ~n16090 ;
  assign n16093 = n39006 & n16092 ;
  assign n39007 = ~n16093 ;
  assign n16094 = n173 & n39007 ;
  assign n15371 = n15340 | n15357 ;
  assign n39008 = ~n15371 ;
  assign n15649 = n39008 & n148 ;
  assign n15650 = n14940 | n15649 ;
  assign n15342 = n14940 & n38659 ;
  assign n39009 = ~n15357 ;
  assign n15370 = n15342 & n39009 ;
  assign n15672 = n15370 & n148 ;
  assign n39010 = ~n15672 ;
  assign n15673 = n15650 & n39010 ;
  assign n16048 = n16028 & n38989 ;
  assign n16049 = n15669 | n16048 ;
  assign n39011 = ~n16030 ;
  assign n16050 = n39011 & n16049 ;
  assign n39012 = ~n16050 ;
  assign n16051 = n171 & n39012 ;
  assign n16052 = n38999 & n16049 ;
  assign n16053 = n15710 | n16052 ;
  assign n39013 = ~n16051 ;
  assign n16054 = n39013 & n16053 ;
  assign n39014 = ~n16054 ;
  assign n16055 = n3631 & n39014 ;
  assign n16056 = n173 | n16055 ;
  assign n39015 = ~n16056 ;
  assign n16111 = n39015 & n16092 ;
  assign n16112 = n15673 | n16111 ;
  assign n39016 = ~n16094 ;
  assign n16113 = n39016 & n16112 ;
  assign n39017 = ~n16113 ;
  assign n16114 = n174 & n39017 ;
  assign n15369 = n15360 | n15361 ;
  assign n39018 = ~n15369 ;
  assign n15641 = n39018 & n148 ;
  assign n15642 = n15021 | n15641 ;
  assign n39019 = ~n15361 ;
  assign n15367 = n15021 & n39019 ;
  assign n15368 = n38665 & n15367 ;
  assign n15645 = n15368 & n148 ;
  assign n39020 = ~n15645 ;
  assign n15646 = n15642 & n39020 ;
  assign n16095 = n174 | n16094 ;
  assign n39021 = ~n16095 ;
  assign n16115 = n39021 & n16112 ;
  assign n16116 = n15646 | n16115 ;
  assign n39022 = ~n16114 ;
  assign n16117 = n39022 & n16116 ;
  assign n39023 = ~n16117 ;
  assign n16118 = n2753 & n39023 ;
  assign n15366 = n15006 & n38675 ;
  assign n39024 = ~n15381 ;
  assign n15394 = n15366 & n39024 ;
  assign n15702 = n15394 & n148 ;
  assign n15395 = n15364 | n15381 ;
  assign n39025 = ~n15395 ;
  assign n15717 = n39025 & n148 ;
  assign n15718 = n15006 | n15717 ;
  assign n39026 = ~n15702 ;
  assign n15719 = n39026 & n15718 ;
  assign n16072 = n16053 & n39005 ;
  assign n16073 = n15751 | n16072 ;
  assign n39027 = ~n16055 ;
  assign n16074 = n39027 & n16073 ;
  assign n39028 = ~n16074 ;
  assign n16075 = n173 & n39028 ;
  assign n16076 = n39015 & n16073 ;
  assign n16077 = n15673 | n16076 ;
  assign n39029 = ~n16075 ;
  assign n16078 = n39029 & n16077 ;
  assign n39030 = ~n16078 ;
  assign n16079 = n174 & n39030 ;
  assign n16080 = n2753 | n16079 ;
  assign n39031 = ~n16080 ;
  assign n16134 = n39031 & n16116 ;
  assign n16135 = n15719 | n16134 ;
  assign n39032 = ~n16118 ;
  assign n16136 = n39032 & n16135 ;
  assign n39033 = ~n16136 ;
  assign n16137 = n176 & n39033 ;
  assign n15393 = n15384 | n15385 ;
  assign n39034 = ~n15393 ;
  assign n15639 = n39034 & n148 ;
  assign n15640 = n15009 | n15639 ;
  assign n39035 = ~n15385 ;
  assign n15391 = n15009 & n39035 ;
  assign n15392 = n38681 & n15391 ;
  assign n15812 = n15392 & n15807 ;
  assign n39036 = ~n15812 ;
  assign n15813 = n15640 & n39036 ;
  assign n16119 = n2431 | n16118 ;
  assign n39037 = ~n16119 ;
  assign n16138 = n39037 & n16135 ;
  assign n16139 = n15813 | n16138 ;
  assign n39038 = ~n16137 ;
  assign n16140 = n39038 & n16139 ;
  assign n39039 = ~n16140 ;
  assign n16141 = n177 & n39039 ;
  assign n15419 = n15388 | n15405 ;
  assign n39040 = ~n15419 ;
  assign n15635 = n39040 & n148 ;
  assign n15636 = n14927 | n15635 ;
  assign n15389 = n14927 & n38691 ;
  assign n39041 = ~n15405 ;
  assign n15418 = n15389 & n39041 ;
  assign n15810 = n15418 & n15807 ;
  assign n39042 = ~n15810 ;
  assign n15811 = n15636 & n39042 ;
  assign n16096 = n16077 & n39021 ;
  assign n16097 = n15646 | n16096 ;
  assign n39043 = ~n16079 ;
  assign n16098 = n39043 & n16097 ;
  assign n39044 = ~n16098 ;
  assign n16099 = n175 & n39044 ;
  assign n16100 = n39031 & n16097 ;
  assign n16101 = n15719 | n16100 ;
  assign n39045 = ~n16099 ;
  assign n16102 = n39045 & n16101 ;
  assign n39046 = ~n16102 ;
  assign n16103 = n2431 & n39046 ;
  assign n16104 = n177 | n16103 ;
  assign n39047 = ~n16104 ;
  assign n16158 = n39047 & n16139 ;
  assign n16159 = n15811 | n16158 ;
  assign n39048 = ~n16141 ;
  assign n16160 = n39048 & n16159 ;
  assign n39049 = ~n16160 ;
  assign n16161 = n178 & n39049 ;
  assign n15417 = n15408 | n15409 ;
  assign n39050 = ~n15417 ;
  assign n15630 = n39050 & n148 ;
  assign n15631 = n14990 | n15630 ;
  assign n39051 = ~n15409 ;
  assign n15415 = n14990 & n39051 ;
  assign n15416 = n38697 & n15415 ;
  assign n15808 = n15416 & n15807 ;
  assign n39052 = ~n15808 ;
  assign n15809 = n15631 & n39052 ;
  assign n16142 = n178 | n16141 ;
  assign n39053 = ~n16142 ;
  assign n16162 = n39053 & n16159 ;
  assign n16163 = n15809 | n16162 ;
  assign n39054 = ~n16161 ;
  assign n16164 = n39054 & n16163 ;
  assign n39055 = ~n16164 ;
  assign n16165 = n1707 & n39055 ;
  assign n15435 = n15412 | n15429 ;
  assign n39056 = ~n15435 ;
  assign n15624 = n39056 & n148 ;
  assign n15625 = n14999 | n15624 ;
  assign n15414 = n14999 & n38707 ;
  assign n39057 = ~n15429 ;
  assign n15434 = n15414 & n39057 ;
  assign n15626 = n15434 & n148 ;
  assign n39058 = ~n15626 ;
  assign n15627 = n15625 & n39058 ;
  assign n16120 = n16101 & n39037 ;
  assign n16121 = n15813 | n16120 ;
  assign n39059 = ~n16103 ;
  assign n16122 = n39059 & n16121 ;
  assign n39060 = ~n16122 ;
  assign n16123 = n177 & n39060 ;
  assign n16124 = n39047 & n16121 ;
  assign n16125 = n15811 | n16124 ;
  assign n39061 = ~n16123 ;
  assign n16126 = n39061 & n16125 ;
  assign n39062 = ~n16126 ;
  assign n16127 = n178 & n39062 ;
  assign n16128 = n1707 | n16127 ;
  assign n39063 = ~n16128 ;
  assign n16172 = n39063 & n16163 ;
  assign n16173 = n15627 | n16172 ;
  assign n39064 = ~n16165 ;
  assign n16174 = n39064 & n16173 ;
  assign n39065 = ~n16174 ;
  assign n16175 = n180 & n39065 ;
  assign n16166 = n1487 | n16165 ;
  assign n39066 = ~n16166 ;
  assign n16176 = n39066 & n16173 ;
  assign n39067 = ~n15433 ;
  assign n15490 = n39067 & n15469 ;
  assign n15491 = n38734 & n15490 ;
  assign n15708 = n15491 & n148 ;
  assign n15445 = n15433 | n15443 ;
  assign n39068 = ~n15445 ;
  assign n15765 = n39068 & n148 ;
  assign n16198 = n15469 | n15765 ;
  assign n39069 = ~n15708 ;
  assign n16199 = n39069 & n16198 ;
  assign n16200 = n16176 | n16199 ;
  assign n39070 = ~n16175 ;
  assign n16201 = n39070 & n16200 ;
  assign n39071 = ~n16201 ;
  assign n16202 = n181 & n39071 ;
  assign n15474 = n15042 & n38723 ;
  assign n39072 = ~n15475 ;
  assign n15488 = n15474 & n39072 ;
  assign n15687 = n15488 & n148 ;
  assign n15489 = n15472 | n15475 ;
  assign n39073 = ~n15489 ;
  assign n15766 = n39073 & n148 ;
  assign n15767 = n15042 | n15766 ;
  assign n39074 = ~n15687 ;
  assign n15768 = n39074 & n15767 ;
  assign n16143 = n16125 & n39053 ;
  assign n16144 = n15809 | n16143 ;
  assign n39075 = ~n16127 ;
  assign n16145 = n39075 & n16144 ;
  assign n39076 = ~n16145 ;
  assign n16146 = n179 & n39076 ;
  assign n16147 = n39063 & n16144 ;
  assign n16148 = n15627 | n16147 ;
  assign n39077 = ~n16146 ;
  assign n16149 = n39077 & n16148 ;
  assign n39078 = ~n16149 ;
  assign n16150 = n1487 & n39078 ;
  assign n16151 = n181 | n16150 ;
  assign n39079 = ~n16151 ;
  assign n16205 = n39079 & n16200 ;
  assign n16206 = n15768 | n16205 ;
  assign n39080 = ~n16202 ;
  assign n16207 = n39080 & n16206 ;
  assign n39081 = ~n16207 ;
  assign n16208 = n182 & n39081 ;
  assign n39082 = ~n15479 ;
  assign n15485 = n15048 & n39082 ;
  assign n15486 = n38729 & n15485 ;
  assign n15711 = n15486 & n148 ;
  assign n15487 = n15478 | n15479 ;
  assign n39083 = ~n15487 ;
  assign n15769 = n39083 & n148 ;
  assign n15770 = n15048 | n15769 ;
  assign n39084 = ~n15711 ;
  assign n15771 = n39084 & n15770 ;
  assign n16203 = n182 | n16202 ;
  assign n39085 = ~n16203 ;
  assign n16209 = n39085 & n16206 ;
  assign n16210 = n15771 | n16209 ;
  assign n39086 = ~n16208 ;
  assign n16211 = n39086 & n16210 ;
  assign n39087 = ~n16211 ;
  assign n16212 = n996 & n39087 ;
  assign n15514 = n15482 | n15500 ;
  assign n39088 = ~n15514 ;
  assign n15683 = n39088 & n148 ;
  assign n15684 = n15050 | n15683 ;
  assign n15484 = n15050 & n38739 ;
  assign n39089 = ~n15500 ;
  assign n15513 = n15484 & n39089 ;
  assign n15772 = n15513 & n148 ;
  assign n39090 = ~n15772 ;
  assign n15773 = n15684 & n39090 ;
  assign n16167 = n16148 & n39066 ;
  assign n16217 = n16167 | n16199 ;
  assign n39091 = ~n16150 ;
  assign n16218 = n39091 & n16217 ;
  assign n39092 = ~n16218 ;
  assign n16219 = n181 & n39092 ;
  assign n16220 = n39079 & n16217 ;
  assign n16221 = n15768 | n16220 ;
  assign n39093 = ~n16219 ;
  assign n16222 = n39093 & n16221 ;
  assign n39094 = ~n16222 ;
  assign n16223 = n182 & n39094 ;
  assign n16224 = n183 | n16223 ;
  assign n39095 = ~n16224 ;
  assign n16225 = n16210 & n39095 ;
  assign n16226 = n15773 | n16225 ;
  assign n39096 = ~n16212 ;
  assign n16227 = n39096 & n16226 ;
  assign n39097 = ~n16227 ;
  assign n16228 = n184 & n39097 ;
  assign n39098 = ~n15504 ;
  assign n15505 = n15054 & n39098 ;
  assign n15506 = n38745 & n15505 ;
  assign n15776 = n15506 & n148 ;
  assign n15507 = n15503 | n15504 ;
  assign n39099 = ~n15507 ;
  assign n15777 = n39099 & n148 ;
  assign n15778 = n15054 | n15777 ;
  assign n39100 = ~n15776 ;
  assign n15779 = n39100 & n15778 ;
  assign n16213 = n838 | n16212 ;
  assign n39101 = ~n16213 ;
  assign n16229 = n39101 & n16226 ;
  assign n16230 = n15779 | n16229 ;
  assign n39102 = ~n16228 ;
  assign n16231 = n39102 & n16230 ;
  assign n39103 = ~n16231 ;
  assign n16232 = n185 & n39103 ;
  assign n15538 = n15510 | n15524 ;
  assign n39104 = ~n15538 ;
  assign n15741 = n39104 & n148 ;
  assign n15742 = n15057 | n15741 ;
  assign n15512 = n15057 & n38755 ;
  assign n39105 = ~n15524 ;
  assign n15537 = n15512 & n39105 ;
  assign n15780 = n15537 & n148 ;
  assign n39106 = ~n15780 ;
  assign n15781 = n15742 & n39106 ;
  assign n16235 = n39085 & n16221 ;
  assign n16236 = n15771 | n16235 ;
  assign n39107 = ~n16223 ;
  assign n16237 = n39107 & n16236 ;
  assign n39108 = ~n16237 ;
  assign n16238 = n183 & n39108 ;
  assign n16239 = n39095 & n16236 ;
  assign n16240 = n15773 | n16239 ;
  assign n39109 = ~n16238 ;
  assign n16241 = n39109 & n16240 ;
  assign n39110 = ~n16241 ;
  assign n16242 = n838 & n39110 ;
  assign n16243 = n185 | n16242 ;
  assign n39111 = ~n16243 ;
  assign n16244 = n16230 & n39111 ;
  assign n16245 = n15781 | n16244 ;
  assign n39112 = ~n16232 ;
  assign n16246 = n39112 & n16245 ;
  assign n39113 = ~n16246 ;
  assign n16247 = n186 & n39113 ;
  assign n39114 = ~n15528 ;
  assign n15534 = n15061 & n39114 ;
  assign n15535 = n38761 & n15534 ;
  assign n15634 = n15535 & n148 ;
  assign n15536 = n15527 | n15528 ;
  assign n39115 = ~n15536 ;
  assign n15782 = n39115 & n148 ;
  assign n15783 = n15061 | n15782 ;
  assign n39116 = ~n15634 ;
  assign n15784 = n39116 & n15783 ;
  assign n16233 = n186 | n16232 ;
  assign n39117 = ~n16233 ;
  assign n16248 = n39117 & n16245 ;
  assign n16249 = n15784 | n16248 ;
  assign n39118 = ~n16247 ;
  assign n16250 = n39118 & n16249 ;
  assign n39119 = ~n16250 ;
  assign n16251 = n528 & n39119 ;
  assign n15562 = n15531 | n15548 ;
  assign n39120 = ~n15562 ;
  assign n15774 = n39120 & n148 ;
  assign n15775 = n15065 | n15774 ;
  assign n15533 = n15065 & n38771 ;
  assign n39121 = ~n15548 ;
  assign n15561 = n15533 & n39121 ;
  assign n15785 = n15561 & n148 ;
  assign n39122 = ~n15785 ;
  assign n15786 = n15775 & n39122 ;
  assign n16254 = n39101 & n16240 ;
  assign n16255 = n15779 | n16254 ;
  assign n39123 = ~n16242 ;
  assign n16256 = n39123 & n16255 ;
  assign n39124 = ~n16256 ;
  assign n16257 = n185 & n39124 ;
  assign n16258 = n39111 & n16255 ;
  assign n16259 = n15781 | n16258 ;
  assign n39125 = ~n16257 ;
  assign n16260 = n39125 & n16259 ;
  assign n39126 = ~n16260 ;
  assign n16261 = n186 & n39126 ;
  assign n16262 = n528 | n16261 ;
  assign n39127 = ~n16262 ;
  assign n16263 = n16249 & n39127 ;
  assign n16264 = n15786 | n16263 ;
  assign n39128 = ~n16251 ;
  assign n16265 = n39128 & n16264 ;
  assign n39129 = ~n16265 ;
  assign n16266 = n188 & n39129 ;
  assign n39130 = ~n15552 ;
  assign n15558 = n15067 & n39130 ;
  assign n15559 = n38777 & n15558 ;
  assign n15787 = n15559 & n148 ;
  assign n15560 = n15551 | n15552 ;
  assign n39131 = ~n15560 ;
  assign n15788 = n39131 & n148 ;
  assign n15789 = n15067 | n15788 ;
  assign n39132 = ~n15787 ;
  assign n15790 = n39132 & n15789 ;
  assign n16252 = n413 | n16251 ;
  assign n39133 = ~n16252 ;
  assign n16267 = n39133 & n16264 ;
  assign n16268 = n15790 | n16267 ;
  assign n39134 = ~n16266 ;
  assign n16269 = n39134 & n16268 ;
  assign n39135 = ~n16269 ;
  assign n16270 = n189 & n39135 ;
  assign n15557 = n15071 & n38787 ;
  assign n39136 = ~n15572 ;
  assign n15583 = n15557 & n39136 ;
  assign n15791 = n15583 & n148 ;
  assign n15584 = n15555 | n15572 ;
  assign n39137 = ~n15584 ;
  assign n15792 = n39137 & n148 ;
  assign n15793 = n15071 | n15792 ;
  assign n39138 = ~n15791 ;
  assign n15794 = n39138 & n15793 ;
  assign n16273 = n39117 & n16259 ;
  assign n16274 = n15784 | n16273 ;
  assign n39139 = ~n16261 ;
  assign n16275 = n39139 & n16274 ;
  assign n39140 = ~n16275 ;
  assign n16276 = n187 & n39140 ;
  assign n16277 = n39127 & n16274 ;
  assign n16278 = n15786 | n16277 ;
  assign n39141 = ~n16276 ;
  assign n16279 = n39141 & n16278 ;
  assign n39142 = ~n16279 ;
  assign n16280 = n413 & n39142 ;
  assign n16281 = n189 | n16280 ;
  assign n39143 = ~n16281 ;
  assign n16282 = n16268 & n39143 ;
  assign n16283 = n15794 | n16282 ;
  assign n39144 = ~n16270 ;
  assign n16284 = n39144 & n16283 ;
  assign n39145 = ~n16284 ;
  assign n16285 = n190 & n39145 ;
  assign n16190 = n38792 & n15590 ;
  assign n39146 = ~n16190 ;
  assign n16191 = n15073 & n39146 ;
  assign n16192 = n38793 & n16191 ;
  assign n16193 = n148 & n16192 ;
  assign n16194 = n15575 | n16190 ;
  assign n39147 = ~n16194 ;
  assign n16195 = n148 & n39147 ;
  assign n16196 = n15073 | n16195 ;
  assign n39148 = ~n16193 ;
  assign n16197 = n39148 & n16196 ;
  assign n16271 = n190 | n16270 ;
  assign n39149 = ~n16271 ;
  assign n16286 = n39149 & n16283 ;
  assign n16287 = n16197 | n16286 ;
  assign n39150 = ~n16285 ;
  assign n16288 = n39150 & n16287 ;
  assign n39151 = ~n16288 ;
  assign n16289 = n287 & n39151 ;
  assign n15582 = n15077 & n38803 ;
  assign n39152 = ~n15594 ;
  assign n15599 = n15582 & n39152 ;
  assign n15707 = n15599 & n148 ;
  assign n15598 = n15579 | n15594 ;
  assign n39153 = ~n15598 ;
  assign n15795 = n39153 & n148 ;
  assign n15796 = n15077 | n15795 ;
  assign n39154 = ~n15707 ;
  assign n15797 = n39154 & n15796 ;
  assign n16292 = n39133 & n16278 ;
  assign n16293 = n15790 | n16292 ;
  assign n39155 = ~n16280 ;
  assign n16294 = n39155 & n16293 ;
  assign n39156 = ~n16294 ;
  assign n16295 = n189 & n39156 ;
  assign n16296 = n39143 & n16293 ;
  assign n16297 = n15794 | n16296 ;
  assign n39157 = ~n16295 ;
  assign n16298 = n39157 & n16297 ;
  assign n39158 = ~n16298 ;
  assign n16299 = n190 & n39158 ;
  assign n16304 = n287 | n16299 ;
  assign n39159 = ~n16304 ;
  assign n16305 = n16287 & n39159 ;
  assign n16306 = n15797 | n16305 ;
  assign n39160 = ~n16289 ;
  assign n16307 = n39160 & n16306 ;
  assign n16308 = n16187 | n16307 ;
  assign n16309 = n31336 & n16308 ;
  assign n15452 = n15078 | n15450 ;
  assign n39161 = ~n15452 ;
  assign n15453 = n14925 & n39161 ;
  assign n15454 = n38826 & n15453 ;
  assign n15606 = n15454 & n38827 ;
  assign n15618 = n15606 & n38828 ;
  assign n15610 = n192 & n15609 ;
  assign n39162 = ~n15079 ;
  assign n15798 = n39162 & n148 ;
  assign n39163 = ~n15798 ;
  assign n15799 = n15608 & n39163 ;
  assign n39164 = ~n15799 ;
  assign n15800 = n15610 & n39164 ;
  assign n15801 = n15618 | n15800 ;
  assign n16290 = n16186 & n39160 ;
  assign n16310 = n16290 & n16306 ;
  assign n16321 = n15801 | n16310 ;
  assign n16322 = n16309 | n16321 ;
  assign n16319 = n16186 | n16307 ;
  assign n16331 = n39149 & n16297 ;
  assign n16332 = n16197 | n16331 ;
  assign n39165 = ~n16299 ;
  assign n16333 = n39165 & n16332 ;
  assign n39166 = ~n16333 ;
  assign n16334 = n191 & n39166 ;
  assign n16300 = n191 | n16299 ;
  assign n39167 = ~n16300 ;
  assign n16335 = n39167 & n16332 ;
  assign n16336 = n15797 | n16335 ;
  assign n39168 = ~n16334 ;
  assign n16337 = n39168 & n16336 ;
  assign n16338 = n16187 | n16337 ;
  assign n16339 = n31336 & n16338 ;
  assign n16340 = n16290 & n16336 ;
  assign n16341 = n15801 | n16340 ;
  assign n147 = n16339 | n16341 ;
  assign n39169 = ~n16319 ;
  assign n16882 = n39169 & n147 ;
  assign n16883 = n16310 | n16882 ;
  assign n16291 = n15797 & n39160 ;
  assign n16301 = n16287 & n39167 ;
  assign n39170 = ~n16301 ;
  assign n16302 = n16291 & n39170 ;
  assign n16374 = n16302 & n147 ;
  assign n16303 = n16289 | n16301 ;
  assign n39171 = ~n16303 ;
  assign n16884 = n39171 & n147 ;
  assign n16885 = n15797 | n16884 ;
  assign n39172 = ~n16374 ;
  assign n16886 = n39172 & n16885 ;
  assign n16887 = n16883 | n16886 ;
  assign n218 = x34 | x35 ;
  assign n39173 = ~x36 ;
  assign n220 = n39173 & n218 ;
  assign n39174 = ~n16322 ;
  assign n16325 = x36 & n39174 ;
  assign n16326 = n220 | n16325 ;
  assign n39175 = ~n16326 ;
  assign n16327 = n15807 & n39175 ;
  assign n219 = x36 | n218 ;
  assign n15457 = n219 & n38825 ;
  assign n15458 = n38826 & n15457 ;
  assign n15607 = n15458 & n38827 ;
  assign n15620 = n15607 & n38828 ;
  assign n16416 = x36 & n147 ;
  assign n39176 = ~n16416 ;
  assign n16417 = n15620 & n39176 ;
  assign n39177 = ~n215 ;
  assign n16402 = n39177 & n147 ;
  assign n16468 = n39173 & n147 ;
  assign n39178 = ~n16468 ;
  assign n16469 = x37 & n39178 ;
  assign n16470 = n16402 | n16469 ;
  assign n16472 = n16417 | n16470 ;
  assign n39179 = ~n16327 ;
  assign n16473 = n39179 & n16472 ;
  assign n39180 = ~n16473 ;
  assign n16474 = n149 & n39180 ;
  assign n39181 = ~n15618 ;
  assign n15803 = n39181 & n148 ;
  assign n39182 = ~n15800 ;
  assign n15804 = n39182 & n15803 ;
  assign n39183 = ~n16310 ;
  assign n16311 = n15804 & n39183 ;
  assign n39184 = ~n16309 ;
  assign n16312 = n39184 & n16311 ;
  assign n16403 = n16312 | n16402 ;
  assign n16404 = x38 & n16403 ;
  assign n16313 = x38 | n16312 ;
  assign n16405 = n16313 | n16402 ;
  assign n39185 = ~n16404 ;
  assign n16406 = n39185 & n16405 ;
  assign n16448 = n219 & n39176 ;
  assign n39186 = ~n16448 ;
  assign n16449 = n148 & n39186 ;
  assign n16450 = n149 | n16449 ;
  assign n39187 = ~n16450 ;
  assign n16476 = n39187 & n16472 ;
  assign n16477 = n16406 | n16476 ;
  assign n39188 = ~n16474 ;
  assign n16478 = n39188 & n16477 ;
  assign n39189 = ~n16478 ;
  assign n16479 = n150 & n39189 ;
  assign n16177 = n15682 | n15820 ;
  assign n39190 = ~n16177 ;
  assign n16370 = n39190 & n147 ;
  assign n16371 = n15720 | n16370 ;
  assign n16178 = n15720 & n39190 ;
  assign n16438 = n16178 & n147 ;
  assign n39191 = ~n16438 ;
  assign n16439 = n16371 & n39191 ;
  assign n16328 = n149 | n16327 ;
  assign n39192 = ~n16328 ;
  assign n16482 = n39192 & n16472 ;
  assign n16483 = n16406 | n16482 ;
  assign n16329 = n148 & n39175 ;
  assign n39193 = ~n16329 ;
  assign n16490 = n39193 & n16472 ;
  assign n39194 = ~n16490 ;
  assign n16491 = n149 & n39194 ;
  assign n16492 = n150 | n16491 ;
  assign n39195 = ~n16492 ;
  assign n16493 = n16483 & n39195 ;
  assign n16494 = n16439 | n16493 ;
  assign n39196 = ~n16479 ;
  assign n16495 = n39196 & n16494 ;
  assign n39197 = ~n16495 ;
  assign n16496 = n13662 & n39197 ;
  assign n16481 = n13662 | n16479 ;
  assign n39198 = ~n16481 ;
  assign n16498 = n39198 & n16494 ;
  assign n39199 = ~n15722 ;
  assign n15727 = n39199 & n15725 ;
  assign n39200 = ~n15729 ;
  assign n15733 = n15727 & n39200 ;
  assign n16421 = n15733 & n147 ;
  assign n15734 = n15722 | n15729 ;
  assign n39201 = ~n15734 ;
  assign n16506 = n39201 & n147 ;
  assign n16507 = n15725 | n16506 ;
  assign n39202 = ~n16421 ;
  assign n16508 = n39202 & n16507 ;
  assign n16509 = n16498 | n16508 ;
  assign n39203 = ~n16496 ;
  assign n16510 = n39203 & n16509 ;
  assign n39204 = ~n16510 ;
  assign n16511 = n152 & n39204 ;
  assign n15829 = n15716 & n38839 ;
  assign n39205 = ~n15731 ;
  assign n15830 = n39205 & n15829 ;
  assign n16395 = n15830 & n147 ;
  assign n15831 = n15731 | n15828 ;
  assign n39206 = ~n15831 ;
  assign n16443 = n39206 & n147 ;
  assign n16444 = n15716 | n16443 ;
  assign n39207 = ~n16395 ;
  assign n16445 = n39207 & n16444 ;
  assign n16497 = n152 | n16496 ;
  assign n39208 = ~n16497 ;
  assign n16512 = n39208 & n16509 ;
  assign n16513 = n16445 | n16512 ;
  assign n39209 = ~n16511 ;
  assign n16514 = n39209 & n16513 ;
  assign n39210 = ~n16514 ;
  assign n16515 = n153 & n39210 ;
  assign n39211 = ~n15833 ;
  assign n15842 = n15740 & n39211 ;
  assign n15843 = n38867 & n15842 ;
  assign n16401 = n15843 & n147 ;
  assign n15844 = n15826 | n15833 ;
  assign n39212 = ~n15844 ;
  assign n16440 = n39212 & n147 ;
  assign n16441 = n15740 | n16440 ;
  assign n39213 = ~n16401 ;
  assign n16442 = n39213 & n16441 ;
  assign n16475 = n150 | n16474 ;
  assign n39214 = ~n16475 ;
  assign n16484 = n39214 & n16483 ;
  assign n16485 = n16439 | n16484 ;
  assign n16486 = n39196 & n16485 ;
  assign n39215 = ~n16486 ;
  assign n16487 = n151 & n39215 ;
  assign n16488 = n39198 & n16485 ;
  assign n16518 = n16488 | n16508 ;
  assign n39216 = ~n16487 ;
  assign n16519 = n39216 & n16518 ;
  assign n39217 = ~n16519 ;
  assign n16520 = n13079 & n39217 ;
  assign n16521 = n153 | n16520 ;
  assign n39218 = ~n16521 ;
  assign n16522 = n16513 & n39218 ;
  assign n16523 = n16442 | n16522 ;
  assign n39219 = ~n16515 ;
  assign n16524 = n39219 & n16523 ;
  assign n39220 = ~n16524 ;
  assign n16525 = n154 & n39220 ;
  assign n15869 = n15695 & n38856 ;
  assign n39221 = ~n15837 ;
  assign n15870 = n39221 & n15869 ;
  assign n16324 = n15870 & n16322 ;
  assign n15868 = n15837 | n15853 ;
  assign n39222 = ~n15868 ;
  assign n16463 = n39222 & n147 ;
  assign n16464 = n15695 | n16463 ;
  assign n39223 = ~n16324 ;
  assign n16465 = n39223 & n16464 ;
  assign n16516 = n154 | n16515 ;
  assign n39224 = ~n16516 ;
  assign n16526 = n39224 & n16523 ;
  assign n16527 = n16465 | n16526 ;
  assign n39225 = ~n16525 ;
  assign n16528 = n39225 & n16527 ;
  assign n39226 = ~n16528 ;
  assign n16529 = n11067 & n39226 ;
  assign n39227 = ~n15855 ;
  assign n15866 = n15698 & n39227 ;
  assign n15867 = n38883 & n15866 ;
  assign n16454 = n15867 & n147 ;
  assign n15865 = n15840 | n15855 ;
  assign n39228 = ~n15865 ;
  assign n16455 = n39228 & n147 ;
  assign n16456 = n15698 | n16455 ;
  assign n39229 = ~n16454 ;
  assign n16457 = n39229 & n16456 ;
  assign n16537 = n39208 & n16518 ;
  assign n16538 = n16445 | n16537 ;
  assign n39230 = ~n16520 ;
  assign n16539 = n39230 & n16538 ;
  assign n39231 = ~n16539 ;
  assign n16540 = n153 & n39231 ;
  assign n16541 = n39218 & n16538 ;
  assign n16542 = n16442 | n16541 ;
  assign n39232 = ~n16540 ;
  assign n16543 = n39232 & n16542 ;
  assign n39233 = ~n16543 ;
  assign n16544 = n154 & n39233 ;
  assign n16545 = n11067 | n16544 ;
  assign n39234 = ~n16545 ;
  assign n16546 = n16527 & n39234 ;
  assign n16547 = n16457 | n16546 ;
  assign n39235 = ~n16529 ;
  assign n16548 = n39235 & n16547 ;
  assign n39236 = ~n16548 ;
  assign n16549 = n156 & n39236 ;
  assign n15893 = n15737 & n38872 ;
  assign n39237 = ~n15859 ;
  assign n15894 = n39237 & n15893 ;
  assign n16407 = n15894 & n147 ;
  assign n15864 = n15858 | n15859 ;
  assign n39238 = ~n15864 ;
  assign n16460 = n39238 & n147 ;
  assign n16461 = n15737 | n16460 ;
  assign n39239 = ~n16407 ;
  assign n16462 = n39239 & n16461 ;
  assign n16530 = n10657 | n16529 ;
  assign n39240 = ~n16530 ;
  assign n16550 = n39240 & n16547 ;
  assign n16551 = n16462 | n16550 ;
  assign n39241 = ~n16549 ;
  assign n16552 = n39241 & n16551 ;
  assign n39242 = ~n16552 ;
  assign n16553 = n157 & n39242 ;
  assign n15892 = n15862 | n15880 ;
  assign n39243 = ~n15892 ;
  assign n16387 = n39243 & n147 ;
  assign n16388 = n15817 | n16387 ;
  assign n39244 = ~n15880 ;
  assign n15890 = n15817 & n39244 ;
  assign n15891 = n38899 & n15890 ;
  assign n16422 = n15891 & n147 ;
  assign n39245 = ~n16422 ;
  assign n16423 = n16388 & n39245 ;
  assign n16561 = n39224 & n16542 ;
  assign n16562 = n16465 | n16561 ;
  assign n39246 = ~n16544 ;
  assign n16563 = n39246 & n16562 ;
  assign n39247 = ~n16563 ;
  assign n16564 = n155 & n39247 ;
  assign n16565 = n39234 & n16562 ;
  assign n16566 = n16457 | n16565 ;
  assign n39248 = ~n16564 ;
  assign n16567 = n39248 & n16566 ;
  assign n39249 = ~n16567 ;
  assign n16568 = n10657 & n39249 ;
  assign n16569 = n157 | n16568 ;
  assign n39250 = ~n16569 ;
  assign n16570 = n16551 & n39250 ;
  assign n16571 = n16423 | n16570 ;
  assign n39251 = ~n16553 ;
  assign n16572 = n39251 & n16571 ;
  assign n39252 = ~n16572 ;
  assign n16573 = n158 & n39252 ;
  assign n16554 = n158 | n16553 ;
  assign n39253 = ~n16554 ;
  assign n16574 = n39253 & n16571 ;
  assign n15917 = n15758 & n38888 ;
  assign n39254 = ~n15884 ;
  assign n15918 = n39254 & n15917 ;
  assign n16434 = n15918 & n147 ;
  assign n15889 = n15883 | n15884 ;
  assign n39255 = ~n15889 ;
  assign n16593 = n39255 & n147 ;
  assign n16594 = n15758 | n16593 ;
  assign n39256 = ~n16434 ;
  assign n16595 = n39256 & n16594 ;
  assign n16596 = n16574 | n16595 ;
  assign n39257 = ~n16573 ;
  assign n16597 = n39257 & n16596 ;
  assign n39258 = ~n16597 ;
  assign n16598 = n8857 & n39258 ;
  assign n16581 = n39240 & n16566 ;
  assign n16582 = n16462 | n16581 ;
  assign n39259 = ~n16568 ;
  assign n16583 = n39259 & n16582 ;
  assign n39260 = ~n16583 ;
  assign n16584 = n157 & n39260 ;
  assign n16585 = n39250 & n16582 ;
  assign n16586 = n16423 | n16585 ;
  assign n39261 = ~n16584 ;
  assign n16587 = n39261 & n16586 ;
  assign n39262 = ~n16587 ;
  assign n16588 = n158 & n39262 ;
  assign n16589 = n8857 | n16588 ;
  assign n39263 = ~n16589 ;
  assign n16600 = n39263 & n16596 ;
  assign n39264 = ~n15904 ;
  assign n15914 = n15677 & n39264 ;
  assign n15915 = n38915 & n15914 ;
  assign n16364 = n15915 & n147 ;
  assign n15916 = n15887 | n15904 ;
  assign n39265 = ~n15916 ;
  assign n16610 = n39265 & n147 ;
  assign n16611 = n15677 | n16610 ;
  assign n39266 = ~n16364 ;
  assign n16612 = n39266 & n16611 ;
  assign n16630 = n16600 | n16612 ;
  assign n39267 = ~n16598 ;
  assign n16631 = n39267 & n16630 ;
  assign n39268 = ~n16631 ;
  assign n16632 = n160 & n39268 ;
  assign n15913 = n15907 | n15908 ;
  assign n39269 = ~n15913 ;
  assign n16354 = n39269 & n147 ;
  assign n16355 = n15756 | n16354 ;
  assign n15941 = n15756 & n38904 ;
  assign n39270 = ~n15908 ;
  assign n15942 = n39270 & n15941 ;
  assign n16504 = n15942 & n147 ;
  assign n39271 = ~n16504 ;
  assign n16505 = n16355 & n39271 ;
  assign n16599 = n160 | n16598 ;
  assign n39272 = ~n16599 ;
  assign n16633 = n39272 & n16630 ;
  assign n16634 = n16505 | n16633 ;
  assign n39273 = ~n16632 ;
  assign n16635 = n39273 & n16634 ;
  assign n39274 = ~n16635 ;
  assign n16636 = n161 & n39274 ;
  assign n39275 = ~n15928 ;
  assign n15938 = n15815 & n39275 ;
  assign n15939 = n38931 & n15938 ;
  assign n16424 = n15939 & n147 ;
  assign n15940 = n15911 | n15928 ;
  assign n39276 = ~n15940 ;
  assign n16451 = n39276 & n147 ;
  assign n16452 = n15815 | n16451 ;
  assign n39277 = ~n16424 ;
  assign n16453 = n39277 & n16452 ;
  assign n16590 = n39253 & n16586 ;
  assign n16604 = n16590 | n16595 ;
  assign n39278 = ~n16588 ;
  assign n16605 = n39278 & n16604 ;
  assign n39279 = ~n16605 ;
  assign n16606 = n159 & n39279 ;
  assign n16607 = n39263 & n16604 ;
  assign n16613 = n16607 | n16612 ;
  assign n39280 = ~n16606 ;
  assign n16614 = n39280 & n16613 ;
  assign n39281 = ~n16614 ;
  assign n16615 = n8534 & n39281 ;
  assign n16616 = n161 | n16615 ;
  assign n39282 = ~n16616 ;
  assign n16648 = n39282 & n16634 ;
  assign n16649 = n16453 | n16648 ;
  assign n39283 = ~n16636 ;
  assign n16650 = n39283 & n16649 ;
  assign n39284 = ~n16650 ;
  assign n16651 = n162 & n39284 ;
  assign n15937 = n15931 | n15932 ;
  assign n39285 = ~n15937 ;
  assign n16393 = n39285 & n147 ;
  assign n16394 = n15754 | n16393 ;
  assign n15964 = n15754 & n38920 ;
  assign n39286 = ~n15932 ;
  assign n15965 = n39286 & n15964 ;
  assign n16458 = n15965 & n147 ;
  assign n39287 = ~n16458 ;
  assign n16459 = n16394 & n39287 ;
  assign n16637 = n162 | n16636 ;
  assign n39288 = ~n16637 ;
  assign n16652 = n39288 & n16649 ;
  assign n16653 = n16459 | n16652 ;
  assign n39289 = ~n16651 ;
  assign n16654 = n39289 & n16653 ;
  assign n39290 = ~n16654 ;
  assign n16655 = n6889 & n39290 ;
  assign n15963 = n15935 | n15952 ;
  assign n39291 = ~n15963 ;
  assign n16391 = n39291 & n147 ;
  assign n16392 = n15764 | n16391 ;
  assign n39292 = ~n15952 ;
  assign n15961 = n15764 & n39292 ;
  assign n15962 = n38947 & n15961 ;
  assign n16432 = n15962 & n147 ;
  assign n39293 = ~n16432 ;
  assign n16433 = n16392 & n39293 ;
  assign n16618 = n39272 & n16613 ;
  assign n16619 = n16505 | n16618 ;
  assign n39294 = ~n16615 ;
  assign n16620 = n39294 & n16619 ;
  assign n39295 = ~n16620 ;
  assign n16621 = n161 & n39295 ;
  assign n16622 = n39282 & n16619 ;
  assign n16623 = n16453 | n16622 ;
  assign n39296 = ~n16621 ;
  assign n16624 = n39296 & n16623 ;
  assign n39297 = ~n16624 ;
  assign n16625 = n162 & n39297 ;
  assign n16626 = n6889 | n16625 ;
  assign n39298 = ~n16626 ;
  assign n16667 = n39298 & n16653 ;
  assign n16668 = n16433 | n16667 ;
  assign n39299 = ~n16655 ;
  assign n16669 = n39299 & n16668 ;
  assign n39300 = ~n16669 ;
  assign n16670 = n164 & n39300 ;
  assign n15989 = n15956 | n15973 ;
  assign n39301 = ~n15989 ;
  assign n16385 = n39301 & n147 ;
  assign n16386 = n15762 | n16385 ;
  assign n15987 = n15762 & n38936 ;
  assign n39302 = ~n15956 ;
  assign n15988 = n39302 & n15987 ;
  assign n16389 = n15988 & n147 ;
  assign n39303 = ~n16389 ;
  assign n16390 = n16386 & n39303 ;
  assign n16656 = n6600 | n16655 ;
  assign n39304 = ~n16656 ;
  assign n16671 = n39304 & n16668 ;
  assign n16672 = n16390 | n16671 ;
  assign n39305 = ~n16670 ;
  assign n16673 = n39305 & n16672 ;
  assign n39306 = ~n16673 ;
  assign n16674 = n165 & n39306 ;
  assign n15986 = n15959 | n15975 ;
  assign n39307 = ~n15986 ;
  assign n16378 = n39307 & n147 ;
  assign n16379 = n15686 | n16378 ;
  assign n39308 = ~n15975 ;
  assign n15984 = n15686 & n39308 ;
  assign n15985 = n38963 & n15984 ;
  assign n16383 = n15985 & n147 ;
  assign n39309 = ~n16383 ;
  assign n16384 = n16379 & n39309 ;
  assign n16638 = n16623 & n39288 ;
  assign n16639 = n16459 | n16638 ;
  assign n39310 = ~n16625 ;
  assign n16640 = n39310 & n16639 ;
  assign n39311 = ~n16640 ;
  assign n16641 = n163 & n39311 ;
  assign n16642 = n39298 & n16639 ;
  assign n16643 = n16433 | n16642 ;
  assign n39312 = ~n16641 ;
  assign n16644 = n39312 & n16643 ;
  assign n39313 = ~n16644 ;
  assign n16645 = n6600 & n39313 ;
  assign n16646 = n165 | n16645 ;
  assign n39314 = ~n16646 ;
  assign n16686 = n39314 & n16672 ;
  assign n16687 = n16384 | n16686 ;
  assign n39315 = ~n16674 ;
  assign n16688 = n39315 & n16687 ;
  assign n39316 = ~n16688 ;
  assign n16689 = n166 & n39316 ;
  assign n16013 = n15979 | n15997 ;
  assign n39317 = ~n16013 ;
  assign n16376 = n39317 & n147 ;
  assign n16377 = n15714 | n16376 ;
  assign n16011 = n15714 & n38952 ;
  assign n39318 = ~n15979 ;
  assign n16012 = n39318 & n16011 ;
  assign n16399 = n16012 & n147 ;
  assign n39319 = ~n16399 ;
  assign n16400 = n16377 & n39319 ;
  assign n16675 = n166 | n16674 ;
  assign n39320 = ~n16675 ;
  assign n16690 = n39320 & n16687 ;
  assign n16691 = n16400 | n16690 ;
  assign n39321 = ~n16689 ;
  assign n16692 = n39321 & n16691 ;
  assign n39322 = ~n16692 ;
  assign n16693 = n5352 & n39322 ;
  assign n16010 = n15982 | n15999 ;
  assign n39323 = ~n16010 ;
  assign n16372 = n39323 & n147 ;
  assign n16373 = n15675 | n16372 ;
  assign n39324 = ~n15999 ;
  assign n16008 = n15675 & n39324 ;
  assign n16009 = n38979 & n16008 ;
  assign n16446 = n16009 & n147 ;
  assign n39325 = ~n16446 ;
  assign n16447 = n16373 & n39325 ;
  assign n16657 = n16643 & n39304 ;
  assign n16658 = n16390 | n16657 ;
  assign n39326 = ~n16645 ;
  assign n16659 = n39326 & n16658 ;
  assign n39327 = ~n16659 ;
  assign n16660 = n165 & n39327 ;
  assign n16661 = n39314 & n16658 ;
  assign n16662 = n16384 | n16661 ;
  assign n39328 = ~n16660 ;
  assign n16663 = n39328 & n16662 ;
  assign n39329 = ~n16663 ;
  assign n16664 = n166 & n39329 ;
  assign n16665 = n5352 | n16664 ;
  assign n39330 = ~n16665 ;
  assign n16705 = n39330 & n16691 ;
  assign n16706 = n16447 | n16705 ;
  assign n39331 = ~n16693 ;
  assign n16707 = n39331 & n16706 ;
  assign n39332 = ~n16707 ;
  assign n16708 = n168 & n39332 ;
  assign n16038 = n16003 | n16021 ;
  assign n39333 = ~n16038 ;
  assign n16358 = n39333 & n147 ;
  assign n16359 = n15665 | n16358 ;
  assign n16036 = n15665 & n38968 ;
  assign n39334 = ~n16003 ;
  assign n16037 = n39334 & n16036 ;
  assign n16365 = n16037 & n147 ;
  assign n39335 = ~n16365 ;
  assign n16366 = n16359 & n39335 ;
  assign n16694 = n4934 | n16693 ;
  assign n39336 = ~n16694 ;
  assign n16709 = n39336 & n16706 ;
  assign n16710 = n16366 | n16709 ;
  assign n39337 = ~n16708 ;
  assign n16711 = n39337 & n16710 ;
  assign n39338 = ~n16711 ;
  assign n16712 = n169 & n39338 ;
  assign n39339 = ~n16023 ;
  assign n16033 = n15744 & n39339 ;
  assign n16034 = n38995 & n16033 ;
  assign n16356 = n16034 & n147 ;
  assign n16035 = n16006 | n16023 ;
  assign n39340 = ~n16035 ;
  assign n16411 = n39340 & n147 ;
  assign n16412 = n15744 | n16411 ;
  assign n39341 = ~n16356 ;
  assign n16413 = n39341 & n16412 ;
  assign n16676 = n16662 & n39320 ;
  assign n16677 = n16400 | n16676 ;
  assign n39342 = ~n16664 ;
  assign n16678 = n39342 & n16677 ;
  assign n39343 = ~n16678 ;
  assign n16679 = n167 & n39343 ;
  assign n16680 = n39330 & n16677 ;
  assign n16681 = n16447 | n16680 ;
  assign n39344 = ~n16679 ;
  assign n16682 = n39344 & n16681 ;
  assign n39345 = ~n16682 ;
  assign n16683 = n4934 & n39345 ;
  assign n16684 = n169 | n16683 ;
  assign n39346 = ~n16684 ;
  assign n16724 = n39346 & n16710 ;
  assign n16725 = n16413 | n16724 ;
  assign n39347 = ~n16712 ;
  assign n16726 = n39347 & n16725 ;
  assign n39348 = ~n16726 ;
  assign n16727 = n170 & n39348 ;
  assign n16061 = n15659 & n38984 ;
  assign n39349 = ~n16027 ;
  assign n16062 = n39349 & n16061 ;
  assign n16360 = n16062 & n147 ;
  assign n16032 = n16026 | n16027 ;
  assign n39350 = ~n16032 ;
  assign n16367 = n39350 & n147 ;
  assign n16368 = n15659 | n16367 ;
  assign n39351 = ~n16360 ;
  assign n16369 = n39351 & n16368 ;
  assign n16713 = n170 | n16712 ;
  assign n39352 = ~n16713 ;
  assign n16728 = n39352 & n16725 ;
  assign n16729 = n16369 | n16728 ;
  assign n39353 = ~n16727 ;
  assign n16730 = n39353 & n16729 ;
  assign n39354 = ~n16730 ;
  assign n16731 = n3940 & n39354 ;
  assign n39355 = ~n16048 ;
  assign n16058 = n15669 & n39355 ;
  assign n16059 = n39011 & n16058 ;
  assign n16353 = n16059 & n147 ;
  assign n16060 = n16030 | n16048 ;
  assign n39356 = ~n16060 ;
  assign n16361 = n39356 & n147 ;
  assign n16362 = n15669 | n16361 ;
  assign n39357 = ~n16353 ;
  assign n16363 = n39357 & n16362 ;
  assign n16695 = n16681 & n39336 ;
  assign n16696 = n16366 | n16695 ;
  assign n39358 = ~n16683 ;
  assign n16697 = n39358 & n16696 ;
  assign n39359 = ~n16697 ;
  assign n16698 = n169 & n39359 ;
  assign n16699 = n39346 & n16696 ;
  assign n16700 = n16413 | n16699 ;
  assign n39360 = ~n16698 ;
  assign n16701 = n39360 & n16700 ;
  assign n39361 = ~n16701 ;
  assign n16702 = n170 & n39361 ;
  assign n16703 = n3940 | n16702 ;
  assign n39362 = ~n16703 ;
  assign n16743 = n39362 & n16729 ;
  assign n16744 = n16363 | n16743 ;
  assign n39363 = ~n16731 ;
  assign n16745 = n39363 & n16744 ;
  assign n39364 = ~n16745 ;
  assign n16746 = n172 & n39364 ;
  assign n16057 = n16051 | n16052 ;
  assign n39365 = ~n16057 ;
  assign n16414 = n39365 & n147 ;
  assign n16415 = n15710 | n16414 ;
  assign n16085 = n15710 & n39000 ;
  assign n39366 = ~n16052 ;
  assign n16086 = n39366 & n16085 ;
  assign n16608 = n16086 & n147 ;
  assign n39367 = ~n16608 ;
  assign n16609 = n16415 & n39367 ;
  assign n16732 = n3631 | n16731 ;
  assign n39368 = ~n16732 ;
  assign n16747 = n39368 & n16744 ;
  assign n16748 = n16609 | n16747 ;
  assign n39369 = ~n16746 ;
  assign n16749 = n39369 & n16748 ;
  assign n39370 = ~n16749 ;
  assign n16750 = n173 & n39370 ;
  assign n16084 = n16055 | n16072 ;
  assign n39371 = ~n16084 ;
  assign n16347 = n39371 & n147 ;
  assign n16348 = n15751 | n16347 ;
  assign n39372 = ~n16072 ;
  assign n16082 = n15751 & n39372 ;
  assign n16083 = n39027 & n16082 ;
  assign n16351 = n16083 & n147 ;
  assign n39373 = ~n16351 ;
  assign n16352 = n16348 & n39373 ;
  assign n16714 = n16700 & n39352 ;
  assign n16715 = n16369 | n16714 ;
  assign n39374 = ~n16702 ;
  assign n16716 = n39374 & n16715 ;
  assign n39375 = ~n16716 ;
  assign n16717 = n171 & n39375 ;
  assign n16718 = n39362 & n16715 ;
  assign n16719 = n16363 | n16718 ;
  assign n39376 = ~n16717 ;
  assign n16720 = n39376 & n16719 ;
  assign n39377 = ~n16720 ;
  assign n16721 = n3631 & n39377 ;
  assign n16722 = n173 | n16721 ;
  assign n39378 = ~n16722 ;
  assign n16762 = n39378 & n16748 ;
  assign n16763 = n16352 | n16762 ;
  assign n39379 = ~n16750 ;
  assign n16764 = n39379 & n16763 ;
  assign n39380 = ~n16764 ;
  assign n16765 = n174 & n39380 ;
  assign n16109 = n15673 & n39016 ;
  assign n39381 = ~n16076 ;
  assign n16110 = n39381 & n16109 ;
  assign n16344 = n16110 & n147 ;
  assign n16081 = n16075 | n16076 ;
  assign n39382 = ~n16081 ;
  assign n16380 = n39382 & n147 ;
  assign n16381 = n15673 | n16380 ;
  assign n39383 = ~n16344 ;
  assign n16382 = n39383 & n16381 ;
  assign n16751 = n174 | n16750 ;
  assign n39384 = ~n16751 ;
  assign n16766 = n39384 & n16763 ;
  assign n16767 = n16382 | n16766 ;
  assign n39385 = ~n16765 ;
  assign n16768 = n39385 & n16767 ;
  assign n39386 = ~n16768 ;
  assign n16769 = n2753 & n39386 ;
  assign n39387 = ~n16096 ;
  assign n16106 = n15646 & n39387 ;
  assign n16107 = n39043 & n16106 ;
  assign n16323 = n16107 & n16322 ;
  assign n16108 = n16079 | n16096 ;
  assign n39388 = ~n16108 ;
  assign n16435 = n39388 & n147 ;
  assign n16436 = n15646 | n16435 ;
  assign n39389 = ~n16323 ;
  assign n16437 = n39389 & n16436 ;
  assign n16733 = n16719 & n39368 ;
  assign n16734 = n16609 | n16733 ;
  assign n39390 = ~n16721 ;
  assign n16735 = n39390 & n16734 ;
  assign n39391 = ~n16735 ;
  assign n16736 = n173 & n39391 ;
  assign n16737 = n39378 & n16734 ;
  assign n16738 = n16352 | n16737 ;
  assign n39392 = ~n16736 ;
  assign n16739 = n39392 & n16738 ;
  assign n39393 = ~n16739 ;
  assign n16740 = n174 & n39393 ;
  assign n16741 = n2753 | n16740 ;
  assign n39394 = ~n16741 ;
  assign n16780 = n39394 & n16767 ;
  assign n16781 = n16437 | n16780 ;
  assign n39395 = ~n16769 ;
  assign n16782 = n39395 & n16781 ;
  assign n39396 = ~n16782 ;
  assign n16783 = n176 & n39396 ;
  assign n16132 = n15719 & n39032 ;
  assign n39397 = ~n16100 ;
  assign n16133 = n39397 & n16132 ;
  assign n16357 = n16133 & n147 ;
  assign n16105 = n16099 | n16100 ;
  assign n39398 = ~n16105 ;
  assign n16396 = n39398 & n147 ;
  assign n16397 = n15719 | n16396 ;
  assign n39399 = ~n16357 ;
  assign n16398 = n39399 & n16397 ;
  assign n16770 = n2431 | n16769 ;
  assign n39400 = ~n16770 ;
  assign n16784 = n39400 & n16781 ;
  assign n16785 = n16398 | n16784 ;
  assign n39401 = ~n16783 ;
  assign n16786 = n39401 & n16785 ;
  assign n39402 = ~n16786 ;
  assign n16787 = n177 & n39402 ;
  assign n39403 = ~n16120 ;
  assign n16129 = n15813 & n39403 ;
  assign n16130 = n39059 & n16129 ;
  assign n16343 = n16130 & n147 ;
  assign n16131 = n16103 | n16120 ;
  assign n39404 = ~n16131 ;
  assign n16408 = n39404 & n147 ;
  assign n16409 = n15813 | n16408 ;
  assign n39405 = ~n16343 ;
  assign n16410 = n39405 & n16409 ;
  assign n16752 = n16738 & n39384 ;
  assign n16753 = n16382 | n16752 ;
  assign n39406 = ~n16740 ;
  assign n16754 = n39406 & n16753 ;
  assign n39407 = ~n16754 ;
  assign n16755 = n175 & n39407 ;
  assign n16756 = n39394 & n16753 ;
  assign n16757 = n16437 | n16756 ;
  assign n39408 = ~n16755 ;
  assign n16758 = n39408 & n16757 ;
  assign n39409 = ~n16758 ;
  assign n16759 = n2431 & n39409 ;
  assign n16760 = n177 | n16759 ;
  assign n39410 = ~n16760 ;
  assign n16790 = n39410 & n16785 ;
  assign n16791 = n16410 | n16790 ;
  assign n39411 = ~n16787 ;
  assign n16792 = n39411 & n16791 ;
  assign n39412 = ~n16792 ;
  assign n16793 = n178 & n39412 ;
  assign n16788 = n178 | n16787 ;
  assign n39413 = ~n16788 ;
  assign n16794 = n39413 & n16791 ;
  assign n16155 = n15811 & n39048 ;
  assign n39414 = ~n16124 ;
  assign n16156 = n39414 & n16155 ;
  assign n16841 = n16156 & n147 ;
  assign n16157 = n16124 | n16141 ;
  assign n39415 = ~n16157 ;
  assign n16842 = n39415 & n147 ;
  assign n16843 = n15811 | n16842 ;
  assign n39416 = ~n16841 ;
  assign n16844 = n39416 & n16843 ;
  assign n16845 = n16794 | n16844 ;
  assign n39417 = ~n16793 ;
  assign n16846 = n39417 & n16845 ;
  assign n39418 = ~n16846 ;
  assign n16847 = n1707 & n39418 ;
  assign n16154 = n16127 | n16143 ;
  assign n39419 = ~n16154 ;
  assign n16419 = n39419 & n147 ;
  assign n16420 = n15809 | n16419 ;
  assign n39420 = ~n16143 ;
  assign n16152 = n15809 & n39420 ;
  assign n16153 = n39075 & n16152 ;
  assign n16466 = n16153 & n147 ;
  assign n39421 = ~n16466 ;
  assign n16467 = n16420 & n39421 ;
  assign n16771 = n16757 & n39400 ;
  assign n16772 = n16398 | n16771 ;
  assign n39422 = ~n16759 ;
  assign n16773 = n39422 & n16772 ;
  assign n39423 = ~n16773 ;
  assign n16774 = n177 & n39423 ;
  assign n16775 = n39410 & n16772 ;
  assign n16776 = n16410 | n16775 ;
  assign n39424 = ~n16774 ;
  assign n16777 = n39424 & n16776 ;
  assign n39425 = ~n16777 ;
  assign n16778 = n178 & n39425 ;
  assign n16779 = n1707 | n16778 ;
  assign n39426 = ~n16779 ;
  assign n16849 = n39426 & n16845 ;
  assign n16850 = n16467 | n16849 ;
  assign n39427 = ~n16847 ;
  assign n16851 = n39427 & n16850 ;
  assign n39428 = ~n16851 ;
  assign n16852 = n180 & n39428 ;
  assign n16171 = n16147 | n16165 ;
  assign n39429 = ~n16171 ;
  assign n16345 = n39429 & n147 ;
  assign n16346 = n15627 | n16345 ;
  assign n16169 = n15627 & n39064 ;
  assign n39430 = ~n16147 ;
  assign n16170 = n39430 & n16169 ;
  assign n16349 = n16170 & n147 ;
  assign n39431 = ~n16349 ;
  assign n16350 = n16346 & n39431 ;
  assign n16848 = n1487 | n16847 ;
  assign n39432 = ~n16848 ;
  assign n16853 = n39432 & n16850 ;
  assign n16854 = n16350 | n16853 ;
  assign n39433 = ~n16852 ;
  assign n16855 = n39433 & n16854 ;
  assign n39434 = ~n16855 ;
  assign n16856 = n181 & n39434 ;
  assign n16789 = n16776 & n39413 ;
  assign n16864 = n16789 | n16844 ;
  assign n39435 = ~n16778 ;
  assign n16865 = n39435 & n16864 ;
  assign n39436 = ~n16865 ;
  assign n16866 = n179 & n39436 ;
  assign n16867 = n39426 & n16864 ;
  assign n16868 = n16467 | n16867 ;
  assign n39437 = ~n16866 ;
  assign n16869 = n39437 & n16868 ;
  assign n39438 = ~n16869 ;
  assign n16870 = n1487 & n39438 ;
  assign n16871 = n181 | n16870 ;
  assign n39439 = ~n16871 ;
  assign n16872 = n16854 & n39439 ;
  assign n39440 = ~n16167 ;
  assign n16215 = n39440 & n16199 ;
  assign n16216 = n39091 & n16215 ;
  assign n16881 = n16216 & n147 ;
  assign n16168 = n16150 | n16167 ;
  assign n39441 = ~n16168 ;
  assign n16431 = n39441 & n147 ;
  assign n16955 = n16199 | n16431 ;
  assign n39442 = ~n16881 ;
  assign n16956 = n39442 & n16955 ;
  assign n16974 = n16872 | n16956 ;
  assign n39443 = ~n16856 ;
  assign n16975 = n39443 & n16974 ;
  assign n39444 = ~n16975 ;
  assign n16976 = n182 & n39444 ;
  assign n16204 = n15768 & n39080 ;
  assign n39445 = ~n16220 ;
  assign n16949 = n16204 & n39445 ;
  assign n16950 = n147 & n16949 ;
  assign n16951 = n16219 | n16220 ;
  assign n39446 = ~n16951 ;
  assign n16952 = n147 & n39446 ;
  assign n16953 = n15768 | n16952 ;
  assign n39447 = ~n16950 ;
  assign n16954 = n39447 & n16953 ;
  assign n16857 = n182 | n16856 ;
  assign n39448 = ~n16857 ;
  assign n16977 = n39448 & n16974 ;
  assign n16978 = n16954 | n16977 ;
  assign n39449 = ~n16976 ;
  assign n16979 = n39449 & n16978 ;
  assign n39450 = ~n16979 ;
  assign n16980 = n996 & n39450 ;
  assign n39451 = ~n16235 ;
  assign n16942 = n15771 & n39451 ;
  assign n16943 = n39107 & n16942 ;
  assign n16944 = n147 & n16943 ;
  assign n16945 = n16223 | n16235 ;
  assign n39452 = ~n16945 ;
  assign n16946 = n147 & n39452 ;
  assign n16947 = n15771 | n16946 ;
  assign n39453 = ~n16944 ;
  assign n16948 = n39453 & n16947 ;
  assign n16876 = n39432 & n16868 ;
  assign n16877 = n16350 | n16876 ;
  assign n39454 = ~n16870 ;
  assign n16878 = n39454 & n16877 ;
  assign n39455 = ~n16878 ;
  assign n16879 = n181 & n39455 ;
  assign n16880 = n39439 & n16877 ;
  assign n16957 = n16880 | n16956 ;
  assign n39456 = ~n16879 ;
  assign n16958 = n39456 & n16957 ;
  assign n39457 = ~n16958 ;
  assign n16959 = n182 & n39457 ;
  assign n16960 = n183 | n16959 ;
  assign n39458 = ~n16960 ;
  assign n16992 = n39458 & n16978 ;
  assign n16993 = n16948 | n16992 ;
  assign n39459 = ~n16980 ;
  assign n16994 = n39459 & n16993 ;
  assign n39460 = ~n16994 ;
  assign n16995 = n184 & n39460 ;
  assign n16214 = n15773 & n39096 ;
  assign n39461 = ~n16239 ;
  assign n16936 = n16214 & n39461 ;
  assign n16937 = n147 & n16936 ;
  assign n16938 = n16238 | n16239 ;
  assign n39462 = ~n16938 ;
  assign n16939 = n147 & n39462 ;
  assign n16940 = n15773 | n16939 ;
  assign n39463 = ~n16937 ;
  assign n16941 = n39463 & n16940 ;
  assign n16981 = n838 | n16980 ;
  assign n39464 = ~n16981 ;
  assign n16996 = n39464 & n16993 ;
  assign n16997 = n16941 | n16996 ;
  assign n39465 = ~n16995 ;
  assign n16998 = n39465 & n16997 ;
  assign n39466 = ~n16998 ;
  assign n16999 = n185 & n39466 ;
  assign n39467 = ~n16254 ;
  assign n16929 = n15779 & n39467 ;
  assign n16930 = n39123 & n16929 ;
  assign n16931 = n16322 & n16930 ;
  assign n16932 = n16242 | n16254 ;
  assign n39468 = ~n16932 ;
  assign n16933 = n147 & n39468 ;
  assign n16934 = n15779 | n16933 ;
  assign n39469 = ~n16931 ;
  assign n16935 = n39469 & n16934 ;
  assign n16962 = n39448 & n16957 ;
  assign n16963 = n16954 | n16962 ;
  assign n39470 = ~n16959 ;
  assign n16964 = n39470 & n16963 ;
  assign n39471 = ~n16964 ;
  assign n16965 = n183 & n39471 ;
  assign n16966 = n39458 & n16963 ;
  assign n16967 = n16948 | n16966 ;
  assign n39472 = ~n16965 ;
  assign n16968 = n39472 & n16967 ;
  assign n39473 = ~n16968 ;
  assign n16969 = n838 & n39473 ;
  assign n16970 = n185 | n16969 ;
  assign n39474 = ~n16970 ;
  assign n17011 = n39474 & n16997 ;
  assign n17012 = n16935 | n17011 ;
  assign n39475 = ~n16999 ;
  assign n17013 = n39475 & n17012 ;
  assign n39476 = ~n17013 ;
  assign n17014 = n186 & n39476 ;
  assign n16234 = n15781 & n39112 ;
  assign n39477 = ~n16258 ;
  assign n16923 = n16234 & n39477 ;
  assign n16924 = n147 & n16923 ;
  assign n16925 = n16257 | n16258 ;
  assign n39478 = ~n16925 ;
  assign n16926 = n147 & n39478 ;
  assign n16927 = n15781 | n16926 ;
  assign n39479 = ~n16924 ;
  assign n16928 = n39479 & n16927 ;
  assign n17000 = n186 | n16999 ;
  assign n39480 = ~n17000 ;
  assign n17015 = n39480 & n17012 ;
  assign n17016 = n16928 | n17015 ;
  assign n39481 = ~n17014 ;
  assign n17017 = n39481 & n17016 ;
  assign n39482 = ~n17017 ;
  assign n17018 = n528 & n39482 ;
  assign n39483 = ~n16273 ;
  assign n16916 = n15784 & n39483 ;
  assign n16917 = n39139 & n16916 ;
  assign n16918 = n147 & n16917 ;
  assign n16919 = n16261 | n16273 ;
  assign n39484 = ~n16919 ;
  assign n16920 = n147 & n39484 ;
  assign n16921 = n15784 | n16920 ;
  assign n39485 = ~n16918 ;
  assign n16922 = n39485 & n16921 ;
  assign n16982 = n16967 & n39464 ;
  assign n16983 = n16941 | n16982 ;
  assign n39486 = ~n16969 ;
  assign n16984 = n39486 & n16983 ;
  assign n39487 = ~n16984 ;
  assign n16985 = n185 & n39487 ;
  assign n16986 = n39474 & n16983 ;
  assign n16987 = n16935 | n16986 ;
  assign n39488 = ~n16985 ;
  assign n16988 = n39488 & n16987 ;
  assign n39489 = ~n16988 ;
  assign n16989 = n186 & n39489 ;
  assign n16990 = n528 | n16989 ;
  assign n39490 = ~n16990 ;
  assign n17030 = n39490 & n17016 ;
  assign n17031 = n16922 | n17030 ;
  assign n39491 = ~n17018 ;
  assign n17032 = n39491 & n17031 ;
  assign n39492 = ~n17032 ;
  assign n17033 = n188 & n39492 ;
  assign n16253 = n15786 & n39128 ;
  assign n39493 = ~n16277 ;
  assign n16910 = n16253 & n39493 ;
  assign n16911 = n147 & n16910 ;
  assign n16912 = n16276 | n16277 ;
  assign n39494 = ~n16912 ;
  assign n16913 = n147 & n39494 ;
  assign n16914 = n15786 | n16913 ;
  assign n39495 = ~n16911 ;
  assign n16915 = n39495 & n16914 ;
  assign n17019 = n413 | n17018 ;
  assign n39496 = ~n17019 ;
  assign n17034 = n39496 & n17031 ;
  assign n17035 = n16915 | n17034 ;
  assign n39497 = ~n17033 ;
  assign n17036 = n39497 & n17035 ;
  assign n39498 = ~n17036 ;
  assign n17037 = n189 & n39498 ;
  assign n39499 = ~n16292 ;
  assign n16903 = n15790 & n39499 ;
  assign n16904 = n39155 & n16903 ;
  assign n16905 = n147 & n16904 ;
  assign n16906 = n16280 | n16292 ;
  assign n39500 = ~n16906 ;
  assign n16907 = n147 & n39500 ;
  assign n16908 = n15790 | n16907 ;
  assign n39501 = ~n16905 ;
  assign n16909 = n39501 & n16908 ;
  assign n17001 = n16987 & n39480 ;
  assign n17002 = n16928 | n17001 ;
  assign n39502 = ~n16989 ;
  assign n17003 = n39502 & n17002 ;
  assign n39503 = ~n17003 ;
  assign n17004 = n187 & n39503 ;
  assign n17005 = n39490 & n17002 ;
  assign n17006 = n16922 | n17005 ;
  assign n39504 = ~n17004 ;
  assign n17007 = n39504 & n17006 ;
  assign n39505 = ~n17007 ;
  assign n17008 = n413 & n39505 ;
  assign n17009 = n189 | n17008 ;
  assign n39506 = ~n17009 ;
  assign n17039 = n39506 & n17035 ;
  assign n17040 = n16909 | n17039 ;
  assign n39507 = ~n17037 ;
  assign n17041 = n39507 & n17040 ;
  assign n39508 = ~n17041 ;
  assign n17042 = n190 & n39508 ;
  assign n16272 = n15794 & n39144 ;
  assign n39509 = ~n16296 ;
  assign n16897 = n16272 & n39509 ;
  assign n16898 = n147 & n16897 ;
  assign n16899 = n16295 | n16296 ;
  assign n39510 = ~n16899 ;
  assign n16900 = n147 & n39510 ;
  assign n16901 = n15794 | n16900 ;
  assign n39511 = ~n16898 ;
  assign n16902 = n39511 & n16901 ;
  assign n17038 = n190 | n17037 ;
  assign n39512 = ~n17038 ;
  assign n17043 = n39512 & n17040 ;
  assign n17044 = n16902 | n17043 ;
  assign n39513 = ~n17042 ;
  assign n17047 = n39513 & n17044 ;
  assign n39514 = ~n17047 ;
  assign n17048 = n287 & n39514 ;
  assign n39515 = ~n16331 ;
  assign n16890 = n16197 & n39515 ;
  assign n16891 = n39165 & n16890 ;
  assign n16892 = n147 & n16891 ;
  assign n16893 = n16299 | n16331 ;
  assign n39516 = ~n16893 ;
  assign n16894 = n147 & n39516 ;
  assign n16895 = n16197 | n16894 ;
  assign n39517 = ~n16892 ;
  assign n16896 = n39517 & n16895 ;
  assign n17020 = n17006 & n39496 ;
  assign n17021 = n16915 | n17020 ;
  assign n39518 = ~n17008 ;
  assign n17022 = n39518 & n17021 ;
  assign n39519 = ~n17022 ;
  assign n17023 = n189 & n39519 ;
  assign n17024 = n39506 & n17021 ;
  assign n17025 = n16909 | n17024 ;
  assign n39520 = ~n17023 ;
  assign n17026 = n39520 & n17025 ;
  assign n39521 = ~n17026 ;
  assign n17027 = n190 & n39521 ;
  assign n17028 = n287 | n17027 ;
  assign n39522 = ~n17028 ;
  assign n17045 = n39522 & n17044 ;
  assign n17052 = n16896 | n17045 ;
  assign n39523 = ~n17048 ;
  assign n17053 = n39523 & n17052 ;
  assign n17054 = n16887 | n17053 ;
  assign n17055 = n31336 & n17054 ;
  assign n16182 = n15618 | n16181 ;
  assign n39524 = ~n16182 ;
  assign n16188 = n39524 & n16185 ;
  assign n16189 = n39182 & n16188 ;
  assign n16314 = n16189 & n39183 ;
  assign n16315 = n39184 & n16314 ;
  assign n16320 = n192 & n16319 ;
  assign n39525 = ~n16186 ;
  assign n16425 = n39525 & n147 ;
  assign n39526 = ~n16425 ;
  assign n16426 = n16307 & n39526 ;
  assign n39527 = ~n16426 ;
  assign n16427 = n16320 & n39527 ;
  assign n16428 = n16315 | n16427 ;
  assign n17050 = n16886 & n39523 ;
  assign n17058 = n17050 & n17052 ;
  assign n17059 = n16428 | n17058 ;
  assign n146 = n17055 | n17059 ;
  assign n221 = x32 | x33 ;
  assign n222 = x34 | n221 ;
  assign n17146 = x34 & n146 ;
  assign n39528 = ~n17146 ;
  assign n17147 = n222 & n39528 ;
  assign n39529 = ~n17147 ;
  assign n17148 = n147 & n39529 ;
  assign n15619 = n222 & n39181 ;
  assign n15802 = n15619 & n39182 ;
  assign n16317 = n15802 & n39183 ;
  assign n16318 = n39184 & n16317 ;
  assign n17212 = n16318 & n39528 ;
  assign n39530 = ~n218 ;
  assign n17080 = n39530 & n146 ;
  assign n39531 = ~x34 ;
  assign n17214 = n39531 & n146 ;
  assign n39532 = ~n17214 ;
  assign n17215 = x35 & n39532 ;
  assign n17216 = n17080 | n17215 ;
  assign n17217 = n17212 | n17216 ;
  assign n39533 = ~n17148 ;
  assign n17219 = n39533 & n17217 ;
  assign n39534 = ~n17219 ;
  assign n17220 = n15807 & n39534 ;
  assign n223 = n39531 & n221 ;
  assign n39535 = ~n146 ;
  assign n17206 = x34 & n39535 ;
  assign n17207 = n223 | n17206 ;
  assign n39536 = ~n17207 ;
  assign n17208 = n16322 & n39536 ;
  assign n17209 = n15807 | n17208 ;
  assign n39537 = ~n17209 ;
  assign n17218 = n39537 & n17217 ;
  assign n39538 = ~n16315 ;
  assign n16330 = n39538 & n16322 ;
  assign n39539 = ~n16427 ;
  assign n16429 = n16330 & n39539 ;
  assign n39540 = ~n17058 ;
  assign n17226 = n16429 & n39540 ;
  assign n39541 = ~n17055 ;
  assign n17227 = n39541 & n17226 ;
  assign n17228 = n17080 | n17227 ;
  assign n17229 = x36 & n17228 ;
  assign n17230 = x36 | n17227 ;
  assign n17231 = n17080 | n17230 ;
  assign n39542 = ~n17229 ;
  assign n17232 = n39542 & n17231 ;
  assign n17233 = n17218 | n17232 ;
  assign n39543 = ~n17220 ;
  assign n17234 = n39543 & n17233 ;
  assign n39544 = ~n17234 ;
  assign n17235 = n149 & n39544 ;
  assign n16418 = n16329 | n16417 ;
  assign n39545 = ~n16418 ;
  assign n17138 = n39545 & n146 ;
  assign n17139 = n16470 | n17138 ;
  assign n16471 = n39545 & n16470 ;
  assign n17210 = n16471 & n146 ;
  assign n39546 = ~n17210 ;
  assign n17211 = n17139 & n39546 ;
  assign n17221 = n149 | n17220 ;
  assign n39547 = ~n17221 ;
  assign n17238 = n39547 & n17233 ;
  assign n17239 = n17211 | n17238 ;
  assign n39548 = ~n17235 ;
  assign n17240 = n39548 & n17239 ;
  assign n39549 = ~n17240 ;
  assign n17241 = n150 & n39549 ;
  assign n39550 = ~n16482 ;
  assign n16489 = n16406 & n39550 ;
  assign n39551 = ~n16491 ;
  assign n16502 = n16489 & n39551 ;
  assign n17102 = n16502 & n146 ;
  assign n16503 = n16482 | n16491 ;
  assign n39552 = ~n16503 ;
  assign n17116 = n39552 & n146 ;
  assign n17117 = n16406 | n17116 ;
  assign n39553 = ~n17102 ;
  assign n17118 = n39553 & n17117 ;
  assign n17236 = n150 | n17235 ;
  assign n39554 = ~n17236 ;
  assign n17242 = n39554 & n17239 ;
  assign n17243 = n17118 | n17242 ;
  assign n39555 = ~n17241 ;
  assign n17244 = n39555 & n17243 ;
  assign n39556 = ~n17244 ;
  assign n17245 = n13662 & n39556 ;
  assign n16501 = n16479 | n16493 ;
  assign n39557 = ~n16501 ;
  assign n17108 = n39557 & n146 ;
  assign n17109 = n16439 | n17108 ;
  assign n16480 = n16439 & n39196 ;
  assign n39558 = ~n16493 ;
  assign n16500 = n16480 & n39558 ;
  assign n17204 = n16500 & n146 ;
  assign n39559 = ~n17204 ;
  assign n17205 = n17109 & n39559 ;
  assign n17222 = n148 & n39534 ;
  assign n17149 = n148 | n17148 ;
  assign n39560 = ~n17149 ;
  assign n17225 = n39560 & n17217 ;
  assign n17254 = n17225 | n17232 ;
  assign n39561 = ~n17222 ;
  assign n17255 = n39561 & n17254 ;
  assign n39562 = ~n17255 ;
  assign n17256 = n149 & n39562 ;
  assign n17257 = n39547 & n17254 ;
  assign n17258 = n17211 | n17257 ;
  assign n39563 = ~n17256 ;
  assign n17259 = n39563 & n17258 ;
  assign n39564 = ~n17259 ;
  assign n17260 = n150 & n39564 ;
  assign n17261 = n151 | n17260 ;
  assign n39565 = ~n17261 ;
  assign n17262 = n17243 & n39565 ;
  assign n17263 = n17205 | n17262 ;
  assign n39566 = ~n17245 ;
  assign n17264 = n39566 & n17263 ;
  assign n39567 = ~n17264 ;
  assign n17265 = n152 & n39567 ;
  assign n16499 = n16496 | n16498 ;
  assign n39568 = ~n16499 ;
  assign n17100 = n39568 & n146 ;
  assign n17101 = n16508 | n17100 ;
  assign n39569 = ~n16498 ;
  assign n16591 = n39569 & n16508 ;
  assign n16592 = n39203 & n16591 ;
  assign n17134 = n16592 & n146 ;
  assign n39570 = ~n17134 ;
  assign n17135 = n17101 & n39570 ;
  assign n17246 = n152 | n17245 ;
  assign n39571 = ~n17246 ;
  assign n17266 = n39571 & n17263 ;
  assign n17267 = n17135 | n17266 ;
  assign n39572 = ~n17265 ;
  assign n17268 = n39572 & n17267 ;
  assign n39573 = ~n17268 ;
  assign n17269 = n153 & n39573 ;
  assign n16517 = n16511 | n16512 ;
  assign n39574 = ~n16517 ;
  assign n17103 = n39574 & n146 ;
  assign n17104 = n16445 | n17103 ;
  assign n16535 = n16445 & n39230 ;
  assign n39575 = ~n16512 ;
  assign n16536 = n39575 & n16535 ;
  assign n17144 = n16536 & n146 ;
  assign n39576 = ~n17144 ;
  assign n17145 = n17104 & n39576 ;
  assign n17277 = n39554 & n17258 ;
  assign n17278 = n17118 | n17277 ;
  assign n39577 = ~n17260 ;
  assign n17279 = n39577 & n17278 ;
  assign n39578 = ~n17279 ;
  assign n17280 = n151 & n39578 ;
  assign n17281 = n39565 & n17278 ;
  assign n17282 = n17205 | n17281 ;
  assign n39579 = ~n17280 ;
  assign n17283 = n39579 & n17282 ;
  assign n39580 = ~n17283 ;
  assign n17284 = n13079 & n39580 ;
  assign n17285 = n153 | n17284 ;
  assign n39581 = ~n17285 ;
  assign n17286 = n17267 & n39581 ;
  assign n17287 = n17145 | n17286 ;
  assign n39582 = ~n17269 ;
  assign n17288 = n39582 & n17287 ;
  assign n39583 = ~n17288 ;
  assign n17289 = n154 & n39583 ;
  assign n39584 = ~n16522 ;
  assign n16532 = n16442 & n39584 ;
  assign n16533 = n39219 & n16532 ;
  assign n17143 = n16533 & n146 ;
  assign n16534 = n16515 | n16522 ;
  assign n39585 = ~n16534 ;
  assign n17153 = n39585 & n146 ;
  assign n17154 = n16442 | n17153 ;
  assign n39586 = ~n17143 ;
  assign n17155 = n39586 & n17154 ;
  assign n17270 = n154 | n17269 ;
  assign n39587 = ~n17270 ;
  assign n17290 = n39587 & n17287 ;
  assign n17291 = n17155 | n17290 ;
  assign n39588 = ~n17289 ;
  assign n17292 = n39588 & n17291 ;
  assign n39589 = ~n17292 ;
  assign n17293 = n11067 & n39589 ;
  assign n16559 = n16465 & n39246 ;
  assign n39590 = ~n16526 ;
  assign n16560 = n39590 & n16559 ;
  assign n17128 = n16560 & n146 ;
  assign n16531 = n16525 | n16526 ;
  assign n39591 = ~n16531 ;
  assign n17160 = n39591 & n146 ;
  assign n17161 = n16465 | n17160 ;
  assign n39592 = ~n17128 ;
  assign n17162 = n39592 & n17161 ;
  assign n17301 = n39571 & n17282 ;
  assign n17302 = n17135 | n17301 ;
  assign n39593 = ~n17284 ;
  assign n17303 = n39593 & n17302 ;
  assign n39594 = ~n17303 ;
  assign n17304 = n153 & n39594 ;
  assign n17305 = n39581 & n17302 ;
  assign n17306 = n17145 | n17305 ;
  assign n39595 = ~n17304 ;
  assign n17307 = n39595 & n17306 ;
  assign n39596 = ~n17307 ;
  assign n17308 = n154 & n39596 ;
  assign n17309 = n11067 | n17308 ;
  assign n39597 = ~n17309 ;
  assign n17310 = n17291 & n39597 ;
  assign n17311 = n17162 | n17310 ;
  assign n39598 = ~n17293 ;
  assign n17312 = n39598 & n17311 ;
  assign n39599 = ~n17312 ;
  assign n17313 = n156 & n39599 ;
  assign n16558 = n16529 | n16546 ;
  assign n39600 = ~n16558 ;
  assign n17168 = n39600 & n146 ;
  assign n17169 = n16457 | n17168 ;
  assign n39601 = ~n16546 ;
  assign n16556 = n16457 & n39601 ;
  assign n16557 = n39235 & n16556 ;
  assign n17172 = n16557 & n146 ;
  assign n39602 = ~n17172 ;
  assign n17173 = n17169 & n39602 ;
  assign n17295 = n10657 | n17293 ;
  assign n39603 = ~n17295 ;
  assign n17314 = n39603 & n17311 ;
  assign n17315 = n17173 | n17314 ;
  assign n39604 = ~n17313 ;
  assign n17316 = n39604 & n17315 ;
  assign n39605 = ~n17316 ;
  assign n17317 = n157 & n39605 ;
  assign n16555 = n16549 | n16550 ;
  assign n39606 = ~n16555 ;
  assign n17110 = n39606 & n146 ;
  assign n17111 = n16462 | n17110 ;
  assign n16579 = n16462 & n39259 ;
  assign n39607 = ~n16550 ;
  assign n16580 = n39607 & n16579 ;
  assign n17179 = n16580 & n146 ;
  assign n39608 = ~n17179 ;
  assign n17180 = n17111 & n39608 ;
  assign n17325 = n39587 & n17306 ;
  assign n17326 = n17155 | n17325 ;
  assign n39609 = ~n17308 ;
  assign n17327 = n39609 & n17326 ;
  assign n39610 = ~n17327 ;
  assign n17328 = n155 & n39610 ;
  assign n17329 = n39597 & n17326 ;
  assign n17330 = n17162 | n17329 ;
  assign n39611 = ~n17328 ;
  assign n17331 = n39611 & n17330 ;
  assign n39612 = ~n17331 ;
  assign n17332 = n10657 & n39612 ;
  assign n17333 = n157 | n17332 ;
  assign n39613 = ~n17333 ;
  assign n17334 = n17315 & n39613 ;
  assign n17335 = n17180 | n17334 ;
  assign n39614 = ~n17317 ;
  assign n17336 = n39614 & n17335 ;
  assign n39615 = ~n17336 ;
  assign n17337 = n158 & n39615 ;
  assign n16578 = n16553 | n16570 ;
  assign n39616 = ~n16578 ;
  assign n17122 = n39616 & n146 ;
  assign n17123 = n16423 | n17122 ;
  assign n39617 = ~n16570 ;
  assign n16576 = n16423 & n39617 ;
  assign n16577 = n39251 & n16576 ;
  assign n17124 = n16577 & n146 ;
  assign n39618 = ~n17124 ;
  assign n17125 = n17123 & n39618 ;
  assign n17318 = n158 | n17317 ;
  assign n39619 = ~n17318 ;
  assign n17338 = n39619 & n17335 ;
  assign n17339 = n17125 | n17338 ;
  assign n39620 = ~n17337 ;
  assign n17340 = n39620 & n17339 ;
  assign n39621 = ~n17340 ;
  assign n17341 = n8857 & n39621 ;
  assign n16575 = n16573 | n16574 ;
  assign n39622 = ~n16575 ;
  assign n17166 = n39622 & n146 ;
  assign n17167 = n16595 | n17166 ;
  assign n16602 = n39278 & n16595 ;
  assign n39623 = ~n16574 ;
  assign n16603 = n39623 & n16602 ;
  assign n17174 = n16603 & n146 ;
  assign n39624 = ~n17174 ;
  assign n17175 = n17167 & n39624 ;
  assign n17349 = n39603 & n17330 ;
  assign n17350 = n17173 | n17349 ;
  assign n39625 = ~n17332 ;
  assign n17351 = n39625 & n17350 ;
  assign n39626 = ~n17351 ;
  assign n17352 = n157 & n39626 ;
  assign n17353 = n39613 & n17350 ;
  assign n17354 = n17180 | n17353 ;
  assign n39627 = ~n17352 ;
  assign n17355 = n39627 & n17354 ;
  assign n39628 = ~n17355 ;
  assign n17356 = n158 & n39628 ;
  assign n17357 = n8857 | n17356 ;
  assign n39629 = ~n17357 ;
  assign n17358 = n17339 & n39629 ;
  assign n17359 = n17175 | n17358 ;
  assign n39630 = ~n17341 ;
  assign n17360 = n39630 & n17359 ;
  assign n39631 = ~n17360 ;
  assign n17361 = n160 & n39631 ;
  assign n39632 = ~n16600 ;
  assign n16628 = n39632 & n16612 ;
  assign n16629 = n39267 & n16628 ;
  assign n17067 = n16629 & n146 ;
  assign n16601 = n16598 | n16600 ;
  assign n39633 = ~n16601 ;
  assign n17150 = n39633 & n146 ;
  assign n17151 = n16612 | n17150 ;
  assign n39634 = ~n17067 ;
  assign n17152 = n39634 & n17151 ;
  assign n17342 = n160 | n17341 ;
  assign n39635 = ~n17342 ;
  assign n17362 = n39635 & n17359 ;
  assign n17363 = n17152 | n17362 ;
  assign n39636 = ~n17361 ;
  assign n17364 = n39636 & n17363 ;
  assign n39637 = ~n17364 ;
  assign n17365 = n161 & n39637 ;
  assign n16617 = n16505 & n39294 ;
  assign n39638 = ~n16633 ;
  assign n16839 = n16617 & n39638 ;
  assign n17084 = n16839 & n146 ;
  assign n16840 = n16632 | n16633 ;
  assign n39639 = ~n16840 ;
  assign n17156 = n39639 & n146 ;
  assign n17157 = n16505 | n17156 ;
  assign n39640 = ~n17084 ;
  assign n17158 = n39640 & n17157 ;
  assign n17373 = n39619 & n17354 ;
  assign n17374 = n17125 | n17373 ;
  assign n39641 = ~n17356 ;
  assign n17375 = n39641 & n17374 ;
  assign n39642 = ~n17375 ;
  assign n17376 = n159 & n39642 ;
  assign n17377 = n39629 & n17374 ;
  assign n17378 = n17175 | n17377 ;
  assign n39643 = ~n17376 ;
  assign n17379 = n39643 & n17378 ;
  assign n39644 = ~n17379 ;
  assign n17380 = n8534 & n39644 ;
  assign n17381 = n161 | n17380 ;
  assign n39645 = ~n17381 ;
  assign n17382 = n17363 & n39645 ;
  assign n17383 = n17158 | n17382 ;
  assign n39646 = ~n17365 ;
  assign n17384 = n39646 & n17383 ;
  assign n39647 = ~n17384 ;
  assign n17385 = n162 & n39647 ;
  assign n39648 = ~n16648 ;
  assign n16836 = n16453 & n39648 ;
  assign n16837 = n39283 & n16836 ;
  assign n17093 = n16837 & n146 ;
  assign n16838 = n16636 | n16648 ;
  assign n39649 = ~n16838 ;
  assign n17097 = n39649 & n146 ;
  assign n17098 = n16453 | n17097 ;
  assign n39650 = ~n17093 ;
  assign n17099 = n39650 & n17098 ;
  assign n17366 = n162 | n17365 ;
  assign n39651 = ~n17366 ;
  assign n17386 = n39651 & n17383 ;
  assign n17387 = n17099 | n17386 ;
  assign n39652 = ~n17385 ;
  assign n17388 = n39652 & n17387 ;
  assign n39653 = ~n17388 ;
  assign n17389 = n6889 & n39653 ;
  assign n16627 = n16459 & n39310 ;
  assign n39654 = ~n16652 ;
  assign n16834 = n16627 & n39654 ;
  assign n17092 = n16834 & n146 ;
  assign n16835 = n16651 | n16652 ;
  assign n39655 = ~n16835 ;
  assign n17163 = n39655 & n146 ;
  assign n17164 = n16459 | n17163 ;
  assign n39656 = ~n17092 ;
  assign n17165 = n39656 & n17164 ;
  assign n17397 = n39635 & n17378 ;
  assign n17398 = n17152 | n17397 ;
  assign n39657 = ~n17380 ;
  assign n17399 = n39657 & n17398 ;
  assign n39658 = ~n17399 ;
  assign n17400 = n161 & n39658 ;
  assign n17401 = n39645 & n17398 ;
  assign n17402 = n17158 | n17401 ;
  assign n39659 = ~n17400 ;
  assign n17403 = n39659 & n17402 ;
  assign n39660 = ~n17403 ;
  assign n17404 = n162 & n39660 ;
  assign n17405 = n6889 | n17404 ;
  assign n39661 = ~n17405 ;
  assign n17406 = n17387 & n39661 ;
  assign n17407 = n17165 | n17406 ;
  assign n39662 = ~n17389 ;
  assign n17408 = n39662 & n17407 ;
  assign n39663 = ~n17408 ;
  assign n17409 = n164 & n39663 ;
  assign n39664 = ~n16667 ;
  assign n16831 = n16433 & n39664 ;
  assign n16832 = n39299 & n16831 ;
  assign n17088 = n16832 & n146 ;
  assign n16833 = n16655 | n16667 ;
  assign n39665 = ~n16833 ;
  assign n17089 = n39665 & n146 ;
  assign n17090 = n16433 | n17089 ;
  assign n39666 = ~n17088 ;
  assign n17091 = n39666 & n17090 ;
  assign n17390 = n6600 | n17389 ;
  assign n39667 = ~n17390 ;
  assign n17410 = n39667 & n17407 ;
  assign n17411 = n17091 | n17410 ;
  assign n39668 = ~n17409 ;
  assign n17412 = n39668 & n17411 ;
  assign n39669 = ~n17412 ;
  assign n17413 = n165 & n39669 ;
  assign n16647 = n16390 & n39326 ;
  assign n39670 = ~n16671 ;
  assign n16829 = n16647 & n39670 ;
  assign n17083 = n16829 & n146 ;
  assign n16830 = n16670 | n16671 ;
  assign n39671 = ~n16830 ;
  assign n17085 = n39671 & n146 ;
  assign n17086 = n16390 | n17085 ;
  assign n39672 = ~n17083 ;
  assign n17087 = n39672 & n17086 ;
  assign n17421 = n39651 & n17402 ;
  assign n17422 = n17099 | n17421 ;
  assign n39673 = ~n17404 ;
  assign n17423 = n39673 & n17422 ;
  assign n39674 = ~n17423 ;
  assign n17424 = n163 & n39674 ;
  assign n17425 = n39661 & n17422 ;
  assign n17426 = n17165 | n17425 ;
  assign n39675 = ~n17424 ;
  assign n17427 = n39675 & n17426 ;
  assign n39676 = ~n17427 ;
  assign n17428 = n6600 & n39676 ;
  assign n17429 = n165 | n17428 ;
  assign n39677 = ~n17429 ;
  assign n17430 = n17411 & n39677 ;
  assign n17431 = n17087 | n17430 ;
  assign n39678 = ~n17413 ;
  assign n17432 = n39678 & n17431 ;
  assign n39679 = ~n17432 ;
  assign n17433 = n166 & n39679 ;
  assign n39680 = ~n16686 ;
  assign n16826 = n16384 & n39680 ;
  assign n16827 = n39315 & n16826 ;
  assign n17076 = n16827 & n146 ;
  assign n16828 = n16674 | n16686 ;
  assign n39681 = ~n16828 ;
  assign n17113 = n39681 & n146 ;
  assign n17114 = n16384 | n17113 ;
  assign n39682 = ~n17076 ;
  assign n17115 = n39682 & n17114 ;
  assign n17414 = n166 | n17413 ;
  assign n39683 = ~n17414 ;
  assign n17434 = n39683 & n17431 ;
  assign n17435 = n17115 | n17434 ;
  assign n39684 = ~n17433 ;
  assign n17436 = n39684 & n17435 ;
  assign n39685 = ~n17436 ;
  assign n17437 = n5352 & n39685 ;
  assign n16825 = n16689 | n16690 ;
  assign n39686 = ~n16825 ;
  assign n17132 = n39686 & n146 ;
  assign n17133 = n16400 | n17132 ;
  assign n16666 = n16400 & n39342 ;
  assign n39687 = ~n16690 ;
  assign n16824 = n16666 & n39687 ;
  assign n17136 = n16824 & n146 ;
  assign n39688 = ~n17136 ;
  assign n17137 = n17133 & n39688 ;
  assign n17445 = n39667 & n17426 ;
  assign n17446 = n17091 | n17445 ;
  assign n39689 = ~n17428 ;
  assign n17447 = n39689 & n17446 ;
  assign n39690 = ~n17447 ;
  assign n17448 = n165 & n39690 ;
  assign n17449 = n39677 & n17446 ;
  assign n17450 = n17087 | n17449 ;
  assign n39691 = ~n17448 ;
  assign n17451 = n39691 & n17450 ;
  assign n39692 = ~n17451 ;
  assign n17452 = n166 & n39692 ;
  assign n17453 = n5352 | n17452 ;
  assign n39693 = ~n17453 ;
  assign n17454 = n17435 & n39693 ;
  assign n17455 = n17137 | n17454 ;
  assign n39694 = ~n17437 ;
  assign n17456 = n39694 & n17455 ;
  assign n39695 = ~n17456 ;
  assign n17457 = n168 & n39695 ;
  assign n39696 = ~n16705 ;
  assign n16821 = n16447 & n39696 ;
  assign n16822 = n39331 & n16821 ;
  assign n17066 = n16822 & n146 ;
  assign n16823 = n16693 | n16705 ;
  assign n39697 = ~n16823 ;
  assign n17129 = n39697 & n146 ;
  assign n17130 = n16447 | n17129 ;
  assign n39698 = ~n17066 ;
  assign n17131 = n39698 & n17130 ;
  assign n17438 = n4934 | n17437 ;
  assign n39699 = ~n17438 ;
  assign n17458 = n39699 & n17455 ;
  assign n17459 = n17131 | n17458 ;
  assign n39700 = ~n17457 ;
  assign n17460 = n39700 & n17459 ;
  assign n39701 = ~n17460 ;
  assign n17461 = n169 & n39701 ;
  assign n16820 = n16708 | n16709 ;
  assign n39702 = ~n16820 ;
  assign n17073 = n39702 & n146 ;
  assign n17074 = n16366 | n17073 ;
  assign n16685 = n16366 & n39358 ;
  assign n39703 = ~n16709 ;
  assign n16819 = n16685 & n39703 ;
  assign n17141 = n16819 & n146 ;
  assign n39704 = ~n17141 ;
  assign n17142 = n17074 & n39704 ;
  assign n17469 = n39683 & n17450 ;
  assign n17470 = n17115 | n17469 ;
  assign n39705 = ~n17452 ;
  assign n17471 = n39705 & n17470 ;
  assign n39706 = ~n17471 ;
  assign n17472 = n167 & n39706 ;
  assign n17473 = n39693 & n17470 ;
  assign n17474 = n17137 | n17473 ;
  assign n39707 = ~n17472 ;
  assign n17475 = n39707 & n17474 ;
  assign n39708 = ~n17475 ;
  assign n17476 = n4934 & n39708 ;
  assign n17477 = n169 | n17476 ;
  assign n39709 = ~n17477 ;
  assign n17478 = n17459 & n39709 ;
  assign n17479 = n17142 | n17478 ;
  assign n39710 = ~n17461 ;
  assign n17480 = n39710 & n17479 ;
  assign n39711 = ~n17480 ;
  assign n17481 = n170 & n39711 ;
  assign n39712 = ~n16724 ;
  assign n16816 = n16413 & n39712 ;
  assign n16817 = n39347 & n16816 ;
  assign n17112 = n16817 & n146 ;
  assign n16818 = n16712 | n16724 ;
  assign n39713 = ~n16818 ;
  assign n17119 = n39713 & n146 ;
  assign n17120 = n16413 | n17119 ;
  assign n39714 = ~n17112 ;
  assign n17121 = n39714 & n17120 ;
  assign n17462 = n170 | n17461 ;
  assign n39715 = ~n17462 ;
  assign n17482 = n39715 & n17479 ;
  assign n17483 = n17121 | n17482 ;
  assign n39716 = ~n17481 ;
  assign n17484 = n39716 & n17483 ;
  assign n39717 = ~n17484 ;
  assign n17485 = n3940 & n39717 ;
  assign n16815 = n16727 | n16728 ;
  assign n39718 = ~n16815 ;
  assign n17081 = n39718 & n146 ;
  assign n17082 = n16369 | n17081 ;
  assign n16704 = n16369 & n39374 ;
  assign n39719 = ~n16728 ;
  assign n16814 = n16704 & n39719 ;
  assign n17170 = n16814 & n146 ;
  assign n39720 = ~n17170 ;
  assign n17171 = n17082 & n39720 ;
  assign n17493 = n39699 & n17474 ;
  assign n17494 = n17131 | n17493 ;
  assign n39721 = ~n17476 ;
  assign n17495 = n39721 & n17494 ;
  assign n39722 = ~n17495 ;
  assign n17496 = n169 & n39722 ;
  assign n17497 = n39709 & n17494 ;
  assign n17498 = n17142 | n17497 ;
  assign n39723 = ~n17496 ;
  assign n17499 = n39723 & n17498 ;
  assign n39724 = ~n17499 ;
  assign n17500 = n170 & n39724 ;
  assign n17501 = n3940 | n17500 ;
  assign n39725 = ~n17501 ;
  assign n17502 = n17483 & n39725 ;
  assign n17503 = n17171 | n17502 ;
  assign n39726 = ~n17485 ;
  assign n17504 = n39726 & n17503 ;
  assign n39727 = ~n17504 ;
  assign n17505 = n172 & n39727 ;
  assign n39728 = ~n16743 ;
  assign n16811 = n16363 & n39728 ;
  assign n16812 = n39363 & n16811 ;
  assign n17075 = n16812 & n146 ;
  assign n16813 = n16731 | n16743 ;
  assign n39729 = ~n16813 ;
  assign n17077 = n39729 & n146 ;
  assign n17078 = n16363 | n17077 ;
  assign n39730 = ~n17075 ;
  assign n17079 = n39730 & n17078 ;
  assign n17487 = n3631 | n17485 ;
  assign n39731 = ~n17487 ;
  assign n17506 = n39731 & n17503 ;
  assign n17507 = n17079 | n17506 ;
  assign n39732 = ~n17505 ;
  assign n17508 = n39732 & n17507 ;
  assign n39733 = ~n17508 ;
  assign n17509 = n173 & n39733 ;
  assign n16723 = n16609 & n39390 ;
  assign n39734 = ~n16747 ;
  assign n16809 = n16723 & n39734 ;
  assign n17069 = n16809 & n146 ;
  assign n16810 = n16746 | n16747 ;
  assign n39735 = ~n16810 ;
  assign n17070 = n39735 & n146 ;
  assign n17071 = n16609 | n17070 ;
  assign n39736 = ~n17069 ;
  assign n17072 = n39736 & n17071 ;
  assign n17517 = n39715 & n17498 ;
  assign n17518 = n17121 | n17517 ;
  assign n39737 = ~n17500 ;
  assign n17519 = n39737 & n17518 ;
  assign n39738 = ~n17519 ;
  assign n17520 = n171 & n39738 ;
  assign n17521 = n39725 & n17518 ;
  assign n17522 = n17171 | n17521 ;
  assign n39739 = ~n17520 ;
  assign n17523 = n39739 & n17522 ;
  assign n39740 = ~n17523 ;
  assign n17524 = n3631 & n39740 ;
  assign n17525 = n173 | n17524 ;
  assign n39741 = ~n17525 ;
  assign n17526 = n17507 & n39741 ;
  assign n17527 = n17072 | n17526 ;
  assign n39742 = ~n17509 ;
  assign n17528 = n39742 & n17527 ;
  assign n39743 = ~n17528 ;
  assign n17529 = n174 & n39743 ;
  assign n39744 = ~n16762 ;
  assign n16806 = n16352 & n39744 ;
  assign n16807 = n39379 & n16806 ;
  assign n17159 = n16807 & n146 ;
  assign n16808 = n16750 | n16762 ;
  assign n39745 = ~n16808 ;
  assign n17176 = n39745 & n146 ;
  assign n17177 = n16352 | n17176 ;
  assign n39746 = ~n17159 ;
  assign n17178 = n39746 & n17177 ;
  assign n17510 = n174 | n17509 ;
  assign n39747 = ~n17510 ;
  assign n17530 = n39747 & n17527 ;
  assign n17533 = n17178 | n17530 ;
  assign n39748 = ~n17529 ;
  assign n17534 = n39748 & n17533 ;
  assign n39749 = ~n17534 ;
  assign n17535 = n2753 & n39749 ;
  assign n16742 = n16382 & n39406 ;
  assign n39750 = ~n16766 ;
  assign n16804 = n16742 & n39750 ;
  assign n17065 = n16804 & n146 ;
  assign n16805 = n16765 | n16766 ;
  assign n39751 = ~n16805 ;
  assign n17105 = n39751 & n146 ;
  assign n17106 = n16382 | n17105 ;
  assign n39752 = ~n17065 ;
  assign n17107 = n39752 & n17106 ;
  assign n17541 = n39731 & n17522 ;
  assign n17542 = n17079 | n17541 ;
  assign n39753 = ~n17524 ;
  assign n17543 = n39753 & n17542 ;
  assign n39754 = ~n17543 ;
  assign n17544 = n173 & n39754 ;
  assign n17545 = n39741 & n17542 ;
  assign n17546 = n17072 | n17545 ;
  assign n39755 = ~n17544 ;
  assign n17547 = n39755 & n17546 ;
  assign n39756 = ~n17547 ;
  assign n17548 = n174 & n39756 ;
  assign n17549 = n2753 | n17548 ;
  assign n39757 = ~n17549 ;
  assign n17550 = n17533 & n39757 ;
  assign n17551 = n17107 | n17550 ;
  assign n39758 = ~n17535 ;
  assign n17552 = n39758 & n17551 ;
  assign n39759 = ~n17552 ;
  assign n17553 = n176 & n39759 ;
  assign n39760 = ~n16780 ;
  assign n16801 = n16437 & n39760 ;
  assign n16802 = n39395 & n16801 ;
  assign n17061 = n16802 & n146 ;
  assign n16803 = n16769 | n16780 ;
  assign n39761 = ~n16803 ;
  assign n17062 = n39761 & n146 ;
  assign n17063 = n16437 | n17062 ;
  assign n39762 = ~n17061 ;
  assign n17064 = n39762 & n17063 ;
  assign n17536 = n2431 | n17535 ;
  assign n39763 = ~n17536 ;
  assign n17554 = n39763 & n17551 ;
  assign n17555 = n17064 | n17554 ;
  assign n39764 = ~n17553 ;
  assign n17556 = n39764 & n17555 ;
  assign n39765 = ~n17556 ;
  assign n17557 = n177 & n39765 ;
  assign n16800 = n16783 | n16784 ;
  assign n39766 = ~n16800 ;
  assign n17181 = n39766 & n146 ;
  assign n17182 = n16398 | n17181 ;
  assign n16761 = n16398 & n39422 ;
  assign n39767 = ~n16784 ;
  assign n16799 = n16761 & n39767 ;
  assign n17183 = n16799 & n146 ;
  assign n39768 = ~n17183 ;
  assign n17184 = n17182 & n39768 ;
  assign n17565 = n39747 & n17546 ;
  assign n17566 = n17178 | n17565 ;
  assign n39769 = ~n17548 ;
  assign n17567 = n39769 & n17566 ;
  assign n39770 = ~n17567 ;
  assign n17568 = n175 & n39770 ;
  assign n17569 = n39757 & n17566 ;
  assign n17570 = n17107 | n17569 ;
  assign n39771 = ~n17568 ;
  assign n17571 = n39771 & n17570 ;
  assign n39772 = ~n17571 ;
  assign n17572 = n2431 & n39772 ;
  assign n17573 = n177 | n17572 ;
  assign n39773 = ~n17573 ;
  assign n17574 = n17555 & n39773 ;
  assign n17575 = n17184 | n17574 ;
  assign n39774 = ~n17557 ;
  assign n17576 = n39774 & n17575 ;
  assign n39775 = ~n17576 ;
  assign n17577 = n178 & n39775 ;
  assign n16798 = n16787 | n16790 ;
  assign n39776 = ~n16798 ;
  assign n17185 = n39776 & n146 ;
  assign n17186 = n16410 | n17185 ;
  assign n39777 = ~n16790 ;
  assign n16796 = n16410 & n39777 ;
  assign n16797 = n39411 & n16796 ;
  assign n17187 = n16797 & n146 ;
  assign n39778 = ~n17187 ;
  assign n17188 = n17186 & n39778 ;
  assign n17558 = n178 | n17557 ;
  assign n39779 = ~n17558 ;
  assign n17578 = n39779 & n17575 ;
  assign n17579 = n17188 | n17578 ;
  assign n39780 = ~n17577 ;
  assign n17580 = n39780 & n17579 ;
  assign n39781 = ~n17580 ;
  assign n17581 = n1707 & n39781 ;
  assign n16862 = n39435 & n16844 ;
  assign n39782 = ~n16794 ;
  assign n16863 = n39782 & n16862 ;
  assign n17140 = n16863 & n146 ;
  assign n16795 = n16793 | n16794 ;
  assign n39783 = ~n16795 ;
  assign n17189 = n39783 & n146 ;
  assign n17190 = n16844 | n17189 ;
  assign n39784 = ~n17140 ;
  assign n17191 = n39784 & n17190 ;
  assign n17589 = n39763 & n17570 ;
  assign n17590 = n17064 | n17589 ;
  assign n39785 = ~n17572 ;
  assign n17591 = n39785 & n17590 ;
  assign n39786 = ~n17591 ;
  assign n17592 = n177 & n39786 ;
  assign n17593 = n39773 & n17590 ;
  assign n17594 = n17184 | n17593 ;
  assign n39787 = ~n17592 ;
  assign n17595 = n39787 & n17594 ;
  assign n39788 = ~n17595 ;
  assign n17596 = n178 & n39788 ;
  assign n17597 = n1707 | n17596 ;
  assign n39789 = ~n17597 ;
  assign n17598 = n17579 & n39789 ;
  assign n17599 = n17191 | n17598 ;
  assign n39790 = ~n17581 ;
  assign n17600 = n39790 & n17599 ;
  assign n39791 = ~n17600 ;
  assign n17601 = n180 & n39791 ;
  assign n39792 = ~n16849 ;
  assign n16859 = n16467 & n39792 ;
  assign n16860 = n39427 & n16859 ;
  assign n17068 = n16860 & n146 ;
  assign n16861 = n16847 | n16849 ;
  assign n39793 = ~n16861 ;
  assign n17094 = n39793 & n146 ;
  assign n17095 = n16467 | n17094 ;
  assign n39794 = ~n17068 ;
  assign n17096 = n39794 & n17095 ;
  assign n17583 = n1487 | n17581 ;
  assign n39795 = ~n17583 ;
  assign n17602 = n39795 & n17599 ;
  assign n17603 = n17096 | n17602 ;
  assign n39796 = ~n17601 ;
  assign n17604 = n39796 & n17603 ;
  assign n39797 = ~n17604 ;
  assign n17605 = n181 & n39797 ;
  assign n16858 = n16852 | n16853 ;
  assign n39798 = ~n16858 ;
  assign n17126 = n39798 & n146 ;
  assign n17127 = n16350 | n17126 ;
  assign n16874 = n16350 & n39454 ;
  assign n39799 = ~n16853 ;
  assign n16875 = n39799 & n16874 ;
  assign n17192 = n16875 & n146 ;
  assign n39800 = ~n17192 ;
  assign n17193 = n17127 & n39800 ;
  assign n17613 = n39779 & n17594 ;
  assign n17614 = n17188 | n17613 ;
  assign n39801 = ~n17596 ;
  assign n17615 = n39801 & n17614 ;
  assign n39802 = ~n17615 ;
  assign n17616 = n179 & n39802 ;
  assign n17617 = n39789 & n17614 ;
  assign n17618 = n17191 | n17617 ;
  assign n39803 = ~n17616 ;
  assign n17619 = n39803 & n17618 ;
  assign n39804 = ~n17619 ;
  assign n17620 = n1487 & n39804 ;
  assign n17621 = n181 | n17620 ;
  assign n39805 = ~n17621 ;
  assign n17622 = n17603 & n39805 ;
  assign n17623 = n17193 | n17622 ;
  assign n39806 = ~n17605 ;
  assign n17624 = n39806 & n17623 ;
  assign n39807 = ~n17624 ;
  assign n17625 = n182 & n39807 ;
  assign n17606 = n182 | n17605 ;
  assign n39808 = ~n17606 ;
  assign n17626 = n39808 & n17623 ;
  assign n39809 = ~n16872 ;
  assign n16972 = n39809 & n16956 ;
  assign n16973 = n39443 & n16972 ;
  assign n17195 = n16973 & n146 ;
  assign n16873 = n16856 | n16872 ;
  assign n39810 = ~n16873 ;
  assign n17194 = n39810 & n146 ;
  assign n17713 = n16956 | n17194 ;
  assign n39811 = ~n17195 ;
  assign n17714 = n39811 & n17713 ;
  assign n17715 = n17626 | n17714 ;
  assign n39812 = ~n17625 ;
  assign n17716 = n39812 & n17715 ;
  assign n39813 = ~n17716 ;
  assign n17717 = n996 & n39813 ;
  assign n16961 = n16954 & n39470 ;
  assign n39814 = ~n16977 ;
  assign n17707 = n16961 & n39814 ;
  assign n17708 = n146 & n17707 ;
  assign n17709 = n16976 | n16977 ;
  assign n39815 = ~n17709 ;
  assign n17710 = n146 & n39815 ;
  assign n17711 = n16954 | n17710 ;
  assign n39816 = ~n17708 ;
  assign n17712 = n39816 & n17711 ;
  assign n17630 = n39795 & n17618 ;
  assign n17631 = n17096 | n17630 ;
  assign n39817 = ~n17620 ;
  assign n17632 = n39817 & n17631 ;
  assign n39818 = ~n17632 ;
  assign n17633 = n181 & n39818 ;
  assign n17634 = n39805 & n17631 ;
  assign n17635 = n17193 | n17634 ;
  assign n39819 = ~n17633 ;
  assign n17636 = n39819 & n17635 ;
  assign n39820 = ~n17636 ;
  assign n17637 = n182 & n39820 ;
  assign n17638 = n183 | n17637 ;
  assign n39821 = ~n17638 ;
  assign n17720 = n39821 & n17715 ;
  assign n17721 = n17712 | n17720 ;
  assign n39822 = ~n17717 ;
  assign n17722 = n39822 & n17721 ;
  assign n39823 = ~n17722 ;
  assign n17723 = n184 & n39823 ;
  assign n39824 = ~n16992 ;
  assign n17700 = n16948 & n39824 ;
  assign n17701 = n39459 & n17700 ;
  assign n17702 = n146 & n17701 ;
  assign n17703 = n16980 | n16992 ;
  assign n39825 = ~n17703 ;
  assign n17704 = n146 & n39825 ;
  assign n17705 = n16948 | n17704 ;
  assign n39826 = ~n17702 ;
  assign n17706 = n39826 & n17705 ;
  assign n17718 = n838 | n17717 ;
  assign n39827 = ~n17718 ;
  assign n17724 = n39827 & n17721 ;
  assign n17725 = n17706 | n17724 ;
  assign n39828 = ~n17723 ;
  assign n17726 = n39828 & n17725 ;
  assign n39829 = ~n17726 ;
  assign n17727 = n185 & n39829 ;
  assign n16971 = n16941 & n39486 ;
  assign n39830 = ~n16996 ;
  assign n17694 = n16971 & n39830 ;
  assign n17695 = n146 & n17694 ;
  assign n17696 = n16995 | n16996 ;
  assign n39831 = ~n17696 ;
  assign n17697 = n146 & n39831 ;
  assign n17698 = n16941 | n17697 ;
  assign n39832 = ~n17695 ;
  assign n17699 = n39832 & n17698 ;
  assign n17640 = n39808 & n17635 ;
  assign n17736 = n17640 | n17714 ;
  assign n39833 = ~n17637 ;
  assign n17737 = n39833 & n17736 ;
  assign n39834 = ~n17737 ;
  assign n17738 = n183 & n39834 ;
  assign n17739 = n39821 & n17736 ;
  assign n17740 = n17712 | n17739 ;
  assign n39835 = ~n17738 ;
  assign n17741 = n39835 & n17740 ;
  assign n39836 = ~n17741 ;
  assign n17742 = n838 & n39836 ;
  assign n17743 = n185 | n17742 ;
  assign n39837 = ~n17743 ;
  assign n17744 = n17725 & n39837 ;
  assign n17745 = n17699 | n17744 ;
  assign n39838 = ~n17727 ;
  assign n17746 = n39838 & n17745 ;
  assign n39839 = ~n17746 ;
  assign n17747 = n186 & n39839 ;
  assign n39840 = ~n17011 ;
  assign n17687 = n16935 & n39840 ;
  assign n17688 = n39475 & n17687 ;
  assign n17689 = n146 & n17688 ;
  assign n17690 = n16999 | n17011 ;
  assign n39841 = ~n17690 ;
  assign n17691 = n146 & n39841 ;
  assign n17692 = n16935 | n17691 ;
  assign n39842 = ~n17689 ;
  assign n17693 = n39842 & n17692 ;
  assign n17728 = n186 | n17727 ;
  assign n39843 = ~n17728 ;
  assign n17748 = n39843 & n17745 ;
  assign n17749 = n17693 | n17748 ;
  assign n39844 = ~n17747 ;
  assign n17750 = n39844 & n17749 ;
  assign n39845 = ~n17750 ;
  assign n17751 = n528 & n39845 ;
  assign n16991 = n16928 & n39502 ;
  assign n39846 = ~n17015 ;
  assign n17681 = n16991 & n39846 ;
  assign n17682 = n146 & n17681 ;
  assign n17683 = n17014 | n17015 ;
  assign n39847 = ~n17683 ;
  assign n17684 = n146 & n39847 ;
  assign n17685 = n16928 | n17684 ;
  assign n39848 = ~n17682 ;
  assign n17686 = n39848 & n17685 ;
  assign n17759 = n39827 & n17740 ;
  assign n17760 = n17706 | n17759 ;
  assign n39849 = ~n17742 ;
  assign n17761 = n39849 & n17760 ;
  assign n39850 = ~n17761 ;
  assign n17762 = n185 & n39850 ;
  assign n17763 = n39837 & n17760 ;
  assign n17764 = n17699 | n17763 ;
  assign n39851 = ~n17762 ;
  assign n17765 = n39851 & n17764 ;
  assign n39852 = ~n17765 ;
  assign n17766 = n186 & n39852 ;
  assign n17767 = n528 | n17766 ;
  assign n39853 = ~n17767 ;
  assign n17768 = n17749 & n39853 ;
  assign n17769 = n17686 | n17768 ;
  assign n39854 = ~n17751 ;
  assign n17770 = n39854 & n17769 ;
  assign n39855 = ~n17770 ;
  assign n17771 = n188 & n39855 ;
  assign n39856 = ~n17030 ;
  assign n17674 = n16922 & n39856 ;
  assign n17675 = n39491 & n17674 ;
  assign n17676 = n146 & n17675 ;
  assign n17677 = n17018 | n17030 ;
  assign n39857 = ~n17677 ;
  assign n17678 = n146 & n39857 ;
  assign n17679 = n16922 | n17678 ;
  assign n39858 = ~n17676 ;
  assign n17680 = n39858 & n17679 ;
  assign n17752 = n413 | n17751 ;
  assign n39859 = ~n17752 ;
  assign n17772 = n39859 & n17769 ;
  assign n17773 = n17680 | n17772 ;
  assign n39860 = ~n17771 ;
  assign n17774 = n39860 & n17773 ;
  assign n39861 = ~n17774 ;
  assign n17775 = n189 & n39861 ;
  assign n17010 = n16915 & n39518 ;
  assign n39862 = ~n17034 ;
  assign n17668 = n17010 & n39862 ;
  assign n17669 = n146 & n17668 ;
  assign n17670 = n17033 | n17034 ;
  assign n39863 = ~n17670 ;
  assign n17671 = n146 & n39863 ;
  assign n17672 = n16915 | n17671 ;
  assign n39864 = ~n17669 ;
  assign n17673 = n39864 & n17672 ;
  assign n17783 = n39843 & n17764 ;
  assign n17784 = n17693 | n17783 ;
  assign n39865 = ~n17766 ;
  assign n17785 = n39865 & n17784 ;
  assign n39866 = ~n17785 ;
  assign n17786 = n187 & n39866 ;
  assign n17787 = n39853 & n17784 ;
  assign n17788 = n17686 | n17787 ;
  assign n39867 = ~n17786 ;
  assign n17789 = n39867 & n17788 ;
  assign n39868 = ~n17789 ;
  assign n17790 = n413 & n39868 ;
  assign n17791 = n189 | n17790 ;
  assign n39869 = ~n17791 ;
  assign n17792 = n17773 & n39869 ;
  assign n17793 = n17673 | n17792 ;
  assign n39870 = ~n17775 ;
  assign n17794 = n39870 & n17793 ;
  assign n39871 = ~n17794 ;
  assign n17795 = n190 & n39871 ;
  assign n39872 = ~n17039 ;
  assign n17661 = n16909 & n39872 ;
  assign n17662 = n39507 & n17661 ;
  assign n17663 = n146 & n17662 ;
  assign n17664 = n17037 | n17039 ;
  assign n39873 = ~n17664 ;
  assign n17665 = n146 & n39873 ;
  assign n17666 = n16909 | n17665 ;
  assign n39874 = ~n17663 ;
  assign n17667 = n39874 & n17666 ;
  assign n17776 = n190 | n17775 ;
  assign n39875 = ~n17776 ;
  assign n17796 = n39875 & n17793 ;
  assign n39876 = ~n17796 ;
  assign n17802 = n17667 & n39876 ;
  assign n39877 = ~n17795 ;
  assign n17803 = n39877 & n17802 ;
  assign n39878 = ~n17045 ;
  assign n17046 = n16896 & n39878 ;
  assign n17049 = n17046 & n39523 ;
  assign n17196 = n17049 & n146 ;
  assign n17051 = n17045 | n17048 ;
  assign n39879 = ~n17051 ;
  assign n17197 = n39879 & n146 ;
  assign n17198 = n16896 | n17197 ;
  assign n39880 = ~n17196 ;
  assign n17199 = n39880 & n17198 ;
  assign n17056 = n16886 | n17053 ;
  assign n39881 = ~n17056 ;
  assign n17203 = n39881 & n146 ;
  assign n17641 = n17058 | n17203 ;
  assign n17642 = n17199 | n17641 ;
  assign n17797 = n17667 | n17796 ;
  assign n17798 = n39877 & n17797 ;
  assign n39882 = ~n17798 ;
  assign n17799 = n287 & n39882 ;
  assign n39883 = ~n17027 ;
  assign n17029 = n16902 & n39883 ;
  assign n39884 = ~n17043 ;
  assign n17655 = n17029 & n39884 ;
  assign n17656 = n146 & n17655 ;
  assign n17657 = n17042 | n17043 ;
  assign n39885 = ~n17657 ;
  assign n17658 = n146 & n39885 ;
  assign n17659 = n16902 | n17658 ;
  assign n39886 = ~n17656 ;
  assign n17660 = n39886 & n17659 ;
  assign n17807 = n39859 & n17788 ;
  assign n17808 = n17680 | n17807 ;
  assign n39887 = ~n17790 ;
  assign n17809 = n39887 & n17808 ;
  assign n39888 = ~n17809 ;
  assign n17810 = n189 & n39888 ;
  assign n17811 = n39869 & n17808 ;
  assign n17812 = n17673 | n17811 ;
  assign n39889 = ~n17810 ;
  assign n17813 = n39889 & n17812 ;
  assign n39890 = ~n17813 ;
  assign n17814 = n190 & n39890 ;
  assign n17815 = n287 | n17814 ;
  assign n39891 = ~n17815 ;
  assign n17816 = n17797 & n39891 ;
  assign n17819 = n17660 | n17816 ;
  assign n39892 = ~n17799 ;
  assign n17820 = n39892 & n17819 ;
  assign n17823 = n17642 | n17820 ;
  assign n17824 = n31336 & n17823 ;
  assign n17057 = n192 & n17056 ;
  assign n39893 = ~n16886 ;
  assign n17200 = n39893 & n146 ;
  assign n39894 = ~n17200 ;
  assign n17201 = n17053 & n39894 ;
  assign n39895 = ~n17201 ;
  assign n17202 = n17057 & n39895 ;
  assign n16375 = n16315 | n16374 ;
  assign n39896 = ~n16375 ;
  assign n16888 = n39896 & n16885 ;
  assign n16889 = n39539 & n16888 ;
  assign n17643 = n16889 & n39540 ;
  assign n17644 = n39541 & n17643 ;
  assign n17645 = n17202 | n17644 ;
  assign n17800 = n17199 & n39892 ;
  assign n17825 = n17800 & n17819 ;
  assign n17826 = n17645 | n17825 ;
  assign n145 = n17824 | n17826 ;
  assign n17885 = n17803 & n145 ;
  assign n18483 = n17796 | n17814 ;
  assign n39897 = ~n18483 ;
  assign n18484 = n145 & n39897 ;
  assign n18485 = n17667 | n18484 ;
  assign n39898 = ~n17885 ;
  assign n18486 = n39898 & n18485 ;
  assign n224 = x30 | x31 ;
  assign n225 = x32 | n224 ;
  assign n17849 = x32 & n145 ;
  assign n39899 = ~n17849 ;
  assign n17930 = n225 & n39899 ;
  assign n39900 = ~n17930 ;
  assign n17931 = n146 & n39900 ;
  assign n16316 = n225 & n39538 ;
  assign n16430 = n16316 & n39539 ;
  assign n17653 = n16430 & n39540 ;
  assign n17654 = n39541 & n17653 ;
  assign n17850 = n17654 & n39899 ;
  assign n39901 = ~n221 ;
  assign n17915 = n39901 & n145 ;
  assign n39902 = ~x32 ;
  assign n18018 = n39902 & n145 ;
  assign n39903 = ~n18018 ;
  assign n18019 = x33 & n39903 ;
  assign n18020 = n17915 | n18019 ;
  assign n18022 = n17850 | n18020 ;
  assign n39904 = ~n17931 ;
  assign n18023 = n39904 & n18022 ;
  assign n39905 = ~n18023 ;
  assign n18024 = n16322 & n39905 ;
  assign n226 = n39902 & n224 ;
  assign n39906 = ~n145 ;
  assign n18009 = x32 & n39906 ;
  assign n18010 = n226 | n18009 ;
  assign n39907 = ~n18010 ;
  assign n18011 = n146 & n39907 ;
  assign n18012 = n16322 | n18011 ;
  assign n39908 = ~n18012 ;
  assign n18027 = n39908 & n18022 ;
  assign n39909 = ~n17644 ;
  assign n17646 = n146 & n39909 ;
  assign n39910 = ~n17202 ;
  assign n17647 = n39910 & n17646 ;
  assign n39911 = ~n17825 ;
  assign n18030 = n17647 & n39911 ;
  assign n39912 = ~n17824 ;
  assign n18031 = n39912 & n18030 ;
  assign n18032 = n17915 | n18031 ;
  assign n18033 = x34 & n18032 ;
  assign n18034 = x34 | n18031 ;
  assign n18035 = n17915 | n18034 ;
  assign n39913 = ~n18033 ;
  assign n18036 = n39913 & n18035 ;
  assign n18037 = n18027 | n18036 ;
  assign n39914 = ~n18024 ;
  assign n18038 = n39914 & n18037 ;
  assign n39915 = ~n18038 ;
  assign n18039 = n15807 & n39915 ;
  assign n17213 = n17208 | n17212 ;
  assign n39916 = ~n17213 ;
  assign n17875 = n39916 & n145 ;
  assign n17876 = n17216 | n17875 ;
  assign n17224 = n39916 & n17216 ;
  assign n17920 = n17224 & n145 ;
  assign n39917 = ~n17920 ;
  assign n17921 = n17876 & n39917 ;
  assign n18025 = n15807 | n18024 ;
  assign n39918 = ~n18025 ;
  assign n18042 = n39918 & n18037 ;
  assign n18043 = n17921 | n18042 ;
  assign n39919 = ~n18039 ;
  assign n18044 = n39919 & n18043 ;
  assign n39920 = ~n18044 ;
  assign n18045 = n149 & n39920 ;
  assign n17223 = n17218 | n17222 ;
  assign n39921 = ~n17223 ;
  assign n17934 = n39921 & n145 ;
  assign n17935 = n17232 | n17934 ;
  assign n39922 = ~n17218 ;
  assign n17252 = n39922 & n17232 ;
  assign n17253 = n39543 & n17252 ;
  assign n18013 = n17253 & n145 ;
  assign n39923 = ~n18013 ;
  assign n18014 = n17935 & n39923 ;
  assign n18040 = n149 | n18039 ;
  assign n39924 = ~n18040 ;
  assign n18046 = n39924 & n18043 ;
  assign n18047 = n18014 | n18046 ;
  assign n39925 = ~n18045 ;
  assign n18048 = n39925 & n18047 ;
  assign n39926 = ~n18048 ;
  assign n18049 = n150 & n39926 ;
  assign n17251 = n17235 | n17238 ;
  assign n39927 = ~n17251 ;
  assign n17899 = n39927 & n145 ;
  assign n17900 = n17211 | n17899 ;
  assign n17237 = n17211 & n39548 ;
  assign n39928 = ~n17238 ;
  assign n17250 = n17237 & n39928 ;
  assign n18016 = n17250 & n145 ;
  assign n39929 = ~n18016 ;
  assign n18017 = n17900 & n39929 ;
  assign n18026 = n147 & n39905 ;
  assign n17932 = n147 | n17931 ;
  assign n39930 = ~n17932 ;
  assign n18029 = n39930 & n18022 ;
  assign n18059 = n18029 | n18036 ;
  assign n39931 = ~n18026 ;
  assign n18060 = n39931 & n18059 ;
  assign n39932 = ~n18060 ;
  assign n18061 = n148 & n39932 ;
  assign n18062 = n39918 & n18059 ;
  assign n18063 = n17921 | n18062 ;
  assign n39933 = ~n18061 ;
  assign n18064 = n39933 & n18063 ;
  assign n39934 = ~n18064 ;
  assign n18065 = n149 & n39934 ;
  assign n18066 = n150 | n18065 ;
  assign n39935 = ~n18066 ;
  assign n18067 = n18047 & n39935 ;
  assign n18068 = n18017 | n18067 ;
  assign n39936 = ~n18049 ;
  assign n18069 = n39936 & n18068 ;
  assign n39937 = ~n18069 ;
  assign n18070 = n151 & n39937 ;
  assign n17276 = n17242 | n17260 ;
  assign n39938 = ~n17276 ;
  assign n17889 = n39938 & n145 ;
  assign n17890 = n17118 | n17889 ;
  assign n39939 = ~n17242 ;
  assign n17248 = n17118 & n39939 ;
  assign n17249 = n39555 & n17248 ;
  assign n17911 = n17249 & n145 ;
  assign n39940 = ~n17911 ;
  assign n17912 = n17890 & n39940 ;
  assign n18050 = n151 | n18049 ;
  assign n39941 = ~n18050 ;
  assign n18071 = n39941 & n18068 ;
  assign n18072 = n17912 | n18071 ;
  assign n39942 = ~n18070 ;
  assign n18073 = n39942 & n18072 ;
  assign n39943 = ~n18073 ;
  assign n18074 = n13079 & n39943 ;
  assign n17275 = n17245 | n17262 ;
  assign n39944 = ~n17275 ;
  assign n17883 = n39944 & n145 ;
  assign n17884 = n17205 | n17883 ;
  assign n17247 = n17205 & n39566 ;
  assign n39945 = ~n17262 ;
  assign n17274 = n17247 & n39945 ;
  assign n17896 = n17274 & n145 ;
  assign n39946 = ~n17896 ;
  assign n17897 = n17884 & n39946 ;
  assign n18082 = n39924 & n18063 ;
  assign n18083 = n18014 | n18082 ;
  assign n39947 = ~n18065 ;
  assign n18084 = n39947 & n18083 ;
  assign n39948 = ~n18084 ;
  assign n18085 = n150 & n39948 ;
  assign n18086 = n39935 & n18083 ;
  assign n18087 = n18017 | n18086 ;
  assign n39949 = ~n18085 ;
  assign n18088 = n39949 & n18087 ;
  assign n39950 = ~n18088 ;
  assign n18089 = n13662 & n39950 ;
  assign n18090 = n152 | n18089 ;
  assign n39951 = ~n18090 ;
  assign n18091 = n18072 & n39951 ;
  assign n18092 = n17897 | n18091 ;
  assign n39952 = ~n18074 ;
  assign n18093 = n39952 & n18092 ;
  assign n39953 = ~n18093 ;
  assign n18094 = n153 & n39953 ;
  assign n17300 = n17266 | n17284 ;
  assign n39954 = ~n17300 ;
  assign n17905 = n39954 & n145 ;
  assign n17906 = n17135 | n17905 ;
  assign n39955 = ~n17266 ;
  assign n17272 = n17135 & n39955 ;
  assign n17273 = n39572 & n17272 ;
  assign n17936 = n17273 & n145 ;
  assign n39956 = ~n17936 ;
  assign n17937 = n17906 & n39956 ;
  assign n18075 = n153 | n18074 ;
  assign n39957 = ~n18075 ;
  assign n18095 = n39957 & n18092 ;
  assign n18096 = n17937 | n18095 ;
  assign n39958 = ~n18094 ;
  assign n18097 = n39958 & n18096 ;
  assign n39959 = ~n18097 ;
  assign n18098 = n154 & n39959 ;
  assign n17271 = n17145 & n39582 ;
  assign n39960 = ~n17286 ;
  assign n17298 = n17271 & n39960 ;
  assign n17891 = n17298 & n145 ;
  assign n17299 = n17269 | n17286 ;
  assign n39961 = ~n17299 ;
  assign n17922 = n39961 & n145 ;
  assign n17923 = n17145 | n17922 ;
  assign n39962 = ~n17891 ;
  assign n17924 = n39962 & n17923 ;
  assign n18106 = n39941 & n18087 ;
  assign n18107 = n17912 | n18106 ;
  assign n39963 = ~n18089 ;
  assign n18108 = n39963 & n18107 ;
  assign n39964 = ~n18108 ;
  assign n18109 = n152 & n39964 ;
  assign n18110 = n39951 & n18107 ;
  assign n18111 = n17897 | n18110 ;
  assign n39965 = ~n18109 ;
  assign n18112 = n39965 & n18111 ;
  assign n39966 = ~n18112 ;
  assign n18113 = n153 & n39966 ;
  assign n18114 = n154 | n18113 ;
  assign n39967 = ~n18114 ;
  assign n18115 = n18096 & n39967 ;
  assign n18116 = n17924 | n18115 ;
  assign n39968 = ~n18098 ;
  assign n18117 = n39968 & n18116 ;
  assign n39969 = ~n18117 ;
  assign n18118 = n155 & n39969 ;
  assign n17324 = n17290 | n17308 ;
  assign n39970 = ~n17324 ;
  assign n17938 = n39970 & n145 ;
  assign n17939 = n17155 | n17938 ;
  assign n39971 = ~n17290 ;
  assign n17296 = n17155 & n39971 ;
  assign n17297 = n39588 & n17296 ;
  assign n17942 = n17297 & n145 ;
  assign n39972 = ~n17942 ;
  assign n17943 = n17939 & n39972 ;
  assign n18099 = n11067 | n18098 ;
  assign n39973 = ~n18099 ;
  assign n18119 = n39973 & n18116 ;
  assign n18120 = n17943 | n18119 ;
  assign n39974 = ~n18118 ;
  assign n18121 = n39974 & n18120 ;
  assign n39975 = ~n18121 ;
  assign n18122 = n10657 & n39975 ;
  assign n17294 = n17162 & n39598 ;
  assign n39976 = ~n17310 ;
  assign n17322 = n17294 & n39976 ;
  assign n17886 = n17322 & n145 ;
  assign n17323 = n17293 | n17310 ;
  assign n39977 = ~n17323 ;
  assign n17944 = n39977 & n145 ;
  assign n17945 = n17162 | n17944 ;
  assign n39978 = ~n17886 ;
  assign n17946 = n39978 & n17945 ;
  assign n18130 = n39957 & n18111 ;
  assign n18131 = n17937 | n18130 ;
  assign n39979 = ~n18113 ;
  assign n18132 = n39979 & n18131 ;
  assign n39980 = ~n18132 ;
  assign n18133 = n154 & n39980 ;
  assign n18134 = n39967 & n18131 ;
  assign n18135 = n17924 | n18134 ;
  assign n39981 = ~n18133 ;
  assign n18136 = n39981 & n18135 ;
  assign n39982 = ~n18136 ;
  assign n18137 = n11067 & n39982 ;
  assign n18138 = n10657 | n18137 ;
  assign n39983 = ~n18138 ;
  assign n18139 = n18120 & n39983 ;
  assign n18140 = n17946 | n18139 ;
  assign n39984 = ~n18122 ;
  assign n18141 = n39984 & n18140 ;
  assign n39985 = ~n18141 ;
  assign n18142 = n157 & n39985 ;
  assign n39986 = ~n17314 ;
  assign n17320 = n17173 & n39986 ;
  assign n17321 = n39604 & n17320 ;
  assign n17902 = n17321 & n145 ;
  assign n17348 = n17314 | n17332 ;
  assign n39987 = ~n17348 ;
  assign n17947 = n39987 & n145 ;
  assign n17948 = n17173 | n17947 ;
  assign n39988 = ~n17902 ;
  assign n17949 = n39988 & n17948 ;
  assign n18123 = n157 | n18122 ;
  assign n39989 = ~n18123 ;
  assign n18143 = n39989 & n18140 ;
  assign n18144 = n17949 | n18143 ;
  assign n39990 = ~n18142 ;
  assign n18145 = n39990 & n18144 ;
  assign n39991 = ~n18145 ;
  assign n18146 = n158 & n39991 ;
  assign n17319 = n17180 & n39614 ;
  assign n39992 = ~n17334 ;
  assign n17346 = n17319 & n39992 ;
  assign n17901 = n17346 & n145 ;
  assign n17347 = n17317 | n17334 ;
  assign n39993 = ~n17347 ;
  assign n17927 = n39993 & n145 ;
  assign n17928 = n17180 | n17927 ;
  assign n39994 = ~n17901 ;
  assign n17929 = n39994 & n17928 ;
  assign n18154 = n39973 & n18135 ;
  assign n18155 = n17943 | n18154 ;
  assign n39995 = ~n18137 ;
  assign n18156 = n39995 & n18155 ;
  assign n39996 = ~n18156 ;
  assign n18157 = n156 & n39996 ;
  assign n18158 = n39983 & n18155 ;
  assign n18159 = n17946 | n18158 ;
  assign n39997 = ~n18157 ;
  assign n18160 = n39997 & n18159 ;
  assign n39998 = ~n18160 ;
  assign n18161 = n157 & n39998 ;
  assign n18162 = n158 | n18161 ;
  assign n39999 = ~n18162 ;
  assign n18163 = n18144 & n39999 ;
  assign n18164 = n17929 | n18163 ;
  assign n40000 = ~n18146 ;
  assign n18165 = n40000 & n18164 ;
  assign n40001 = ~n18165 ;
  assign n18166 = n159 & n40001 ;
  assign n40002 = ~n17338 ;
  assign n17344 = n17125 & n40002 ;
  assign n17345 = n39620 & n17344 ;
  assign n17898 = n17345 & n145 ;
  assign n17372 = n17338 | n17356 ;
  assign n40003 = ~n17372 ;
  assign n17954 = n40003 & n145 ;
  assign n17955 = n17125 | n17954 ;
  assign n40004 = ~n17898 ;
  assign n17956 = n40004 & n17955 ;
  assign n18147 = n8857 | n18146 ;
  assign n40005 = ~n18147 ;
  assign n18167 = n40005 & n18164 ;
  assign n18171 = n17956 | n18167 ;
  assign n40006 = ~n18166 ;
  assign n18172 = n40006 & n18171 ;
  assign n40007 = ~n18172 ;
  assign n18173 = n8534 & n40007 ;
  assign n17371 = n17341 | n17358 ;
  assign n40008 = ~n17371 ;
  assign n17916 = n40008 & n145 ;
  assign n17917 = n17175 | n17916 ;
  assign n17343 = n17175 & n39630 ;
  assign n40009 = ~n17358 ;
  assign n17370 = n17343 & n40009 ;
  assign n17925 = n17370 & n145 ;
  assign n40010 = ~n17925 ;
  assign n17926 = n17917 & n40010 ;
  assign n18178 = n39989 & n18159 ;
  assign n18179 = n17949 | n18178 ;
  assign n40011 = ~n18161 ;
  assign n18180 = n40011 & n18179 ;
  assign n40012 = ~n18180 ;
  assign n18181 = n158 & n40012 ;
  assign n18182 = n39999 & n18179 ;
  assign n18183 = n17929 | n18182 ;
  assign n40013 = ~n18181 ;
  assign n18184 = n40013 & n18183 ;
  assign n40014 = ~n18184 ;
  assign n18185 = n8857 & n40014 ;
  assign n18186 = n160 | n18185 ;
  assign n40015 = ~n18186 ;
  assign n18187 = n18171 & n40015 ;
  assign n18188 = n17926 | n18187 ;
  assign n40016 = ~n18173 ;
  assign n18189 = n40016 & n18188 ;
  assign n40017 = ~n18189 ;
  assign n18190 = n161 & n40017 ;
  assign n40018 = ~n17362 ;
  assign n17368 = n17152 & n40018 ;
  assign n17369 = n39636 & n17368 ;
  assign n17864 = n17369 & n145 ;
  assign n17396 = n17362 | n17380 ;
  assign n40019 = ~n17396 ;
  assign n17951 = n40019 & n145 ;
  assign n17952 = n17152 | n17951 ;
  assign n40020 = ~n17864 ;
  assign n17953 = n40020 & n17952 ;
  assign n18174 = n161 | n18173 ;
  assign n40021 = ~n18174 ;
  assign n18191 = n40021 & n18188 ;
  assign n18192 = n17953 | n18191 ;
  assign n40022 = ~n18190 ;
  assign n18193 = n40022 & n18192 ;
  assign n40023 = ~n18193 ;
  assign n18194 = n162 & n40023 ;
  assign n17367 = n17158 & n39646 ;
  assign n40024 = ~n17382 ;
  assign n17394 = n17367 & n40024 ;
  assign n17867 = n17394 & n145 ;
  assign n17395 = n17365 | n17382 ;
  assign n40025 = ~n17395 ;
  assign n17877 = n40025 & n145 ;
  assign n17878 = n17158 | n17877 ;
  assign n40026 = ~n17867 ;
  assign n17879 = n40026 & n17878 ;
  assign n18202 = n40005 & n18183 ;
  assign n18203 = n17956 | n18202 ;
  assign n40027 = ~n18185 ;
  assign n18204 = n40027 & n18203 ;
  assign n40028 = ~n18204 ;
  assign n18205 = n160 & n40028 ;
  assign n18206 = n40015 & n18203 ;
  assign n18207 = n17926 | n18206 ;
  assign n40029 = ~n18205 ;
  assign n18208 = n40029 & n18207 ;
  assign n40030 = ~n18208 ;
  assign n18209 = n161 & n40030 ;
  assign n18210 = n162 | n18209 ;
  assign n40031 = ~n18210 ;
  assign n18211 = n18192 & n40031 ;
  assign n18212 = n17879 | n18211 ;
  assign n40032 = ~n18194 ;
  assign n18213 = n40032 & n18212 ;
  assign n40033 = ~n18213 ;
  assign n18214 = n163 & n40033 ;
  assign n17420 = n17386 | n17404 ;
  assign n40034 = ~n17420 ;
  assign n17873 = n40034 & n145 ;
  assign n17874 = n17099 | n17873 ;
  assign n40035 = ~n17386 ;
  assign n17392 = n17099 & n40035 ;
  assign n17393 = n39652 & n17392 ;
  assign n17903 = n17393 & n145 ;
  assign n40036 = ~n17903 ;
  assign n17904 = n17874 & n40036 ;
  assign n18196 = n6889 | n18194 ;
  assign n40037 = ~n18196 ;
  assign n18215 = n40037 & n18212 ;
  assign n18216 = n17904 | n18215 ;
  assign n40038 = ~n18214 ;
  assign n18217 = n40038 & n18216 ;
  assign n40039 = ~n18217 ;
  assign n18218 = n6600 & n40039 ;
  assign n17419 = n17389 | n17406 ;
  assign n40040 = ~n17419 ;
  assign n17871 = n40040 & n145 ;
  assign n17872 = n17165 | n17871 ;
  assign n17391 = n17165 & n39662 ;
  assign n40041 = ~n17406 ;
  assign n17418 = n17391 & n40041 ;
  assign n17887 = n17418 & n145 ;
  assign n40042 = ~n17887 ;
  assign n17888 = n17872 & n40042 ;
  assign n18226 = n40021 & n18207 ;
  assign n18227 = n17953 | n18226 ;
  assign n40043 = ~n18209 ;
  assign n18228 = n40043 & n18227 ;
  assign n40044 = ~n18228 ;
  assign n18229 = n162 & n40044 ;
  assign n18230 = n40031 & n18227 ;
  assign n18231 = n17879 | n18230 ;
  assign n40045 = ~n18229 ;
  assign n18232 = n40045 & n18231 ;
  assign n40046 = ~n18232 ;
  assign n18233 = n6889 & n40046 ;
  assign n18234 = n6600 | n18233 ;
  assign n40047 = ~n18234 ;
  assign n18235 = n18216 & n40047 ;
  assign n18236 = n17888 | n18235 ;
  assign n40048 = ~n18218 ;
  assign n18237 = n40048 & n18236 ;
  assign n40049 = ~n18237 ;
  assign n18238 = n165 & n40049 ;
  assign n17444 = n17410 | n17428 ;
  assign n40050 = ~n17444 ;
  assign n17865 = n40050 & n145 ;
  assign n17866 = n17091 | n17865 ;
  assign n40051 = ~n17410 ;
  assign n17416 = n17091 & n40051 ;
  assign n17417 = n39668 & n17416 ;
  assign n17918 = n17417 & n145 ;
  assign n40052 = ~n17918 ;
  assign n17919 = n17866 & n40052 ;
  assign n18219 = n165 | n18218 ;
  assign n40053 = ~n18219 ;
  assign n18239 = n40053 & n18236 ;
  assign n18240 = n17919 | n18239 ;
  assign n40054 = ~n18238 ;
  assign n18241 = n40054 & n18240 ;
  assign n40055 = ~n18241 ;
  assign n18242 = n166 & n40055 ;
  assign n17443 = n17413 | n17430 ;
  assign n40056 = ~n17443 ;
  assign n17854 = n40056 & n145 ;
  assign n17855 = n17087 | n17854 ;
  assign n17415 = n17087 & n39678 ;
  assign n40057 = ~n17430 ;
  assign n17442 = n17415 & n40057 ;
  assign n17907 = n17442 & n145 ;
  assign n40058 = ~n17907 ;
  assign n17908 = n17855 & n40058 ;
  assign n18250 = n40037 & n18231 ;
  assign n18251 = n17904 | n18250 ;
  assign n40059 = ~n18233 ;
  assign n18252 = n40059 & n18251 ;
  assign n40060 = ~n18252 ;
  assign n18253 = n164 & n40060 ;
  assign n18254 = n40047 & n18251 ;
  assign n18255 = n17888 | n18254 ;
  assign n40061 = ~n18253 ;
  assign n18256 = n40061 & n18255 ;
  assign n40062 = ~n18256 ;
  assign n18257 = n165 & n40062 ;
  assign n18258 = n166 | n18257 ;
  assign n40063 = ~n18258 ;
  assign n18259 = n18240 & n40063 ;
  assign n18260 = n17908 | n18259 ;
  assign n40064 = ~n18242 ;
  assign n18261 = n40064 & n18260 ;
  assign n40065 = ~n18261 ;
  assign n18262 = n167 & n40065 ;
  assign n40066 = ~n17434 ;
  assign n17440 = n17115 & n40066 ;
  assign n17441 = n39684 & n17440 ;
  assign n17844 = n17441 & n145 ;
  assign n17468 = n17434 | n17452 ;
  assign n40067 = ~n17468 ;
  assign n17845 = n40067 & n145 ;
  assign n17846 = n17115 | n17845 ;
  assign n40068 = ~n17844 ;
  assign n17847 = n40068 & n17846 ;
  assign n18243 = n5352 | n18242 ;
  assign n40069 = ~n18243 ;
  assign n18263 = n40069 & n18260 ;
  assign n18264 = n17847 | n18263 ;
  assign n40070 = ~n18262 ;
  assign n18265 = n40070 & n18264 ;
  assign n40071 = ~n18265 ;
  assign n18266 = n4934 & n40071 ;
  assign n17439 = n17137 & n39694 ;
  assign n40072 = ~n17454 ;
  assign n17466 = n17439 & n40072 ;
  assign n17835 = n17466 & n145 ;
  assign n17467 = n17437 | n17454 ;
  assign n40073 = ~n17467 ;
  assign n17861 = n40073 & n145 ;
  assign n17862 = n17137 | n17861 ;
  assign n40074 = ~n17835 ;
  assign n17863 = n40074 & n17862 ;
  assign n18274 = n40053 & n18255 ;
  assign n18275 = n17919 | n18274 ;
  assign n40075 = ~n18257 ;
  assign n18276 = n40075 & n18275 ;
  assign n40076 = ~n18276 ;
  assign n18277 = n166 & n40076 ;
  assign n18278 = n40063 & n18275 ;
  assign n18279 = n17908 | n18278 ;
  assign n40077 = ~n18277 ;
  assign n18280 = n40077 & n18279 ;
  assign n40078 = ~n18280 ;
  assign n18281 = n5352 & n40078 ;
  assign n18282 = n4934 | n18281 ;
  assign n40079 = ~n18282 ;
  assign n18283 = n18264 & n40079 ;
  assign n18284 = n17863 | n18283 ;
  assign n40080 = ~n18266 ;
  assign n18285 = n40080 & n18284 ;
  assign n40081 = ~n18285 ;
  assign n18286 = n169 & n40081 ;
  assign n40082 = ~n17458 ;
  assign n17464 = n17131 & n40082 ;
  assign n17465 = n39700 & n17464 ;
  assign n17838 = n17465 & n145 ;
  assign n17492 = n17458 | n17476 ;
  assign n40083 = ~n17492 ;
  assign n17841 = n40083 & n145 ;
  assign n17842 = n17131 | n17841 ;
  assign n40084 = ~n17838 ;
  assign n17843 = n40084 & n17842 ;
  assign n18267 = n169 | n18266 ;
  assign n40085 = ~n18267 ;
  assign n18287 = n40085 & n18284 ;
  assign n18288 = n17843 | n18287 ;
  assign n40086 = ~n18286 ;
  assign n18289 = n40086 & n18288 ;
  assign n40087 = ~n18289 ;
  assign n18290 = n170 & n40087 ;
  assign n17463 = n17142 & n39710 ;
  assign n40088 = ~n17478 ;
  assign n17490 = n17463 & n40088 ;
  assign n17829 = n17490 & n145 ;
  assign n17491 = n17461 | n17478 ;
  assign n40089 = ~n17491 ;
  assign n17832 = n40089 & n145 ;
  assign n17833 = n17142 | n17832 ;
  assign n40090 = ~n17829 ;
  assign n17834 = n40090 & n17833 ;
  assign n18298 = n40069 & n18279 ;
  assign n18299 = n17847 | n18298 ;
  assign n40091 = ~n18281 ;
  assign n18300 = n40091 & n18299 ;
  assign n40092 = ~n18300 ;
  assign n18301 = n168 & n40092 ;
  assign n18302 = n40079 & n18299 ;
  assign n18303 = n17863 | n18302 ;
  assign n40093 = ~n18301 ;
  assign n18304 = n40093 & n18303 ;
  assign n40094 = ~n18304 ;
  assign n18305 = n169 & n40094 ;
  assign n18306 = n170 | n18305 ;
  assign n40095 = ~n18306 ;
  assign n18307 = n18288 & n40095 ;
  assign n18308 = n17834 | n18307 ;
  assign n40096 = ~n18290 ;
  assign n18309 = n40096 & n18308 ;
  assign n40097 = ~n18309 ;
  assign n18310 = n171 & n40097 ;
  assign n17516 = n17482 | n17500 ;
  assign n40098 = ~n17516 ;
  assign n17859 = n40098 & n145 ;
  assign n17860 = n17121 | n17859 ;
  assign n40099 = ~n17482 ;
  assign n17488 = n17121 & n40099 ;
  assign n17489 = n39716 & n17488 ;
  assign n17869 = n17489 & n145 ;
  assign n40100 = ~n17869 ;
  assign n17870 = n17860 & n40100 ;
  assign n18291 = n3940 | n18290 ;
  assign n40101 = ~n18291 ;
  assign n18311 = n40101 & n18308 ;
  assign n18312 = n17870 | n18311 ;
  assign n40102 = ~n18310 ;
  assign n18313 = n40102 & n18312 ;
  assign n40103 = ~n18313 ;
  assign n18314 = n3631 & n40103 ;
  assign n17515 = n17485 | n17502 ;
  assign n40104 = ~n17515 ;
  assign n17892 = n40104 & n145 ;
  assign n17893 = n17171 | n17892 ;
  assign n17486 = n17171 & n39726 ;
  assign n40105 = ~n17502 ;
  assign n17514 = n17486 & n40105 ;
  assign n17940 = n17514 & n145 ;
  assign n40106 = ~n17940 ;
  assign n17941 = n17893 & n40106 ;
  assign n18322 = n40085 & n18303 ;
  assign n18323 = n17843 | n18322 ;
  assign n40107 = ~n18305 ;
  assign n18324 = n40107 & n18323 ;
  assign n40108 = ~n18324 ;
  assign n18325 = n170 & n40108 ;
  assign n18326 = n40095 & n18323 ;
  assign n18327 = n17834 | n18326 ;
  assign n40109 = ~n18325 ;
  assign n18328 = n40109 & n18327 ;
  assign n40110 = ~n18328 ;
  assign n18329 = n3940 & n40110 ;
  assign n18330 = n3631 | n18329 ;
  assign n40111 = ~n18330 ;
  assign n18331 = n18312 & n40111 ;
  assign n18332 = n17941 | n18331 ;
  assign n40112 = ~n18314 ;
  assign n18333 = n40112 & n18332 ;
  assign n40113 = ~n18333 ;
  assign n18334 = n173 & n40113 ;
  assign n40114 = ~n17506 ;
  assign n17512 = n17079 & n40114 ;
  assign n17513 = n39732 & n17512 ;
  assign n17828 = n17513 & n145 ;
  assign n17540 = n17506 | n17524 ;
  assign n40115 = ~n17540 ;
  assign n17851 = n40115 & n145 ;
  assign n17852 = n17079 | n17851 ;
  assign n40116 = ~n17828 ;
  assign n17853 = n40116 & n17852 ;
  assign n18315 = n173 | n18314 ;
  assign n40117 = ~n18315 ;
  assign n18335 = n40117 & n18332 ;
  assign n18336 = n17853 | n18335 ;
  assign n40118 = ~n18334 ;
  assign n18337 = n40118 & n18336 ;
  assign n40119 = ~n18337 ;
  assign n18338 = n174 & n40119 ;
  assign n17511 = n17072 & n39742 ;
  assign n40120 = ~n17526 ;
  assign n17538 = n17511 & n40120 ;
  assign n17848 = n17538 & n145 ;
  assign n17539 = n17509 | n17526 ;
  assign n40121 = ~n17539 ;
  assign n17880 = n40121 & n145 ;
  assign n17881 = n17072 | n17880 ;
  assign n40122 = ~n17848 ;
  assign n17882 = n40122 & n17881 ;
  assign n18346 = n40101 & n18327 ;
  assign n18347 = n17870 | n18346 ;
  assign n40123 = ~n18329 ;
  assign n18348 = n40123 & n18347 ;
  assign n40124 = ~n18348 ;
  assign n18349 = n172 & n40124 ;
  assign n18350 = n40111 & n18347 ;
  assign n18351 = n17941 | n18350 ;
  assign n40125 = ~n18349 ;
  assign n18352 = n40125 & n18351 ;
  assign n40126 = ~n18352 ;
  assign n18353 = n173 & n40126 ;
  assign n18354 = n174 | n18353 ;
  assign n40127 = ~n18354 ;
  assign n18355 = n18336 & n40127 ;
  assign n18356 = n17882 | n18355 ;
  assign n40128 = ~n18338 ;
  assign n18357 = n40128 & n18356 ;
  assign n40129 = ~n18357 ;
  assign n18358 = n175 & n40129 ;
  assign n40130 = ~n17530 ;
  assign n17531 = n17178 & n40130 ;
  assign n17532 = n39748 & n17531 ;
  assign n17836 = n17532 & n145 ;
  assign n17564 = n17530 | n17548 ;
  assign n40131 = ~n17564 ;
  assign n17856 = n40131 & n145 ;
  assign n17857 = n17178 | n17856 ;
  assign n40132 = ~n17836 ;
  assign n17858 = n40132 & n17857 ;
  assign n18339 = n2753 | n18338 ;
  assign n40133 = ~n18339 ;
  assign n18359 = n40133 & n18356 ;
  assign n18360 = n17858 | n18359 ;
  assign n40134 = ~n18358 ;
  assign n18361 = n40134 & n18360 ;
  assign n40135 = ~n18361 ;
  assign n18362 = n2431 & n40135 ;
  assign n17563 = n17535 | n17550 ;
  assign n40136 = ~n17563 ;
  assign n17839 = n40136 & n145 ;
  assign n17840 = n17107 | n17839 ;
  assign n17537 = n17107 & n39758 ;
  assign n40137 = ~n17550 ;
  assign n17562 = n17537 & n40137 ;
  assign n17957 = n17562 & n145 ;
  assign n40138 = ~n17957 ;
  assign n17958 = n17840 & n40138 ;
  assign n18370 = n40117 & n18351 ;
  assign n18371 = n17853 | n18370 ;
  assign n40139 = ~n18353 ;
  assign n18372 = n40139 & n18371 ;
  assign n40140 = ~n18372 ;
  assign n18373 = n174 & n40140 ;
  assign n18374 = n40127 & n18371 ;
  assign n18375 = n17882 | n18374 ;
  assign n40141 = ~n18373 ;
  assign n18376 = n40141 & n18375 ;
  assign n40142 = ~n18376 ;
  assign n18377 = n2753 & n40142 ;
  assign n18378 = n2431 | n18377 ;
  assign n40143 = ~n18378 ;
  assign n18379 = n18360 & n40143 ;
  assign n18380 = n17958 | n18379 ;
  assign n40144 = ~n18362 ;
  assign n18381 = n40144 & n18380 ;
  assign n40145 = ~n18381 ;
  assign n18382 = n177 & n40145 ;
  assign n17588 = n17554 | n17572 ;
  assign n40146 = ~n17588 ;
  assign n17961 = n40146 & n145 ;
  assign n17962 = n17064 | n17961 ;
  assign n40147 = ~n17554 ;
  assign n17560 = n17064 & n40147 ;
  assign n17561 = n39764 & n17560 ;
  assign n17963 = n17561 & n145 ;
  assign n40148 = ~n17963 ;
  assign n17964 = n17962 & n40148 ;
  assign n18363 = n177 | n18362 ;
  assign n40149 = ~n18363 ;
  assign n18383 = n40149 & n18380 ;
  assign n18384 = n17964 | n18383 ;
  assign n40150 = ~n18382 ;
  assign n18385 = n40150 & n18384 ;
  assign n40151 = ~n18385 ;
  assign n18386 = n178 & n40151 ;
  assign n17587 = n17557 | n17574 ;
  assign n40152 = ~n17587 ;
  assign n17965 = n40152 & n145 ;
  assign n17966 = n17184 | n17965 ;
  assign n17559 = n17184 & n39774 ;
  assign n40153 = ~n17574 ;
  assign n17586 = n17559 & n40153 ;
  assign n17967 = n17586 & n145 ;
  assign n40154 = ~n17967 ;
  assign n17968 = n17966 & n40154 ;
  assign n18394 = n40133 & n18375 ;
  assign n18395 = n17858 | n18394 ;
  assign n40155 = ~n18377 ;
  assign n18396 = n40155 & n18395 ;
  assign n40156 = ~n18396 ;
  assign n18397 = n176 & n40156 ;
  assign n18398 = n40143 & n18395 ;
  assign n18399 = n17958 | n18398 ;
  assign n40157 = ~n18397 ;
  assign n18400 = n40157 & n18399 ;
  assign n40158 = ~n18400 ;
  assign n18401 = n177 & n40158 ;
  assign n18402 = n178 | n18401 ;
  assign n40159 = ~n18402 ;
  assign n18403 = n18384 & n40159 ;
  assign n18404 = n17968 | n18403 ;
  assign n40160 = ~n18386 ;
  assign n18405 = n40160 & n18404 ;
  assign n40161 = ~n18405 ;
  assign n18406 = n179 & n40161 ;
  assign n17612 = n17578 | n17596 ;
  assign n40162 = ~n17612 ;
  assign n17969 = n40162 & n145 ;
  assign n17970 = n17188 | n17969 ;
  assign n40163 = ~n17578 ;
  assign n17584 = n17188 & n40163 ;
  assign n17585 = n39780 & n17584 ;
  assign n17971 = n17585 & n145 ;
  assign n40164 = ~n17971 ;
  assign n17972 = n17970 & n40164 ;
  assign n18387 = n1707 | n18386 ;
  assign n40165 = ~n18387 ;
  assign n18407 = n40165 & n18404 ;
  assign n18411 = n17972 | n18407 ;
  assign n40166 = ~n18406 ;
  assign n18412 = n40166 & n18411 ;
  assign n40167 = ~n18412 ;
  assign n18413 = n1487 & n40167 ;
  assign n17611 = n17581 | n17598 ;
  assign n40168 = ~n17611 ;
  assign n17973 = n40168 & n145 ;
  assign n17974 = n17191 | n17973 ;
  assign n17582 = n17191 & n39790 ;
  assign n40169 = ~n17598 ;
  assign n17610 = n17582 & n40169 ;
  assign n17975 = n17610 & n145 ;
  assign n40170 = ~n17975 ;
  assign n17976 = n17974 & n40170 ;
  assign n18418 = n40149 & n18399 ;
  assign n18419 = n17964 | n18418 ;
  assign n40171 = ~n18401 ;
  assign n18420 = n40171 & n18419 ;
  assign n40172 = ~n18420 ;
  assign n18421 = n178 & n40172 ;
  assign n18422 = n40159 & n18419 ;
  assign n18423 = n17968 | n18422 ;
  assign n40173 = ~n18421 ;
  assign n18424 = n40173 & n18423 ;
  assign n40174 = ~n18424 ;
  assign n18425 = n1707 & n40174 ;
  assign n18426 = n1487 | n18425 ;
  assign n40175 = ~n18426 ;
  assign n18427 = n18411 & n40175 ;
  assign n18428 = n17976 | n18427 ;
  assign n40176 = ~n18413 ;
  assign n18429 = n40176 & n18428 ;
  assign n40177 = ~n18429 ;
  assign n18430 = n181 & n40177 ;
  assign n17629 = n17602 | n17620 ;
  assign n40178 = ~n17629 ;
  assign n17909 = n40178 & n145 ;
  assign n17910 = n17096 | n17909 ;
  assign n40179 = ~n17602 ;
  assign n17608 = n17096 & n40179 ;
  assign n17609 = n39796 & n17608 ;
  assign n17977 = n17609 & n145 ;
  assign n40180 = ~n17977 ;
  assign n17978 = n17910 & n40180 ;
  assign n18414 = n181 | n18413 ;
  assign n40181 = ~n18414 ;
  assign n18431 = n40181 & n18428 ;
  assign n18432 = n17978 | n18431 ;
  assign n40182 = ~n18430 ;
  assign n18433 = n40182 & n18432 ;
  assign n40183 = ~n18433 ;
  assign n18434 = n182 & n40183 ;
  assign n17607 = n17193 & n39806 ;
  assign n40184 = ~n17622 ;
  assign n17627 = n17607 & n40184 ;
  assign n17868 = n17627 & n145 ;
  assign n17628 = n17605 | n17622 ;
  assign n40185 = ~n17628 ;
  assign n17979 = n40185 & n145 ;
  assign n17980 = n17193 | n17979 ;
  assign n40186 = ~n17868 ;
  assign n17981 = n40186 & n17980 ;
  assign n18442 = n40165 & n18423 ;
  assign n18443 = n17972 | n18442 ;
  assign n40187 = ~n18425 ;
  assign n18444 = n40187 & n18443 ;
  assign n40188 = ~n18444 ;
  assign n18445 = n180 & n40188 ;
  assign n18446 = n40175 & n18443 ;
  assign n18447 = n17976 | n18446 ;
  assign n40189 = ~n18445 ;
  assign n18448 = n40189 & n18447 ;
  assign n40190 = ~n18448 ;
  assign n18449 = n181 & n40190 ;
  assign n18450 = n182 | n18449 ;
  assign n40191 = ~n18450 ;
  assign n18451 = n18432 & n40191 ;
  assign n18452 = n17981 | n18451 ;
  assign n40192 = ~n18434 ;
  assign n18453 = n40192 & n18452 ;
  assign n40193 = ~n18453 ;
  assign n18454 = n183 & n40193 ;
  assign n18435 = n183 | n18434 ;
  assign n40194 = ~n18435 ;
  assign n18455 = n40194 & n18452 ;
  assign n40195 = ~n17626 ;
  assign n17734 = n40195 & n17714 ;
  assign n17735 = n39812 & n17734 ;
  assign n17983 = n17735 & n145 ;
  assign n17639 = n17626 | n17637 ;
  assign n40196 = ~n17639 ;
  assign n17982 = n40196 & n145 ;
  assign n18487 = n17714 | n17982 ;
  assign n40197 = ~n17983 ;
  assign n18488 = n40197 & n18487 ;
  assign n18489 = n18455 | n18488 ;
  assign n40198 = ~n18454 ;
  assign n18490 = n40198 & n18489 ;
  assign n40199 = ~n18490 ;
  assign n18491 = n838 & n40199 ;
  assign n17733 = n17717 | n17720 ;
  assign n40200 = ~n17733 ;
  assign n17986 = n40200 & n145 ;
  assign n17987 = n17712 | n17986 ;
  assign n17719 = n17712 & n39822 ;
  assign n40201 = ~n17720 ;
  assign n17732 = n17719 & n40201 ;
  assign n17990 = n17732 & n145 ;
  assign n40202 = ~n17990 ;
  assign n17991 = n17987 & n40202 ;
  assign n18459 = n40181 & n18447 ;
  assign n18460 = n17978 | n18459 ;
  assign n40203 = ~n18449 ;
  assign n18461 = n40203 & n18460 ;
  assign n40204 = ~n18461 ;
  assign n18462 = n182 & n40204 ;
  assign n18463 = n40191 & n18460 ;
  assign n18464 = n17981 | n18463 ;
  assign n40205 = ~n18462 ;
  assign n18465 = n40205 & n18464 ;
  assign n40206 = ~n18465 ;
  assign n18466 = n996 & n40206 ;
  assign n18467 = n838 | n18466 ;
  assign n40207 = ~n18467 ;
  assign n18494 = n40207 & n18489 ;
  assign n18495 = n17991 | n18494 ;
  assign n40208 = ~n18491 ;
  assign n18496 = n40208 & n18495 ;
  assign n40209 = ~n18496 ;
  assign n18497 = n185 & n40209 ;
  assign n17758 = n17724 | n17742 ;
  assign n40210 = ~n17758 ;
  assign n17894 = n40210 & n145 ;
  assign n17895 = n17706 | n17894 ;
  assign n40211 = ~n17724 ;
  assign n17730 = n17706 & n40211 ;
  assign n17731 = n39828 & n17730 ;
  assign n17984 = n17731 & n145 ;
  assign n40212 = ~n17984 ;
  assign n17985 = n17895 & n40212 ;
  assign n18492 = n185 | n18491 ;
  assign n40213 = ~n18492 ;
  assign n18498 = n40213 & n18495 ;
  assign n18499 = n17985 | n18498 ;
  assign n40214 = ~n18497 ;
  assign n18500 = n40214 & n18499 ;
  assign n40215 = ~n18500 ;
  assign n18501 = n186 & n40215 ;
  assign n17756 = n17727 | n17744 ;
  assign n40216 = ~n17756 ;
  assign n17988 = n40216 & n145 ;
  assign n17989 = n17699 | n17988 ;
  assign n17729 = n17699 & n39838 ;
  assign n40217 = ~n17744 ;
  assign n17757 = n17729 & n40217 ;
  assign n17992 = n17757 & n145 ;
  assign n40218 = ~n17992 ;
  assign n17993 = n17989 & n40218 ;
  assign n18468 = n40194 & n18464 ;
  assign n18511 = n18468 | n18488 ;
  assign n40219 = ~n18466 ;
  assign n18512 = n40219 & n18511 ;
  assign n40220 = ~n18512 ;
  assign n18513 = n184 & n40220 ;
  assign n18514 = n40207 & n18511 ;
  assign n18515 = n17991 | n18514 ;
  assign n40221 = ~n18513 ;
  assign n18516 = n40221 & n18515 ;
  assign n40222 = ~n18516 ;
  assign n18517 = n185 & n40222 ;
  assign n18518 = n186 | n18517 ;
  assign n40223 = ~n18518 ;
  assign n18519 = n18499 & n40223 ;
  assign n18520 = n17993 | n18519 ;
  assign n40224 = ~n18501 ;
  assign n18521 = n40224 & n18520 ;
  assign n40225 = ~n18521 ;
  assign n18522 = n187 & n40225 ;
  assign n40226 = ~n17748 ;
  assign n17754 = n17693 & n40226 ;
  assign n17755 = n39844 & n17754 ;
  assign n17950 = n17755 & n145 ;
  assign n17782 = n17748 | n17766 ;
  assign n40227 = ~n17782 ;
  assign n17994 = n40227 & n145 ;
  assign n17995 = n17693 | n17994 ;
  assign n40228 = ~n17950 ;
  assign n17996 = n40228 & n17995 ;
  assign n18502 = n528 | n18501 ;
  assign n40229 = ~n18502 ;
  assign n18523 = n40229 & n18520 ;
  assign n18524 = n17996 | n18523 ;
  assign n40230 = ~n18522 ;
  assign n18525 = n40230 & n18524 ;
  assign n40231 = ~n18525 ;
  assign n18526 = n413 & n40231 ;
  assign n17780 = n17751 | n17768 ;
  assign n40232 = ~n17780 ;
  assign n17959 = n40232 & n145 ;
  assign n17960 = n17686 | n17959 ;
  assign n17753 = n17686 & n39854 ;
  assign n40233 = ~n17768 ;
  assign n17781 = n17753 & n40233 ;
  assign n17998 = n17781 & n145 ;
  assign n40234 = ~n17998 ;
  assign n17999 = n17960 & n40234 ;
  assign n18534 = n40213 & n18515 ;
  assign n18535 = n17985 | n18534 ;
  assign n40235 = ~n18517 ;
  assign n18536 = n40235 & n18535 ;
  assign n40236 = ~n18536 ;
  assign n18537 = n186 & n40236 ;
  assign n18538 = n40223 & n18535 ;
  assign n18539 = n17993 | n18538 ;
  assign n40237 = ~n18537 ;
  assign n18540 = n40237 & n18539 ;
  assign n40238 = ~n18540 ;
  assign n18541 = n528 & n40238 ;
  assign n18542 = n413 | n18541 ;
  assign n40239 = ~n18542 ;
  assign n18543 = n18524 & n40239 ;
  assign n18544 = n17999 | n18543 ;
  assign n40240 = ~n18526 ;
  assign n18545 = n40240 & n18544 ;
  assign n40241 = ~n18545 ;
  assign n18546 = n189 & n40241 ;
  assign n17806 = n17772 | n17790 ;
  assign n40242 = ~n17806 ;
  assign n17830 = n40242 & n145 ;
  assign n17831 = n17680 | n17830 ;
  assign n40243 = ~n17772 ;
  assign n17778 = n17680 & n40243 ;
  assign n17779 = n39860 & n17778 ;
  assign n17913 = n17779 & n145 ;
  assign n40244 = ~n17913 ;
  assign n17914 = n17831 & n40244 ;
  assign n18528 = n189 | n18526 ;
  assign n40245 = ~n18528 ;
  assign n18547 = n40245 & n18544 ;
  assign n18548 = n17914 | n18547 ;
  assign n40246 = ~n18546 ;
  assign n18549 = n40246 & n18548 ;
  assign n40247 = ~n18549 ;
  assign n18550 = n190 & n40247 ;
  assign n18552 = n287 | n18550 ;
  assign n17777 = n17673 & n39870 ;
  assign n40248 = ~n17792 ;
  assign n17804 = n17777 & n40248 ;
  assign n17837 = n17804 & n145 ;
  assign n17805 = n17775 | n17792 ;
  assign n40249 = ~n17805 ;
  assign n18000 = n40249 & n145 ;
  assign n18001 = n17673 | n18000 ;
  assign n40250 = ~n17837 ;
  assign n18002 = n40250 & n18001 ;
  assign n18556 = n40229 & n18539 ;
  assign n18557 = n17996 | n18556 ;
  assign n40251 = ~n18541 ;
  assign n18558 = n40251 & n18557 ;
  assign n40252 = ~n18558 ;
  assign n18559 = n188 & n40252 ;
  assign n18560 = n40239 & n18557 ;
  assign n18561 = n17999 | n18560 ;
  assign n40253 = ~n18559 ;
  assign n18562 = n40253 & n18561 ;
  assign n40254 = ~n18562 ;
  assign n18563 = n189 & n40254 ;
  assign n18564 = n190 | n18563 ;
  assign n40255 = ~n18564 ;
  assign n18565 = n18548 & n40255 ;
  assign n18566 = n18002 | n18565 ;
  assign n40256 = ~n18552 ;
  assign n18567 = n40256 & n18566 ;
  assign n18568 = n18486 | n18567 ;
  assign n17801 = n17660 & n39892 ;
  assign n40257 = ~n17816 ;
  assign n17817 = n17801 & n40257 ;
  assign n17997 = n17817 & n145 ;
  assign n17818 = n17799 | n17816 ;
  assign n40258 = ~n17818 ;
  assign n18003 = n40258 & n145 ;
  assign n18004 = n17660 | n18003 ;
  assign n40259 = ~n17997 ;
  assign n18005 = n40259 & n18004 ;
  assign n40260 = ~n18550 ;
  assign n18571 = n40260 & n18566 ;
  assign n40261 = ~n18571 ;
  assign n18572 = n191 & n40261 ;
  assign n40262 = ~n18572 ;
  assign n18573 = n18005 & n40262 ;
  assign n18574 = n18568 & n18573 ;
  assign n18579 = n18568 & n40262 ;
  assign n18580 = n18005 | n18579 ;
  assign n17821 = n17199 | n17820 ;
  assign n40263 = ~n17821 ;
  assign n18015 = n40263 & n145 ;
  assign n18469 = n17825 | n18015 ;
  assign n18470 = n18005 | n18469 ;
  assign n18551 = n191 | n18550 ;
  assign n40264 = ~n18551 ;
  assign n18582 = n40264 & n18566 ;
  assign n18583 = n18486 | n18582 ;
  assign n18584 = n40262 & n18583 ;
  assign n18585 = n18470 | n18584 ;
  assign n18586 = n31336 & n18585 ;
  assign n17822 = n192 & n17821 ;
  assign n40265 = ~n17199 ;
  assign n18006 = n40265 & n145 ;
  assign n40266 = ~n18006 ;
  assign n18007 = n17820 & n40266 ;
  assign n40267 = ~n18007 ;
  assign n18008 = n17822 & n40267 ;
  assign n17648 = n17196 | n17644 ;
  assign n40268 = ~n17648 ;
  assign n17649 = n17198 & n40268 ;
  assign n17650 = n39910 & n17649 ;
  assign n18471 = n17650 & n39911 ;
  assign n18472 = n39912 & n18471 ;
  assign n18473 = n18008 | n18472 ;
  assign n18592 = n18573 & n18583 ;
  assign n18593 = n18473 | n18592 ;
  assign n144 = n18586 | n18593 ;
  assign n40269 = ~n18580 ;
  assign n18779 = n40269 & n144 ;
  assign n18780 = n18574 | n18779 ;
  assign n40270 = ~n18582 ;
  assign n19265 = n18486 & n40270 ;
  assign n19266 = n40262 & n19265 ;
  assign n19267 = n144 & n19266 ;
  assign n19269 = n18572 | n18582 ;
  assign n40271 = ~n19269 ;
  assign n19270 = n144 & n40271 ;
  assign n19271 = n18486 | n19270 ;
  assign n40272 = ~n19267 ;
  assign n19272 = n40272 & n19271 ;
  assign n19273 = n18780 | n19272 ;
  assign n227 = x28 | x29 ;
  assign n228 = x30 | n227 ;
  assign n18611 = x30 & n144 ;
  assign n40273 = ~n18611 ;
  assign n18612 = n228 & n40273 ;
  assign n40274 = ~n18612 ;
  assign n18613 = n145 & n40274 ;
  assign n18614 = n146 | n18613 ;
  assign n17651 = n228 & n39909 ;
  assign n17652 = n39910 & n17651 ;
  assign n18481 = n17652 & n39911 ;
  assign n18482 = n39912 & n18481 ;
  assign n18675 = n18482 & n40273 ;
  assign n40275 = ~n224 ;
  assign n18681 = n40275 & n144 ;
  assign n40276 = ~x30 ;
  assign n18683 = n40276 & n144 ;
  assign n40277 = ~n18683 ;
  assign n18684 = x31 & n40277 ;
  assign n18694 = n18681 | n18684 ;
  assign n18695 = n18675 | n18694 ;
  assign n40278 = ~n18614 ;
  assign n18696 = n40278 & n18695 ;
  assign n40279 = ~n18472 ;
  assign n18474 = n145 & n40279 ;
  assign n40280 = ~n18008 ;
  assign n18475 = n40280 & n18474 ;
  assign n40281 = ~n18574 ;
  assign n18576 = n18475 & n40281 ;
  assign n40282 = ~n18586 ;
  assign n18587 = n18576 & n40282 ;
  assign n18588 = x32 | n18587 ;
  assign n18682 = n18588 | n18681 ;
  assign n18697 = n18587 | n18681 ;
  assign n18698 = x32 & n18697 ;
  assign n40283 = ~n18698 ;
  assign n18699 = n18682 & n40283 ;
  assign n18700 = n18696 | n18699 ;
  assign n229 = n40276 & n227 ;
  assign n18575 = n18473 | n18574 ;
  assign n18795 = n18470 | n18579 ;
  assign n18796 = n31336 & n18795 ;
  assign n18797 = n18575 | n18796 ;
  assign n40284 = ~n18797 ;
  assign n18798 = x30 & n40284 ;
  assign n18799 = n229 | n18798 ;
  assign n40285 = ~n18799 ;
  assign n18800 = n145 & n40285 ;
  assign n40286 = ~n18800 ;
  assign n18801 = n18695 & n40286 ;
  assign n40287 = ~n18801 ;
  assign n18802 = n146 & n40287 ;
  assign n40288 = ~n18802 ;
  assign n18803 = n18700 & n40288 ;
  assign n40289 = ~n18803 ;
  assign n18804 = n16322 & n40289 ;
  assign n17933 = n17850 | n17931 ;
  assign n40290 = ~n17933 ;
  assign n18021 = n40290 & n18020 ;
  assign n18705 = n18021 & n144 ;
  assign n18709 = n40290 & n144 ;
  assign n18710 = n18020 | n18709 ;
  assign n40291 = ~n18705 ;
  assign n18711 = n40291 & n18710 ;
  assign n40292 = ~n18613 ;
  assign n18701 = n40292 & n18695 ;
  assign n40293 = ~n18701 ;
  assign n18702 = n146 & n40293 ;
  assign n18703 = n16322 | n18702 ;
  assign n18811 = n146 | n18800 ;
  assign n40294 = ~n18811 ;
  assign n18812 = n18695 & n40294 ;
  assign n18813 = n18699 | n18812 ;
  assign n40295 = ~n18703 ;
  assign n18814 = n40295 & n18813 ;
  assign n18815 = n18711 | n18814 ;
  assign n40296 = ~n18804 ;
  assign n18816 = n40296 & n18815 ;
  assign n40297 = ~n18816 ;
  assign n18817 = n15807 & n40297 ;
  assign n40298 = ~n18027 ;
  assign n18057 = n40298 & n18036 ;
  assign n18058 = n39931 & n18057 ;
  assign n18743 = n18058 & n144 ;
  assign n18028 = n18026 | n18027 ;
  assign n40299 = ~n18028 ;
  assign n18744 = n40299 & n144 ;
  assign n18745 = n18036 | n18744 ;
  assign n40300 = ~n18743 ;
  assign n18746 = n40300 & n18745 ;
  assign n18805 = n15807 | n18804 ;
  assign n40301 = ~n18805 ;
  assign n18819 = n40301 & n18815 ;
  assign n18820 = n18746 | n18819 ;
  assign n40302 = ~n18817 ;
  assign n18821 = n40302 & n18820 ;
  assign n40303 = ~n18821 ;
  assign n18822 = n149 & n40303 ;
  assign n18056 = n18039 | n18042 ;
  assign n40304 = ~n18056 ;
  assign n18679 = n40304 & n144 ;
  assign n18680 = n17921 | n18679 ;
  assign n18041 = n17921 & n39919 ;
  assign n40305 = ~n18042 ;
  assign n18055 = n18041 & n40305 ;
  assign n18724 = n18055 & n144 ;
  assign n40306 = ~n18724 ;
  assign n18725 = n18680 & n40306 ;
  assign n18818 = n149 | n18817 ;
  assign n40307 = ~n18818 ;
  assign n18823 = n40307 & n18820 ;
  assign n18824 = n18725 | n18823 ;
  assign n40308 = ~n18822 ;
  assign n18825 = n40308 & n18824 ;
  assign n40309 = ~n18825 ;
  assign n18826 = n150 & n40309 ;
  assign n18054 = n18045 | n18046 ;
  assign n40310 = ~n18054 ;
  assign n18660 = n40310 & n144 ;
  assign n18661 = n18014 | n18660 ;
  assign n40311 = ~n18046 ;
  assign n18052 = n18014 & n40311 ;
  assign n18053 = n39925 & n18052 ;
  assign n18692 = n18053 & n144 ;
  assign n40312 = ~n18692 ;
  assign n18693 = n18661 & n40312 ;
  assign n18806 = n147 & n40289 ;
  assign n18808 = n147 | n18802 ;
  assign n40313 = ~n18808 ;
  assign n18831 = n40313 & n18813 ;
  assign n18832 = n18711 | n18831 ;
  assign n40314 = ~n18806 ;
  assign n18833 = n40314 & n18832 ;
  assign n40315 = ~n18833 ;
  assign n18834 = n148 & n40315 ;
  assign n18835 = n40301 & n18832 ;
  assign n18836 = n18746 | n18835 ;
  assign n40316 = ~n18834 ;
  assign n18837 = n40316 & n18836 ;
  assign n40317 = ~n18837 ;
  assign n18838 = n149 & n40317 ;
  assign n18839 = n150 | n18838 ;
  assign n40318 = ~n18839 ;
  assign n18840 = n18824 & n40318 ;
  assign n18841 = n18693 | n18840 ;
  assign n40319 = ~n18826 ;
  assign n18842 = n40319 & n18841 ;
  assign n40320 = ~n18842 ;
  assign n18843 = n151 & n40320 ;
  assign n18051 = n18017 & n39936 ;
  assign n40321 = ~n18067 ;
  assign n18080 = n18051 & n40321 ;
  assign n18597 = n18080 & n144 ;
  assign n18081 = n18049 | n18067 ;
  assign n40322 = ~n18081 ;
  assign n18636 = n40322 & n144 ;
  assign n18637 = n18017 | n18636 ;
  assign n40323 = ~n18597 ;
  assign n18638 = n40323 & n18637 ;
  assign n18827 = n151 | n18826 ;
  assign n40324 = ~n18827 ;
  assign n18844 = n40324 & n18841 ;
  assign n18845 = n18638 | n18844 ;
  assign n40325 = ~n18843 ;
  assign n18846 = n40325 & n18845 ;
  assign n40326 = ~n18846 ;
  assign n18847 = n13079 & n40326 ;
  assign n40327 = ~n18071 ;
  assign n18077 = n17912 & n40327 ;
  assign n18078 = n39942 & n18077 ;
  assign n18596 = n18078 & n144 ;
  assign n18079 = n18070 | n18071 ;
  assign n40328 = ~n18079 ;
  assign n18706 = n40328 & n144 ;
  assign n18707 = n17912 | n18706 ;
  assign n40329 = ~n18596 ;
  assign n18708 = n40329 & n18707 ;
  assign n18856 = n40307 & n18836 ;
  assign n18857 = n18725 | n18856 ;
  assign n40330 = ~n18838 ;
  assign n18858 = n40330 & n18857 ;
  assign n40331 = ~n18858 ;
  assign n18859 = n150 & n40331 ;
  assign n18860 = n40318 & n18857 ;
  assign n18861 = n18693 | n18860 ;
  assign n40332 = ~n18859 ;
  assign n18862 = n40332 & n18861 ;
  assign n40333 = ~n18862 ;
  assign n18863 = n13662 & n40333 ;
  assign n18864 = n152 | n18863 ;
  assign n40334 = ~n18864 ;
  assign n18865 = n18845 & n40334 ;
  assign n18866 = n18708 | n18865 ;
  assign n40335 = ~n18847 ;
  assign n18867 = n40335 & n18866 ;
  assign n40336 = ~n18867 ;
  assign n18868 = n153 & n40336 ;
  assign n18105 = n18074 | n18091 ;
  assign n40337 = ~n18105 ;
  assign n18658 = n40337 & n144 ;
  assign n18659 = n17897 | n18658 ;
  assign n18076 = n17897 & n39952 ;
  assign n40338 = ~n18091 ;
  assign n18104 = n18076 & n40338 ;
  assign n18717 = n18104 & n144 ;
  assign n40339 = ~n18717 ;
  assign n18718 = n18659 & n40339 ;
  assign n18848 = n153 | n18847 ;
  assign n40340 = ~n18848 ;
  assign n18869 = n40340 & n18866 ;
  assign n18870 = n18718 | n18869 ;
  assign n40341 = ~n18868 ;
  assign n18871 = n40341 & n18870 ;
  assign n40342 = ~n18871 ;
  assign n18872 = n154 & n40342 ;
  assign n18103 = n18094 | n18095 ;
  assign n40343 = ~n18103 ;
  assign n18608 = n40343 & n144 ;
  assign n18609 = n17937 | n18608 ;
  assign n40344 = ~n18095 ;
  assign n18101 = n17937 & n40344 ;
  assign n18102 = n39958 & n18101 ;
  assign n18650 = n18102 & n144 ;
  assign n40345 = ~n18650 ;
  assign n18651 = n18609 & n40345 ;
  assign n18880 = n40324 & n18861 ;
  assign n18881 = n18638 | n18880 ;
  assign n40346 = ~n18863 ;
  assign n18882 = n40346 & n18881 ;
  assign n40347 = ~n18882 ;
  assign n18883 = n152 & n40347 ;
  assign n18884 = n40334 & n18881 ;
  assign n18885 = n18708 | n18884 ;
  assign n40348 = ~n18883 ;
  assign n18886 = n40348 & n18885 ;
  assign n40349 = ~n18886 ;
  assign n18887 = n153 & n40349 ;
  assign n18888 = n154 | n18887 ;
  assign n40350 = ~n18888 ;
  assign n18889 = n18870 & n40350 ;
  assign n18890 = n18651 | n18889 ;
  assign n40351 = ~n18872 ;
  assign n18891 = n40351 & n18890 ;
  assign n40352 = ~n18891 ;
  assign n18892 = n155 & n40352 ;
  assign n18129 = n18098 | n18115 ;
  assign n40353 = ~n18129 ;
  assign n18617 = n40353 & n144 ;
  assign n18618 = n17924 | n18617 ;
  assign n18100 = n17924 & n39968 ;
  assign n40354 = ~n18115 ;
  assign n18128 = n18100 & n40354 ;
  assign n18786 = n18128 & n144 ;
  assign n40355 = ~n18786 ;
  assign n18787 = n18618 & n40355 ;
  assign n18873 = n11067 | n18872 ;
  assign n40356 = ~n18873 ;
  assign n18893 = n40356 & n18890 ;
  assign n18894 = n18787 | n18893 ;
  assign n40357 = ~n18892 ;
  assign n18895 = n40357 & n18894 ;
  assign n40358 = ~n18895 ;
  assign n18896 = n10657 & n40358 ;
  assign n40359 = ~n18119 ;
  assign n18125 = n17943 & n40359 ;
  assign n18126 = n39974 & n18125 ;
  assign n18664 = n18126 & n144 ;
  assign n18127 = n18118 | n18119 ;
  assign n40360 = ~n18127 ;
  assign n18740 = n40360 & n144 ;
  assign n18741 = n17943 | n18740 ;
  assign n40361 = ~n18664 ;
  assign n18742 = n40361 & n18741 ;
  assign n18904 = n40340 & n18885 ;
  assign n18905 = n18718 | n18904 ;
  assign n40362 = ~n18887 ;
  assign n18906 = n40362 & n18905 ;
  assign n40363 = ~n18906 ;
  assign n18907 = n154 & n40363 ;
  assign n18908 = n40350 & n18905 ;
  assign n18909 = n18651 | n18908 ;
  assign n40364 = ~n18907 ;
  assign n18910 = n40364 & n18909 ;
  assign n40365 = ~n18910 ;
  assign n18911 = n11067 & n40365 ;
  assign n18912 = n10657 | n18911 ;
  assign n40366 = ~n18912 ;
  assign n18913 = n18894 & n40366 ;
  assign n18914 = n18742 | n18913 ;
  assign n40367 = ~n18896 ;
  assign n18915 = n40367 & n18914 ;
  assign n40368 = ~n18915 ;
  assign n18916 = n157 & n40368 ;
  assign n18124 = n17946 & n39984 ;
  assign n40369 = ~n18139 ;
  assign n18152 = n18124 & n40369 ;
  assign n18595 = n18152 & n144 ;
  assign n18153 = n18122 | n18139 ;
  assign n40370 = ~n18153 ;
  assign n18670 = n40370 & n144 ;
  assign n18671 = n17946 | n18670 ;
  assign n40371 = ~n18595 ;
  assign n18672 = n40371 & n18671 ;
  assign n18897 = n157 | n18896 ;
  assign n40372 = ~n18897 ;
  assign n18917 = n40372 & n18914 ;
  assign n18918 = n18672 | n18917 ;
  assign n40373 = ~n18916 ;
  assign n18919 = n40373 & n18918 ;
  assign n40374 = ~n18919 ;
  assign n18920 = n158 & n40374 ;
  assign n18151 = n18142 | n18143 ;
  assign n40375 = ~n18151 ;
  assign n18662 = n40375 & n144 ;
  assign n18663 = n17949 | n18662 ;
  assign n40376 = ~n18143 ;
  assign n18149 = n17949 & n40376 ;
  assign n18150 = n39990 & n18149 ;
  assign n18715 = n18150 & n144 ;
  assign n40377 = ~n18715 ;
  assign n18716 = n18663 & n40377 ;
  assign n18928 = n40356 & n18909 ;
  assign n18929 = n18787 | n18928 ;
  assign n40378 = ~n18911 ;
  assign n18930 = n40378 & n18929 ;
  assign n40379 = ~n18930 ;
  assign n18931 = n156 & n40379 ;
  assign n18932 = n40366 & n18929 ;
  assign n18933 = n18742 | n18932 ;
  assign n40380 = ~n18931 ;
  assign n18934 = n40380 & n18933 ;
  assign n40381 = ~n18934 ;
  assign n18935 = n157 & n40381 ;
  assign n18936 = n158 | n18935 ;
  assign n40382 = ~n18936 ;
  assign n18937 = n18918 & n40382 ;
  assign n18938 = n18716 | n18937 ;
  assign n40383 = ~n18920 ;
  assign n18939 = n40383 & n18938 ;
  assign n40384 = ~n18939 ;
  assign n18940 = n159 & n40384 ;
  assign n18148 = n17929 & n40000 ;
  assign n40385 = ~n18163 ;
  assign n18176 = n18148 & n40385 ;
  assign n18704 = n18176 & n144 ;
  assign n18177 = n18146 | n18163 ;
  assign n40386 = ~n18177 ;
  assign n18712 = n40386 & n144 ;
  assign n18713 = n17929 | n18712 ;
  assign n40387 = ~n18704 ;
  assign n18714 = n40387 & n18713 ;
  assign n18921 = n8857 | n18920 ;
  assign n40388 = ~n18921 ;
  assign n18941 = n40388 & n18938 ;
  assign n18942 = n18714 | n18941 ;
  assign n40389 = ~n18940 ;
  assign n18943 = n40389 & n18942 ;
  assign n40390 = ~n18943 ;
  assign n18944 = n8534 & n40390 ;
  assign n18170 = n18166 | n18167 ;
  assign n40391 = ~n18170 ;
  assign n18722 = n40391 & n144 ;
  assign n18723 = n17956 | n18722 ;
  assign n40392 = ~n18167 ;
  assign n18168 = n17956 & n40392 ;
  assign n18169 = n40006 & n18168 ;
  assign n18774 = n18169 & n144 ;
  assign n40393 = ~n18774 ;
  assign n18775 = n18723 & n40393 ;
  assign n18952 = n40372 & n18933 ;
  assign n18953 = n18672 | n18952 ;
  assign n40394 = ~n18935 ;
  assign n18954 = n40394 & n18953 ;
  assign n40395 = ~n18954 ;
  assign n18955 = n158 & n40395 ;
  assign n18956 = n40382 & n18953 ;
  assign n18957 = n18716 | n18956 ;
  assign n40396 = ~n18955 ;
  assign n18958 = n40396 & n18957 ;
  assign n40397 = ~n18958 ;
  assign n18959 = n8857 & n40397 ;
  assign n18960 = n160 | n18959 ;
  assign n40398 = ~n18960 ;
  assign n18961 = n18942 & n40398 ;
  assign n18962 = n18775 | n18961 ;
  assign n40399 = ~n18944 ;
  assign n18963 = n40399 & n18962 ;
  assign n40400 = ~n18963 ;
  assign n18964 = n161 & n40400 ;
  assign n18175 = n17926 & n40016 ;
  assign n40401 = ~n18187 ;
  assign n18200 = n18175 & n40401 ;
  assign n18626 = n18200 & n144 ;
  assign n18201 = n18173 | n18187 ;
  assign n40402 = ~n18201 ;
  assign n18757 = n40402 & n144 ;
  assign n18758 = n17926 | n18757 ;
  assign n40403 = ~n18626 ;
  assign n18759 = n40403 & n18758 ;
  assign n18945 = n161 | n18944 ;
  assign n40404 = ~n18945 ;
  assign n18965 = n40404 & n18962 ;
  assign n18966 = n18759 | n18965 ;
  assign n40405 = ~n18964 ;
  assign n18967 = n40405 & n18966 ;
  assign n40406 = ~n18967 ;
  assign n18968 = n162 & n40406 ;
  assign n18199 = n18190 | n18191 ;
  assign n40407 = ~n18199 ;
  assign n18656 = n40407 & n144 ;
  assign n18657 = n17953 | n18656 ;
  assign n40408 = ~n18191 ;
  assign n18197 = n17953 & n40408 ;
  assign n18198 = n40022 & n18197 ;
  assign n18755 = n18198 & n144 ;
  assign n40409 = ~n18755 ;
  assign n18756 = n18657 & n40409 ;
  assign n18976 = n40388 & n18957 ;
  assign n18977 = n18714 | n18976 ;
  assign n40410 = ~n18959 ;
  assign n18978 = n40410 & n18977 ;
  assign n40411 = ~n18978 ;
  assign n18979 = n160 & n40411 ;
  assign n18980 = n40398 & n18977 ;
  assign n18981 = n18775 | n18980 ;
  assign n40412 = ~n18979 ;
  assign n18982 = n40412 & n18981 ;
  assign n40413 = ~n18982 ;
  assign n18983 = n161 & n40413 ;
  assign n18984 = n162 | n18983 ;
  assign n40414 = ~n18984 ;
  assign n18985 = n18966 & n40414 ;
  assign n18986 = n18756 | n18985 ;
  assign n40415 = ~n18968 ;
  assign n18987 = n40415 & n18986 ;
  assign n40416 = ~n18987 ;
  assign n18988 = n163 & n40416 ;
  assign n18195 = n17879 & n40032 ;
  assign n40417 = ~n18211 ;
  assign n18224 = n18195 & n40417 ;
  assign n18615 = n18224 & n144 ;
  assign n18225 = n18194 | n18211 ;
  assign n40418 = ~n18225 ;
  assign n18665 = n40418 & n144 ;
  assign n18666 = n17879 | n18665 ;
  assign n40419 = ~n18615 ;
  assign n18667 = n40419 & n18666 ;
  assign n18969 = n6889 | n18968 ;
  assign n40420 = ~n18969 ;
  assign n18989 = n40420 & n18986 ;
  assign n18990 = n18667 | n18989 ;
  assign n40421 = ~n18988 ;
  assign n18991 = n40421 & n18990 ;
  assign n40422 = ~n18991 ;
  assign n18992 = n6600 & n40422 ;
  assign n18223 = n18214 | n18215 ;
  assign n40423 = ~n18223 ;
  assign n18690 = n40423 & n144 ;
  assign n18691 = n17904 | n18690 ;
  assign n40424 = ~n18215 ;
  assign n18221 = n17904 & n40424 ;
  assign n18222 = n40038 & n18221 ;
  assign n18760 = n18222 & n144 ;
  assign n40425 = ~n18760 ;
  assign n18761 = n18691 & n40425 ;
  assign n18999 = n40404 & n18981 ;
  assign n19000 = n18759 | n18999 ;
  assign n40426 = ~n18983 ;
  assign n19001 = n40426 & n19000 ;
  assign n40427 = ~n19001 ;
  assign n19002 = n162 & n40427 ;
  assign n19003 = n40414 & n19000 ;
  assign n19004 = n18756 | n19003 ;
  assign n40428 = ~n19002 ;
  assign n19005 = n40428 & n19004 ;
  assign n40429 = ~n19005 ;
  assign n19006 = n6889 & n40429 ;
  assign n19007 = n6600 | n19006 ;
  assign n40430 = ~n19007 ;
  assign n19008 = n18990 & n40430 ;
  assign n19009 = n18761 | n19008 ;
  assign n40431 = ~n18992 ;
  assign n19010 = n40431 & n19009 ;
  assign n40432 = ~n19010 ;
  assign n19011 = n165 & n40432 ;
  assign n18220 = n17888 & n40048 ;
  assign n40433 = ~n18235 ;
  assign n18248 = n18220 & n40433 ;
  assign n18735 = n18248 & n144 ;
  assign n18249 = n18218 | n18235 ;
  assign n40434 = ~n18249 ;
  assign n18737 = n40434 & n144 ;
  assign n18738 = n17888 | n18737 ;
  assign n40435 = ~n18735 ;
  assign n18739 = n40435 & n18738 ;
  assign n18993 = n165 | n18992 ;
  assign n40436 = ~n18993 ;
  assign n19012 = n40436 & n19009 ;
  assign n19013 = n18739 | n19012 ;
  assign n40437 = ~n19011 ;
  assign n19014 = n40437 & n19013 ;
  assign n40438 = ~n19014 ;
  assign n19015 = n166 & n40438 ;
  assign n40439 = ~n18239 ;
  assign n18245 = n17919 & n40439 ;
  assign n18246 = n40054 & n18245 ;
  assign n18749 = n18246 & n144 ;
  assign n18247 = n18238 | n18239 ;
  assign n40440 = ~n18247 ;
  assign n18771 = n40440 & n144 ;
  assign n18772 = n17919 | n18771 ;
  assign n40441 = ~n18749 ;
  assign n18773 = n40441 & n18772 ;
  assign n19024 = n40420 & n19004 ;
  assign n19025 = n18667 | n19024 ;
  assign n40442 = ~n19006 ;
  assign n19026 = n40442 & n19025 ;
  assign n40443 = ~n19026 ;
  assign n19027 = n164 & n40443 ;
  assign n19028 = n40430 & n19025 ;
  assign n19029 = n18761 | n19028 ;
  assign n40444 = ~n19027 ;
  assign n19030 = n40444 & n19029 ;
  assign n40445 = ~n19030 ;
  assign n19031 = n165 & n40445 ;
  assign n19032 = n166 | n19031 ;
  assign n40446 = ~n19032 ;
  assign n19033 = n19013 & n40446 ;
  assign n19034 = n18773 | n19033 ;
  assign n40447 = ~n19015 ;
  assign n19035 = n40447 & n19034 ;
  assign n40448 = ~n19035 ;
  assign n19036 = n167 & n40448 ;
  assign n18244 = n17908 & n40064 ;
  assign n40449 = ~n18259 ;
  assign n18272 = n18244 & n40449 ;
  assign n18736 = n18272 & n144 ;
  assign n18273 = n18242 | n18259 ;
  assign n40450 = ~n18273 ;
  assign n18783 = n40450 & n144 ;
  assign n18784 = n17908 | n18783 ;
  assign n40451 = ~n18736 ;
  assign n18785 = n40451 & n18784 ;
  assign n19016 = n5352 | n19015 ;
  assign n40452 = ~n19016 ;
  assign n19037 = n40452 & n19034 ;
  assign n19038 = n18785 | n19037 ;
  assign n40453 = ~n19036 ;
  assign n19039 = n40453 & n19038 ;
  assign n40454 = ~n19039 ;
  assign n19040 = n4934 & n40454 ;
  assign n18271 = n18262 | n18263 ;
  assign n40455 = ~n18271 ;
  assign n18765 = n40455 & n144 ;
  assign n18766 = n17847 | n18765 ;
  assign n40456 = ~n18263 ;
  assign n18269 = n17847 & n40456 ;
  assign n18270 = n40070 & n18269 ;
  assign n18788 = n18270 & n144 ;
  assign n40457 = ~n18788 ;
  assign n18789 = n18766 & n40457 ;
  assign n19048 = n40436 & n19029 ;
  assign n19049 = n18739 | n19048 ;
  assign n40458 = ~n19031 ;
  assign n19050 = n40458 & n19049 ;
  assign n40459 = ~n19050 ;
  assign n19051 = n166 & n40459 ;
  assign n19052 = n40446 & n19049 ;
  assign n19053 = n18773 | n19052 ;
  assign n40460 = ~n19051 ;
  assign n19054 = n40460 & n19053 ;
  assign n40461 = ~n19054 ;
  assign n19055 = n5352 & n40461 ;
  assign n19056 = n4934 | n19055 ;
  assign n40462 = ~n19056 ;
  assign n19057 = n19038 & n40462 ;
  assign n19058 = n18789 | n19057 ;
  assign n40463 = ~n19040 ;
  assign n19059 = n40463 & n19058 ;
  assign n40464 = ~n19059 ;
  assign n19060 = n169 & n40464 ;
  assign n18268 = n17863 & n40080 ;
  assign n40465 = ~n18283 ;
  assign n18296 = n18268 & n40465 ;
  assign n18673 = n18296 & n144 ;
  assign n18297 = n18266 | n18283 ;
  assign n40466 = ~n18297 ;
  assign n18776 = n40466 & n144 ;
  assign n18777 = n17863 | n18776 ;
  assign n40467 = ~n18673 ;
  assign n18778 = n40467 & n18777 ;
  assign n19041 = n169 | n19040 ;
  assign n40468 = ~n19041 ;
  assign n19061 = n40468 & n19058 ;
  assign n19062 = n18778 | n19061 ;
  assign n40469 = ~n19060 ;
  assign n19063 = n40469 & n19062 ;
  assign n40470 = ~n19063 ;
  assign n19064 = n170 & n40470 ;
  assign n18295 = n18286 | n18287 ;
  assign n40471 = ~n18295 ;
  assign n18598 = n40471 & n144 ;
  assign n18599 = n17843 | n18598 ;
  assign n40472 = ~n18287 ;
  assign n18293 = n17843 & n40472 ;
  assign n18294 = n40086 & n18293 ;
  assign n18677 = n18294 & n144 ;
  assign n40473 = ~n18677 ;
  assign n18678 = n18599 & n40473 ;
  assign n19072 = n40452 & n19053 ;
  assign n19073 = n18785 | n19072 ;
  assign n40474 = ~n19055 ;
  assign n19074 = n40474 & n19073 ;
  assign n40475 = ~n19074 ;
  assign n19075 = n168 & n40475 ;
  assign n19076 = n40462 & n19073 ;
  assign n19077 = n18789 | n19076 ;
  assign n40476 = ~n19075 ;
  assign n19078 = n40476 & n19077 ;
  assign n40477 = ~n19078 ;
  assign n19079 = n169 & n40477 ;
  assign n19080 = n170 | n19079 ;
  assign n40478 = ~n19080 ;
  assign n19081 = n19062 & n40478 ;
  assign n19082 = n18678 | n19081 ;
  assign n40479 = ~n19064 ;
  assign n19083 = n40479 & n19082 ;
  assign n40480 = ~n19083 ;
  assign n19084 = n171 & n40480 ;
  assign n18292 = n17834 & n40096 ;
  assign n40481 = ~n18307 ;
  assign n18320 = n18292 & n40481 ;
  assign n18674 = n18320 & n144 ;
  assign n18321 = n18290 | n18307 ;
  assign n40482 = ~n18321 ;
  assign n18790 = n40482 & n144 ;
  assign n18791 = n17834 | n18790 ;
  assign n40483 = ~n18674 ;
  assign n18792 = n40483 & n18791 ;
  assign n19065 = n3940 | n19064 ;
  assign n40484 = ~n19065 ;
  assign n19085 = n40484 & n19082 ;
  assign n19086 = n18792 | n19085 ;
  assign n40485 = ~n19084 ;
  assign n19087 = n40485 & n19086 ;
  assign n40486 = ~n19087 ;
  assign n19088 = n3631 & n40486 ;
  assign n18319 = n18310 | n18311 ;
  assign n40487 = ~n18319 ;
  assign n18769 = n40487 & n144 ;
  assign n18770 = n17870 | n18769 ;
  assign n40488 = ~n18311 ;
  assign n18317 = n17870 & n40488 ;
  assign n18318 = n40102 & n18317 ;
  assign n18781 = n18318 & n144 ;
  assign n40489 = ~n18781 ;
  assign n18782 = n18770 & n40489 ;
  assign n19095 = n40468 & n19077 ;
  assign n19096 = n18778 | n19095 ;
  assign n40490 = ~n19079 ;
  assign n19097 = n40490 & n19096 ;
  assign n40491 = ~n19097 ;
  assign n19098 = n170 & n40491 ;
  assign n19099 = n40478 & n19096 ;
  assign n19100 = n18678 | n19099 ;
  assign n40492 = ~n19098 ;
  assign n19101 = n40492 & n19100 ;
  assign n40493 = ~n19101 ;
  assign n19102 = n3940 & n40493 ;
  assign n19103 = n3631 | n19102 ;
  assign n40494 = ~n19103 ;
  assign n19104 = n19086 & n40494 ;
  assign n19105 = n18782 | n19104 ;
  assign n40495 = ~n19088 ;
  assign n19106 = n40495 & n19105 ;
  assign n40496 = ~n19106 ;
  assign n19107 = n173 & n40496 ;
  assign n18345 = n18314 | n18331 ;
  assign n40497 = ~n18345 ;
  assign n18668 = n40497 & n144 ;
  assign n18669 = n17941 | n18668 ;
  assign n18316 = n17941 & n40112 ;
  assign n40498 = ~n18331 ;
  assign n18344 = n18316 & n40498 ;
  assign n18793 = n18344 & n144 ;
  assign n40499 = ~n18793 ;
  assign n18794 = n18669 & n40499 ;
  assign n19089 = n173 | n19088 ;
  assign n40500 = ~n19089 ;
  assign n19108 = n40500 & n19105 ;
  assign n19109 = n18794 | n19108 ;
  assign n40501 = ~n19107 ;
  assign n19110 = n40501 & n19109 ;
  assign n40502 = ~n19110 ;
  assign n19111 = n174 & n40502 ;
  assign n18343 = n18334 | n18335 ;
  assign n40503 = ~n18343 ;
  assign n18652 = n40503 & n144 ;
  assign n18653 = n17853 | n18652 ;
  assign n40504 = ~n18335 ;
  assign n18341 = n17853 & n40504 ;
  assign n18342 = n40118 & n18341 ;
  assign n18654 = n18342 & n144 ;
  assign n40505 = ~n18654 ;
  assign n18655 = n18653 & n40505 ;
  assign n19120 = n40484 & n19100 ;
  assign n19121 = n18792 | n19120 ;
  assign n40506 = ~n19102 ;
  assign n19122 = n40506 & n19121 ;
  assign n40507 = ~n19122 ;
  assign n19123 = n172 & n40507 ;
  assign n19124 = n40494 & n19121 ;
  assign n19125 = n18782 | n19124 ;
  assign n40508 = ~n19123 ;
  assign n19126 = n40508 & n19125 ;
  assign n40509 = ~n19126 ;
  assign n19127 = n173 & n40509 ;
  assign n19128 = n174 | n19127 ;
  assign n40510 = ~n19128 ;
  assign n19129 = n19109 & n40510 ;
  assign n19130 = n18655 | n19129 ;
  assign n40511 = ~n19111 ;
  assign n19131 = n40511 & n19130 ;
  assign n40512 = ~n19131 ;
  assign n19132 = n175 & n40512 ;
  assign n18369 = n18338 | n18355 ;
  assign n40513 = ~n18369 ;
  assign n18646 = n40513 & n144 ;
  assign n18647 = n17882 | n18646 ;
  assign n18340 = n17882 & n40128 ;
  assign n40514 = ~n18355 ;
  assign n18368 = n18340 & n40514 ;
  assign n18648 = n18368 & n144 ;
  assign n40515 = ~n18648 ;
  assign n18649 = n18647 & n40515 ;
  assign n19112 = n2753 | n19111 ;
  assign n40516 = ~n19112 ;
  assign n19133 = n40516 & n19130 ;
  assign n19134 = n18649 | n19133 ;
  assign n40517 = ~n19132 ;
  assign n19135 = n40517 & n19134 ;
  assign n40518 = ~n19135 ;
  assign n19136 = n2431 & n40518 ;
  assign n18367 = n18358 | n18359 ;
  assign n40519 = ~n18367 ;
  assign n18641 = n40519 & n144 ;
  assign n18642 = n17858 | n18641 ;
  assign n40520 = ~n18359 ;
  assign n18365 = n17858 & n40520 ;
  assign n18366 = n40134 & n18365 ;
  assign n18643 = n18366 & n144 ;
  assign n40521 = ~n18643 ;
  assign n18644 = n18642 & n40521 ;
  assign n19144 = n40500 & n19125 ;
  assign n19145 = n18794 | n19144 ;
  assign n40522 = ~n19127 ;
  assign n19146 = n40522 & n19145 ;
  assign n40523 = ~n19146 ;
  assign n19147 = n174 & n40523 ;
  assign n19148 = n40510 & n19145 ;
  assign n19149 = n18655 | n19148 ;
  assign n40524 = ~n19147 ;
  assign n19150 = n40524 & n19149 ;
  assign n40525 = ~n19150 ;
  assign n19151 = n2753 & n40525 ;
  assign n19152 = n2431 | n19151 ;
  assign n40526 = ~n19152 ;
  assign n19153 = n19134 & n40526 ;
  assign n19154 = n18644 | n19153 ;
  assign n40527 = ~n19136 ;
  assign n19155 = n40527 & n19154 ;
  assign n40528 = ~n19155 ;
  assign n19156 = n177 & n40528 ;
  assign n18393 = n18362 | n18379 ;
  assign n40529 = ~n18393 ;
  assign n18604 = n40529 & n144 ;
  assign n18605 = n17958 | n18604 ;
  assign n18364 = n17958 & n40144 ;
  assign n40530 = ~n18379 ;
  assign n18392 = n18364 & n40530 ;
  assign n18634 = n18392 & n144 ;
  assign n40531 = ~n18634 ;
  assign n18635 = n18605 & n40531 ;
  assign n19137 = n177 | n19136 ;
  assign n40532 = ~n19137 ;
  assign n19157 = n40532 & n19154 ;
  assign n19158 = n18635 | n19157 ;
  assign n40533 = ~n19156 ;
  assign n19159 = n40533 & n19158 ;
  assign n40534 = ~n19159 ;
  assign n19160 = n178 & n40534 ;
  assign n40535 = ~n18383 ;
  assign n18389 = n17964 & n40535 ;
  assign n18390 = n40150 & n18389 ;
  assign n18676 = n18390 & n144 ;
  assign n18391 = n18382 | n18383 ;
  assign n40536 = ~n18391 ;
  assign n18719 = n40536 & n144 ;
  assign n18720 = n17964 | n18719 ;
  assign n40537 = ~n18676 ;
  assign n18721 = n40537 & n18720 ;
  assign n19168 = n40516 & n19149 ;
  assign n19169 = n18649 | n19168 ;
  assign n40538 = ~n19151 ;
  assign n19170 = n40538 & n19169 ;
  assign n40539 = ~n19170 ;
  assign n19171 = n176 & n40539 ;
  assign n19172 = n40526 & n19169 ;
  assign n19173 = n18644 | n19172 ;
  assign n40540 = ~n19171 ;
  assign n19174 = n40540 & n19173 ;
  assign n40541 = ~n19174 ;
  assign n19175 = n177 & n40541 ;
  assign n19176 = n178 | n19175 ;
  assign n40542 = ~n19176 ;
  assign n19177 = n19158 & n40542 ;
  assign n19178 = n18721 | n19177 ;
  assign n40543 = ~n19160 ;
  assign n19179 = n40543 & n19178 ;
  assign n40544 = ~n19179 ;
  assign n19180 = n179 & n40544 ;
  assign n18417 = n18386 | n18403 ;
  assign n40545 = ~n18417 ;
  assign n18630 = n40545 & n144 ;
  assign n18631 = n17968 | n18630 ;
  assign n18388 = n17968 & n40160 ;
  assign n40546 = ~n18403 ;
  assign n18416 = n18388 & n40546 ;
  assign n18632 = n18416 & n144 ;
  assign n40547 = ~n18632 ;
  assign n18633 = n18631 & n40547 ;
  assign n19161 = n1707 | n19160 ;
  assign n40548 = ~n19161 ;
  assign n19181 = n40548 & n19178 ;
  assign n19182 = n18633 | n19181 ;
  assign n40549 = ~n19180 ;
  assign n19183 = n40549 & n19182 ;
  assign n40550 = ~n19183 ;
  assign n19184 = n1487 & n40550 ;
  assign n18410 = n18406 | n18407 ;
  assign n40551 = ~n18410 ;
  assign n18747 = n40551 & n144 ;
  assign n18748 = n17972 | n18747 ;
  assign n40552 = ~n18407 ;
  assign n18408 = n17972 & n40552 ;
  assign n18409 = n40166 & n18408 ;
  assign n18753 = n18409 & n144 ;
  assign n40553 = ~n18753 ;
  assign n18754 = n18748 & n40553 ;
  assign n19192 = n40532 & n19173 ;
  assign n19193 = n18635 | n19192 ;
  assign n40554 = ~n19175 ;
  assign n19194 = n40554 & n19193 ;
  assign n40555 = ~n19194 ;
  assign n19195 = n178 & n40555 ;
  assign n19196 = n40542 & n19193 ;
  assign n19197 = n18721 | n19196 ;
  assign n40556 = ~n19195 ;
  assign n19198 = n40556 & n19197 ;
  assign n40557 = ~n19198 ;
  assign n19199 = n1707 & n40557 ;
  assign n19200 = n1487 | n19199 ;
  assign n40558 = ~n19200 ;
  assign n19201 = n19182 & n40558 ;
  assign n19202 = n18754 | n19201 ;
  assign n40559 = ~n19184 ;
  assign n19203 = n40559 & n19202 ;
  assign n40560 = ~n19203 ;
  assign n19204 = n181 & n40560 ;
  assign n18415 = n17976 & n40176 ;
  assign n40561 = ~n18427 ;
  assign n18440 = n18415 & n40561 ;
  assign n18629 = n18440 & n144 ;
  assign n18441 = n18413 | n18427 ;
  assign n40562 = ~n18441 ;
  assign n18762 = n40562 & n144 ;
  assign n18763 = n17976 | n18762 ;
  assign n40563 = ~n18629 ;
  assign n18764 = n40563 & n18763 ;
  assign n19185 = n181 | n19184 ;
  assign n40564 = ~n19185 ;
  assign n19205 = n40564 & n19202 ;
  assign n19206 = n18764 | n19205 ;
  assign n40565 = ~n19204 ;
  assign n19207 = n40565 & n19206 ;
  assign n40566 = ~n19207 ;
  assign n19208 = n182 & n40566 ;
  assign n18439 = n18430 | n18431 ;
  assign n40567 = ~n18439 ;
  assign n18624 = n40567 & n144 ;
  assign n18625 = n17978 | n18624 ;
  assign n40568 = ~n18431 ;
  assign n18437 = n17978 & n40568 ;
  assign n18438 = n40182 & n18437 ;
  assign n18627 = n18438 & n144 ;
  assign n40569 = ~n18627 ;
  assign n18628 = n18625 & n40569 ;
  assign n19216 = n40548 & n19197 ;
  assign n19217 = n18633 | n19216 ;
  assign n40570 = ~n19199 ;
  assign n19218 = n40570 & n19217 ;
  assign n40571 = ~n19218 ;
  assign n19219 = n180 & n40571 ;
  assign n19220 = n40558 & n19217 ;
  assign n19221 = n18754 | n19220 ;
  assign n40572 = ~n19219 ;
  assign n19222 = n40572 & n19221 ;
  assign n40573 = ~n19222 ;
  assign n19223 = n181 & n40573 ;
  assign n19224 = n182 | n19223 ;
  assign n40574 = ~n19224 ;
  assign n19225 = n19206 & n40574 ;
  assign n19226 = n18628 | n19225 ;
  assign n40575 = ~n19208 ;
  assign n19227 = n40575 & n19226 ;
  assign n40576 = ~n19227 ;
  assign n19228 = n183 & n40576 ;
  assign n18436 = n17981 & n40192 ;
  assign n40577 = ~n18451 ;
  assign n18457 = n18436 & n40577 ;
  assign n18616 = n18457 & n144 ;
  assign n18458 = n18434 | n18451 ;
  assign n40578 = ~n18458 ;
  assign n18687 = n40578 & n144 ;
  assign n18688 = n17981 | n18687 ;
  assign n40579 = ~n18616 ;
  assign n18689 = n40579 & n18688 ;
  assign n19209 = n183 | n19208 ;
  assign n40580 = ~n19209 ;
  assign n19229 = n40580 & n19226 ;
  assign n19230 = n18689 | n19229 ;
  assign n40581 = ~n19228 ;
  assign n19231 = n40581 & n19230 ;
  assign n40582 = ~n19231 ;
  assign n19232 = n838 & n40582 ;
  assign n19240 = n40564 & n19221 ;
  assign n19241 = n18764 | n19240 ;
  assign n40583 = ~n19223 ;
  assign n19242 = n40583 & n19241 ;
  assign n40584 = ~n19242 ;
  assign n19243 = n182 & n40584 ;
  assign n19244 = n40574 & n19241 ;
  assign n19245 = n18628 | n19244 ;
  assign n40585 = ~n19243 ;
  assign n19246 = n40585 & n19245 ;
  assign n40586 = ~n19246 ;
  assign n19247 = n996 & n40586 ;
  assign n19248 = n838 | n19247 ;
  assign n40587 = ~n19248 ;
  assign n19249 = n19230 & n40587 ;
  assign n40588 = ~n18455 ;
  assign n18509 = n40588 & n18488 ;
  assign n18510 = n40198 & n18509 ;
  assign n18610 = n18510 & n144 ;
  assign n18456 = n18454 | n18455 ;
  assign n40589 = ~n18456 ;
  assign n18645 = n40589 & n144 ;
  assign n19284 = n18488 | n18645 ;
  assign n40590 = ~n18610 ;
  assign n19285 = n40590 & n19284 ;
  assign n19303 = n19249 | n19285 ;
  assign n40591 = ~n19232 ;
  assign n19304 = n40591 & n19303 ;
  assign n40592 = ~n19304 ;
  assign n19305 = n185 & n40592 ;
  assign n18508 = n18491 | n18494 ;
  assign n40593 = ~n18508 ;
  assign n18622 = n40593 & n144 ;
  assign n18623 = n17991 | n18622 ;
  assign n18493 = n17991 & n40208 ;
  assign n40594 = ~n18494 ;
  assign n18507 = n18493 & n40594 ;
  assign n18767 = n18507 & n144 ;
  assign n40595 = ~n18767 ;
  assign n18768 = n18623 & n40595 ;
  assign n19233 = n185 | n19232 ;
  assign n40596 = ~n19233 ;
  assign n19306 = n40596 & n19303 ;
  assign n19309 = n18768 | n19306 ;
  assign n40597 = ~n19305 ;
  assign n19310 = n40597 & n19309 ;
  assign n40598 = ~n19310 ;
  assign n19311 = n186 & n40598 ;
  assign n18506 = n18497 | n18498 ;
  assign n40599 = ~n18506 ;
  assign n18602 = n40599 & n144 ;
  assign n18603 = n17985 | n18602 ;
  assign n40600 = ~n18498 ;
  assign n18504 = n17985 & n40600 ;
  assign n18505 = n40214 & n18504 ;
  assign n18606 = n18505 & n144 ;
  assign n40601 = ~n18606 ;
  assign n18607 = n18603 & n40601 ;
  assign n19253 = n40580 & n19245 ;
  assign n19254 = n18689 | n19253 ;
  assign n40602 = ~n19247 ;
  assign n19255 = n40602 & n19254 ;
  assign n40603 = ~n19255 ;
  assign n19256 = n184 & n40603 ;
  assign n19257 = n40587 & n19254 ;
  assign n19286 = n19257 | n19285 ;
  assign n40604 = ~n19256 ;
  assign n19287 = n40604 & n19286 ;
  assign n40605 = ~n19287 ;
  assign n19288 = n185 & n40605 ;
  assign n19289 = n186 | n19288 ;
  assign n40606 = ~n19289 ;
  assign n19323 = n40606 & n19309 ;
  assign n19324 = n18607 | n19323 ;
  assign n40607 = ~n19311 ;
  assign n19325 = n40607 & n19324 ;
  assign n40608 = ~n19325 ;
  assign n19326 = n187 & n40608 ;
  assign n18503 = n17993 & n40224 ;
  assign n40609 = ~n18519 ;
  assign n18532 = n18503 & n40609 ;
  assign n18601 = n18532 & n144 ;
  assign n18533 = n18501 | n18519 ;
  assign n40610 = ~n18533 ;
  assign n18619 = n40610 & n144 ;
  assign n18620 = n17993 | n18619 ;
  assign n40611 = ~n18601 ;
  assign n18621 = n40611 & n18620 ;
  assign n19312 = n528 | n19311 ;
  assign n40612 = ~n19312 ;
  assign n19327 = n40612 & n19324 ;
  assign n19328 = n18621 | n19327 ;
  assign n40613 = ~n19326 ;
  assign n19329 = n40613 & n19328 ;
  assign n40614 = ~n19329 ;
  assign n19330 = n413 & n40614 ;
  assign n40615 = ~n18523 ;
  assign n18529 = n17996 & n40615 ;
  assign n18530 = n40230 & n18529 ;
  assign n18600 = n18530 & n144 ;
  assign n18531 = n18522 | n18523 ;
  assign n40616 = ~n18531 ;
  assign n18750 = n40616 & n144 ;
  assign n18751 = n17996 | n18750 ;
  assign n40617 = ~n18600 ;
  assign n18752 = n40617 & n18751 ;
  assign n19291 = n40596 & n19286 ;
  assign n19292 = n18768 | n19291 ;
  assign n40618 = ~n19288 ;
  assign n19293 = n40618 & n19292 ;
  assign n40619 = ~n19293 ;
  assign n19294 = n186 & n40619 ;
  assign n19295 = n40606 & n19292 ;
  assign n19296 = n18607 | n19295 ;
  assign n40620 = ~n19294 ;
  assign n19297 = n40620 & n19296 ;
  assign n40621 = ~n19297 ;
  assign n19298 = n528 & n40621 ;
  assign n19299 = n413 | n19298 ;
  assign n40622 = ~n19299 ;
  assign n19342 = n40622 & n19328 ;
  assign n19343 = n18752 | n19342 ;
  assign n40623 = ~n19330 ;
  assign n19344 = n40623 & n19343 ;
  assign n40624 = ~n19344 ;
  assign n19345 = n189 & n40624 ;
  assign n18555 = n18526 | n18543 ;
  assign n40625 = ~n18555 ;
  assign n18685 = n40625 & n144 ;
  assign n18686 = n17999 | n18685 ;
  assign n18527 = n17999 & n40240 ;
  assign n40626 = ~n18543 ;
  assign n18554 = n18527 & n40626 ;
  assign n18726 = n18554 & n144 ;
  assign n40627 = ~n18726 ;
  assign n18727 = n18686 & n40627 ;
  assign n19331 = n189 | n19330 ;
  assign n40628 = ~n19331 ;
  assign n19346 = n40628 & n19343 ;
  assign n19347 = n18727 | n19346 ;
  assign n40629 = ~n19345 ;
  assign n19348 = n40629 & n19347 ;
  assign n40630 = ~n19348 ;
  assign n19349 = n190 & n40630 ;
  assign n19276 = n40245 & n18561 ;
  assign n40631 = ~n19276 ;
  assign n19277 = n17914 & n40631 ;
  assign n19278 = n40246 & n19277 ;
  assign n19279 = n144 & n19278 ;
  assign n19280 = n18546 | n19276 ;
  assign n40632 = ~n19280 ;
  assign n19281 = n144 & n40632 ;
  assign n19282 = n17914 | n19281 ;
  assign n40633 = ~n19279 ;
  assign n19283 = n40633 & n19282 ;
  assign n19313 = n19296 & n40612 ;
  assign n19314 = n18621 | n19313 ;
  assign n40634 = ~n19298 ;
  assign n19315 = n40634 & n19314 ;
  assign n40635 = ~n19315 ;
  assign n19316 = n188 & n40635 ;
  assign n19317 = n40622 & n19314 ;
  assign n19318 = n18752 | n19317 ;
  assign n40636 = ~n19316 ;
  assign n19319 = n40636 & n19318 ;
  assign n40637 = ~n19319 ;
  assign n19320 = n189 & n40637 ;
  assign n19321 = n190 | n19320 ;
  assign n40638 = ~n19321 ;
  assign n19387 = n40638 & n19347 ;
  assign n19388 = n19283 | n19387 ;
  assign n40639 = ~n19349 ;
  assign n19389 = n40639 & n19388 ;
  assign n40640 = ~n19389 ;
  assign n19390 = n191 & n40640 ;
  assign n18570 = n18550 | n18565 ;
  assign n40641 = ~n18570 ;
  assign n18639 = n40641 & n144 ;
  assign n18640 = n18002 | n18639 ;
  assign n18553 = n18002 & n40260 ;
  assign n40642 = ~n18565 ;
  assign n18569 = n18553 & n40642 ;
  assign n19263 = n18569 & n18797 ;
  assign n40643 = ~n19263 ;
  assign n19264 = n18640 & n40643 ;
  assign n19350 = n191 | n19349 ;
  assign n40644 = ~n19350 ;
  assign n19391 = n40644 & n19388 ;
  assign n19392 = n19264 | n19391 ;
  assign n40645 = ~n19390 ;
  assign n19393 = n40645 & n19392 ;
  assign n19394 = n19273 | n19393 ;
  assign n19395 = n31336 & n19394 ;
  assign n18476 = n17997 | n18472 ;
  assign n40646 = ~n18476 ;
  assign n18477 = n18004 & n40646 ;
  assign n18478 = n40280 & n18477 ;
  assign n18577 = n18478 & n40281 ;
  assign n18589 = n18577 & n40282 ;
  assign n18581 = n192 & n18580 ;
  assign n40647 = ~n18005 ;
  assign n18729 = n40647 & n144 ;
  assign n40648 = ~n18729 ;
  assign n18730 = n18579 & n40648 ;
  assign n40649 = ~n18730 ;
  assign n18731 = n18581 & n40649 ;
  assign n18732 = n18589 | n18731 ;
  assign n19332 = n19318 & n40628 ;
  assign n19333 = n18727 | n19332 ;
  assign n40650 = ~n19320 ;
  assign n19334 = n40650 & n19333 ;
  assign n40651 = ~n19334 ;
  assign n19335 = n190 & n40651 ;
  assign n19336 = n40638 & n19333 ;
  assign n19337 = n19283 | n19336 ;
  assign n40652 = ~n19335 ;
  assign n19338 = n40652 & n19337 ;
  assign n40653 = ~n19338 ;
  assign n19339 = n287 & n40653 ;
  assign n40654 = ~n19339 ;
  assign n19340 = n19272 & n40654 ;
  assign n19396 = n19340 & n19392 ;
  assign n19397 = n18732 | n19396 ;
  assign n143 = n19395 | n19397 ;
  assign n19354 = n287 | n19349 ;
  assign n40655 = ~n19354 ;
  assign n19355 = n19337 & n40655 ;
  assign n19356 = n19264 | n19355 ;
  assign n19360 = n19340 & n19356 ;
  assign n19357 = n40654 & n19356 ;
  assign n19385 = n19272 | n19357 ;
  assign n40656 = ~n19385 ;
  assign n19604 = n40656 & n143 ;
  assign n19605 = n19360 | n19604 ;
  assign n19341 = n19264 & n40654 ;
  assign n19351 = n19337 & n40644 ;
  assign n40657 = ~n19351 ;
  assign n19352 = n19341 & n40657 ;
  assign n20032 = n19352 & n143 ;
  assign n19353 = n19339 | n19351 ;
  assign n40658 = ~n19353 ;
  assign n20066 = n40658 & n143 ;
  assign n20067 = n19264 | n20066 ;
  assign n40659 = ~n20032 ;
  assign n20068 = n40659 & n20067 ;
  assign n20069 = n19605 | n20068 ;
  assign n40660 = ~n19387 ;
  assign n20072 = n19283 & n40660 ;
  assign n20073 = n40639 & n20072 ;
  assign n20074 = n143 & n20073 ;
  assign n20075 = n19349 | n19387 ;
  assign n40661 = ~n20075 ;
  assign n20076 = n143 & n40661 ;
  assign n20077 = n19283 | n20076 ;
  assign n40662 = ~n20074 ;
  assign n20078 = n40662 & n20077 ;
  assign n230 = x26 | x27 ;
  assign n40663 = ~x28 ;
  assign n232 = n40663 & n230 ;
  assign n19358 = n19273 | n19357 ;
  assign n19359 = n31336 & n19358 ;
  assign n19361 = n18732 | n19360 ;
  assign n19362 = n19359 | n19361 ;
  assign n40664 = ~n19362 ;
  assign n19371 = x28 & n40664 ;
  assign n19372 = n232 | n19371 ;
  assign n40665 = ~n19372 ;
  assign n19373 = n18797 & n40665 ;
  assign n231 = x28 | n230 ;
  assign n18479 = n231 & n40279 ;
  assign n18480 = n40280 & n18479 ;
  assign n18578 = n18480 & n40281 ;
  assign n18591 = n18578 & n40282 ;
  assign n19435 = x28 & n143 ;
  assign n40666 = ~n19435 ;
  assign n19436 = n18591 & n40666 ;
  assign n19503 = n40663 & n143 ;
  assign n40667 = ~n19503 ;
  assign n19504 = x29 & n40667 ;
  assign n40668 = ~n227 ;
  assign n19510 = n40668 & n143 ;
  assign n19523 = n19504 | n19510 ;
  assign n19525 = n19436 | n19523 ;
  assign n40669 = ~n19373 ;
  assign n19526 = n40669 & n19525 ;
  assign n40670 = ~n19526 ;
  assign n19527 = n145 & n40670 ;
  assign n19486 = n231 & n40666 ;
  assign n40671 = ~n19486 ;
  assign n19487 = n144 & n40671 ;
  assign n19488 = n145 | n19487 ;
  assign n40672 = ~n19488 ;
  assign n19529 = n40672 & n19525 ;
  assign n40673 = ~n18589 ;
  assign n18728 = n40673 & n144 ;
  assign n40674 = ~n18731 ;
  assign n18733 = n18728 & n40674 ;
  assign n40675 = ~n19360 ;
  assign n19376 = n18733 & n40675 ;
  assign n40676 = ~n19359 ;
  assign n19377 = n40676 & n19376 ;
  assign n19378 = x30 | n19377 ;
  assign n19511 = n19378 | n19510 ;
  assign n19530 = n19377 | n19510 ;
  assign n19531 = x30 & n19530 ;
  assign n40677 = ~n19531 ;
  assign n19532 = n19511 & n40677 ;
  assign n19533 = n19529 | n19532 ;
  assign n40678 = ~n19527 ;
  assign n19534 = n40678 & n19533 ;
  assign n40679 = ~n19534 ;
  assign n19535 = n146 & n40679 ;
  assign n18809 = n18675 | n18800 ;
  assign n40680 = ~n18809 ;
  assign n19465 = n40680 & n143 ;
  assign n19466 = n18694 | n19465 ;
  assign n18810 = n18694 & n40680 ;
  assign n19481 = n18810 & n143 ;
  assign n40681 = ~n19481 ;
  assign n19482 = n19466 & n40681 ;
  assign n19528 = n146 | n19527 ;
  assign n19374 = n145 | n19373 ;
  assign n40682 = ~n19374 ;
  assign n19538 = n40682 & n19525 ;
  assign n19545 = n19532 | n19538 ;
  assign n40683 = ~n19528 ;
  assign n19564 = n40683 & n19545 ;
  assign n19565 = n19482 | n19564 ;
  assign n40684 = ~n19535 ;
  assign n19566 = n40684 & n19565 ;
  assign n40685 = ~n19566 ;
  assign n19567 = n147 & n40685 ;
  assign n19262 = n18702 | n18812 ;
  assign n40686 = ~n19262 ;
  assign n19426 = n40686 & n143 ;
  assign n19427 = n18699 | n19426 ;
  assign n40687 = ~n18812 ;
  assign n19260 = n18699 & n40687 ;
  assign n40688 = ~n18702 ;
  assign n19261 = n40688 & n19260 ;
  assign n19491 = n19261 & n143 ;
  assign n40689 = ~n19491 ;
  assign n19492 = n19427 & n40689 ;
  assign n19537 = n16322 | n19535 ;
  assign n40690 = ~n19537 ;
  assign n19568 = n40690 & n19565 ;
  assign n19569 = n19492 | n19568 ;
  assign n40691 = ~n19567 ;
  assign n19570 = n40691 & n19569 ;
  assign n40692 = ~n19570 ;
  assign n19571 = n15807 & n40692 ;
  assign n19259 = n18806 | n18814 ;
  assign n40693 = ~n19259 ;
  assign n19454 = n40693 & n143 ;
  assign n19455 = n18711 | n19454 ;
  assign n18807 = n18711 & n40314 ;
  assign n40694 = ~n18814 ;
  assign n19258 = n18807 & n40694 ;
  assign n19479 = n19258 & n143 ;
  assign n40695 = ~n19479 ;
  assign n19480 = n19455 & n40695 ;
  assign n19375 = n144 & n40665 ;
  assign n40696 = ~n19375 ;
  assign n19539 = n40696 & n19525 ;
  assign n40697 = ~n19539 ;
  assign n19540 = n145 & n40697 ;
  assign n19541 = n146 | n19540 ;
  assign n40698 = ~n19541 ;
  assign n19546 = n40698 & n19545 ;
  assign n19547 = n19482 | n19546 ;
  assign n19548 = n40684 & n19547 ;
  assign n40699 = ~n19548 ;
  assign n19549 = n16322 & n40699 ;
  assign n19550 = n148 | n19549 ;
  assign n40700 = ~n19550 ;
  assign n19584 = n40700 & n19569 ;
  assign n19585 = n19480 | n19584 ;
  assign n40701 = ~n19571 ;
  assign n19586 = n40701 & n19585 ;
  assign n40702 = ~n19586 ;
  assign n19587 = n149 & n40702 ;
  assign n40703 = ~n18819 ;
  assign n18828 = n18746 & n40703 ;
  assign n18829 = n40302 & n18828 ;
  assign n19369 = n18829 & n19362 ;
  assign n18830 = n18817 | n18819 ;
  assign n40704 = ~n18830 ;
  assign n19451 = n40704 & n143 ;
  assign n19452 = n18746 | n19451 ;
  assign n40705 = ~n19369 ;
  assign n19453 = n40705 & n19452 ;
  assign n19572 = n149 | n19571 ;
  assign n40706 = ~n19572 ;
  assign n19588 = n40706 & n19585 ;
  assign n19589 = n19453 | n19588 ;
  assign n40707 = ~n19587 ;
  assign n19590 = n40707 & n19589 ;
  assign n40708 = ~n19590 ;
  assign n19591 = n150 & n40708 ;
  assign n19551 = n40690 & n19547 ;
  assign n19552 = n19492 | n19551 ;
  assign n40709 = ~n19549 ;
  assign n19553 = n40709 & n19552 ;
  assign n40710 = ~n19553 ;
  assign n19554 = n148 & n40710 ;
  assign n19555 = n40700 & n19552 ;
  assign n19556 = n19480 | n19555 ;
  assign n40711 = ~n19554 ;
  assign n19557 = n40711 & n19556 ;
  assign n40712 = ~n19557 ;
  assign n19558 = n149 & n40712 ;
  assign n19559 = n150 | n19558 ;
  assign n40713 = ~n19559 ;
  assign n19593 = n40713 & n19589 ;
  assign n18854 = n18725 & n40330 ;
  assign n40714 = ~n18823 ;
  assign n18855 = n40714 & n18854 ;
  assign n19368 = n18855 & n19362 ;
  assign n18853 = n18823 | n18838 ;
  assign n40715 = ~n18853 ;
  assign n19613 = n40715 & n143 ;
  assign n19614 = n18725 | n19613 ;
  assign n40716 = ~n19368 ;
  assign n19615 = n40716 & n19614 ;
  assign n19616 = n19593 | n19615 ;
  assign n40717 = ~n19591 ;
  assign n19617 = n40717 & n19616 ;
  assign n40718 = ~n19617 ;
  assign n19618 = n151 & n40718 ;
  assign n18852 = n18826 | n18840 ;
  assign n40719 = ~n18852 ;
  assign n19402 = n40719 & n143 ;
  assign n19403 = n18693 | n19402 ;
  assign n40720 = ~n18840 ;
  assign n18850 = n18693 & n40720 ;
  assign n18851 = n40319 & n18850 ;
  assign n19469 = n18851 & n143 ;
  assign n40721 = ~n19469 ;
  assign n19470 = n19403 & n40721 ;
  assign n19592 = n151 | n19591 ;
  assign n40722 = ~n19592 ;
  assign n19619 = n40722 & n19616 ;
  assign n19620 = n19470 | n19619 ;
  assign n40723 = ~n19618 ;
  assign n19621 = n40723 & n19620 ;
  assign n40724 = ~n19621 ;
  assign n19622 = n13079 & n40724 ;
  assign n18849 = n18843 | n18844 ;
  assign n40725 = ~n18849 ;
  assign n19508 = n40725 & n143 ;
  assign n19509 = n18638 | n19508 ;
  assign n18878 = n18638 & n40346 ;
  assign n40726 = ~n18844 ;
  assign n18879 = n40726 & n18878 ;
  assign n19609 = n18879 & n143 ;
  assign n40727 = ~n19609 ;
  assign n19610 = n19509 & n40727 ;
  assign n19573 = n19556 & n40706 ;
  assign n19574 = n19453 | n19573 ;
  assign n40728 = ~n19558 ;
  assign n19575 = n40728 & n19574 ;
  assign n40729 = ~n19575 ;
  assign n19576 = n150 & n40729 ;
  assign n19577 = n40713 & n19574 ;
  assign n19625 = n19577 | n19615 ;
  assign n40730 = ~n19576 ;
  assign n19626 = n40730 & n19625 ;
  assign n40731 = ~n19626 ;
  assign n19627 = n13662 & n40731 ;
  assign n19628 = n152 | n19627 ;
  assign n40732 = ~n19628 ;
  assign n19629 = n19620 & n40732 ;
  assign n19630 = n19610 | n19629 ;
  assign n40733 = ~n19622 ;
  assign n19631 = n40733 & n19630 ;
  assign n40734 = ~n19631 ;
  assign n19632 = n153 & n40734 ;
  assign n40735 = ~n18865 ;
  assign n18875 = n18708 & n40735 ;
  assign n18876 = n40335 & n18875 ;
  assign n19432 = n18876 & n143 ;
  assign n18877 = n18847 | n18865 ;
  assign n40736 = ~n18877 ;
  assign n19516 = n40736 & n143 ;
  assign n19517 = n18708 | n19516 ;
  assign n40737 = ~n19432 ;
  assign n19518 = n40737 & n19517 ;
  assign n19623 = n153 | n19622 ;
  assign n40738 = ~n19623 ;
  assign n19633 = n40738 & n19630 ;
  assign n19634 = n19518 | n19633 ;
  assign n40739 = ~n19632 ;
  assign n19635 = n40739 & n19634 ;
  assign n40740 = ~n19635 ;
  assign n19636 = n154 & n40740 ;
  assign n18874 = n18868 | n18869 ;
  assign n40741 = ~n18874 ;
  assign n19498 = n40741 & n143 ;
  assign n19499 = n18718 | n19498 ;
  assign n18902 = n18718 & n40362 ;
  assign n40742 = ~n18869 ;
  assign n18903 = n40742 & n18902 ;
  assign n19519 = n18903 & n143 ;
  assign n40743 = ~n19519 ;
  assign n19520 = n19499 & n40743 ;
  assign n19639 = n40722 & n19625 ;
  assign n19640 = n19470 | n19639 ;
  assign n40744 = ~n19627 ;
  assign n19641 = n40744 & n19640 ;
  assign n40745 = ~n19641 ;
  assign n19642 = n152 & n40745 ;
  assign n19643 = n40732 & n19640 ;
  assign n19644 = n19610 | n19643 ;
  assign n40746 = ~n19642 ;
  assign n19645 = n40746 & n19644 ;
  assign n40747 = ~n19645 ;
  assign n19646 = n153 & n40747 ;
  assign n19647 = n154 | n19646 ;
  assign n40748 = ~n19647 ;
  assign n19648 = n19634 & n40748 ;
  assign n19649 = n19520 | n19648 ;
  assign n40749 = ~n19636 ;
  assign n19650 = n40749 & n19649 ;
  assign n40750 = ~n19650 ;
  assign n19651 = n155 & n40750 ;
  assign n40751 = ~n18889 ;
  assign n18899 = n18651 & n40751 ;
  assign n18900 = n40351 & n18899 ;
  assign n19367 = n18900 & n19362 ;
  assign n18901 = n18872 | n18889 ;
  assign n40752 = ~n18901 ;
  assign n19606 = n40752 & n143 ;
  assign n19607 = n18651 | n19606 ;
  assign n40753 = ~n19367 ;
  assign n19608 = n40753 & n19607 ;
  assign n19637 = n11067 | n19636 ;
  assign n40754 = ~n19637 ;
  assign n19652 = n40754 & n19649 ;
  assign n19653 = n19608 | n19652 ;
  assign n40755 = ~n19651 ;
  assign n19654 = n40755 & n19653 ;
  assign n40756 = ~n19654 ;
  assign n19655 = n10657 & n40756 ;
  assign n18898 = n18892 | n18893 ;
  assign n40757 = ~n18898 ;
  assign n19493 = n40757 & n143 ;
  assign n19494 = n18787 | n19493 ;
  assign n18926 = n18787 & n40378 ;
  assign n40758 = ~n18893 ;
  assign n18927 = n40758 & n18926 ;
  assign n19611 = n18927 & n143 ;
  assign n40759 = ~n19611 ;
  assign n19612 = n19494 & n40759 ;
  assign n19658 = n40738 & n19644 ;
  assign n19659 = n19518 | n19658 ;
  assign n40760 = ~n19646 ;
  assign n19660 = n40760 & n19659 ;
  assign n40761 = ~n19660 ;
  assign n19661 = n154 & n40761 ;
  assign n19662 = n40748 & n19659 ;
  assign n19663 = n19520 | n19662 ;
  assign n40762 = ~n19661 ;
  assign n19664 = n40762 & n19663 ;
  assign n40763 = ~n19664 ;
  assign n19665 = n11067 & n40763 ;
  assign n19666 = n10657 | n19665 ;
  assign n40764 = ~n19666 ;
  assign n19667 = n19653 & n40764 ;
  assign n19668 = n19612 | n19667 ;
  assign n40765 = ~n19655 ;
  assign n19669 = n40765 & n19668 ;
  assign n40766 = ~n19669 ;
  assign n19670 = n157 & n40766 ;
  assign n18925 = n18896 | n18913 ;
  assign n40767 = ~n18925 ;
  assign n19447 = n40767 & n143 ;
  assign n19448 = n18742 | n19447 ;
  assign n40768 = ~n18913 ;
  assign n18923 = n18742 & n40768 ;
  assign n18924 = n40367 & n18923 ;
  assign n19514 = n18924 & n143 ;
  assign n40769 = ~n19514 ;
  assign n19515 = n19448 & n40769 ;
  assign n19656 = n157 | n19655 ;
  assign n40770 = ~n19656 ;
  assign n19671 = n40770 & n19668 ;
  assign n19672 = n19515 | n19671 ;
  assign n40771 = ~n19670 ;
  assign n19673 = n40771 & n19672 ;
  assign n40772 = ~n19673 ;
  assign n19674 = n158 & n40772 ;
  assign n18950 = n18672 & n40394 ;
  assign n40773 = ~n18917 ;
  assign n18951 = n40773 & n18950 ;
  assign n19366 = n18951 & n19362 ;
  assign n18922 = n18916 | n18917 ;
  assign n40774 = ~n18922 ;
  assign n19416 = n40774 & n143 ;
  assign n19417 = n18672 | n19416 ;
  assign n40775 = ~n19366 ;
  assign n19418 = n40775 & n19417 ;
  assign n19677 = n40754 & n19663 ;
  assign n19678 = n19608 | n19677 ;
  assign n40776 = ~n19665 ;
  assign n19679 = n40776 & n19678 ;
  assign n40777 = ~n19679 ;
  assign n19680 = n156 & n40777 ;
  assign n19681 = n40764 & n19678 ;
  assign n19682 = n19612 | n19681 ;
  assign n40778 = ~n19680 ;
  assign n19683 = n40778 & n19682 ;
  assign n40779 = ~n19683 ;
  assign n19684 = n157 & n40779 ;
  assign n19685 = n158 | n19684 ;
  assign n40780 = ~n19685 ;
  assign n19686 = n19672 & n40780 ;
  assign n19687 = n19418 | n19686 ;
  assign n40781 = ~n19674 ;
  assign n19688 = n40781 & n19687 ;
  assign n40782 = ~n19688 ;
  assign n19689 = n159 & n40782 ;
  assign n19675 = n8857 | n19674 ;
  assign n40783 = ~n19675 ;
  assign n19690 = n40783 & n19687 ;
  assign n40784 = ~n18937 ;
  assign n18947 = n18716 & n40784 ;
  assign n18948 = n40383 & n18947 ;
  assign n19724 = n18948 & n143 ;
  assign n18949 = n18920 | n18937 ;
  assign n40785 = ~n18949 ;
  assign n19725 = n40785 & n143 ;
  assign n19726 = n18716 | n19725 ;
  assign n40786 = ~n19724 ;
  assign n19727 = n40786 & n19726 ;
  assign n19728 = n19690 | n19727 ;
  assign n40787 = ~n19689 ;
  assign n19729 = n40787 & n19728 ;
  assign n40788 = ~n19729 ;
  assign n19730 = n8534 & n40788 ;
  assign n18946 = n18940 | n18941 ;
  assign n40789 = ~n18946 ;
  assign n19458 = n40789 & n143 ;
  assign n19459 = n18714 | n19458 ;
  assign n18974 = n18714 & n40410 ;
  assign n40790 = ~n18941 ;
  assign n18975 = n40790 & n18974 ;
  assign n19460 = n18975 & n143 ;
  assign n40791 = ~n19460 ;
  assign n19461 = n19459 & n40791 ;
  assign n19691 = n40770 & n19682 ;
  assign n19692 = n19515 | n19691 ;
  assign n40792 = ~n19684 ;
  assign n19693 = n40792 & n19692 ;
  assign n40793 = ~n19693 ;
  assign n19694 = n158 & n40793 ;
  assign n19695 = n40780 & n19692 ;
  assign n19696 = n19418 | n19695 ;
  assign n40794 = ~n19694 ;
  assign n19697 = n40794 & n19696 ;
  assign n40795 = ~n19697 ;
  assign n19698 = n8857 & n40795 ;
  assign n19699 = n160 | n19698 ;
  assign n40796 = ~n19699 ;
  assign n19733 = n40796 & n19728 ;
  assign n19734 = n19461 | n19733 ;
  assign n40797 = ~n19730 ;
  assign n19735 = n40797 & n19734 ;
  assign n40798 = ~n19735 ;
  assign n19736 = n161 & n40798 ;
  assign n18973 = n18944 | n18961 ;
  assign n40799 = ~n18973 ;
  assign n19443 = n40799 & n143 ;
  assign n19444 = n18775 | n19443 ;
  assign n40800 = ~n18961 ;
  assign n18971 = n18775 & n40800 ;
  assign n18972 = n40399 & n18971 ;
  assign n19445 = n18972 & n143 ;
  assign n40801 = ~n19445 ;
  assign n19446 = n19444 & n40801 ;
  assign n19731 = n161 | n19730 ;
  assign n40802 = ~n19731 ;
  assign n19737 = n40802 & n19734 ;
  assign n19738 = n19446 | n19737 ;
  assign n40803 = ~n19736 ;
  assign n19739 = n40803 & n19738 ;
  assign n40804 = ~n19739 ;
  assign n19740 = n162 & n40804 ;
  assign n18970 = n18964 | n18965 ;
  assign n40805 = ~n18970 ;
  assign n19439 = n40805 & n143 ;
  assign n19440 = n18759 | n19439 ;
  assign n18997 = n18759 & n40426 ;
  assign n40806 = ~n18965 ;
  assign n18998 = n40806 & n18997 ;
  assign n19441 = n18998 & n143 ;
  assign n40807 = ~n19441 ;
  assign n19442 = n19440 & n40807 ;
  assign n19700 = n40783 & n19696 ;
  assign n19743 = n19700 | n19727 ;
  assign n40808 = ~n19698 ;
  assign n19744 = n40808 & n19743 ;
  assign n40809 = ~n19744 ;
  assign n19745 = n160 & n40809 ;
  assign n19746 = n40796 & n19743 ;
  assign n19747 = n19461 | n19746 ;
  assign n40810 = ~n19745 ;
  assign n19748 = n40810 & n19747 ;
  assign n40811 = ~n19748 ;
  assign n19749 = n161 & n40811 ;
  assign n19750 = n162 | n19749 ;
  assign n40812 = ~n19750 ;
  assign n19751 = n19738 & n40812 ;
  assign n19752 = n19442 | n19751 ;
  assign n40813 = ~n19740 ;
  assign n19753 = n40813 & n19752 ;
  assign n40814 = ~n19753 ;
  assign n19754 = n163 & n40814 ;
  assign n18994 = n18968 | n18985 ;
  assign n40815 = ~n18994 ;
  assign n19433 = n40815 & n143 ;
  assign n19434 = n18756 | n19433 ;
  assign n40816 = ~n18985 ;
  assign n18995 = n18756 & n40816 ;
  assign n18996 = n40415 & n18995 ;
  assign n19467 = n18996 & n143 ;
  assign n40817 = ~n19467 ;
  assign n19468 = n19434 & n40817 ;
  assign n19741 = n6889 | n19740 ;
  assign n40818 = ~n19741 ;
  assign n19755 = n40818 & n19752 ;
  assign n19756 = n19468 | n19755 ;
  assign n40819 = ~n19754 ;
  assign n19757 = n40819 & n19756 ;
  assign n40820 = ~n19757 ;
  assign n19758 = n6600 & n40820 ;
  assign n19023 = n18989 | n19006 ;
  assign n40821 = ~n19023 ;
  assign n19521 = n40821 & n143 ;
  assign n19522 = n18667 | n19521 ;
  assign n19021 = n18667 & n40442 ;
  assign n40822 = ~n18989 ;
  assign n19022 = n40822 & n19021 ;
  assign n19599 = n19022 & n143 ;
  assign n40823 = ~n19599 ;
  assign n19600 = n19522 & n40823 ;
  assign n19761 = n40802 & n19747 ;
  assign n19762 = n19446 | n19761 ;
  assign n40824 = ~n19749 ;
  assign n19763 = n40824 & n19762 ;
  assign n40825 = ~n19763 ;
  assign n19764 = n162 & n40825 ;
  assign n19765 = n40812 & n19762 ;
  assign n19766 = n19442 | n19765 ;
  assign n40826 = ~n19764 ;
  assign n19767 = n40826 & n19766 ;
  assign n40827 = ~n19767 ;
  assign n19768 = n6889 & n40827 ;
  assign n19769 = n6600 | n19768 ;
  assign n40828 = ~n19769 ;
  assign n19770 = n19756 & n40828 ;
  assign n19771 = n19600 | n19770 ;
  assign n40829 = ~n19758 ;
  assign n19772 = n40829 & n19771 ;
  assign n40830 = ~n19772 ;
  assign n19773 = n165 & n40830 ;
  assign n40831 = ~n19008 ;
  assign n19018 = n18761 & n40831 ;
  assign n19019 = n40431 & n19018 ;
  assign n19431 = n19019 & n143 ;
  assign n19020 = n18992 | n19008 ;
  assign n40832 = ~n19020 ;
  assign n19462 = n40832 & n143 ;
  assign n19463 = n18761 | n19462 ;
  assign n40833 = ~n19431 ;
  assign n19464 = n40833 & n19463 ;
  assign n19759 = n165 | n19758 ;
  assign n40834 = ~n19759 ;
  assign n19774 = n40834 & n19771 ;
  assign n19775 = n19464 | n19774 ;
  assign n40835 = ~n19773 ;
  assign n19776 = n40835 & n19775 ;
  assign n40836 = ~n19776 ;
  assign n19777 = n166 & n40836 ;
  assign n19046 = n18739 & n40458 ;
  assign n40837 = ~n19012 ;
  assign n19047 = n40837 & n19046 ;
  assign n19365 = n19047 & n19362 ;
  assign n19017 = n19011 | n19012 ;
  assign n40838 = ~n19017 ;
  assign n19423 = n40838 & n143 ;
  assign n19424 = n18739 | n19423 ;
  assign n40839 = ~n19365 ;
  assign n19425 = n40839 & n19424 ;
  assign n19780 = n40818 & n19766 ;
  assign n19781 = n19468 | n19780 ;
  assign n40840 = ~n19768 ;
  assign n19782 = n40840 & n19781 ;
  assign n40841 = ~n19782 ;
  assign n19783 = n164 & n40841 ;
  assign n19784 = n40828 & n19781 ;
  assign n19787 = n19600 | n19784 ;
  assign n40842 = ~n19783 ;
  assign n19788 = n40842 & n19787 ;
  assign n40843 = ~n19788 ;
  assign n19789 = n165 & n40843 ;
  assign n19790 = n166 | n19789 ;
  assign n40844 = ~n19790 ;
  assign n19791 = n19775 & n40844 ;
  assign n19792 = n19425 | n19791 ;
  assign n40845 = ~n19777 ;
  assign n19793 = n40845 & n19792 ;
  assign n40846 = ~n19793 ;
  assign n19794 = n167 & n40846 ;
  assign n40847 = ~n19033 ;
  assign n19043 = n18773 & n40847 ;
  assign n19044 = n40447 & n19043 ;
  assign n19422 = n19044 & n143 ;
  assign n19045 = n19015 | n19033 ;
  assign n40848 = ~n19045 ;
  assign n19495 = n40848 & n143 ;
  assign n19496 = n18773 | n19495 ;
  assign n40849 = ~n19422 ;
  assign n19497 = n40849 & n19496 ;
  assign n19778 = n5352 | n19777 ;
  assign n40850 = ~n19778 ;
  assign n19795 = n40850 & n19792 ;
  assign n19796 = n19497 | n19795 ;
  assign n40851 = ~n19794 ;
  assign n19797 = n40851 & n19796 ;
  assign n40852 = ~n19797 ;
  assign n19798 = n4934 & n40852 ;
  assign n19070 = n18785 & n40474 ;
  assign n40853 = ~n19037 ;
  assign n19071 = n40853 & n19070 ;
  assign n19421 = n19071 & n143 ;
  assign n19042 = n19036 | n19037 ;
  assign n40854 = ~n19042 ;
  assign n19428 = n40854 & n143 ;
  assign n19429 = n18785 | n19428 ;
  assign n40855 = ~n19421 ;
  assign n19430 = n40855 & n19429 ;
  assign n19801 = n40834 & n19787 ;
  assign n19802 = n19464 | n19801 ;
  assign n40856 = ~n19789 ;
  assign n19803 = n40856 & n19802 ;
  assign n40857 = ~n19803 ;
  assign n19804 = n166 & n40857 ;
  assign n19805 = n40844 & n19802 ;
  assign n19806 = n19425 | n19805 ;
  assign n40858 = ~n19804 ;
  assign n19807 = n40858 & n19806 ;
  assign n40859 = ~n19807 ;
  assign n19808 = n5352 & n40859 ;
  assign n19809 = n4934 | n19808 ;
  assign n40860 = ~n19809 ;
  assign n19810 = n19796 & n40860 ;
  assign n19811 = n19430 | n19810 ;
  assign n40861 = ~n19798 ;
  assign n19812 = n40861 & n19811 ;
  assign n40862 = ~n19812 ;
  assign n19813 = n169 & n40862 ;
  assign n19069 = n19040 | n19057 ;
  assign n40863 = ~n19069 ;
  assign n19419 = n40863 & n143 ;
  assign n19420 = n18789 | n19419 ;
  assign n40864 = ~n19057 ;
  assign n19067 = n18789 & n40864 ;
  assign n19068 = n40463 & n19067 ;
  assign n19506 = n19068 & n143 ;
  assign n40865 = ~n19506 ;
  assign n19507 = n19420 & n40865 ;
  assign n19799 = n169 | n19798 ;
  assign n40866 = ~n19799 ;
  assign n19814 = n40866 & n19811 ;
  assign n19815 = n19507 | n19814 ;
  assign n40867 = ~n19813 ;
  assign n19816 = n40867 & n19815 ;
  assign n40868 = ~n19816 ;
  assign n19817 = n170 & n40868 ;
  assign n19066 = n19060 | n19061 ;
  assign n40869 = ~n19066 ;
  assign n19449 = n40869 & n143 ;
  assign n19450 = n18778 | n19449 ;
  assign n19093 = n18778 & n40490 ;
  assign n40870 = ~n19061 ;
  assign n19094 = n40870 & n19093 ;
  assign n19471 = n19094 & n143 ;
  assign n40871 = ~n19471 ;
  assign n19472 = n19450 & n40871 ;
  assign n19820 = n40850 & n19806 ;
  assign n19821 = n19497 | n19820 ;
  assign n40872 = ~n19808 ;
  assign n19822 = n40872 & n19821 ;
  assign n40873 = ~n19822 ;
  assign n19823 = n168 & n40873 ;
  assign n19824 = n40860 & n19821 ;
  assign n19825 = n19430 | n19824 ;
  assign n40874 = ~n19823 ;
  assign n19826 = n40874 & n19825 ;
  assign n40875 = ~n19826 ;
  assign n19827 = n169 & n40875 ;
  assign n19828 = n170 | n19827 ;
  assign n40876 = ~n19828 ;
  assign n19829 = n19815 & n40876 ;
  assign n19830 = n19472 | n19829 ;
  assign n40877 = ~n19817 ;
  assign n19831 = n40877 & n19830 ;
  assign n40878 = ~n19831 ;
  assign n19832 = n171 & n40878 ;
  assign n19092 = n19064 | n19081 ;
  assign n40879 = ~n19092 ;
  assign n19412 = n40879 & n143 ;
  assign n19413 = n18678 | n19412 ;
  assign n40880 = ~n19081 ;
  assign n19090 = n18678 & n40880 ;
  assign n19091 = n40479 & n19090 ;
  assign n19456 = n19091 & n143 ;
  assign n40881 = ~n19456 ;
  assign n19457 = n19413 & n40881 ;
  assign n19818 = n3940 | n19817 ;
  assign n40882 = ~n19818 ;
  assign n19833 = n40882 & n19830 ;
  assign n19834 = n19457 | n19833 ;
  assign n40883 = ~n19832 ;
  assign n19835 = n40883 & n19834 ;
  assign n40884 = ~n19835 ;
  assign n19836 = n3631 & n40884 ;
  assign n19117 = n18792 & n40506 ;
  assign n40885 = ~n19085 ;
  assign n19118 = n40885 & n19117 ;
  assign n19408 = n19118 & n143 ;
  assign n19119 = n19085 | n19102 ;
  assign n40886 = ~n19119 ;
  assign n19596 = n40886 & n143 ;
  assign n19597 = n18792 | n19596 ;
  assign n40887 = ~n19408 ;
  assign n19598 = n40887 & n19597 ;
  assign n19839 = n40866 & n19825 ;
  assign n19840 = n19507 | n19839 ;
  assign n40888 = ~n19827 ;
  assign n19841 = n40888 & n19840 ;
  assign n40889 = ~n19841 ;
  assign n19842 = n170 & n40889 ;
  assign n19843 = n40876 & n19840 ;
  assign n19844 = n19472 | n19843 ;
  assign n40890 = ~n19842 ;
  assign n19845 = n40890 & n19844 ;
  assign n40891 = ~n19845 ;
  assign n19846 = n3940 & n40891 ;
  assign n19847 = n3631 | n19846 ;
  assign n40892 = ~n19847 ;
  assign n19848 = n19834 & n40892 ;
  assign n19849 = n19598 | n19848 ;
  assign n40893 = ~n19836 ;
  assign n19850 = n40893 & n19849 ;
  assign n40894 = ~n19850 ;
  assign n19851 = n173 & n40894 ;
  assign n19116 = n19088 | n19104 ;
  assign n40895 = ~n19116 ;
  assign n19404 = n40895 & n143 ;
  assign n19405 = n18782 | n19404 ;
  assign n40896 = ~n19104 ;
  assign n19114 = n18782 & n40896 ;
  assign n19115 = n40495 & n19114 ;
  assign n19406 = n19115 & n143 ;
  assign n40897 = ~n19406 ;
  assign n19407 = n19405 & n40897 ;
  assign n19837 = n173 | n19836 ;
  assign n40898 = ~n19837 ;
  assign n19852 = n40898 & n19849 ;
  assign n19853 = n19407 | n19852 ;
  assign n40899 = ~n19851 ;
  assign n19854 = n40899 & n19853 ;
  assign n40900 = ~n19854 ;
  assign n19855 = n174 & n40900 ;
  assign n19113 = n19107 | n19108 ;
  assign n40901 = ~n19113 ;
  assign n19400 = n40901 & n143 ;
  assign n19401 = n18794 | n19400 ;
  assign n19142 = n18794 & n40522 ;
  assign n40902 = ~n19108 ;
  assign n19143 = n40902 & n19142 ;
  assign n19414 = n19143 & n143 ;
  assign n40903 = ~n19414 ;
  assign n19415 = n19401 & n40903 ;
  assign n19858 = n40882 & n19844 ;
  assign n19859 = n19457 | n19858 ;
  assign n40904 = ~n19846 ;
  assign n19860 = n40904 & n19859 ;
  assign n40905 = ~n19860 ;
  assign n19861 = n172 & n40905 ;
  assign n19862 = n40892 & n19859 ;
  assign n19863 = n19598 | n19862 ;
  assign n40906 = ~n19861 ;
  assign n19864 = n40906 & n19863 ;
  assign n40907 = ~n19864 ;
  assign n19865 = n173 & n40907 ;
  assign n19866 = n174 | n19865 ;
  assign n40908 = ~n19866 ;
  assign n19867 = n19853 & n40908 ;
  assign n19868 = n19415 | n19867 ;
  assign n40909 = ~n19855 ;
  assign n19869 = n40909 & n19868 ;
  assign n40910 = ~n19869 ;
  assign n19870 = n175 & n40910 ;
  assign n40911 = ~n19129 ;
  assign n19139 = n18655 & n40911 ;
  assign n19140 = n40511 & n19139 ;
  assign n19399 = n19140 & n143 ;
  assign n19141 = n19111 | n19129 ;
  assign n40912 = ~n19141 ;
  assign n19483 = n40912 & n143 ;
  assign n19484 = n18655 | n19483 ;
  assign n40913 = ~n19399 ;
  assign n19485 = n40913 & n19484 ;
  assign n19856 = n2753 | n19855 ;
  assign n40914 = ~n19856 ;
  assign n19871 = n40914 & n19868 ;
  assign n19872 = n19485 | n19871 ;
  assign n40915 = ~n19870 ;
  assign n19873 = n40915 & n19872 ;
  assign n40916 = ~n19873 ;
  assign n19874 = n2431 & n40916 ;
  assign n19876 = n40898 & n19863 ;
  assign n19877 = n19407 | n19876 ;
  assign n40917 = ~n19865 ;
  assign n19878 = n40917 & n19877 ;
  assign n40918 = ~n19878 ;
  assign n19879 = n174 & n40918 ;
  assign n19880 = n40908 & n19877 ;
  assign n19881 = n19415 | n19880 ;
  assign n40919 = ~n19879 ;
  assign n19882 = n40919 & n19881 ;
  assign n40920 = ~n19882 ;
  assign n19883 = n2753 & n40920 ;
  assign n19884 = n2431 | n19883 ;
  assign n40921 = ~n19884 ;
  assign n19885 = n19872 & n40921 ;
  assign n19166 = n18649 & n40538 ;
  assign n40922 = ~n19133 ;
  assign n19167 = n40922 & n19166 ;
  assign n19505 = n19167 & n143 ;
  assign n19138 = n19132 | n19133 ;
  assign n40923 = ~n19138 ;
  assign n19932 = n40923 & n143 ;
  assign n19933 = n18649 | n19932 ;
  assign n40924 = ~n19505 ;
  assign n19934 = n40924 & n19933 ;
  assign n19943 = n19885 | n19934 ;
  assign n40925 = ~n19874 ;
  assign n19944 = n40925 & n19943 ;
  assign n40926 = ~n19944 ;
  assign n19945 = n177 & n40926 ;
  assign n19875 = n177 | n19874 ;
  assign n40927 = ~n19875 ;
  assign n19946 = n40927 & n19943 ;
  assign n40928 = ~n19153 ;
  assign n19163 = n18644 & n40928 ;
  assign n19164 = n40527 & n19163 ;
  assign n19950 = n19164 & n143 ;
  assign n19165 = n19136 | n19153 ;
  assign n40929 = ~n19165 ;
  assign n19951 = n40929 & n143 ;
  assign n19952 = n18644 | n19951 ;
  assign n40930 = ~n19950 ;
  assign n19953 = n40930 & n19952 ;
  assign n19954 = n19946 | n19953 ;
  assign n40931 = ~n19945 ;
  assign n19955 = n40931 & n19954 ;
  assign n40932 = ~n19955 ;
  assign n19956 = n178 & n40932 ;
  assign n19190 = n18635 & n40554 ;
  assign n40933 = ~n19157 ;
  assign n19191 = n40933 & n19190 ;
  assign n19364 = n19191 & n19362 ;
  assign n19162 = n19156 | n19157 ;
  assign n40934 = ~n19162 ;
  assign n19601 = n40934 & n143 ;
  assign n19602 = n18635 | n19601 ;
  assign n40935 = ~n19364 ;
  assign n19603 = n40935 & n19602 ;
  assign n19886 = n40914 & n19881 ;
  assign n19887 = n19485 | n19886 ;
  assign n40936 = ~n19883 ;
  assign n19888 = n40936 & n19887 ;
  assign n40937 = ~n19888 ;
  assign n19889 = n176 & n40937 ;
  assign n19890 = n40921 & n19887 ;
  assign n19935 = n19890 | n19934 ;
  assign n40938 = ~n19889 ;
  assign n19936 = n40938 & n19935 ;
  assign n40939 = ~n19936 ;
  assign n19937 = n177 & n40939 ;
  assign n19938 = n178 | n19937 ;
  assign n40940 = ~n19938 ;
  assign n19959 = n40940 & n19954 ;
  assign n19960 = n19603 | n19959 ;
  assign n40941 = ~n19956 ;
  assign n19961 = n40941 & n19960 ;
  assign n40942 = ~n19961 ;
  assign n19962 = n179 & n40942 ;
  assign n40943 = ~n19177 ;
  assign n19187 = n18721 & n40943 ;
  assign n19188 = n40543 & n19187 ;
  assign n19363 = n19188 & n19362 ;
  assign n19189 = n19160 | n19177 ;
  assign n40944 = ~n19189 ;
  assign n19500 = n40944 & n143 ;
  assign n19501 = n18721 | n19500 ;
  assign n40945 = ~n19363 ;
  assign n19502 = n40945 & n19501 ;
  assign n19957 = n1707 | n19956 ;
  assign n40946 = ~n19957 ;
  assign n19963 = n40946 & n19960 ;
  assign n19964 = n19502 | n19963 ;
  assign n40947 = ~n19962 ;
  assign n19965 = n40947 & n19964 ;
  assign n40948 = ~n19965 ;
  assign n19966 = n1487 & n40948 ;
  assign n19939 = n40927 & n19935 ;
  assign n19970 = n19939 | n19953 ;
  assign n40949 = ~n19937 ;
  assign n19971 = n40949 & n19970 ;
  assign n40950 = ~n19971 ;
  assign n19972 = n178 & n40950 ;
  assign n19973 = n40940 & n19970 ;
  assign n19974 = n19603 | n19973 ;
  assign n40951 = ~n19972 ;
  assign n19975 = n40951 & n19974 ;
  assign n40952 = ~n19975 ;
  assign n19976 = n1707 & n40952 ;
  assign n19977 = n1487 | n19976 ;
  assign n40953 = ~n19977 ;
  assign n19978 = n19964 & n40953 ;
  assign n19214 = n18633 & n40570 ;
  assign n40954 = ~n19181 ;
  assign n19215 = n40954 & n19214 ;
  assign n19990 = n19215 & n143 ;
  assign n19186 = n19180 | n19181 ;
  assign n40955 = ~n19186 ;
  assign n19991 = n40955 & n143 ;
  assign n19992 = n18633 | n19991 ;
  assign n40956 = ~n19990 ;
  assign n19993 = n40956 & n19992 ;
  assign n20002 = n19978 | n19993 ;
  assign n40957 = ~n19966 ;
  assign n20003 = n40957 & n20002 ;
  assign n40958 = ~n20003 ;
  assign n20004 = n181 & n40958 ;
  assign n19967 = n181 | n19966 ;
  assign n40959 = ~n19967 ;
  assign n20005 = n40959 & n20002 ;
  assign n19211 = n19184 | n19201 ;
  assign n40960 = ~n19211 ;
  assign n19512 = n40960 & n143 ;
  assign n19513 = n18754 | n19512 ;
  assign n40961 = ~n19201 ;
  assign n19212 = n18754 & n40961 ;
  assign n19213 = n40559 & n19212 ;
  assign n20006 = n19213 & n143 ;
  assign n40962 = ~n20006 ;
  assign n20007 = n19513 & n40962 ;
  assign n20008 = n20005 | n20007 ;
  assign n40963 = ~n20004 ;
  assign n20009 = n40963 & n20008 ;
  assign n40964 = ~n20009 ;
  assign n20010 = n182 & n40964 ;
  assign n19238 = n18764 & n40583 ;
  assign n40965 = ~n19205 ;
  assign n19239 = n40965 & n19238 ;
  assign n19438 = n19239 & n143 ;
  assign n19210 = n19204 | n19205 ;
  assign n40966 = ~n19210 ;
  assign n19947 = n40966 & n143 ;
  assign n19948 = n18764 | n19947 ;
  assign n40967 = ~n19438 ;
  assign n19949 = n40967 & n19948 ;
  assign n19979 = n40946 & n19974 ;
  assign n19980 = n19502 | n19979 ;
  assign n40968 = ~n19976 ;
  assign n19981 = n40968 & n19980 ;
  assign n40969 = ~n19981 ;
  assign n19982 = n180 & n40969 ;
  assign n19983 = n40953 & n19980 ;
  assign n19994 = n19983 | n19993 ;
  assign n40970 = ~n19982 ;
  assign n19995 = n40970 & n19994 ;
  assign n40971 = ~n19995 ;
  assign n19996 = n181 & n40971 ;
  assign n19997 = n182 | n19996 ;
  assign n40972 = ~n19997 ;
  assign n20013 = n40972 & n20008 ;
  assign n20014 = n19949 | n20013 ;
  assign n40973 = ~n20010 ;
  assign n20015 = n40973 & n20014 ;
  assign n40974 = ~n20015 ;
  assign n20016 = n183 & n40974 ;
  assign n20011 = n183 | n20010 ;
  assign n40975 = ~n20011 ;
  assign n20017 = n40975 & n20014 ;
  assign n40976 = ~n19225 ;
  assign n19235 = n18628 & n40976 ;
  assign n19236 = n40575 & n19235 ;
  assign n20034 = n19236 & n143 ;
  assign n19237 = n19208 | n19225 ;
  assign n40977 = ~n19237 ;
  assign n20035 = n40977 & n143 ;
  assign n20036 = n18628 | n20035 ;
  assign n40978 = ~n20034 ;
  assign n20037 = n40978 & n20036 ;
  assign n20038 = n20017 | n20037 ;
  assign n40979 = ~n20016 ;
  assign n20039 = n40979 & n20038 ;
  assign n40980 = ~n20039 ;
  assign n20040 = n838 & n40980 ;
  assign n19998 = n40959 & n19994 ;
  assign n20020 = n19998 | n20007 ;
  assign n40981 = ~n19996 ;
  assign n20021 = n40981 & n20020 ;
  assign n40982 = ~n20021 ;
  assign n20022 = n182 & n40982 ;
  assign n20023 = n40972 & n20020 ;
  assign n20024 = n19949 | n20023 ;
  assign n40983 = ~n20022 ;
  assign n20025 = n40983 & n20024 ;
  assign n40984 = ~n20025 ;
  assign n20026 = n996 & n40984 ;
  assign n20027 = n838 | n20026 ;
  assign n40985 = ~n20027 ;
  assign n20042 = n40985 & n20038 ;
  assign n19234 = n19228 | n19229 ;
  assign n40986 = ~n19234 ;
  assign n19489 = n40986 & n143 ;
  assign n19490 = n18689 | n19489 ;
  assign n19251 = n18689 & n40602 ;
  assign n40987 = ~n19229 ;
  assign n19252 = n40987 & n19251 ;
  assign n20050 = n19252 & n143 ;
  assign n40988 = ~n20050 ;
  assign n20051 = n19490 & n40988 ;
  assign n20060 = n20042 | n20051 ;
  assign n40989 = ~n20040 ;
  assign n20061 = n40989 & n20060 ;
  assign n40990 = ~n20061 ;
  assign n20062 = n185 & n40990 ;
  assign n20041 = n185 | n20040 ;
  assign n40991 = ~n20041 ;
  assign n20063 = n40991 & n20060 ;
  assign n40992 = ~n19249 ;
  assign n19301 = n40992 & n19285 ;
  assign n19302 = n40591 & n19301 ;
  assign n20064 = n19302 & n143 ;
  assign n19250 = n19232 | n19249 ;
  assign n40993 = ~n19250 ;
  assign n20065 = n40993 & n143 ;
  assign n20105 = n19285 | n20065 ;
  assign n40994 = ~n20064 ;
  assign n20106 = n40994 & n20105 ;
  assign n20107 = n20063 | n20106 ;
  assign n40995 = ~n20062 ;
  assign n20108 = n40995 & n20107 ;
  assign n40996 = ~n20108 ;
  assign n20109 = n186 & n40996 ;
  assign n19290 = n18768 & n40618 ;
  assign n40997 = ~n19306 ;
  assign n19307 = n19290 & n40997 ;
  assign n19370 = n19307 & n19362 ;
  assign n19308 = n19305 | n19306 ;
  assign n40998 = ~n19308 ;
  assign n19409 = n40998 & n143 ;
  assign n19410 = n18768 | n19409 ;
  assign n40999 = ~n19370 ;
  assign n19411 = n40999 & n19410 ;
  assign n20028 = n40975 & n20024 ;
  assign n20045 = n20028 | n20037 ;
  assign n41000 = ~n20026 ;
  assign n20046 = n41000 & n20045 ;
  assign n41001 = ~n20046 ;
  assign n20047 = n184 & n41001 ;
  assign n20048 = n40985 & n20045 ;
  assign n20052 = n20048 | n20051 ;
  assign n41002 = ~n20047 ;
  assign n20053 = n41002 & n20052 ;
  assign n41003 = ~n20053 ;
  assign n20054 = n185 & n41003 ;
  assign n20055 = n186 | n20054 ;
  assign n41004 = ~n20055 ;
  assign n20112 = n41004 & n20107 ;
  assign n20113 = n19411 | n20112 ;
  assign n41005 = ~n20109 ;
  assign n20114 = n41005 & n20113 ;
  assign n41006 = ~n20114 ;
  assign n20115 = n187 & n41006 ;
  assign n41007 = ~n19323 ;
  assign n20098 = n18607 & n41007 ;
  assign n20099 = n40607 & n20098 ;
  assign n20100 = n143 & n20099 ;
  assign n20101 = n19311 | n19323 ;
  assign n41008 = ~n20101 ;
  assign n20102 = n143 & n41008 ;
  assign n20103 = n18607 | n20102 ;
  assign n41009 = ~n20100 ;
  assign n20104 = n41009 & n20103 ;
  assign n20110 = n528 | n20109 ;
  assign n41010 = ~n20110 ;
  assign n20116 = n41010 & n20113 ;
  assign n20117 = n20104 | n20116 ;
  assign n41011 = ~n20115 ;
  assign n20118 = n41011 & n20117 ;
  assign n41012 = ~n20118 ;
  assign n20119 = n413 & n41012 ;
  assign n19300 = n18621 & n40634 ;
  assign n41013 = ~n19327 ;
  assign n20092 = n19300 & n41013 ;
  assign n20093 = n143 & n20092 ;
  assign n20094 = n19326 | n19327 ;
  assign n41014 = ~n20094 ;
  assign n20095 = n143 & n41014 ;
  assign n20096 = n18621 | n20095 ;
  assign n41015 = ~n20093 ;
  assign n20097 = n41015 & n20096 ;
  assign n20056 = n40991 & n20052 ;
  assign n20124 = n20056 | n20106 ;
  assign n41016 = ~n20054 ;
  assign n20125 = n41016 & n20124 ;
  assign n41017 = ~n20125 ;
  assign n20126 = n186 & n41017 ;
  assign n20127 = n41004 & n20124 ;
  assign n20128 = n19411 | n20127 ;
  assign n41018 = ~n20126 ;
  assign n20129 = n41018 & n20128 ;
  assign n41019 = ~n20129 ;
  assign n20130 = n528 & n41019 ;
  assign n20131 = n413 | n20130 ;
  assign n41020 = ~n20131 ;
  assign n20132 = n20117 & n41020 ;
  assign n20133 = n20097 | n20132 ;
  assign n41021 = ~n20119 ;
  assign n20134 = n41021 & n20133 ;
  assign n41022 = ~n20134 ;
  assign n20135 = n189 & n41022 ;
  assign n41023 = ~n19342 ;
  assign n20085 = n18752 & n41023 ;
  assign n20086 = n40623 & n20085 ;
  assign n20087 = n143 & n20086 ;
  assign n20088 = n19330 | n19342 ;
  assign n41024 = ~n20088 ;
  assign n20089 = n143 & n41024 ;
  assign n20090 = n18752 | n20089 ;
  assign n41025 = ~n20087 ;
  assign n20091 = n41025 & n20090 ;
  assign n20120 = n189 | n20119 ;
  assign n41026 = ~n20120 ;
  assign n20136 = n41026 & n20133 ;
  assign n20137 = n20091 | n20136 ;
  assign n41027 = ~n20135 ;
  assign n20138 = n41027 & n20137 ;
  assign n41028 = ~n20138 ;
  assign n20139 = n190 & n41028 ;
  assign n20140 = n287 | n20139 ;
  assign n19322 = n18727 & n40650 ;
  assign n41029 = ~n19346 ;
  assign n20079 = n19322 & n41029 ;
  assign n20080 = n143 & n20079 ;
  assign n20081 = n19345 | n19346 ;
  assign n41030 = ~n20081 ;
  assign n20082 = n143 & n41030 ;
  assign n20083 = n18727 | n20082 ;
  assign n41031 = ~n20080 ;
  assign n20084 = n41031 & n20083 ;
  assign n20142 = n41010 & n20128 ;
  assign n20143 = n20104 | n20142 ;
  assign n41032 = ~n20130 ;
  assign n20144 = n41032 & n20143 ;
  assign n41033 = ~n20144 ;
  assign n20145 = n188 & n41033 ;
  assign n20146 = n41020 & n20143 ;
  assign n20147 = n20097 | n20146 ;
  assign n41034 = ~n20145 ;
  assign n20148 = n41034 & n20147 ;
  assign n41035 = ~n20148 ;
  assign n20149 = n189 & n41035 ;
  assign n20150 = n190 | n20149 ;
  assign n20151 = n41026 & n20147 ;
  assign n20152 = n20091 | n20151 ;
  assign n41036 = ~n20150 ;
  assign n20155 = n41036 & n20152 ;
  assign n20156 = n20084 | n20155 ;
  assign n41037 = ~n20140 ;
  assign n20157 = n41037 & n20156 ;
  assign n20159 = n20078 | n20157 ;
  assign n41038 = ~n20149 ;
  assign n20153 = n41038 & n20152 ;
  assign n41039 = ~n20153 ;
  assign n20154 = n190 & n41039 ;
  assign n41040 = ~n20154 ;
  assign n20160 = n41040 & n20156 ;
  assign n41041 = ~n20160 ;
  assign n20161 = n287 & n41041 ;
  assign n41042 = ~n20161 ;
  assign n20162 = n20159 & n41042 ;
  assign n20163 = n20069 | n20162 ;
  assign n20164 = n31336 & n20163 ;
  assign n19268 = n18589 | n19267 ;
  assign n41043 = ~n19268 ;
  assign n19274 = n41043 & n19271 ;
  assign n19275 = n40674 & n19274 ;
  assign n19379 = n19275 & n40675 ;
  assign n19380 = n40676 & n19379 ;
  assign n19386 = n192 & n19385 ;
  assign n41044 = ~n19272 ;
  assign n19473 = n41044 & n143 ;
  assign n41045 = ~n19473 ;
  assign n19474 = n19357 & n41045 ;
  assign n41046 = ~n19474 ;
  assign n19475 = n19386 & n41046 ;
  assign n19476 = n19380 | n19475 ;
  assign n20167 = n20068 & n41042 ;
  assign n20168 = n20159 & n20167 ;
  assign n20169 = n19476 | n20168 ;
  assign n142 = n20164 | n20169 ;
  assign n20165 = n20068 | n20162 ;
  assign n20166 = n192 & n20165 ;
  assign n41047 = ~n20068 ;
  assign n20332 = n41047 & n142 ;
  assign n41048 = ~n20332 ;
  assign n20333 = n20162 & n41048 ;
  assign n41049 = ~n20333 ;
  assign n20334 = n20166 & n41049 ;
  assign n20033 = n19380 | n20032 ;
  assign n41050 = ~n20033 ;
  assign n20070 = n41050 & n20067 ;
  assign n41051 = ~n19475 ;
  assign n20071 = n41051 & n20070 ;
  assign n41052 = ~n20168 ;
  assign n20876 = n20071 & n41052 ;
  assign n41053 = ~n20164 ;
  assign n20877 = n41053 & n20876 ;
  assign n20878 = n20334 | n20877 ;
  assign n41054 = ~n20157 ;
  assign n20158 = n20078 & n41054 ;
  assign n20885 = n20158 & n41042 ;
  assign n20886 = n142 & n20885 ;
  assign n20888 = n20157 | n20161 ;
  assign n41055 = ~n20888 ;
  assign n20889 = n142 & n41055 ;
  assign n20890 = n20078 | n20889 ;
  assign n41056 = ~n20886 ;
  assign n20891 = n41056 & n20890 ;
  assign n233 = x24 | x25 ;
  assign n234 = x26 | n233 ;
  assign n20261 = x26 & n142 ;
  assign n41057 = ~n20261 ;
  assign n20262 = n234 & n41057 ;
  assign n41058 = ~n20262 ;
  assign n20263 = n143 & n41058 ;
  assign n18590 = n234 & n40673 ;
  assign n18734 = n18590 & n40674 ;
  assign n19383 = n18734 & n40675 ;
  assign n19384 = n40676 & n19383 ;
  assign n20335 = n19384 & n41057 ;
  assign n41059 = ~n230 ;
  assign n20221 = n41059 & n142 ;
  assign n41060 = ~x26 ;
  assign n20352 = n41060 & n142 ;
  assign n41061 = ~n20352 ;
  assign n20353 = x27 & n41061 ;
  assign n20354 = n20221 | n20353 ;
  assign n20355 = n20335 | n20354 ;
  assign n41062 = ~n20263 ;
  assign n20358 = n41062 & n20355 ;
  assign n41063 = ~n20358 ;
  assign n20359 = n18797 & n41063 ;
  assign n235 = n41060 & n233 ;
  assign n41064 = ~n142 ;
  assign n20340 = x26 & n41064 ;
  assign n20341 = n235 | n20340 ;
  assign n41065 = ~n20341 ;
  assign n20342 = n19362 & n41065 ;
  assign n20343 = n18797 | n20342 ;
  assign n41066 = ~n20343 ;
  assign n20356 = n41066 & n20355 ;
  assign n41067 = ~n19380 ;
  assign n19381 = n19362 & n41067 ;
  assign n19477 = n19381 & n41051 ;
  assign n20364 = n19477 & n41052 ;
  assign n20365 = n41053 & n20364 ;
  assign n20366 = n20221 | n20365 ;
  assign n20367 = x28 & n20366 ;
  assign n20368 = x28 | n20365 ;
  assign n20369 = n20221 | n20368 ;
  assign n41068 = ~n20367 ;
  assign n20370 = n41068 & n20369 ;
  assign n20371 = n20356 | n20370 ;
  assign n41069 = ~n20359 ;
  assign n20372 = n41069 & n20371 ;
  assign n41070 = ~n20372 ;
  assign n20373 = n145 & n41070 ;
  assign n19437 = n19375 | n19436 ;
  assign n41071 = ~n19437 ;
  assign n19524 = n41071 & n19523 ;
  assign n20338 = n19524 & n142 ;
  assign n20345 = n41071 & n142 ;
  assign n20346 = n19523 | n20345 ;
  assign n41072 = ~n20338 ;
  assign n20347 = n41072 & n20346 ;
  assign n20360 = n145 | n20359 ;
  assign n41073 = ~n20360 ;
  assign n20376 = n41073 & n20371 ;
  assign n20377 = n20347 | n20376 ;
  assign n41074 = ~n20373 ;
  assign n20378 = n41074 & n20377 ;
  assign n41075 = ~n20378 ;
  assign n20379 = n146 & n41075 ;
  assign n41076 = ~n19538 ;
  assign n19543 = n19532 & n41076 ;
  assign n41077 = ~n19540 ;
  assign n19544 = n41077 & n19543 ;
  assign n20339 = n19544 & n142 ;
  assign n19542 = n19538 | n19540 ;
  assign n41078 = ~n19542 ;
  assign n20348 = n41078 & n142 ;
  assign n20349 = n19532 | n20348 ;
  assign n41079 = ~n20339 ;
  assign n20350 = n41079 & n20349 ;
  assign n20374 = n146 | n20373 ;
  assign n41080 = ~n20374 ;
  assign n20380 = n41080 & n20377 ;
  assign n20381 = n20350 | n20380 ;
  assign n41081 = ~n20379 ;
  assign n20382 = n41081 & n20381 ;
  assign n41082 = ~n20382 ;
  assign n20383 = n16322 & n41082 ;
  assign n19595 = n19535 | n19546 ;
  assign n41083 = ~n19595 ;
  assign n20330 = n41083 & n142 ;
  assign n20331 = n19482 | n20330 ;
  assign n19536 = n19482 & n40684 ;
  assign n41084 = ~n19546 ;
  assign n19594 = n19536 & n41084 ;
  assign n20336 = n19594 & n142 ;
  assign n41085 = ~n20336 ;
  assign n20337 = n20331 & n41085 ;
  assign n20361 = n144 & n41063 ;
  assign n20264 = n144 | n20263 ;
  assign n41086 = ~n20264 ;
  assign n20363 = n41086 & n20355 ;
  assign n20392 = n20363 | n20370 ;
  assign n41087 = ~n20361 ;
  assign n20393 = n41087 & n20392 ;
  assign n41088 = ~n20393 ;
  assign n20394 = n145 & n41088 ;
  assign n20395 = n41073 & n20392 ;
  assign n20396 = n20347 | n20395 ;
  assign n41089 = ~n20394 ;
  assign n20397 = n41089 & n20396 ;
  assign n41090 = ~n20397 ;
  assign n20398 = n146 & n41090 ;
  assign n20399 = n147 | n20398 ;
  assign n41091 = ~n20399 ;
  assign n20400 = n20381 & n41091 ;
  assign n20401 = n20337 | n20400 ;
  assign n41092 = ~n20383 ;
  assign n20402 = n41092 & n20401 ;
  assign n41093 = ~n20402 ;
  assign n20403 = n148 & n41093 ;
  assign n19563 = n19549 | n19551 ;
  assign n41094 = ~n19563 ;
  assign n20241 = n41094 & n142 ;
  assign n20242 = n19492 | n20241 ;
  assign n41095 = ~n19551 ;
  assign n19561 = n19492 & n41095 ;
  assign n19562 = n40709 & n19561 ;
  assign n20290 = n19562 & n142 ;
  assign n41096 = ~n20290 ;
  assign n20291 = n20242 & n41096 ;
  assign n20384 = n148 | n20383 ;
  assign n41097 = ~n20384 ;
  assign n20404 = n41097 & n20401 ;
  assign n20405 = n20291 | n20404 ;
  assign n41098 = ~n20403 ;
  assign n20406 = n41098 & n20405 ;
  assign n41099 = ~n20406 ;
  assign n20407 = n149 & n41099 ;
  assign n19582 = n19480 & n40701 ;
  assign n41100 = ~n19555 ;
  assign n19583 = n41100 & n19582 ;
  assign n20199 = n19583 & n142 ;
  assign n19560 = n19554 | n19555 ;
  assign n41101 = ~n19560 ;
  assign n20258 = n41101 & n142 ;
  assign n20259 = n19480 | n20258 ;
  assign n41102 = ~n20199 ;
  assign n20260 = n41102 & n20259 ;
  assign n20415 = n41080 & n20396 ;
  assign n20416 = n20350 | n20415 ;
  assign n41103 = ~n20398 ;
  assign n20417 = n41103 & n20416 ;
  assign n41104 = ~n20417 ;
  assign n20418 = n147 & n41104 ;
  assign n20419 = n41091 & n20416 ;
  assign n20420 = n20337 | n20419 ;
  assign n41105 = ~n20418 ;
  assign n20421 = n41105 & n20420 ;
  assign n41106 = ~n20421 ;
  assign n20422 = n15807 & n41106 ;
  assign n20423 = n149 | n20422 ;
  assign n41107 = ~n20423 ;
  assign n20424 = n20405 & n41107 ;
  assign n20425 = n20260 | n20424 ;
  assign n41108 = ~n20407 ;
  assign n20426 = n41108 & n20425 ;
  assign n41109 = ~n20426 ;
  assign n20427 = n150 & n41109 ;
  assign n41110 = ~n19573 ;
  assign n19579 = n19453 & n41110 ;
  assign n19580 = n40728 & n19579 ;
  assign n20220 = n19580 & n142 ;
  assign n19581 = n19558 | n19573 ;
  assign n41111 = ~n19581 ;
  assign n20248 = n41111 & n142 ;
  assign n20249 = n19453 | n20248 ;
  assign n41112 = ~n20220 ;
  assign n20250 = n41112 & n20249 ;
  assign n20408 = n150 | n20407 ;
  assign n41113 = ~n20408 ;
  assign n20428 = n41113 & n20425 ;
  assign n20429 = n20250 | n20428 ;
  assign n41114 = ~n20427 ;
  assign n20430 = n41114 & n20429 ;
  assign n41115 = ~n20430 ;
  assign n20431 = n13662 & n41115 ;
  assign n19722 = n40717 & n19615 ;
  assign n41116 = ~n19577 ;
  assign n19723 = n41116 & n19722 ;
  assign n20219 = n19723 & n142 ;
  assign n19578 = n19576 | n19577 ;
  assign n41117 = ~n19578 ;
  assign n20226 = n41117 & n142 ;
  assign n20227 = n19615 | n20226 ;
  assign n41118 = ~n20219 ;
  assign n20228 = n41118 & n20227 ;
  assign n20439 = n41097 & n20420 ;
  assign n20440 = n20291 | n20439 ;
  assign n41119 = ~n20422 ;
  assign n20441 = n41119 & n20440 ;
  assign n41120 = ~n20441 ;
  assign n20442 = n149 & n41120 ;
  assign n20443 = n41107 & n20440 ;
  assign n20444 = n20260 | n20443 ;
  assign n41121 = ~n20442 ;
  assign n20445 = n41121 & n20444 ;
  assign n41122 = ~n20445 ;
  assign n20446 = n150 & n41122 ;
  assign n20447 = n151 | n20446 ;
  assign n41123 = ~n20447 ;
  assign n20448 = n20429 & n41123 ;
  assign n20449 = n20228 | n20448 ;
  assign n41124 = ~n20431 ;
  assign n20450 = n41124 & n20449 ;
  assign n41125 = ~n20450 ;
  assign n20451 = n152 & n41125 ;
  assign n19721 = n19627 | n19639 ;
  assign n41126 = ~n19721 ;
  assign n20231 = n41126 & n142 ;
  assign n20232 = n19470 | n20231 ;
  assign n41127 = ~n19639 ;
  assign n19719 = n19470 & n41127 ;
  assign n19720 = n40744 & n19719 ;
  assign n20251 = n19720 & n142 ;
  assign n41128 = ~n20251 ;
  assign n20252 = n20232 & n41128 ;
  assign n20432 = n152 | n20431 ;
  assign n41129 = ~n20432 ;
  assign n20452 = n41129 & n20449 ;
  assign n20453 = n20252 | n20452 ;
  assign n41130 = ~n20451 ;
  assign n20454 = n41130 & n20453 ;
  assign n41131 = ~n20454 ;
  assign n20455 = n153 & n41131 ;
  assign n19717 = n19642 | n19643 ;
  assign n41132 = ~n19717 ;
  assign n20268 = n41132 & n142 ;
  assign n20269 = n19610 | n20268 ;
  assign n19624 = n19610 & n40733 ;
  assign n41133 = ~n19643 ;
  assign n19718 = n19624 & n41133 ;
  assign n20275 = n19718 & n142 ;
  assign n41134 = ~n20275 ;
  assign n20276 = n20269 & n41134 ;
  assign n20463 = n41113 & n20444 ;
  assign n20464 = n20250 | n20463 ;
  assign n41135 = ~n20446 ;
  assign n20465 = n41135 & n20464 ;
  assign n41136 = ~n20465 ;
  assign n20466 = n151 & n41136 ;
  assign n20467 = n41123 & n20464 ;
  assign n20468 = n20228 | n20467 ;
  assign n41137 = ~n20466 ;
  assign n20469 = n41137 & n20468 ;
  assign n41138 = ~n20469 ;
  assign n20470 = n13079 & n41138 ;
  assign n20471 = n153 | n20470 ;
  assign n41139 = ~n20471 ;
  assign n20472 = n20453 & n41139 ;
  assign n20473 = n20276 | n20472 ;
  assign n41140 = ~n20455 ;
  assign n20474 = n41140 & n20473 ;
  assign n41141 = ~n20474 ;
  assign n20475 = n154 & n41141 ;
  assign n41142 = ~n19658 ;
  assign n19714 = n19518 & n41142 ;
  assign n19715 = n40760 & n19714 ;
  assign n20222 = n19715 & n142 ;
  assign n19716 = n19646 | n19658 ;
  assign n41143 = ~n19716 ;
  assign n20255 = n41143 & n142 ;
  assign n20256 = n19518 | n20255 ;
  assign n41144 = ~n20222 ;
  assign n20257 = n41144 & n20256 ;
  assign n20456 = n154 | n20455 ;
  assign n41145 = ~n20456 ;
  assign n20476 = n41145 & n20473 ;
  assign n20477 = n20257 | n20476 ;
  assign n41146 = ~n20475 ;
  assign n20478 = n41146 & n20477 ;
  assign n41147 = ~n20478 ;
  assign n20479 = n11067 & n41147 ;
  assign n19638 = n19520 & n40749 ;
  assign n41148 = ~n19662 ;
  assign n19712 = n19638 & n41148 ;
  assign n20243 = n19712 & n142 ;
  assign n19713 = n19661 | n19662 ;
  assign n41149 = ~n19713 ;
  assign n20277 = n41149 & n142 ;
  assign n20278 = n19520 | n20277 ;
  assign n41150 = ~n20243 ;
  assign n20279 = n41150 & n20278 ;
  assign n20487 = n41129 & n20468 ;
  assign n20488 = n20252 | n20487 ;
  assign n41151 = ~n20470 ;
  assign n20489 = n41151 & n20488 ;
  assign n41152 = ~n20489 ;
  assign n20490 = n153 & n41152 ;
  assign n20491 = n41139 & n20488 ;
  assign n20492 = n20276 | n20491 ;
  assign n41153 = ~n20490 ;
  assign n20493 = n41153 & n20492 ;
  assign n41154 = ~n20493 ;
  assign n20494 = n154 & n41154 ;
  assign n20495 = n11067 | n20494 ;
  assign n41155 = ~n20495 ;
  assign n20496 = n20477 & n41155 ;
  assign n20497 = n20279 | n20496 ;
  assign n41156 = ~n20479 ;
  assign n20498 = n41156 & n20497 ;
  assign n41157 = ~n20498 ;
  assign n20499 = n156 & n41157 ;
  assign n41158 = ~n19677 ;
  assign n19709 = n19608 & n41158 ;
  assign n19710 = n40776 & n19709 ;
  assign n20233 = n19710 & n142 ;
  assign n19711 = n19665 | n19677 ;
  assign n41159 = ~n19711 ;
  assign n20244 = n41159 & n142 ;
  assign n20245 = n19608 | n20244 ;
  assign n41160 = ~n20233 ;
  assign n20246 = n41160 & n20245 ;
  assign n20480 = n10657 | n20479 ;
  assign n41161 = ~n20480 ;
  assign n20500 = n41161 & n20497 ;
  assign n20501 = n20246 | n20500 ;
  assign n41162 = ~n20499 ;
  assign n20502 = n41162 & n20501 ;
  assign n41163 = ~n20502 ;
  assign n20503 = n157 & n41163 ;
  assign n19708 = n19680 | n19681 ;
  assign n41164 = ~n19708 ;
  assign n20282 = n41164 & n142 ;
  assign n20283 = n19612 | n20282 ;
  assign n19657 = n19612 & n40765 ;
  assign n41165 = ~n19681 ;
  assign n19707 = n19657 & n41165 ;
  assign n20288 = n19707 & n142 ;
  assign n41166 = ~n20288 ;
  assign n20289 = n20283 & n41166 ;
  assign n20511 = n41145 & n20492 ;
  assign n20512 = n20257 | n20511 ;
  assign n41167 = ~n20494 ;
  assign n20513 = n41167 & n20512 ;
  assign n41168 = ~n20513 ;
  assign n20514 = n155 & n41168 ;
  assign n20515 = n41155 & n20512 ;
  assign n20516 = n20279 | n20515 ;
  assign n41169 = ~n20514 ;
  assign n20517 = n41169 & n20516 ;
  assign n41170 = ~n20517 ;
  assign n20518 = n10657 & n41170 ;
  assign n20519 = n157 | n20518 ;
  assign n41171 = ~n20519 ;
  assign n20520 = n20501 & n41171 ;
  assign n20521 = n20289 | n20520 ;
  assign n41172 = ~n20503 ;
  assign n20522 = n41172 & n20521 ;
  assign n41173 = ~n20522 ;
  assign n20523 = n158 & n41173 ;
  assign n19704 = n19684 | n19691 ;
  assign n41174 = ~n19704 ;
  assign n20253 = n41174 & n142 ;
  assign n20254 = n19515 | n20253 ;
  assign n41175 = ~n19691 ;
  assign n19705 = n19515 & n41175 ;
  assign n19706 = n40792 & n19705 ;
  assign n20280 = n19706 & n142 ;
  assign n41176 = ~n20280 ;
  assign n20281 = n20254 & n41176 ;
  assign n20504 = n158 | n20503 ;
  assign n41177 = ~n20504 ;
  assign n20524 = n41177 & n20521 ;
  assign n20525 = n20281 | n20524 ;
  assign n41178 = ~n20523 ;
  assign n20526 = n41178 & n20525 ;
  assign n41179 = ~n20526 ;
  assign n20527 = n8857 & n41179 ;
  assign n19676 = n19418 & n40781 ;
  assign n41180 = ~n19695 ;
  assign n19702 = n19676 & n41180 ;
  assign n20204 = n19702 & n142 ;
  assign n19703 = n19694 | n19695 ;
  assign n41181 = ~n19703 ;
  assign n20223 = n41181 & n142 ;
  assign n20224 = n19418 | n20223 ;
  assign n41182 = ~n20204 ;
  assign n20225 = n41182 & n20224 ;
  assign n20535 = n41161 & n20516 ;
  assign n20536 = n20246 | n20535 ;
  assign n41183 = ~n20518 ;
  assign n20537 = n41183 & n20536 ;
  assign n41184 = ~n20537 ;
  assign n20538 = n157 & n41184 ;
  assign n20539 = n41171 & n20536 ;
  assign n20540 = n20289 | n20539 ;
  assign n41185 = ~n20538 ;
  assign n20541 = n41185 & n20540 ;
  assign n41186 = ~n20541 ;
  assign n20542 = n158 & n41186 ;
  assign n20543 = n8857 | n20542 ;
  assign n41187 = ~n20543 ;
  assign n20544 = n20525 & n41187 ;
  assign n20545 = n20225 | n20544 ;
  assign n41188 = ~n20527 ;
  assign n20546 = n41188 & n20545 ;
  assign n41189 = ~n20546 ;
  assign n20547 = n160 & n41189 ;
  assign n41190 = ~n19700 ;
  assign n19930 = n41190 & n19727 ;
  assign n19931 = n40808 & n19930 ;
  assign n20247 = n19931 & n142 ;
  assign n19701 = n19698 | n19700 ;
  assign n41191 = ~n19701 ;
  assign n20272 = n41191 & n142 ;
  assign n20273 = n19727 | n20272 ;
  assign n41192 = ~n20247 ;
  assign n20274 = n41192 & n20273 ;
  assign n20528 = n160 | n20527 ;
  assign n41193 = ~n20528 ;
  assign n20548 = n41193 & n20545 ;
  assign n20549 = n20274 | n20548 ;
  assign n41194 = ~n20547 ;
  assign n20550 = n41194 & n20549 ;
  assign n41195 = ~n20550 ;
  assign n20551 = n161 & n41195 ;
  assign n19929 = n19745 | n19746 ;
  assign n41196 = ~n19929 ;
  assign n20239 = n41196 & n142 ;
  assign n20240 = n19461 | n20239 ;
  assign n19732 = n19461 & n40797 ;
  assign n41197 = ~n19746 ;
  assign n19928 = n19732 & n41197 ;
  assign n20284 = n19928 & n142 ;
  assign n41198 = ~n20284 ;
  assign n20285 = n20240 & n41198 ;
  assign n20559 = n41177 & n20540 ;
  assign n20560 = n20281 | n20559 ;
  assign n41199 = ~n20542 ;
  assign n20561 = n41199 & n20560 ;
  assign n41200 = ~n20561 ;
  assign n20562 = n159 & n41200 ;
  assign n20563 = n41187 & n20560 ;
  assign n20564 = n20225 | n20563 ;
  assign n41201 = ~n20562 ;
  assign n20565 = n41201 & n20564 ;
  assign n41202 = ~n20565 ;
  assign n20566 = n8534 & n41202 ;
  assign n20567 = n161 | n20566 ;
  assign n41203 = ~n20567 ;
  assign n20568 = n20549 & n41203 ;
  assign n20569 = n20285 | n20568 ;
  assign n41204 = ~n20551 ;
  assign n20570 = n41204 & n20569 ;
  assign n41205 = ~n20570 ;
  assign n20571 = n162 & n41205 ;
  assign n19927 = n19749 | n19761 ;
  assign n41206 = ~n19927 ;
  assign n20193 = n41206 & n142 ;
  assign n20194 = n19446 | n20193 ;
  assign n41207 = ~n19761 ;
  assign n19925 = n19446 & n41207 ;
  assign n19926 = n40824 & n19925 ;
  assign n20217 = n19926 & n142 ;
  assign n41208 = ~n20217 ;
  assign n20218 = n20194 & n41208 ;
  assign n20552 = n162 | n20551 ;
  assign n41209 = ~n20552 ;
  assign n20572 = n41209 & n20569 ;
  assign n20573 = n20218 | n20572 ;
  assign n41210 = ~n20571 ;
  assign n20574 = n41210 & n20573 ;
  assign n41211 = ~n20574 ;
  assign n20575 = n6889 & n41211 ;
  assign n19742 = n19442 & n40813 ;
  assign n41212 = ~n19765 ;
  assign n19923 = n19742 & n41212 ;
  assign n20209 = n19923 & n142 ;
  assign n19924 = n19764 | n19765 ;
  assign n41213 = ~n19924 ;
  assign n20212 = n41213 & n142 ;
  assign n20213 = n19442 | n20212 ;
  assign n41214 = ~n20209 ;
  assign n20214 = n41214 & n20213 ;
  assign n20583 = n41193 & n20564 ;
  assign n20584 = n20274 | n20583 ;
  assign n41215 = ~n20566 ;
  assign n20585 = n41215 & n20584 ;
  assign n41216 = ~n20585 ;
  assign n20586 = n161 & n41216 ;
  assign n20587 = n41203 & n20584 ;
  assign n20588 = n20285 | n20587 ;
  assign n41217 = ~n20586 ;
  assign n20589 = n41217 & n20588 ;
  assign n41218 = ~n20589 ;
  assign n20590 = n162 & n41218 ;
  assign n20591 = n6889 | n20590 ;
  assign n41219 = ~n20591 ;
  assign n20592 = n20573 & n41219 ;
  assign n20593 = n20214 | n20592 ;
  assign n41220 = ~n20575 ;
  assign n20594 = n41220 & n20593 ;
  assign n41221 = ~n20594 ;
  assign n20595 = n164 & n41221 ;
  assign n19922 = n19768 | n19780 ;
  assign n41222 = ~n19922 ;
  assign n20207 = n41222 & n142 ;
  assign n20208 = n19468 | n20207 ;
  assign n41223 = ~n19780 ;
  assign n19920 = n19468 & n41223 ;
  assign n19921 = n40840 & n19920 ;
  assign n20237 = n19921 & n142 ;
  assign n41224 = ~n20237 ;
  assign n20238 = n20208 & n41224 ;
  assign n20576 = n6600 | n20575 ;
  assign n41225 = ~n20576 ;
  assign n20596 = n41225 & n20593 ;
  assign n20597 = n20238 | n20596 ;
  assign n41226 = ~n20595 ;
  assign n20598 = n41226 & n20597 ;
  assign n41227 = ~n20598 ;
  assign n20599 = n165 & n41227 ;
  assign n19786 = n19783 | n19784 ;
  assign n41228 = ~n19786 ;
  assign n20205 = n41228 & n142 ;
  assign n20206 = n19600 | n20205 ;
  assign n19760 = n19600 & n40829 ;
  assign n41229 = ~n19784 ;
  assign n19785 = n19760 & n41229 ;
  assign n20270 = n19785 & n142 ;
  assign n41230 = ~n20270 ;
  assign n20271 = n20206 & n41230 ;
  assign n20607 = n41209 & n20588 ;
  assign n20608 = n20218 | n20607 ;
  assign n41231 = ~n20590 ;
  assign n20609 = n41231 & n20608 ;
  assign n41232 = ~n20609 ;
  assign n20610 = n163 & n41232 ;
  assign n20611 = n41219 & n20608 ;
  assign n20612 = n20214 | n20611 ;
  assign n41233 = ~n20610 ;
  assign n20613 = n41233 & n20612 ;
  assign n41234 = ~n20613 ;
  assign n20614 = n6600 & n41234 ;
  assign n20615 = n165 | n20614 ;
  assign n41235 = ~n20615 ;
  assign n20616 = n20597 & n41235 ;
  assign n20617 = n20271 | n20616 ;
  assign n41236 = ~n20599 ;
  assign n20618 = n41236 & n20617 ;
  assign n41237 = ~n20618 ;
  assign n20619 = n166 & n41237 ;
  assign n41238 = ~n19801 ;
  assign n19917 = n19464 & n41238 ;
  assign n19918 = n40856 & n19917 ;
  assign n20200 = n19918 & n142 ;
  assign n19919 = n19789 | n19801 ;
  assign n41239 = ~n19919 ;
  assign n20201 = n41239 & n142 ;
  assign n20202 = n19464 | n20201 ;
  assign n41240 = ~n20200 ;
  assign n20203 = n41240 & n20202 ;
  assign n20600 = n166 | n20599 ;
  assign n41241 = ~n20600 ;
  assign n20620 = n41241 & n20617 ;
  assign n20621 = n20203 | n20620 ;
  assign n41242 = ~n20619 ;
  assign n20622 = n41242 & n20621 ;
  assign n41243 = ~n20622 ;
  assign n20623 = n5352 & n41243 ;
  assign n19916 = n19804 | n19805 ;
  assign n41244 = ~n19916 ;
  assign n20197 = n41244 & n142 ;
  assign n20198 = n19425 | n20197 ;
  assign n19779 = n19425 & n40845 ;
  assign n41245 = ~n19805 ;
  assign n19915 = n19779 & n41245 ;
  assign n20229 = n19915 & n142 ;
  assign n41246 = ~n20229 ;
  assign n20230 = n20198 & n41246 ;
  assign n20631 = n41225 & n20612 ;
  assign n20632 = n20238 | n20631 ;
  assign n41247 = ~n20614 ;
  assign n20633 = n41247 & n20632 ;
  assign n41248 = ~n20633 ;
  assign n20634 = n165 & n41248 ;
  assign n20635 = n41235 & n20632 ;
  assign n20636 = n20271 | n20635 ;
  assign n41249 = ~n20634 ;
  assign n20637 = n41249 & n20636 ;
  assign n41250 = ~n20637 ;
  assign n20638 = n166 & n41250 ;
  assign n20639 = n5352 | n20638 ;
  assign n41251 = ~n20639 ;
  assign n20640 = n20621 & n41251 ;
  assign n20641 = n20230 | n20640 ;
  assign n41252 = ~n20623 ;
  assign n20642 = n41252 & n20641 ;
  assign n41253 = ~n20642 ;
  assign n20643 = n168 & n41253 ;
  assign n41254 = ~n19820 ;
  assign n19913 = n19497 & n41254 ;
  assign n19914 = n40872 & n19913 ;
  assign n20187 = n19914 & n142 ;
  assign n19912 = n19808 | n19820 ;
  assign n41255 = ~n19912 ;
  assign n20188 = n41255 & n142 ;
  assign n20189 = n19497 | n20188 ;
  assign n41256 = ~n20187 ;
  assign n20190 = n41256 & n20189 ;
  assign n20624 = n4934 | n20623 ;
  assign n41257 = ~n20624 ;
  assign n20644 = n41257 & n20641 ;
  assign n20645 = n20190 | n20644 ;
  assign n41258 = ~n20643 ;
  assign n20646 = n41258 & n20645 ;
  assign n41259 = ~n20646 ;
  assign n20647 = n169 & n41259 ;
  assign n19911 = n19823 | n19824 ;
  assign n41260 = ~n19911 ;
  assign n20175 = n41260 & n142 ;
  assign n20176 = n19430 | n20175 ;
  assign n19800 = n19430 & n40861 ;
  assign n41261 = ~n19824 ;
  assign n19910 = n19800 & n41261 ;
  assign n20185 = n19910 & n142 ;
  assign n41262 = ~n20185 ;
  assign n20186 = n20176 & n41262 ;
  assign n20655 = n41241 & n20636 ;
  assign n20656 = n20203 | n20655 ;
  assign n41263 = ~n20638 ;
  assign n20657 = n41263 & n20656 ;
  assign n41264 = ~n20657 ;
  assign n20658 = n167 & n41264 ;
  assign n20659 = n41251 & n20656 ;
  assign n20660 = n20230 | n20659 ;
  assign n41265 = ~n20658 ;
  assign n20661 = n41265 & n20660 ;
  assign n41266 = ~n20661 ;
  assign n20662 = n4934 & n41266 ;
  assign n20663 = n169 | n20662 ;
  assign n41267 = ~n20663 ;
  assign n20664 = n20645 & n41267 ;
  assign n20665 = n20186 | n20664 ;
  assign n41268 = ~n20647 ;
  assign n20666 = n41268 & n20665 ;
  assign n41269 = ~n20666 ;
  assign n20667 = n170 & n41269 ;
  assign n19909 = n19827 | n19839 ;
  assign n41270 = ~n19909 ;
  assign n20183 = n41270 & n142 ;
  assign n20184 = n19507 | n20183 ;
  assign n41271 = ~n19839 ;
  assign n19907 = n19507 & n41271 ;
  assign n19908 = n40888 & n19907 ;
  assign n20292 = n19908 & n142 ;
  assign n41272 = ~n20292 ;
  assign n20293 = n20184 & n41272 ;
  assign n20648 = n170 | n20647 ;
  assign n41273 = ~n20648 ;
  assign n20668 = n41273 & n20665 ;
  assign n20669 = n20293 | n20668 ;
  assign n41274 = ~n20667 ;
  assign n20670 = n41274 & n20669 ;
  assign n41275 = ~n20670 ;
  assign n20671 = n3940 & n41275 ;
  assign n19819 = n19472 & n40877 ;
  assign n41276 = ~n19843 ;
  assign n19905 = n19819 & n41276 ;
  assign n20179 = n19905 & n142 ;
  assign n19906 = n19842 | n19843 ;
  assign n41277 = ~n19906 ;
  assign n20180 = n41277 & n142 ;
  assign n20181 = n19472 | n20180 ;
  assign n41278 = ~n20179 ;
  assign n20182 = n41278 & n20181 ;
  assign n20679 = n41257 & n20660 ;
  assign n20680 = n20190 | n20679 ;
  assign n41279 = ~n20662 ;
  assign n20681 = n41279 & n20680 ;
  assign n41280 = ~n20681 ;
  assign n20682 = n169 & n41280 ;
  assign n20683 = n41267 & n20680 ;
  assign n20684 = n20186 | n20683 ;
  assign n41281 = ~n20682 ;
  assign n20685 = n41281 & n20684 ;
  assign n41282 = ~n20685 ;
  assign n20686 = n170 & n41282 ;
  assign n20687 = n3940 | n20686 ;
  assign n41283 = ~n20687 ;
  assign n20688 = n20669 & n41283 ;
  assign n20689 = n20182 | n20688 ;
  assign n41284 = ~n20671 ;
  assign n20690 = n41284 & n20689 ;
  assign n41285 = ~n20690 ;
  assign n20691 = n172 & n41285 ;
  assign n41286 = ~n19858 ;
  assign n19902 = n19457 & n41286 ;
  assign n19903 = n40904 & n19902 ;
  assign n20192 = n19903 & n142 ;
  assign n19904 = n19846 | n19858 ;
  assign n41287 = ~n19904 ;
  assign n20265 = n41287 & n142 ;
  assign n20266 = n19457 | n20265 ;
  assign n41288 = ~n20192 ;
  assign n20267 = n41288 & n20266 ;
  assign n20672 = n3631 | n20671 ;
  assign n41289 = ~n20672 ;
  assign n20692 = n41289 & n20689 ;
  assign n20693 = n20267 | n20692 ;
  assign n41290 = ~n20691 ;
  assign n20694 = n41290 & n20693 ;
  assign n41291 = ~n20694 ;
  assign n20695 = n173 & n41291 ;
  assign n19901 = n19861 | n19862 ;
  assign n41292 = ~n19901 ;
  assign n20177 = n41292 & n142 ;
  assign n20178 = n19598 | n20177 ;
  assign n19838 = n19598 & n40893 ;
  assign n41293 = ~n19862 ;
  assign n19900 = n19838 & n41293 ;
  assign n20215 = n19900 & n142 ;
  assign n41294 = ~n20215 ;
  assign n20216 = n20178 & n41294 ;
  assign n20703 = n41273 & n20684 ;
  assign n20704 = n20293 | n20703 ;
  assign n41295 = ~n20686 ;
  assign n20705 = n41295 & n20704 ;
  assign n41296 = ~n20705 ;
  assign n20706 = n171 & n41296 ;
  assign n20707 = n41283 & n20704 ;
  assign n20708 = n20182 | n20707 ;
  assign n41297 = ~n20706 ;
  assign n20709 = n41297 & n20708 ;
  assign n41298 = ~n20709 ;
  assign n20710 = n3631 & n41298 ;
  assign n20711 = n173 | n20710 ;
  assign n41299 = ~n20711 ;
  assign n20712 = n20693 & n41299 ;
  assign n20713 = n20216 | n20712 ;
  assign n41300 = ~n20695 ;
  assign n20714 = n41300 & n20713 ;
  assign n41301 = ~n20714 ;
  assign n20715 = n174 & n41301 ;
  assign n41302 = ~n19876 ;
  assign n19898 = n19407 & n41302 ;
  assign n19899 = n40917 & n19898 ;
  assign n20171 = n19899 & n142 ;
  assign n19897 = n19865 | n19876 ;
  assign n41303 = ~n19897 ;
  assign n20172 = n41303 & n142 ;
  assign n20173 = n19407 | n20172 ;
  assign n41304 = ~n20171 ;
  assign n20174 = n41304 & n20173 ;
  assign n20696 = n174 | n20695 ;
  assign n41305 = ~n20696 ;
  assign n20716 = n41305 & n20713 ;
  assign n20717 = n20174 | n20716 ;
  assign n41306 = ~n20715 ;
  assign n20718 = n41306 & n20717 ;
  assign n41307 = ~n20718 ;
  assign n20719 = n2753 & n41307 ;
  assign n19896 = n19879 | n19880 ;
  assign n41308 = ~n19896 ;
  assign n20195 = n41308 & n142 ;
  assign n20196 = n19415 | n20195 ;
  assign n19857 = n19415 & n40909 ;
  assign n41309 = ~n19880 ;
  assign n19895 = n19857 & n41309 ;
  assign n20210 = n19895 & n142 ;
  assign n41310 = ~n20210 ;
  assign n20211 = n20196 & n41310 ;
  assign n20727 = n41289 & n20708 ;
  assign n20728 = n20267 | n20727 ;
  assign n41311 = ~n20710 ;
  assign n20729 = n41311 & n20728 ;
  assign n41312 = ~n20729 ;
  assign n20730 = n173 & n41312 ;
  assign n20731 = n41299 & n20728 ;
  assign n20732 = n20216 | n20731 ;
  assign n41313 = ~n20730 ;
  assign n20733 = n41313 & n20732 ;
  assign n41314 = ~n20733 ;
  assign n20734 = n174 & n41314 ;
  assign n20735 = n2753 | n20734 ;
  assign n41315 = ~n20735 ;
  assign n20736 = n20717 & n41315 ;
  assign n20737 = n20211 | n20736 ;
  assign n41316 = ~n20719 ;
  assign n20738 = n41316 & n20737 ;
  assign n41317 = ~n20738 ;
  assign n20739 = n176 & n41317 ;
  assign n19892 = n19883 | n19886 ;
  assign n41318 = ~n19892 ;
  assign n20294 = n41318 & n142 ;
  assign n20295 = n19485 | n20294 ;
  assign n41319 = ~n19886 ;
  assign n19893 = n19485 & n41319 ;
  assign n19894 = n40936 & n19893 ;
  assign n20297 = n19894 & n142 ;
  assign n41320 = ~n20297 ;
  assign n20298 = n20295 & n41320 ;
  assign n20720 = n2431 | n20719 ;
  assign n41321 = ~n20720 ;
  assign n20740 = n41321 & n20737 ;
  assign n20743 = n20298 | n20740 ;
  assign n41322 = ~n20739 ;
  assign n20744 = n41322 & n20743 ;
  assign n41323 = ~n20744 ;
  assign n20745 = n177 & n41323 ;
  assign n19891 = n19889 | n19890 ;
  assign n41324 = ~n19891 ;
  assign n20299 = n41324 & n142 ;
  assign n20300 = n19934 | n20299 ;
  assign n19941 = n40925 & n19934 ;
  assign n41325 = ~n19890 ;
  assign n19942 = n41325 & n19941 ;
  assign n20303 = n19942 & n142 ;
  assign n41326 = ~n20303 ;
  assign n20304 = n20300 & n41326 ;
  assign n20751 = n41305 & n20732 ;
  assign n20752 = n20174 | n20751 ;
  assign n41327 = ~n20734 ;
  assign n20753 = n41327 & n20752 ;
  assign n41328 = ~n20753 ;
  assign n20754 = n175 & n41328 ;
  assign n20755 = n41315 & n20752 ;
  assign n20756 = n20211 | n20755 ;
  assign n41329 = ~n20754 ;
  assign n20757 = n41329 & n20756 ;
  assign n41330 = ~n20757 ;
  assign n20758 = n2431 & n41330 ;
  assign n20759 = n177 | n20758 ;
  assign n41331 = ~n20759 ;
  assign n20760 = n20743 & n41331 ;
  assign n20761 = n20304 | n20760 ;
  assign n41332 = ~n20745 ;
  assign n20762 = n41332 & n20761 ;
  assign n41333 = ~n20762 ;
  assign n20763 = n178 & n41333 ;
  assign n19940 = n19937 | n19939 ;
  assign n41334 = ~n19940 ;
  assign n20308 = n41334 & n142 ;
  assign n20309 = n19953 | n20308 ;
  assign n41335 = ~n19939 ;
  assign n19968 = n41335 & n19953 ;
  assign n19969 = n40949 & n19968 ;
  assign n20311 = n19969 & n142 ;
  assign n41336 = ~n20311 ;
  assign n20312 = n20309 & n41336 ;
  assign n20746 = n178 | n20745 ;
  assign n41337 = ~n20746 ;
  assign n20764 = n41337 & n20761 ;
  assign n20767 = n20312 | n20764 ;
  assign n41338 = ~n20763 ;
  assign n20768 = n41338 & n20767 ;
  assign n41339 = ~n20768 ;
  assign n20769 = n1707 & n41339 ;
  assign n19989 = n19972 | n19973 ;
  assign n41340 = ~n19989 ;
  assign n20286 = n41340 & n142 ;
  assign n20287 = n19603 | n20286 ;
  assign n19958 = n19603 & n40941 ;
  assign n41341 = ~n19973 ;
  assign n19988 = n19958 & n41341 ;
  assign n20313 = n19988 & n142 ;
  assign n41342 = ~n20313 ;
  assign n20314 = n20287 & n41342 ;
  assign n20775 = n41321 & n20756 ;
  assign n20776 = n20298 | n20775 ;
  assign n41343 = ~n20758 ;
  assign n20777 = n41343 & n20776 ;
  assign n41344 = ~n20777 ;
  assign n20778 = n177 & n41344 ;
  assign n20779 = n41331 & n20776 ;
  assign n20780 = n20304 | n20779 ;
  assign n41345 = ~n20778 ;
  assign n20781 = n41345 & n20780 ;
  assign n41346 = ~n20781 ;
  assign n20782 = n178 & n41346 ;
  assign n20783 = n1707 | n20782 ;
  assign n41347 = ~n20783 ;
  assign n20784 = n20767 & n41347 ;
  assign n20785 = n20314 | n20784 ;
  assign n41348 = ~n20769 ;
  assign n20786 = n41348 & n20785 ;
  assign n41349 = ~n20786 ;
  assign n20787 = n180 & n41349 ;
  assign n19987 = n19976 | n19979 ;
  assign n41350 = ~n19987 ;
  assign n20315 = n41350 & n142 ;
  assign n20316 = n19502 | n20315 ;
  assign n41351 = ~n19979 ;
  assign n19985 = n19502 & n41351 ;
  assign n19986 = n40968 & n19985 ;
  assign n20317 = n19986 & n142 ;
  assign n41352 = ~n20317 ;
  assign n20318 = n20316 & n41352 ;
  assign n20770 = n1487 | n20769 ;
  assign n41353 = ~n20770 ;
  assign n20788 = n41353 & n20785 ;
  assign n20789 = n20318 | n20788 ;
  assign n41354 = ~n20787 ;
  assign n20790 = n41354 & n20789 ;
  assign n41355 = ~n20790 ;
  assign n20791 = n181 & n41355 ;
  assign n19984 = n19982 | n19983 ;
  assign n41356 = ~n19984 ;
  assign n20319 = n41356 & n142 ;
  assign n20320 = n19993 | n20319 ;
  assign n20000 = n40957 & n19993 ;
  assign n41357 = ~n19983 ;
  assign n20001 = n41357 & n20000 ;
  assign n20321 = n20001 & n142 ;
  assign n41358 = ~n20321 ;
  assign n20322 = n20320 & n41358 ;
  assign n20799 = n41337 & n20780 ;
  assign n20800 = n20312 | n20799 ;
  assign n41359 = ~n20782 ;
  assign n20801 = n41359 & n20800 ;
  assign n41360 = ~n20801 ;
  assign n20802 = n179 & n41360 ;
  assign n20803 = n41347 & n20800 ;
  assign n20804 = n20314 | n20803 ;
  assign n41361 = ~n20802 ;
  assign n20805 = n41361 & n20804 ;
  assign n41362 = ~n20805 ;
  assign n20806 = n1487 & n41362 ;
  assign n20807 = n181 | n20806 ;
  assign n41363 = ~n20807 ;
  assign n20808 = n20789 & n41363 ;
  assign n20809 = n20322 | n20808 ;
  assign n41364 = ~n20791 ;
  assign n20810 = n41364 & n20809 ;
  assign n41365 = ~n20810 ;
  assign n20811 = n182 & n41365 ;
  assign n41366 = ~n19998 ;
  assign n20018 = n41366 & n20007 ;
  assign n20019 = n40981 & n20018 ;
  assign n20310 = n20019 & n142 ;
  assign n19999 = n19996 | n19998 ;
  assign n41367 = ~n19999 ;
  assign n20323 = n41367 & n142 ;
  assign n20324 = n20007 | n20323 ;
  assign n41368 = ~n20310 ;
  assign n20325 = n41368 & n20324 ;
  assign n20792 = n182 | n20791 ;
  assign n41369 = ~n20792 ;
  assign n20812 = n41369 & n20809 ;
  assign n20815 = n20325 | n20812 ;
  assign n41370 = ~n20811 ;
  assign n20816 = n41370 & n20815 ;
  assign n41371 = ~n20816 ;
  assign n20817 = n996 & n41371 ;
  assign n20012 = n19949 & n40973 ;
  assign n41372 = ~n20023 ;
  assign n20030 = n20012 & n41372 ;
  assign n20191 = n20030 & n142 ;
  assign n20031 = n20022 | n20023 ;
  assign n41373 = ~n20031 ;
  assign n20234 = n41373 & n142 ;
  assign n20235 = n19949 | n20234 ;
  assign n41374 = ~n20191 ;
  assign n20236 = n41374 & n20235 ;
  assign n20823 = n41353 & n20804 ;
  assign n20824 = n20318 | n20823 ;
  assign n41375 = ~n20806 ;
  assign n20825 = n41375 & n20824 ;
  assign n41376 = ~n20825 ;
  assign n20826 = n181 & n41376 ;
  assign n20827 = n41363 & n20824 ;
  assign n20828 = n20322 | n20827 ;
  assign n41377 = ~n20826 ;
  assign n20829 = n41377 & n20828 ;
  assign n41378 = ~n20829 ;
  assign n20830 = n182 & n41378 ;
  assign n20831 = n183 | n20830 ;
  assign n41379 = ~n20831 ;
  assign n20832 = n20815 & n41379 ;
  assign n20833 = n20236 | n20832 ;
  assign n41380 = ~n20817 ;
  assign n20834 = n41380 & n20833 ;
  assign n41381 = ~n20834 ;
  assign n20835 = n184 & n41381 ;
  assign n41382 = ~n20028 ;
  assign n20043 = n41382 & n20037 ;
  assign n20044 = n41000 & n20043 ;
  assign n20296 = n20044 & n142 ;
  assign n20029 = n20026 | n20028 ;
  assign n41383 = ~n20029 ;
  assign n20305 = n41383 & n142 ;
  assign n20306 = n20037 | n20305 ;
  assign n41384 = ~n20296 ;
  assign n20307 = n41384 & n20306 ;
  assign n20818 = n838 | n20817 ;
  assign n41385 = ~n20818 ;
  assign n20836 = n41385 & n20833 ;
  assign n20839 = n20307 | n20836 ;
  assign n41386 = ~n20835 ;
  assign n20840 = n41386 & n20839 ;
  assign n41387 = ~n20840 ;
  assign n20841 = n185 & n41387 ;
  assign n20049 = n20047 | n20048 ;
  assign n41388 = ~n20049 ;
  assign n20301 = n41388 & n142 ;
  assign n20302 = n20051 | n20301 ;
  assign n20058 = n40989 & n20051 ;
  assign n41389 = ~n20048 ;
  assign n20059 = n41389 & n20058 ;
  assign n20326 = n20059 & n142 ;
  assign n41390 = ~n20326 ;
  assign n20327 = n20302 & n41390 ;
  assign n20847 = n41369 & n20828 ;
  assign n20848 = n20325 | n20847 ;
  assign n41391 = ~n20830 ;
  assign n20849 = n41391 & n20848 ;
  assign n41392 = ~n20849 ;
  assign n20850 = n183 & n41392 ;
  assign n20851 = n41379 & n20848 ;
  assign n20852 = n20236 | n20851 ;
  assign n41393 = ~n20850 ;
  assign n20853 = n41393 & n20852 ;
  assign n41394 = ~n20853 ;
  assign n20854 = n838 & n41394 ;
  assign n20855 = n185 | n20854 ;
  assign n41395 = ~n20855 ;
  assign n20856 = n20839 & n41395 ;
  assign n20857 = n20327 | n20856 ;
  assign n41396 = ~n20841 ;
  assign n20858 = n41396 & n20857 ;
  assign n41397 = ~n20858 ;
  assign n20859 = n186 & n41397 ;
  assign n20842 = n186 | n20841 ;
  assign n41398 = ~n20842 ;
  assign n20860 = n41398 & n20857 ;
  assign n41399 = ~n20056 ;
  assign n20122 = n41399 & n20106 ;
  assign n20123 = n41016 & n20122 ;
  assign n20329 = n20123 & n142 ;
  assign n20057 = n20054 | n20056 ;
  assign n41400 = ~n20057 ;
  assign n20328 = n41400 & n142 ;
  assign n20927 = n20106 | n20328 ;
  assign n41401 = ~n20329 ;
  assign n20928 = n41401 & n20927 ;
  assign n20929 = n20860 | n20928 ;
  assign n41402 = ~n20859 ;
  assign n20930 = n41402 & n20929 ;
  assign n41403 = ~n20930 ;
  assign n20931 = n528 & n41403 ;
  assign n20111 = n19411 & n41005 ;
  assign n41404 = ~n20127 ;
  assign n20921 = n20111 & n41404 ;
  assign n20922 = n142 & n20921 ;
  assign n20923 = n20126 | n20127 ;
  assign n41405 = ~n20923 ;
  assign n20924 = n142 & n41405 ;
  assign n20925 = n19411 | n20924 ;
  assign n41406 = ~n20922 ;
  assign n20926 = n41406 & n20925 ;
  assign n20864 = n41385 & n20852 ;
  assign n20865 = n20307 | n20864 ;
  assign n41407 = ~n20854 ;
  assign n20866 = n41407 & n20865 ;
  assign n41408 = ~n20866 ;
  assign n20867 = n185 & n41408 ;
  assign n20868 = n41395 & n20865 ;
  assign n20869 = n20327 | n20868 ;
  assign n41409 = ~n20867 ;
  assign n20870 = n41409 & n20869 ;
  assign n41410 = ~n20870 ;
  assign n20871 = n186 & n41410 ;
  assign n20872 = n528 | n20871 ;
  assign n41411 = ~n20872 ;
  assign n20934 = n41411 & n20929 ;
  assign n20935 = n20926 | n20934 ;
  assign n41412 = ~n20931 ;
  assign n20936 = n41412 & n20935 ;
  assign n41413 = ~n20936 ;
  assign n20937 = n188 & n41413 ;
  assign n41414 = ~n20142 ;
  assign n20914 = n20104 & n41414 ;
  assign n20915 = n41032 & n20914 ;
  assign n20916 = n142 & n20915 ;
  assign n20917 = n20130 | n20142 ;
  assign n41415 = ~n20917 ;
  assign n20918 = n142 & n41415 ;
  assign n20919 = n20104 | n20918 ;
  assign n41416 = ~n20916 ;
  assign n20920 = n41416 & n20919 ;
  assign n20932 = n413 | n20931 ;
  assign n41417 = ~n20932 ;
  assign n20938 = n41417 & n20935 ;
  assign n20939 = n20920 | n20938 ;
  assign n41418 = ~n20937 ;
  assign n20940 = n41418 & n20939 ;
  assign n41419 = ~n20940 ;
  assign n20941 = n189 & n41419 ;
  assign n20121 = n20097 & n41021 ;
  assign n41420 = ~n20146 ;
  assign n20908 = n20121 & n41420 ;
  assign n20909 = n142 & n20908 ;
  assign n20910 = n20145 | n20146 ;
  assign n41421 = ~n20910 ;
  assign n20911 = n142 & n41421 ;
  assign n20912 = n20097 | n20911 ;
  assign n41422 = ~n20909 ;
  assign n20913 = n41422 & n20912 ;
  assign n20874 = n41398 & n20869 ;
  assign n20950 = n20874 | n20928 ;
  assign n41423 = ~n20871 ;
  assign n20951 = n41423 & n20950 ;
  assign n41424 = ~n20951 ;
  assign n20952 = n187 & n41424 ;
  assign n20953 = n41411 & n20950 ;
  assign n20954 = n20926 | n20953 ;
  assign n41425 = ~n20952 ;
  assign n20955 = n41425 & n20954 ;
  assign n41426 = ~n20955 ;
  assign n20956 = n413 & n41426 ;
  assign n20957 = n189 | n20956 ;
  assign n41427 = ~n20957 ;
  assign n20958 = n20939 & n41427 ;
  assign n20959 = n20913 | n20958 ;
  assign n41428 = ~n20941 ;
  assign n20960 = n41428 & n20959 ;
  assign n41429 = ~n20960 ;
  assign n20961 = n190 & n41429 ;
  assign n20901 = n20149 | n20151 ;
  assign n41430 = ~n20901 ;
  assign n20902 = n142 & n41430 ;
  assign n20903 = n20091 | n20902 ;
  assign n41431 = ~n20151 ;
  assign n20904 = n20091 & n41431 ;
  assign n20905 = n41038 & n20904 ;
  assign n20906 = n142 & n20905 ;
  assign n41432 = ~n20906 ;
  assign n20907 = n20903 & n41432 ;
  assign n20942 = n190 | n20941 ;
  assign n41433 = ~n20942 ;
  assign n20962 = n41433 & n20959 ;
  assign n20963 = n20907 | n20962 ;
  assign n41434 = ~n20961 ;
  assign n20964 = n41434 & n20963 ;
  assign n41435 = ~n20964 ;
  assign n20965 = n287 & n41435 ;
  assign n41436 = ~n20965 ;
  assign n20967 = n20891 & n41436 ;
  assign n41437 = ~n20139 ;
  assign n20141 = n20084 & n41437 ;
  assign n41438 = ~n20155 ;
  assign n20895 = n20141 & n41438 ;
  assign n20896 = n142 & n20895 ;
  assign n20897 = n20154 | n20155 ;
  assign n41439 = ~n20897 ;
  assign n20898 = n142 & n41439 ;
  assign n20899 = n20084 | n20898 ;
  assign n41440 = ~n20896 ;
  assign n20900 = n41440 & n20899 ;
  assign n20973 = n41417 & n20954 ;
  assign n20974 = n20920 | n20973 ;
  assign n41441 = ~n20956 ;
  assign n20975 = n41441 & n20974 ;
  assign n41442 = ~n20975 ;
  assign n20976 = n189 & n41442 ;
  assign n20977 = n41427 & n20974 ;
  assign n20978 = n20913 | n20977 ;
  assign n41443 = ~n20976 ;
  assign n20979 = n41443 & n20978 ;
  assign n41444 = ~n20979 ;
  assign n20980 = n190 & n41444 ;
  assign n20981 = n287 | n20980 ;
  assign n41445 = ~n20981 ;
  assign n20982 = n20963 & n41445 ;
  assign n20983 = n20900 | n20982 ;
  assign n20984 = n20967 & n20983 ;
  assign n20985 = n20878 | n20984 ;
  assign n41446 = ~n20165 ;
  assign n20351 = n41446 & n142 ;
  assign n20875 = n20168 | n20351 ;
  assign n20892 = n20875 | n20891 ;
  assign n20988 = n41436 & n20983 ;
  assign n20989 = n20892 | n20988 ;
  assign n20990 = n31336 & n20989 ;
  assign n141 = n20985 | n20990 ;
  assign n41447 = ~n20891 ;
  assign n21186 = n41447 & n141 ;
  assign n41448 = ~n21186 ;
  assign n21187 = n20988 & n41448 ;
  assign n21208 = n20891 | n20988 ;
  assign n21210 = n192 & n21208 ;
  assign n41449 = ~n21187 ;
  assign n21211 = n41449 & n21210 ;
  assign n20887 = n20877 | n20886 ;
  assign n41450 = ~n20887 ;
  assign n20893 = n41450 & n20890 ;
  assign n41451 = ~n20334 ;
  assign n20894 = n41451 & n20893 ;
  assign n41452 = ~n20984 ;
  assign n21749 = n20894 & n41452 ;
  assign n41453 = ~n20990 ;
  assign n21750 = n41453 & n21749 ;
  assign n21751 = n21211 | n21750 ;
  assign n41454 = ~n20962 ;
  assign n20968 = n20907 & n41454 ;
  assign n20969 = n41434 & n20968 ;
  assign n21185 = n20969 & n141 ;
  assign n21761 = n20962 | n20980 ;
  assign n41455 = ~n21761 ;
  assign n21762 = n141 & n41455 ;
  assign n21763 = n20907 | n21762 ;
  assign n41456 = ~n21185 ;
  assign n21764 = n41456 & n21763 ;
  assign n236 = x22 | x23 ;
  assign n237 = x24 | n236 ;
  assign n21065 = x24 & n141 ;
  assign n41457 = ~n21065 ;
  assign n21088 = n237 & n41457 ;
  assign n41458 = ~n21088 ;
  assign n21089 = n142 & n41458 ;
  assign n19382 = n237 & n41067 ;
  assign n19478 = n19382 & n41051 ;
  assign n20883 = n19478 & n41052 ;
  assign n20884 = n41053 & n20883 ;
  assign n21066 = n20884 & n41457 ;
  assign n41459 = ~n233 ;
  assign n21064 = n41459 & n141 ;
  assign n41460 = ~x24 ;
  assign n21196 = n41460 & n141 ;
  assign n41461 = ~n21196 ;
  assign n21197 = x25 & n41461 ;
  assign n21198 = n21064 | n21197 ;
  assign n21199 = n21066 | n21198 ;
  assign n41462 = ~n21089 ;
  assign n21200 = n41462 & n21199 ;
  assign n41463 = ~n21200 ;
  assign n21201 = n19362 & n41463 ;
  assign n238 = n41460 & n236 ;
  assign n41464 = ~n141 ;
  assign n21188 = x24 & n41464 ;
  assign n21189 = n238 | n21188 ;
  assign n41465 = ~n21189 ;
  assign n21190 = n142 & n41465 ;
  assign n21191 = n19362 | n21190 ;
  assign n41466 = ~n21191 ;
  assign n21205 = n41466 & n21199 ;
  assign n41467 = ~n20877 ;
  assign n20879 = n142 & n41467 ;
  assign n20880 = n41451 & n20879 ;
  assign n21212 = n20880 & n41452 ;
  assign n21213 = n41453 & n21212 ;
  assign n21214 = n21064 | n21213 ;
  assign n21215 = x26 & n21214 ;
  assign n21216 = x26 | n21213 ;
  assign n21217 = n21064 | n21216 ;
  assign n41468 = ~n21215 ;
  assign n21218 = n41468 & n21217 ;
  assign n21219 = n21205 | n21218 ;
  assign n41469 = ~n21201 ;
  assign n21220 = n41469 & n21219 ;
  assign n41470 = ~n21220 ;
  assign n21221 = n18797 & n41470 ;
  assign n20344 = n20335 | n20342 ;
  assign n41471 = ~n20344 ;
  assign n21082 = n41471 & n141 ;
  assign n21083 = n20354 | n21082 ;
  assign n20357 = n41471 & n20354 ;
  assign n21086 = n20357 & n141 ;
  assign n41472 = ~n21086 ;
  assign n21087 = n21083 & n41472 ;
  assign n21202 = n18797 | n21201 ;
  assign n41473 = ~n21202 ;
  assign n21224 = n41473 & n21219 ;
  assign n21225 = n21087 | n21224 ;
  assign n41474 = ~n21221 ;
  assign n21226 = n41474 & n21225 ;
  assign n41475 = ~n21226 ;
  assign n21227 = n145 & n41475 ;
  assign n20362 = n20356 | n20361 ;
  assign n41476 = ~n20362 ;
  assign n21084 = n41476 & n141 ;
  assign n21085 = n20370 | n21084 ;
  assign n41477 = ~n20356 ;
  assign n20390 = n41477 & n20370 ;
  assign n20391 = n41069 & n20390 ;
  assign n21192 = n20391 & n141 ;
  assign n41478 = ~n21192 ;
  assign n21193 = n21085 & n41478 ;
  assign n21222 = n145 | n21221 ;
  assign n41479 = ~n21222 ;
  assign n21228 = n41479 & n21225 ;
  assign n21229 = n21193 | n21228 ;
  assign n41480 = ~n21227 ;
  assign n21230 = n41480 & n21229 ;
  assign n41481 = ~n21230 ;
  assign n21231 = n146 & n41481 ;
  assign n20389 = n20373 | n20376 ;
  assign n41482 = ~n20389 ;
  assign n21058 = n41482 & n141 ;
  assign n21059 = n20347 | n21058 ;
  assign n20375 = n20347 & n41074 ;
  assign n41483 = ~n20376 ;
  assign n20388 = n20375 & n41483 ;
  assign n21194 = n20388 & n141 ;
  assign n41484 = ~n21194 ;
  assign n21195 = n21059 & n41484 ;
  assign n21203 = n143 & n41463 ;
  assign n21090 = n143 | n21089 ;
  assign n41485 = ~n21090 ;
  assign n21207 = n41485 & n21199 ;
  assign n21241 = n21207 | n21218 ;
  assign n41486 = ~n21203 ;
  assign n21242 = n41486 & n21241 ;
  assign n41487 = ~n21242 ;
  assign n21243 = n144 & n41487 ;
  assign n21244 = n41473 & n21241 ;
  assign n21245 = n21087 | n21244 ;
  assign n41488 = ~n21243 ;
  assign n21246 = n41488 & n21245 ;
  assign n41489 = ~n21246 ;
  assign n21247 = n145 & n41489 ;
  assign n21248 = n146 | n21247 ;
  assign n41490 = ~n21248 ;
  assign n21249 = n21229 & n41490 ;
  assign n21250 = n21195 | n21249 ;
  assign n41491 = ~n21231 ;
  assign n21251 = n41491 & n21250 ;
  assign n41492 = ~n21251 ;
  assign n21252 = n147 & n41492 ;
  assign n20414 = n20380 | n20398 ;
  assign n41493 = ~n20414 ;
  assign n21060 = n41493 & n141 ;
  assign n21061 = n20350 | n21060 ;
  assign n41494 = ~n20380 ;
  assign n20386 = n20350 & n41494 ;
  assign n20387 = n41081 & n20386 ;
  assign n21062 = n20387 & n141 ;
  assign n41495 = ~n21062 ;
  assign n21063 = n21061 & n41495 ;
  assign n21232 = n147 | n21231 ;
  assign n41496 = ~n21232 ;
  assign n21253 = n41496 & n21250 ;
  assign n21254 = n21063 | n21253 ;
  assign n41497 = ~n21252 ;
  assign n21255 = n41497 & n21254 ;
  assign n41498 = ~n21255 ;
  assign n21256 = n15807 & n41498 ;
  assign n20413 = n20383 | n20400 ;
  assign n41499 = ~n20413 ;
  assign n21001 = n41499 & n141 ;
  assign n21002 = n20337 | n21001 ;
  assign n20385 = n20337 & n41092 ;
  assign n41500 = ~n20400 ;
  assign n20412 = n20385 & n41500 ;
  assign n21098 = n20412 & n141 ;
  assign n41501 = ~n21098 ;
  assign n21099 = n21002 & n41501 ;
  assign n21264 = n41479 & n21245 ;
  assign n21265 = n21193 | n21264 ;
  assign n41502 = ~n21247 ;
  assign n21266 = n41502 & n21265 ;
  assign n41503 = ~n21266 ;
  assign n21267 = n146 & n41503 ;
  assign n21268 = n41490 & n21265 ;
  assign n21269 = n21195 | n21268 ;
  assign n41504 = ~n21267 ;
  assign n21270 = n41504 & n21269 ;
  assign n41505 = ~n21270 ;
  assign n21271 = n16322 & n41505 ;
  assign n21272 = n148 | n21271 ;
  assign n41506 = ~n21272 ;
  assign n21273 = n21254 & n41506 ;
  assign n21274 = n21099 | n21273 ;
  assign n41507 = ~n21256 ;
  assign n21275 = n41507 & n21274 ;
  assign n41508 = ~n21275 ;
  assign n21276 = n149 & n41508 ;
  assign n20438 = n20404 | n20422 ;
  assign n41509 = ~n20438 ;
  assign n21056 = n41509 & n141 ;
  assign n21057 = n20291 | n21056 ;
  assign n41510 = ~n20404 ;
  assign n20410 = n20291 & n41510 ;
  assign n20411 = n41098 & n20410 ;
  assign n21092 = n20411 & n141 ;
  assign n41511 = ~n21092 ;
  assign n21093 = n21057 & n41511 ;
  assign n21257 = n149 | n21256 ;
  assign n41512 = ~n21257 ;
  assign n21277 = n41512 & n21274 ;
  assign n21278 = n21093 | n21277 ;
  assign n41513 = ~n21276 ;
  assign n21279 = n41513 & n21278 ;
  assign n41514 = ~n21279 ;
  assign n21280 = n150 & n41514 ;
  assign n20437 = n20407 | n20424 ;
  assign n41515 = ~n20437 ;
  assign n21008 = n41515 & n141 ;
  assign n21009 = n20260 | n21008 ;
  assign n20409 = n20260 & n41108 ;
  assign n41516 = ~n20424 ;
  assign n20436 = n20409 & n41516 ;
  assign n21080 = n20436 & n141 ;
  assign n41517 = ~n21080 ;
  assign n21081 = n21009 & n41517 ;
  assign n21288 = n41496 & n21269 ;
  assign n21289 = n21063 | n21288 ;
  assign n41518 = ~n21271 ;
  assign n21290 = n41518 & n21289 ;
  assign n41519 = ~n21290 ;
  assign n21291 = n148 & n41519 ;
  assign n21292 = n41506 & n21289 ;
  assign n21293 = n21099 | n21292 ;
  assign n41520 = ~n21291 ;
  assign n21294 = n41520 & n21293 ;
  assign n41521 = ~n21294 ;
  assign n21295 = n149 & n41521 ;
  assign n21296 = n150 | n21295 ;
  assign n41522 = ~n21296 ;
  assign n21297 = n21278 & n41522 ;
  assign n21298 = n21081 | n21297 ;
  assign n41523 = ~n21280 ;
  assign n21299 = n41523 & n21298 ;
  assign n41524 = ~n21299 ;
  assign n21300 = n151 & n41524 ;
  assign n41525 = ~n20428 ;
  assign n20434 = n20250 & n41525 ;
  assign n20435 = n41114 & n20434 ;
  assign n21094 = n20435 & n141 ;
  assign n20462 = n20428 | n20446 ;
  assign n41526 = ~n20462 ;
  assign n21103 = n41526 & n141 ;
  assign n21104 = n20250 | n21103 ;
  assign n41527 = ~n21094 ;
  assign n21105 = n41527 & n21104 ;
  assign n21281 = n151 | n21280 ;
  assign n41528 = ~n21281 ;
  assign n21301 = n41528 & n21298 ;
  assign n21302 = n21105 | n21301 ;
  assign n41529 = ~n21300 ;
  assign n21303 = n41529 & n21302 ;
  assign n41530 = ~n21303 ;
  assign n21304 = n13079 & n41530 ;
  assign n20433 = n20228 & n41124 ;
  assign n41531 = ~n20448 ;
  assign n20460 = n20433 & n41531 ;
  assign n21069 = n20460 & n141 ;
  assign n20461 = n20431 | n20448 ;
  assign n41532 = ~n20461 ;
  assign n21073 = n41532 & n141 ;
  assign n21074 = n20228 | n21073 ;
  assign n41533 = ~n21069 ;
  assign n21075 = n41533 & n21074 ;
  assign n21312 = n41512 & n21293 ;
  assign n21313 = n21093 | n21312 ;
  assign n41534 = ~n21295 ;
  assign n21314 = n41534 & n21313 ;
  assign n41535 = ~n21314 ;
  assign n21315 = n150 & n41535 ;
  assign n21316 = n41522 & n21313 ;
  assign n21317 = n21081 | n21316 ;
  assign n41536 = ~n21315 ;
  assign n21318 = n41536 & n21317 ;
  assign n41537 = ~n21318 ;
  assign n21319 = n13662 & n41537 ;
  assign n21320 = n152 | n21319 ;
  assign n41538 = ~n21320 ;
  assign n21321 = n21302 & n41538 ;
  assign n21322 = n21075 | n21321 ;
  assign n41539 = ~n21304 ;
  assign n21323 = n41539 & n21322 ;
  assign n41540 = ~n21323 ;
  assign n21324 = n153 & n41540 ;
  assign n20486 = n20452 | n20470 ;
  assign n41541 = ~n20486 ;
  assign n21031 = n41541 & n141 ;
  assign n21032 = n20252 | n21031 ;
  assign n41542 = ~n20452 ;
  assign n20458 = n20252 & n41542 ;
  assign n20459 = n41130 & n20458 ;
  assign n21109 = n20459 & n141 ;
  assign n41543 = ~n21109 ;
  assign n21110 = n21032 & n41543 ;
  assign n21305 = n153 | n21304 ;
  assign n41544 = ~n21305 ;
  assign n21325 = n41544 & n21322 ;
  assign n21326 = n21110 | n21325 ;
  assign n41545 = ~n21324 ;
  assign n21327 = n41545 & n21326 ;
  assign n41546 = ~n21327 ;
  assign n21328 = n154 & n41546 ;
  assign n20485 = n20455 | n20472 ;
  assign n41547 = ~n20485 ;
  assign n21067 = n41547 & n141 ;
  assign n21068 = n20276 | n21067 ;
  assign n20457 = n20276 & n41140 ;
  assign n41548 = ~n20472 ;
  assign n20484 = n20457 & n41548 ;
  assign n21123 = n20484 & n141 ;
  assign n41549 = ~n21123 ;
  assign n21124 = n21068 & n41549 ;
  assign n21336 = n41528 & n21317 ;
  assign n21337 = n21105 | n21336 ;
  assign n41550 = ~n21319 ;
  assign n21338 = n41550 & n21337 ;
  assign n41551 = ~n21338 ;
  assign n21339 = n152 & n41551 ;
  assign n21340 = n41538 & n21337 ;
  assign n21341 = n21075 | n21340 ;
  assign n41552 = ~n21339 ;
  assign n21342 = n41552 & n21341 ;
  assign n41553 = ~n21342 ;
  assign n21343 = n153 & n41553 ;
  assign n21344 = n154 | n21343 ;
  assign n41554 = ~n21344 ;
  assign n21345 = n21326 & n41554 ;
  assign n21346 = n21124 | n21345 ;
  assign n41555 = ~n21328 ;
  assign n21347 = n41555 & n21346 ;
  assign n41556 = ~n21347 ;
  assign n21348 = n155 & n41556 ;
  assign n20510 = n20476 | n20494 ;
  assign n41557 = ~n20510 ;
  assign n21033 = n41557 & n141 ;
  assign n21034 = n20257 | n21033 ;
  assign n41558 = ~n20476 ;
  assign n20482 = n20257 & n41558 ;
  assign n20483 = n41146 & n20482 ;
  assign n21127 = n20483 & n141 ;
  assign n41559 = ~n21127 ;
  assign n21128 = n21034 & n41559 ;
  assign n21329 = n11067 | n21328 ;
  assign n41560 = ~n21329 ;
  assign n21349 = n41560 & n21346 ;
  assign n21350 = n21128 | n21349 ;
  assign n41561 = ~n21348 ;
  assign n21351 = n41561 & n21350 ;
  assign n41562 = ~n21351 ;
  assign n21352 = n10657 & n41562 ;
  assign n20481 = n20279 & n41156 ;
  assign n41563 = ~n20496 ;
  assign n20508 = n20481 & n41563 ;
  assign n21010 = n20508 & n141 ;
  assign n20509 = n20479 | n20496 ;
  assign n41564 = ~n20509 ;
  assign n21095 = n41564 & n141 ;
  assign n21096 = n20279 | n21095 ;
  assign n41565 = ~n21010 ;
  assign n21097 = n41565 & n21096 ;
  assign n21360 = n41544 & n21341 ;
  assign n21361 = n21110 | n21360 ;
  assign n41566 = ~n21343 ;
  assign n21362 = n41566 & n21361 ;
  assign n41567 = ~n21362 ;
  assign n21363 = n154 & n41567 ;
  assign n21364 = n41554 & n21361 ;
  assign n21365 = n21124 | n21364 ;
  assign n41568 = ~n21363 ;
  assign n21366 = n41568 & n21365 ;
  assign n41569 = ~n21366 ;
  assign n21367 = n11067 & n41569 ;
  assign n21368 = n10657 | n21367 ;
  assign n41570 = ~n21368 ;
  assign n21369 = n21350 & n41570 ;
  assign n21370 = n21097 | n21369 ;
  assign n41571 = ~n21352 ;
  assign n21371 = n41571 & n21370 ;
  assign n41572 = ~n21371 ;
  assign n21372 = n157 & n41572 ;
  assign n41573 = ~n20500 ;
  assign n20506 = n20246 & n41573 ;
  assign n20507 = n41162 & n20506 ;
  assign n21044 = n20507 & n141 ;
  assign n20534 = n20500 | n20518 ;
  assign n41574 = ~n20534 ;
  assign n21070 = n41574 & n141 ;
  assign n21071 = n20246 | n21070 ;
  assign n41575 = ~n21044 ;
  assign n21072 = n41575 & n21071 ;
  assign n21353 = n157 | n21352 ;
  assign n41576 = ~n21353 ;
  assign n21373 = n41576 & n21370 ;
  assign n21374 = n21072 | n21373 ;
  assign n41577 = ~n21372 ;
  assign n21375 = n41577 & n21374 ;
  assign n41578 = ~n21375 ;
  assign n21376 = n158 & n41578 ;
  assign n20505 = n20289 & n41172 ;
  assign n41579 = ~n20520 ;
  assign n20532 = n20505 & n41579 ;
  assign n21050 = n20532 & n141 ;
  assign n20533 = n20503 | n20520 ;
  assign n41580 = ~n20533 ;
  assign n21106 = n41580 & n141 ;
  assign n21107 = n20289 | n21106 ;
  assign n41581 = ~n21050 ;
  assign n21108 = n41581 & n21107 ;
  assign n21384 = n41560 & n21365 ;
  assign n21385 = n21128 | n21384 ;
  assign n41582 = ~n21367 ;
  assign n21386 = n41582 & n21385 ;
  assign n41583 = ~n21386 ;
  assign n21387 = n156 & n41583 ;
  assign n21388 = n41570 & n21385 ;
  assign n21389 = n21097 | n21388 ;
  assign n41584 = ~n21387 ;
  assign n21390 = n41584 & n21389 ;
  assign n41585 = ~n21390 ;
  assign n21391 = n157 & n41585 ;
  assign n21392 = n158 | n21391 ;
  assign n41586 = ~n21392 ;
  assign n21393 = n21374 & n41586 ;
  assign n21394 = n21108 | n21393 ;
  assign n41587 = ~n21376 ;
  assign n21395 = n41587 & n21394 ;
  assign n41588 = ~n21395 ;
  assign n21396 = n159 & n41588 ;
  assign n20558 = n20524 | n20542 ;
  assign n41589 = ~n20558 ;
  assign n21042 = n41589 & n141 ;
  assign n21043 = n20281 | n21042 ;
  assign n41590 = ~n20524 ;
  assign n20530 = n20281 & n41590 ;
  assign n20531 = n41178 & n20530 ;
  assign n21051 = n20531 & n141 ;
  assign n41591 = ~n21051 ;
  assign n21052 = n21043 & n41591 ;
  assign n21377 = n8857 | n21376 ;
  assign n41592 = ~n21377 ;
  assign n21397 = n41592 & n21394 ;
  assign n21401 = n21052 | n21397 ;
  assign n41593 = ~n21396 ;
  assign n21402 = n41593 & n21401 ;
  assign n41594 = ~n21402 ;
  assign n21403 = n8534 & n41594 ;
  assign n20529 = n20225 & n41188 ;
  assign n41595 = ~n20544 ;
  assign n20556 = n20529 & n41595 ;
  assign n21021 = n20556 & n141 ;
  assign n20557 = n20527 | n20544 ;
  assign n41596 = ~n20557 ;
  assign n21028 = n41596 & n141 ;
  assign n21029 = n20225 | n21028 ;
  assign n41597 = ~n21021 ;
  assign n21030 = n41597 & n21029 ;
  assign n21408 = n41576 & n21389 ;
  assign n21409 = n21072 | n21408 ;
  assign n41598 = ~n21391 ;
  assign n21410 = n41598 & n21409 ;
  assign n41599 = ~n21410 ;
  assign n21411 = n158 & n41599 ;
  assign n21412 = n41586 & n21409 ;
  assign n21413 = n21108 | n21412 ;
  assign n41600 = ~n21411 ;
  assign n21414 = n41600 & n21413 ;
  assign n41601 = ~n21414 ;
  assign n21415 = n8857 & n41601 ;
  assign n21416 = n160 | n21415 ;
  assign n41602 = ~n21416 ;
  assign n21417 = n21401 & n41602 ;
  assign n21418 = n21030 | n21417 ;
  assign n41603 = ~n21403 ;
  assign n21419 = n41603 & n21418 ;
  assign n41604 = ~n21419 ;
  assign n21420 = n161 & n41604 ;
  assign n41605 = ~n20548 ;
  assign n20554 = n20274 & n41605 ;
  assign n20555 = n41194 & n20554 ;
  assign n21007 = n20555 & n141 ;
  assign n20582 = n20548 | n20566 ;
  assign n41606 = ~n20582 ;
  assign n21100 = n41606 & n141 ;
  assign n21101 = n20274 | n21100 ;
  assign n41607 = ~n21007 ;
  assign n21102 = n41607 & n21101 ;
  assign n21404 = n161 | n21403 ;
  assign n41608 = ~n21404 ;
  assign n21421 = n41608 & n21418 ;
  assign n21422 = n21102 | n21421 ;
  assign n41609 = ~n21420 ;
  assign n21423 = n41609 & n21422 ;
  assign n41610 = ~n21423 ;
  assign n21424 = n162 & n41610 ;
  assign n20553 = n20285 & n41204 ;
  assign n41611 = ~n20568 ;
  assign n20580 = n20553 & n41611 ;
  assign n21016 = n20580 & n141 ;
  assign n20581 = n20551 | n20568 ;
  assign n41612 = ~n20581 ;
  assign n21118 = n41612 & n141 ;
  assign n21119 = n20285 | n21118 ;
  assign n41613 = ~n21016 ;
  assign n21120 = n41613 & n21119 ;
  assign n21432 = n41592 & n21413 ;
  assign n21433 = n21052 | n21432 ;
  assign n41614 = ~n21415 ;
  assign n21434 = n41614 & n21433 ;
  assign n41615 = ~n21434 ;
  assign n21435 = n160 & n41615 ;
  assign n21436 = n41602 & n21433 ;
  assign n21437 = n21030 | n21436 ;
  assign n41616 = ~n21435 ;
  assign n21438 = n41616 & n21437 ;
  assign n41617 = ~n21438 ;
  assign n21439 = n161 & n41617 ;
  assign n21440 = n162 | n21439 ;
  assign n41618 = ~n21440 ;
  assign n21441 = n21422 & n41618 ;
  assign n21442 = n21120 | n21441 ;
  assign n41619 = ~n21424 ;
  assign n21443 = n41619 & n21442 ;
  assign n41620 = ~n21443 ;
  assign n21444 = n163 & n41620 ;
  assign n20606 = n20572 | n20590 ;
  assign n41621 = ~n20606 ;
  assign n21022 = n41621 & n141 ;
  assign n21023 = n20218 | n21022 ;
  assign n41622 = ~n20572 ;
  assign n20578 = n20218 & n41622 ;
  assign n20579 = n41210 & n20578 ;
  assign n21038 = n20579 & n141 ;
  assign n41623 = ~n21038 ;
  assign n21039 = n21023 & n41623 ;
  assign n21425 = n6889 | n21424 ;
  assign n41624 = ~n21425 ;
  assign n21445 = n41624 & n21442 ;
  assign n21446 = n21039 | n21445 ;
  assign n41625 = ~n21444 ;
  assign n21447 = n41625 & n21446 ;
  assign n41626 = ~n21447 ;
  assign n21448 = n6600 & n41626 ;
  assign n20605 = n20575 | n20592 ;
  assign n41627 = ~n20605 ;
  assign n21014 = n41627 & n141 ;
  assign n21015 = n20214 | n21014 ;
  assign n20577 = n20214 & n41220 ;
  assign n41628 = ~n20592 ;
  assign n20604 = n20577 & n41628 ;
  assign n21078 = n20604 & n141 ;
  assign n41629 = ~n21078 ;
  assign n21079 = n21015 & n41629 ;
  assign n21456 = n41608 & n21437 ;
  assign n21457 = n21102 | n21456 ;
  assign n41630 = ~n21439 ;
  assign n21458 = n41630 & n21457 ;
  assign n41631 = ~n21458 ;
  assign n21459 = n162 & n41631 ;
  assign n21460 = n41618 & n21457 ;
  assign n21461 = n21120 | n21460 ;
  assign n41632 = ~n21459 ;
  assign n21462 = n41632 & n21461 ;
  assign n41633 = ~n21462 ;
  assign n21463 = n6889 & n41633 ;
  assign n21464 = n6600 | n21463 ;
  assign n41634 = ~n21464 ;
  assign n21465 = n21446 & n41634 ;
  assign n21466 = n21079 | n21465 ;
  assign n41635 = ~n21448 ;
  assign n21467 = n41635 & n21466 ;
  assign n41636 = ~n21467 ;
  assign n21468 = n165 & n41636 ;
  assign n41637 = ~n20596 ;
  assign n20602 = n20238 & n41637 ;
  assign n20603 = n41226 & n20602 ;
  assign n21006 = n20603 & n141 ;
  assign n20630 = n20596 | n20614 ;
  assign n41638 = ~n20630 ;
  assign n21011 = n41638 & n141 ;
  assign n21012 = n20238 | n21011 ;
  assign n41639 = ~n21006 ;
  assign n21013 = n41639 & n21012 ;
  assign n21449 = n165 | n21448 ;
  assign n41640 = ~n21449 ;
  assign n21469 = n41640 & n21466 ;
  assign n21470 = n21013 | n21469 ;
  assign n41641 = ~n21468 ;
  assign n21471 = n41641 & n21470 ;
  assign n41642 = ~n21471 ;
  assign n21472 = n166 & n41642 ;
  assign n20629 = n20599 | n20616 ;
  assign n41643 = ~n20629 ;
  assign n21040 = n41643 & n141 ;
  assign n21041 = n20271 | n21040 ;
  assign n20601 = n20271 & n41236 ;
  assign n41644 = ~n20616 ;
  assign n20628 = n20601 & n41644 ;
  assign n21116 = n20628 & n141 ;
  assign n41645 = ~n21116 ;
  assign n21117 = n21041 & n41645 ;
  assign n21480 = n41624 & n21461 ;
  assign n21481 = n21039 | n21480 ;
  assign n41646 = ~n21463 ;
  assign n21482 = n41646 & n21481 ;
  assign n41647 = ~n21482 ;
  assign n21483 = n164 & n41647 ;
  assign n21484 = n41634 & n21481 ;
  assign n21485 = n21079 | n21484 ;
  assign n41648 = ~n21483 ;
  assign n21486 = n41648 & n21485 ;
  assign n41649 = ~n21486 ;
  assign n21487 = n165 & n41649 ;
  assign n21488 = n166 | n21487 ;
  assign n41650 = ~n21488 ;
  assign n21489 = n21470 & n41650 ;
  assign n21490 = n21117 | n21489 ;
  assign n41651 = ~n21472 ;
  assign n21491 = n41651 & n21490 ;
  assign n41652 = ~n21491 ;
  assign n21492 = n167 & n41652 ;
  assign n41653 = ~n20620 ;
  assign n20626 = n20203 & n41653 ;
  assign n20627 = n41242 & n20626 ;
  assign n20998 = n20627 & n141 ;
  assign n20654 = n20620 | n20638 ;
  assign n41654 = ~n20654 ;
  assign n21003 = n41654 & n141 ;
  assign n21004 = n20203 | n21003 ;
  assign n41655 = ~n20998 ;
  assign n21005 = n41655 & n21004 ;
  assign n21473 = n5352 | n21472 ;
  assign n41656 = ~n21473 ;
  assign n21493 = n41656 & n21490 ;
  assign n21494 = n21005 | n21493 ;
  assign n41657 = ~n21492 ;
  assign n21495 = n41657 & n21494 ;
  assign n41658 = ~n21495 ;
  assign n21496 = n4934 & n41658 ;
  assign n20653 = n20623 | n20640 ;
  assign n41659 = ~n20653 ;
  assign n20996 = n41659 & n141 ;
  assign n20997 = n20230 | n20996 ;
  assign n20625 = n20230 & n41252 ;
  assign n41660 = ~n20640 ;
  assign n20652 = n20625 & n41660 ;
  assign n21131 = n20652 & n141 ;
  assign n41661 = ~n21131 ;
  assign n21132 = n20997 & n41661 ;
  assign n21504 = n41640 & n21485 ;
  assign n21505 = n21013 | n21504 ;
  assign n41662 = ~n21487 ;
  assign n21506 = n41662 & n21505 ;
  assign n41663 = ~n21506 ;
  assign n21507 = n166 & n41663 ;
  assign n21508 = n41650 & n21505 ;
  assign n21509 = n21117 | n21508 ;
  assign n41664 = ~n21507 ;
  assign n21510 = n41664 & n21509 ;
  assign n41665 = ~n21510 ;
  assign n21511 = n5352 & n41665 ;
  assign n21512 = n4934 | n21511 ;
  assign n41666 = ~n21512 ;
  assign n21513 = n21494 & n41666 ;
  assign n21514 = n21132 | n21513 ;
  assign n41667 = ~n21496 ;
  assign n21515 = n41667 & n21514 ;
  assign n41668 = ~n21515 ;
  assign n21516 = n169 & n41668 ;
  assign n41669 = ~n20644 ;
  assign n20650 = n20190 & n41669 ;
  assign n20651 = n41258 & n20650 ;
  assign n20995 = n20651 & n141 ;
  assign n20678 = n20644 | n20662 ;
  assign n41670 = ~n20678 ;
  assign n21035 = n41670 & n141 ;
  assign n21036 = n20190 | n21035 ;
  assign n41671 = ~n20995 ;
  assign n21037 = n41671 & n21036 ;
  assign n21497 = n169 | n21496 ;
  assign n41672 = ~n21497 ;
  assign n21517 = n41672 & n21514 ;
  assign n21518 = n21037 | n21517 ;
  assign n41673 = ~n21516 ;
  assign n21519 = n41673 & n21518 ;
  assign n41674 = ~n21519 ;
  assign n21520 = n170 & n41674 ;
  assign n20649 = n20186 & n41268 ;
  assign n41675 = ~n20664 ;
  assign n20676 = n20649 & n41675 ;
  assign n20994 = n20676 & n141 ;
  assign n20677 = n20647 | n20664 ;
  assign n41676 = ~n20677 ;
  assign n21045 = n41676 & n141 ;
  assign n21046 = n20186 | n21045 ;
  assign n41677 = ~n20994 ;
  assign n21047 = n41677 & n21046 ;
  assign n21528 = n41656 & n21509 ;
  assign n21529 = n21005 | n21528 ;
  assign n41678 = ~n21511 ;
  assign n21530 = n41678 & n21529 ;
  assign n41679 = ~n21530 ;
  assign n21531 = n168 & n41679 ;
  assign n21532 = n41666 & n21529 ;
  assign n21533 = n21132 | n21532 ;
  assign n41680 = ~n21531 ;
  assign n21534 = n41680 & n21533 ;
  assign n41681 = ~n21534 ;
  assign n21535 = n169 & n41681 ;
  assign n21536 = n170 | n21535 ;
  assign n41682 = ~n21536 ;
  assign n21537 = n21518 & n41682 ;
  assign n21538 = n21047 | n21537 ;
  assign n41683 = ~n21520 ;
  assign n21539 = n41683 & n21538 ;
  assign n41684 = ~n21539 ;
  assign n21540 = n171 & n41684 ;
  assign n20702 = n20668 | n20686 ;
  assign n41685 = ~n20702 ;
  assign n20999 = n41685 & n141 ;
  assign n21000 = n20293 | n20999 ;
  assign n41686 = ~n20668 ;
  assign n20674 = n20293 & n41686 ;
  assign n20675 = n41274 & n20674 ;
  assign n21017 = n20675 & n141 ;
  assign n41687 = ~n21017 ;
  assign n21018 = n21000 & n41687 ;
  assign n21521 = n3940 | n21520 ;
  assign n41688 = ~n21521 ;
  assign n21541 = n41688 & n21538 ;
  assign n21542 = n21018 | n21541 ;
  assign n41689 = ~n21540 ;
  assign n21543 = n41689 & n21542 ;
  assign n41690 = ~n21543 ;
  assign n21544 = n3631 & n41690 ;
  assign n20701 = n20671 | n20688 ;
  assign n41691 = ~n20701 ;
  assign n20992 = n41691 & n141 ;
  assign n20993 = n20182 | n20992 ;
  assign n20673 = n20182 & n41284 ;
  assign n41692 = ~n20688 ;
  assign n20700 = n20673 & n41692 ;
  assign n21133 = n20700 & n141 ;
  assign n41693 = ~n21133 ;
  assign n21134 = n20993 & n41693 ;
  assign n21552 = n41672 & n21533 ;
  assign n21553 = n21037 | n21552 ;
  assign n41694 = ~n21535 ;
  assign n21554 = n41694 & n21553 ;
  assign n41695 = ~n21554 ;
  assign n21555 = n170 & n41695 ;
  assign n21556 = n41682 & n21553 ;
  assign n21557 = n21047 | n21556 ;
  assign n41696 = ~n21555 ;
  assign n21558 = n41696 & n21557 ;
  assign n41697 = ~n21558 ;
  assign n21559 = n3940 & n41697 ;
  assign n21560 = n3631 | n21559 ;
  assign n41698 = ~n21560 ;
  assign n21561 = n21542 & n41698 ;
  assign n21562 = n21134 | n21561 ;
  assign n41699 = ~n21544 ;
  assign n21563 = n41699 & n21562 ;
  assign n41700 = ~n21563 ;
  assign n21564 = n173 & n41700 ;
  assign n20726 = n20692 | n20710 ;
  assign n41701 = ~n20726 ;
  assign n21019 = n41701 & n141 ;
  assign n21020 = n20267 | n21019 ;
  assign n41702 = ~n20692 ;
  assign n20698 = n20267 & n41702 ;
  assign n20699 = n41290 & n20698 ;
  assign n21137 = n20699 & n141 ;
  assign n41703 = ~n21137 ;
  assign n21138 = n21020 & n41703 ;
  assign n21545 = n173 | n21544 ;
  assign n41704 = ~n21545 ;
  assign n21565 = n41704 & n21562 ;
  assign n21566 = n21138 | n21565 ;
  assign n41705 = ~n21564 ;
  assign n21567 = n41705 & n21566 ;
  assign n41706 = ~n21567 ;
  assign n21568 = n174 & n41706 ;
  assign n20697 = n20216 & n41300 ;
  assign n41707 = ~n20712 ;
  assign n20724 = n20697 & n41707 ;
  assign n21053 = n20724 & n141 ;
  assign n20725 = n20695 | n20712 ;
  assign n41708 = ~n20725 ;
  assign n21111 = n41708 & n141 ;
  assign n21112 = n20216 | n21111 ;
  assign n41709 = ~n21053 ;
  assign n21113 = n41709 & n21112 ;
  assign n21576 = n41688 & n21557 ;
  assign n21577 = n21018 | n21576 ;
  assign n41710 = ~n21559 ;
  assign n21578 = n41710 & n21577 ;
  assign n41711 = ~n21578 ;
  assign n21579 = n172 & n41711 ;
  assign n21580 = n41698 & n21577 ;
  assign n21581 = n21134 | n21580 ;
  assign n41712 = ~n21579 ;
  assign n21582 = n41712 & n21581 ;
  assign n41713 = ~n21582 ;
  assign n21583 = n173 & n41713 ;
  assign n21584 = n174 | n21583 ;
  assign n41714 = ~n21584 ;
  assign n21585 = n21566 & n41714 ;
  assign n21586 = n21113 | n21585 ;
  assign n41715 = ~n21568 ;
  assign n21587 = n41715 & n21586 ;
  assign n41716 = ~n21587 ;
  assign n21588 = n175 & n41716 ;
  assign n20750 = n20716 | n20734 ;
  assign n41717 = ~n20750 ;
  assign n21076 = n41717 & n141 ;
  assign n21077 = n20174 | n21076 ;
  assign n41718 = ~n20716 ;
  assign n20722 = n20174 & n41718 ;
  assign n20723 = n41306 & n20722 ;
  assign n21139 = n20723 & n141 ;
  assign n41719 = ~n21139 ;
  assign n21140 = n21077 & n41719 ;
  assign n21569 = n2753 | n21568 ;
  assign n41720 = ~n21569 ;
  assign n21589 = n41720 & n21586 ;
  assign n21590 = n21140 | n21589 ;
  assign n41721 = ~n21588 ;
  assign n21591 = n41721 & n21590 ;
  assign n41722 = ~n21591 ;
  assign n21592 = n2431 & n41722 ;
  assign n20749 = n20719 | n20736 ;
  assign n41723 = ~n20749 ;
  assign n21141 = n41723 & n141 ;
  assign n21142 = n20211 | n21141 ;
  assign n20721 = n20211 & n41316 ;
  assign n41724 = ~n20736 ;
  assign n20748 = n20721 & n41724 ;
  assign n21143 = n20748 & n141 ;
  assign n41725 = ~n21143 ;
  assign n21144 = n21142 & n41725 ;
  assign n21600 = n41704 & n21581 ;
  assign n21601 = n21138 | n21600 ;
  assign n41726 = ~n21583 ;
  assign n21602 = n41726 & n21601 ;
  assign n41727 = ~n21602 ;
  assign n21603 = n174 & n41727 ;
  assign n21604 = n41714 & n21601 ;
  assign n21605 = n21113 | n21604 ;
  assign n41728 = ~n21603 ;
  assign n21606 = n41728 & n21605 ;
  assign n41729 = ~n21606 ;
  assign n21607 = n2753 & n41729 ;
  assign n21608 = n2431 | n21607 ;
  assign n41730 = ~n21608 ;
  assign n21609 = n21590 & n41730 ;
  assign n21610 = n21144 | n21609 ;
  assign n41731 = ~n21592 ;
  assign n21611 = n41731 & n21610 ;
  assign n41732 = ~n21611 ;
  assign n21612 = n177 & n41732 ;
  assign n20774 = n20740 | n20758 ;
  assign n41733 = ~n20774 ;
  assign n21145 = n41733 & n141 ;
  assign n21146 = n20298 | n21145 ;
  assign n41734 = ~n20740 ;
  assign n20741 = n20298 & n41734 ;
  assign n20742 = n41322 & n20741 ;
  assign n21147 = n20742 & n141 ;
  assign n41735 = ~n21147 ;
  assign n21148 = n21146 & n41735 ;
  assign n21593 = n177 | n21592 ;
  assign n41736 = ~n21593 ;
  assign n21613 = n41736 & n21610 ;
  assign n21614 = n21148 | n21613 ;
  assign n41737 = ~n21612 ;
  assign n21615 = n41737 & n21614 ;
  assign n41738 = ~n21615 ;
  assign n21616 = n178 & n41738 ;
  assign n20773 = n20745 | n20760 ;
  assign n41739 = ~n20773 ;
  assign n21149 = n41739 & n141 ;
  assign n21150 = n20304 | n21149 ;
  assign n20747 = n20304 & n41332 ;
  assign n41740 = ~n20760 ;
  assign n20772 = n20747 & n41740 ;
  assign n21151 = n20772 & n141 ;
  assign n41741 = ~n21151 ;
  assign n21152 = n21150 & n41741 ;
  assign n21624 = n41720 & n21605 ;
  assign n21625 = n21140 | n21624 ;
  assign n41742 = ~n21607 ;
  assign n21626 = n41742 & n21625 ;
  assign n41743 = ~n21626 ;
  assign n21627 = n176 & n41743 ;
  assign n21628 = n41730 & n21625 ;
  assign n21629 = n21144 | n21628 ;
  assign n41744 = ~n21627 ;
  assign n21630 = n41744 & n21629 ;
  assign n41745 = ~n21630 ;
  assign n21631 = n177 & n41745 ;
  assign n21632 = n178 | n21631 ;
  assign n41746 = ~n21632 ;
  assign n21633 = n21614 & n41746 ;
  assign n21634 = n21152 | n21633 ;
  assign n41747 = ~n21616 ;
  assign n21635 = n41747 & n21634 ;
  assign n41748 = ~n21635 ;
  assign n21636 = n179 & n41748 ;
  assign n20798 = n20764 | n20782 ;
  assign n41749 = ~n20798 ;
  assign n21135 = n41749 & n141 ;
  assign n21136 = n20312 | n21135 ;
  assign n41750 = ~n20764 ;
  assign n20765 = n20312 & n41750 ;
  assign n20766 = n41338 & n20765 ;
  assign n21154 = n20766 & n141 ;
  assign n41751 = ~n21154 ;
  assign n21155 = n21136 & n41751 ;
  assign n21617 = n1707 | n21616 ;
  assign n41752 = ~n21617 ;
  assign n21637 = n41752 & n21634 ;
  assign n21638 = n21155 | n21637 ;
  assign n41753 = ~n21636 ;
  assign n21639 = n41753 & n21638 ;
  assign n41754 = ~n21639 ;
  assign n21640 = n1487 & n41754 ;
  assign n20771 = n20314 & n41348 ;
  assign n41755 = ~n20784 ;
  assign n20796 = n20771 & n41755 ;
  assign n21156 = n20796 & n141 ;
  assign n20797 = n20769 | n20784 ;
  assign n41756 = ~n20797 ;
  assign n21158 = n41756 & n141 ;
  assign n21159 = n20314 | n21158 ;
  assign n41757 = ~n21156 ;
  assign n21160 = n41757 & n21159 ;
  assign n21648 = n41736 & n21629 ;
  assign n21649 = n21148 | n21648 ;
  assign n41758 = ~n21631 ;
  assign n21650 = n41758 & n21649 ;
  assign n41759 = ~n21650 ;
  assign n21651 = n178 & n41759 ;
  assign n21652 = n41746 & n21649 ;
  assign n21653 = n21152 | n21652 ;
  assign n41760 = ~n21651 ;
  assign n21654 = n41760 & n21653 ;
  assign n41761 = ~n21654 ;
  assign n21655 = n1707 & n41761 ;
  assign n21656 = n1487 | n21655 ;
  assign n41762 = ~n21656 ;
  assign n21657 = n21638 & n41762 ;
  assign n21658 = n21160 | n21657 ;
  assign n41763 = ~n21640 ;
  assign n21659 = n41763 & n21658 ;
  assign n41764 = ~n21659 ;
  assign n21660 = n181 & n41764 ;
  assign n20822 = n20788 | n20806 ;
  assign n41765 = ~n20822 ;
  assign n21161 = n41765 & n141 ;
  assign n21162 = n20318 | n21161 ;
  assign n41766 = ~n20788 ;
  assign n20794 = n20318 & n41766 ;
  assign n20795 = n41354 & n20794 ;
  assign n21163 = n20795 & n141 ;
  assign n41767 = ~n21163 ;
  assign n21164 = n21162 & n41767 ;
  assign n21641 = n181 | n21640 ;
  assign n41768 = ~n21641 ;
  assign n21661 = n41768 & n21658 ;
  assign n21662 = n21164 | n21661 ;
  assign n41769 = ~n21660 ;
  assign n21663 = n41769 & n21662 ;
  assign n41770 = ~n21663 ;
  assign n21664 = n182 & n41770 ;
  assign n20820 = n20791 | n20808 ;
  assign n41771 = ~n20820 ;
  assign n21024 = n41771 & n141 ;
  assign n21025 = n20322 | n21024 ;
  assign n20793 = n20322 & n41364 ;
  assign n41772 = ~n20808 ;
  assign n20821 = n20793 & n41772 ;
  assign n21165 = n20821 & n141 ;
  assign n41773 = ~n21165 ;
  assign n21166 = n21025 & n41773 ;
  assign n21670 = n41752 & n21653 ;
  assign n21671 = n21155 | n21670 ;
  assign n41774 = ~n21655 ;
  assign n21672 = n41774 & n21671 ;
  assign n41775 = ~n21672 ;
  assign n21673 = n180 & n41775 ;
  assign n21674 = n41762 & n21671 ;
  assign n21675 = n21160 | n21674 ;
  assign n41776 = ~n21673 ;
  assign n21676 = n41776 & n21675 ;
  assign n41777 = ~n21676 ;
  assign n21677 = n181 & n41777 ;
  assign n21678 = n182 | n21677 ;
  assign n41778 = ~n21678 ;
  assign n21679 = n21662 & n41778 ;
  assign n21680 = n21166 | n21679 ;
  assign n41779 = ~n21664 ;
  assign n21681 = n41779 & n21680 ;
  assign n41780 = ~n21681 ;
  assign n21682 = n183 & n41780 ;
  assign n41781 = ~n20812 ;
  assign n20813 = n20325 & n41781 ;
  assign n20814 = n41370 & n20813 ;
  assign n21153 = n20814 & n141 ;
  assign n20846 = n20812 | n20830 ;
  assign n41782 = ~n20846 ;
  assign n21167 = n41782 & n141 ;
  assign n21168 = n20325 | n21167 ;
  assign n41783 = ~n21153 ;
  assign n21169 = n41783 & n21168 ;
  assign n21666 = n183 | n21664 ;
  assign n41784 = ~n21666 ;
  assign n21683 = n41784 & n21680 ;
  assign n21684 = n21169 | n21683 ;
  assign n41785 = ~n21682 ;
  assign n21685 = n41785 & n21684 ;
  assign n41786 = ~n21685 ;
  assign n21686 = n838 & n41786 ;
  assign n20845 = n20817 | n20832 ;
  assign n41787 = ~n20845 ;
  assign n21170 = n41787 & n141 ;
  assign n21171 = n20236 | n21170 ;
  assign n20819 = n20236 & n41380 ;
  assign n41788 = ~n20832 ;
  assign n20844 = n20819 & n41788 ;
  assign n21173 = n20844 & n141 ;
  assign n41789 = ~n21173 ;
  assign n21174 = n21171 & n41789 ;
  assign n21696 = n41768 & n21675 ;
  assign n21697 = n21164 | n21696 ;
  assign n41790 = ~n21677 ;
  assign n21698 = n41790 & n21697 ;
  assign n41791 = ~n21698 ;
  assign n21699 = n182 & n41791 ;
  assign n21700 = n41778 & n21697 ;
  assign n21701 = n21166 | n21700 ;
  assign n41792 = ~n21699 ;
  assign n21702 = n41792 & n21701 ;
  assign n41793 = ~n21702 ;
  assign n21703 = n996 & n41793 ;
  assign n21704 = n838 | n21703 ;
  assign n41794 = ~n21704 ;
  assign n21705 = n21684 & n41794 ;
  assign n21706 = n21174 | n21705 ;
  assign n41795 = ~n21686 ;
  assign n21707 = n41795 & n21706 ;
  assign n41796 = ~n21707 ;
  assign n21708 = n185 & n41796 ;
  assign n20863 = n20836 | n20854 ;
  assign n41797 = ~n20863 ;
  assign n21125 = n41797 & n141 ;
  assign n21126 = n20307 | n21125 ;
  assign n41798 = ~n20836 ;
  assign n20837 = n20307 & n41798 ;
  assign n20838 = n41386 & n20837 ;
  assign n21175 = n20838 & n141 ;
  assign n41799 = ~n21175 ;
  assign n21176 = n21126 & n41799 ;
  assign n21687 = n185 | n21686 ;
  assign n41800 = ~n21687 ;
  assign n21709 = n41800 & n21706 ;
  assign n21710 = n21176 | n21709 ;
  assign n41801 = ~n21708 ;
  assign n21711 = n41801 & n21710 ;
  assign n41802 = ~n21711 ;
  assign n21712 = n186 & n41802 ;
  assign n20862 = n20841 | n20856 ;
  assign n41803 = ~n20862 ;
  assign n21114 = n41803 & n141 ;
  assign n21115 = n20327 | n21114 ;
  assign n20843 = n20327 & n41396 ;
  assign n41804 = ~n20856 ;
  assign n20861 = n20843 & n41804 ;
  assign n21177 = n20861 & n141 ;
  assign n41805 = ~n21177 ;
  assign n21178 = n21115 & n41805 ;
  assign n21720 = n41784 & n21701 ;
  assign n21721 = n21169 | n21720 ;
  assign n41806 = ~n21703 ;
  assign n21722 = n41806 & n21721 ;
  assign n41807 = ~n21722 ;
  assign n21723 = n184 & n41807 ;
  assign n21724 = n41794 & n21721 ;
  assign n21725 = n21174 | n21724 ;
  assign n41808 = ~n21723 ;
  assign n21726 = n41808 & n21725 ;
  assign n41809 = ~n21726 ;
  assign n21727 = n185 & n41809 ;
  assign n21728 = n186 | n21727 ;
  assign n41810 = ~n21728 ;
  assign n21729 = n21710 & n41810 ;
  assign n21730 = n21178 | n21729 ;
  assign n41811 = ~n21712 ;
  assign n21731 = n41811 & n21730 ;
  assign n41812 = ~n21731 ;
  assign n21732 = n187 & n41812 ;
  assign n21713 = n528 | n21712 ;
  assign n41813 = ~n21713 ;
  assign n21733 = n41813 & n21730 ;
  assign n41814 = ~n20860 ;
  assign n20948 = n41814 & n20928 ;
  assign n20949 = n41402 & n20948 ;
  assign n21157 = n20949 & n141 ;
  assign n20873 = n20860 | n20871 ;
  assign n41815 = ~n20873 ;
  assign n21179 = n41815 & n141 ;
  assign n21765 = n20928 | n21179 ;
  assign n41816 = ~n21157 ;
  assign n21766 = n41816 & n21765 ;
  assign n21767 = n21733 | n21766 ;
  assign n41817 = ~n21732 ;
  assign n21768 = n41817 & n21767 ;
  assign n41818 = ~n21768 ;
  assign n21769 = n413 & n41818 ;
  assign n20933 = n20926 & n41412 ;
  assign n41819 = ~n20934 ;
  assign n20946 = n20933 & n41819 ;
  assign n21172 = n20946 & n141 ;
  assign n20947 = n20931 | n20934 ;
  assign n41820 = ~n20947 ;
  assign n21180 = n41820 & n141 ;
  assign n21181 = n20926 | n21180 ;
  assign n41821 = ~n21172 ;
  assign n21182 = n41821 & n21181 ;
  assign n21737 = n41800 & n21725 ;
  assign n21738 = n21176 | n21737 ;
  assign n41822 = ~n21727 ;
  assign n21739 = n41822 & n21738 ;
  assign n41823 = ~n21739 ;
  assign n21740 = n186 & n41823 ;
  assign n21741 = n41810 & n21738 ;
  assign n21742 = n21178 | n21741 ;
  assign n41824 = ~n21740 ;
  assign n21743 = n41824 & n21742 ;
  assign n41825 = ~n21743 ;
  assign n21744 = n528 & n41825 ;
  assign n21745 = n413 | n21744 ;
  assign n41826 = ~n21745 ;
  assign n21772 = n41826 & n21767 ;
  assign n21773 = n21182 | n21772 ;
  assign n41827 = ~n21769 ;
  assign n21774 = n41827 & n21773 ;
  assign n41828 = ~n21774 ;
  assign n21775 = n189 & n41828 ;
  assign n20972 = n20938 | n20956 ;
  assign n41829 = ~n20972 ;
  assign n21121 = n41829 & n141 ;
  assign n21122 = n20920 | n21121 ;
  assign n41830 = ~n20938 ;
  assign n20944 = n20920 & n41830 ;
  assign n20945 = n41418 & n20944 ;
  assign n21183 = n20945 & n141 ;
  assign n41831 = ~n21183 ;
  assign n21184 = n21122 & n41831 ;
  assign n21771 = n189 | n21769 ;
  assign n41832 = ~n21771 ;
  assign n21776 = n41832 & n21773 ;
  assign n21777 = n21184 | n21776 ;
  assign n41833 = ~n21775 ;
  assign n21778 = n41833 & n21777 ;
  assign n41834 = ~n21778 ;
  assign n21779 = n190 & n41834 ;
  assign n21781 = n287 | n21779 ;
  assign n20971 = n20941 | n20958 ;
  assign n41835 = ~n20971 ;
  assign n21048 = n41835 & n141 ;
  assign n21049 = n20913 | n21048 ;
  assign n20943 = n20913 & n41428 ;
  assign n41836 = ~n20958 ;
  assign n20970 = n20943 & n41836 ;
  assign n21054 = n20970 & n141 ;
  assign n41837 = ~n21054 ;
  assign n21055 = n21049 & n41837 ;
  assign n21746 = n41813 & n21742 ;
  assign n21787 = n21746 | n21766 ;
  assign n41838 = ~n21744 ;
  assign n21788 = n41838 & n21787 ;
  assign n41839 = ~n21788 ;
  assign n21789 = n188 & n41839 ;
  assign n21790 = n41826 & n21787 ;
  assign n21791 = n21182 | n21790 ;
  assign n41840 = ~n21789 ;
  assign n21792 = n41840 & n21791 ;
  assign n41841 = ~n21792 ;
  assign n21793 = n189 & n41841 ;
  assign n21794 = n190 | n21793 ;
  assign n41842 = ~n21794 ;
  assign n21795 = n21777 & n41842 ;
  assign n21796 = n21055 | n21795 ;
  assign n41843 = ~n21781 ;
  assign n21797 = n41843 & n21796 ;
  assign n21798 = n21764 | n21797 ;
  assign n20987 = n20965 | n20982 ;
  assign n41844 = ~n20987 ;
  assign n21026 = n41844 & n141 ;
  assign n21027 = n20900 | n21026 ;
  assign n20966 = n20900 & n41436 ;
  assign n41845 = ~n20982 ;
  assign n20986 = n20966 & n41845 ;
  assign n21129 = n20986 & n141 ;
  assign n41846 = ~n21129 ;
  assign n21130 = n21027 & n41846 ;
  assign n41847 = ~n21779 ;
  assign n21801 = n41847 & n21796 ;
  assign n41848 = ~n21801 ;
  assign n21802 = n191 & n41848 ;
  assign n41849 = ~n21802 ;
  assign n21803 = n21130 & n41849 ;
  assign n21804 = n21798 & n21803 ;
  assign n21805 = n21751 | n21804 ;
  assign n41850 = ~n21208 ;
  assign n21209 = n141 & n41850 ;
  assign n21747 = n20984 | n21209 ;
  assign n21748 = n21130 | n21747 ;
  assign n21809 = n21798 & n41849 ;
  assign n22028 = n21748 | n21809 ;
  assign n22029 = n31336 & n22028 ;
  assign n22030 = n21805 | n22029 ;
  assign n21810 = n21130 | n21809 ;
  assign n21780 = n191 | n21779 ;
  assign n41851 = ~n21780 ;
  assign n21812 = n41851 & n21796 ;
  assign n21813 = n21764 | n21812 ;
  assign n21814 = n41849 & n21813 ;
  assign n21815 = n21748 | n21814 ;
  assign n21816 = n31336 & n21815 ;
  assign n21822 = n21803 & n21813 ;
  assign n21823 = n21751 | n21822 ;
  assign n140 = n21816 | n21823 ;
  assign n41852 = ~n21810 ;
  assign n22012 = n41852 & n140 ;
  assign n22013 = n21804 | n22012 ;
  assign n41853 = ~n21812 ;
  assign n22604 = n21764 & n41853 ;
  assign n22605 = n41849 & n22604 ;
  assign n22606 = n140 & n22605 ;
  assign n22608 = n21802 | n21812 ;
  assign n41854 = ~n22608 ;
  assign n22609 = n140 & n41854 ;
  assign n22610 = n21764 | n22609 ;
  assign n41855 = ~n22606 ;
  assign n22611 = n41855 & n22610 ;
  assign n22612 = n22013 | n22611 ;
  assign n41856 = ~n21750 ;
  assign n21752 = n141 & n41856 ;
  assign n41857 = ~n21211 ;
  assign n21753 = n41857 & n21752 ;
  assign n41858 = ~n21804 ;
  assign n21806 = n21753 & n41858 ;
  assign n41859 = ~n21816 ;
  assign n21817 = n21806 & n41859 ;
  assign n21818 = x24 | n21817 ;
  assign n41860 = ~n236 ;
  assign n21917 = n41860 & n140 ;
  assign n21918 = n21818 | n21917 ;
  assign n21919 = n21817 | n21917 ;
  assign n21920 = x24 & n21919 ;
  assign n41861 = ~n21920 ;
  assign n21921 = n21918 & n41861 ;
  assign n239 = x20 | x21 ;
  assign n240 = x22 | n239 ;
  assign n21901 = x22 & n140 ;
  assign n41862 = ~n21901 ;
  assign n21922 = n240 & n41862 ;
  assign n41863 = ~n21922 ;
  assign n21923 = n141 & n41863 ;
  assign n21924 = n142 | n21923 ;
  assign n20881 = n240 & n41467 ;
  assign n20882 = n41451 & n20881 ;
  assign n21759 = n20882 & n41452 ;
  assign n21760 = n41453 & n21759 ;
  assign n21902 = n21760 & n41862 ;
  assign n41864 = ~x22 ;
  assign n21939 = n41864 & n140 ;
  assign n41865 = ~n21939 ;
  assign n21940 = x23 & n41865 ;
  assign n21941 = n21917 | n21940 ;
  assign n21942 = n21902 | n21941 ;
  assign n41866 = ~n21924 ;
  assign n21943 = n41866 & n21942 ;
  assign n21944 = n21921 | n21943 ;
  assign n241 = n41864 & n239 ;
  assign n41867 = ~n22030 ;
  assign n22037 = x22 & n41867 ;
  assign n22038 = n241 | n22037 ;
  assign n41868 = ~n22038 ;
  assign n22039 = n141 & n41868 ;
  assign n41869 = ~n22039 ;
  assign n22040 = n21942 & n41869 ;
  assign n41870 = ~n22040 ;
  assign n22041 = n142 & n41870 ;
  assign n41871 = ~n22041 ;
  assign n22042 = n21944 & n41871 ;
  assign n41872 = ~n22042 ;
  assign n22061 = n143 & n41872 ;
  assign n21091 = n21066 | n21089 ;
  assign n41873 = ~n21091 ;
  assign n21204 = n41873 & n21198 ;
  assign n21952 = n21204 & n140 ;
  assign n21971 = n41873 & n140 ;
  assign n21972 = n21198 | n21971 ;
  assign n41874 = ~n21952 ;
  assign n21973 = n41874 & n21972 ;
  assign n22065 = n143 | n22041 ;
  assign n41875 = ~n22065 ;
  assign n22066 = n21944 & n41875 ;
  assign n22067 = n21973 | n22066 ;
  assign n41876 = ~n22061 ;
  assign n22068 = n41876 & n22067 ;
  assign n41877 = ~n22068 ;
  assign n22069 = n144 & n41877 ;
  assign n41878 = ~n21205 ;
  assign n21239 = n41878 & n21218 ;
  assign n21240 = n41486 & n21239 ;
  assign n21908 = n21240 & n140 ;
  assign n21206 = n21203 | n21205 ;
  assign n41879 = ~n21206 ;
  assign n21911 = n41879 & n140 ;
  assign n21912 = n21218 | n21911 ;
  assign n41880 = ~n21908 ;
  assign n21913 = n41880 & n21912 ;
  assign n22043 = n19362 & n41872 ;
  assign n22047 = n18797 | n22043 ;
  assign n41881 = ~n22047 ;
  assign n22070 = n41881 & n22067 ;
  assign n22071 = n21913 | n22070 ;
  assign n41882 = ~n22069 ;
  assign n22072 = n41882 & n22071 ;
  assign n41883 = ~n22072 ;
  assign n22073 = n145 & n41883 ;
  assign n21223 = n21087 & n41474 ;
  assign n41884 = ~n21224 ;
  assign n21237 = n21223 & n41884 ;
  assign n21895 = n21237 & n140 ;
  assign n21238 = n21221 | n21224 ;
  assign n41885 = ~n21238 ;
  assign n21959 = n41885 & n140 ;
  assign n21960 = n21087 | n21959 ;
  assign n41886 = ~n21895 ;
  assign n21961 = n41886 & n21960 ;
  assign n41887 = ~n21923 ;
  assign n21946 = n41887 & n21942 ;
  assign n41888 = ~n21946 ;
  assign n21947 = n142 & n41888 ;
  assign n21948 = n19362 | n21947 ;
  assign n41889 = ~n21948 ;
  assign n21949 = n21944 & n41889 ;
  assign n21974 = n21949 | n21973 ;
  assign n41890 = ~n22043 ;
  assign n22044 = n21974 & n41890 ;
  assign n41891 = ~n22044 ;
  assign n22045 = n18797 & n41891 ;
  assign n22046 = n145 | n22045 ;
  assign n41892 = ~n22046 ;
  assign n22090 = n41892 & n22071 ;
  assign n22091 = n21961 | n22090 ;
  assign n41893 = ~n22073 ;
  assign n22092 = n41893 & n22091 ;
  assign n41894 = ~n22092 ;
  assign n22093 = n146 & n41894 ;
  assign n21236 = n21227 | n21228 ;
  assign n41895 = ~n21236 ;
  assign n21879 = n41895 & n140 ;
  assign n21880 = n21193 | n21879 ;
  assign n41896 = ~n21228 ;
  assign n21234 = n21193 & n41896 ;
  assign n21235 = n41480 & n21234 ;
  assign n21889 = n21235 & n140 ;
  assign n41897 = ~n21889 ;
  assign n21890 = n21880 & n41897 ;
  assign n22074 = n146 | n22073 ;
  assign n41898 = ~n22074 ;
  assign n22094 = n41898 & n22091 ;
  assign n22095 = n21890 | n22094 ;
  assign n41899 = ~n22093 ;
  assign n22096 = n41899 & n22095 ;
  assign n41900 = ~n22096 ;
  assign n22097 = n16322 & n41900 ;
  assign n21263 = n21231 | n21249 ;
  assign n41901 = ~n21263 ;
  assign n21896 = n41901 & n140 ;
  assign n21897 = n21195 | n21896 ;
  assign n21233 = n21195 & n41491 ;
  assign n41902 = ~n21249 ;
  assign n21262 = n21233 & n41902 ;
  assign n21934 = n21262 & n140 ;
  assign n41903 = ~n21934 ;
  assign n21935 = n21897 & n41903 ;
  assign n22048 = n21974 & n41881 ;
  assign n22049 = n21913 | n22048 ;
  assign n41904 = ~n22045 ;
  assign n22050 = n41904 & n22049 ;
  assign n41905 = ~n22050 ;
  assign n22051 = n145 & n41905 ;
  assign n22052 = n41892 & n22049 ;
  assign n22053 = n21961 | n22052 ;
  assign n41906 = ~n22051 ;
  assign n22054 = n41906 & n22053 ;
  assign n41907 = ~n22054 ;
  assign n22055 = n146 & n41907 ;
  assign n22056 = n147 | n22055 ;
  assign n41908 = ~n22056 ;
  assign n22113 = n41908 & n22095 ;
  assign n22114 = n21935 | n22113 ;
  assign n41909 = ~n22097 ;
  assign n22115 = n41909 & n22114 ;
  assign n41910 = ~n22115 ;
  assign n22116 = n148 & n41910 ;
  assign n41911 = ~n21253 ;
  assign n21259 = n21063 & n41911 ;
  assign n21260 = n41497 & n21259 ;
  assign n21955 = n21260 & n140 ;
  assign n21261 = n21252 | n21253 ;
  assign n41912 = ~n21261 ;
  assign n21956 = n41912 & n140 ;
  assign n21957 = n21063 | n21956 ;
  assign n41913 = ~n21955 ;
  assign n21958 = n41913 & n21957 ;
  assign n22098 = n148 | n22097 ;
  assign n41914 = ~n22098 ;
  assign n22117 = n41914 & n22114 ;
  assign n22118 = n21958 | n22117 ;
  assign n41915 = ~n22116 ;
  assign n22119 = n41915 & n22118 ;
  assign n41916 = ~n22119 ;
  assign n22120 = n149 & n41916 ;
  assign n21258 = n21099 & n41507 ;
  assign n41917 = ~n21273 ;
  assign n21286 = n21258 & n41917 ;
  assign n21881 = n21286 & n140 ;
  assign n21287 = n21256 | n21273 ;
  assign n41918 = ~n21287 ;
  assign n21903 = n41918 & n140 ;
  assign n21904 = n21099 | n21903 ;
  assign n41919 = ~n21881 ;
  assign n21905 = n41919 & n21904 ;
  assign n22075 = n22053 & n41898 ;
  assign n22076 = n21890 | n22075 ;
  assign n41920 = ~n22055 ;
  assign n22077 = n41920 & n22076 ;
  assign n41921 = ~n22077 ;
  assign n22078 = n147 & n41921 ;
  assign n22079 = n41908 & n22076 ;
  assign n22080 = n21935 | n22079 ;
  assign n41922 = ~n22078 ;
  assign n22081 = n41922 & n22080 ;
  assign n41923 = ~n22081 ;
  assign n22082 = n15807 & n41923 ;
  assign n22083 = n149 | n22082 ;
  assign n41924 = ~n22083 ;
  assign n22134 = n41924 & n22118 ;
  assign n22135 = n21905 | n22134 ;
  assign n41925 = ~n22120 ;
  assign n22136 = n41925 & n22135 ;
  assign n41926 = ~n22136 ;
  assign n22137 = n150 & n41926 ;
  assign n21285 = n21276 | n21277 ;
  assign n41927 = ~n21285 ;
  assign n21932 = n41927 & n140 ;
  assign n21933 = n21093 | n21932 ;
  assign n41928 = ~n21277 ;
  assign n21283 = n21093 & n41928 ;
  assign n21284 = n41513 & n21283 ;
  assign n21966 = n21284 & n140 ;
  assign n41929 = ~n21966 ;
  assign n21967 = n21933 & n41929 ;
  assign n22121 = n150 | n22120 ;
  assign n41930 = ~n22121 ;
  assign n22138 = n41930 & n22135 ;
  assign n22139 = n21967 | n22138 ;
  assign n41931 = ~n22137 ;
  assign n22140 = n41931 & n22139 ;
  assign n41932 = ~n22140 ;
  assign n22141 = n13662 & n41932 ;
  assign n22099 = n22080 & n41914 ;
  assign n22100 = n21958 | n22099 ;
  assign n41933 = ~n22082 ;
  assign n22101 = n41933 & n22100 ;
  assign n41934 = ~n22101 ;
  assign n22102 = n149 & n41934 ;
  assign n22103 = n41924 & n22100 ;
  assign n22104 = n21905 | n22103 ;
  assign n41935 = ~n22102 ;
  assign n22105 = n41935 & n22104 ;
  assign n41936 = ~n22105 ;
  assign n22106 = n150 & n41936 ;
  assign n22107 = n151 | n22106 ;
  assign n41937 = ~n22107 ;
  assign n22143 = n41937 & n22139 ;
  assign n21311 = n21280 | n21297 ;
  assign n41938 = ~n21311 ;
  assign n21930 = n41938 & n140 ;
  assign n21931 = n21081 | n21930 ;
  assign n21282 = n21081 & n41523 ;
  assign n41939 = ~n21297 ;
  assign n21310 = n21282 & n41939 ;
  assign n22150 = n21310 & n22030 ;
  assign n41940 = ~n22150 ;
  assign n22151 = n21931 & n41940 ;
  assign n22152 = n22143 | n22151 ;
  assign n41941 = ~n22141 ;
  assign n22153 = n41941 & n22152 ;
  assign n41942 = ~n22153 ;
  assign n22154 = n152 & n41942 ;
  assign n41943 = ~n21301 ;
  assign n21307 = n21105 & n41943 ;
  assign n21308 = n41529 & n21307 ;
  assign n21891 = n21308 & n140 ;
  assign n21309 = n21300 | n21301 ;
  assign n41944 = ~n21309 ;
  assign n21936 = n41944 & n140 ;
  assign n21937 = n21105 | n21936 ;
  assign n41945 = ~n21891 ;
  assign n21938 = n41945 & n21937 ;
  assign n22142 = n152 | n22141 ;
  assign n41946 = ~n22142 ;
  assign n22155 = n41946 & n22152 ;
  assign n22156 = n21938 | n22155 ;
  assign n41947 = ~n22154 ;
  assign n22157 = n41947 & n22156 ;
  assign n41948 = ~n22157 ;
  assign n22158 = n153 & n41948 ;
  assign n21335 = n21304 | n21321 ;
  assign n41949 = ~n21335 ;
  assign n21875 = n41949 & n140 ;
  assign n21876 = n21075 | n21875 ;
  assign n21306 = n21075 & n41539 ;
  assign n41950 = ~n21321 ;
  assign n21334 = n21306 & n41950 ;
  assign n21882 = n21334 & n140 ;
  assign n41951 = ~n21882 ;
  assign n21883 = n21876 & n41951 ;
  assign n22122 = n22104 & n41930 ;
  assign n22123 = n21967 | n22122 ;
  assign n41952 = ~n22106 ;
  assign n22124 = n41952 & n22123 ;
  assign n41953 = ~n22124 ;
  assign n22125 = n151 & n41953 ;
  assign n22126 = n41937 & n22123 ;
  assign n22161 = n22126 | n22151 ;
  assign n41954 = ~n22125 ;
  assign n22162 = n41954 & n22161 ;
  assign n41955 = ~n22162 ;
  assign n22163 = n13079 & n41955 ;
  assign n22164 = n153 | n22163 ;
  assign n41956 = ~n22164 ;
  assign n22165 = n22156 & n41956 ;
  assign n22166 = n21883 | n22165 ;
  assign n41957 = ~n22158 ;
  assign n22167 = n41957 & n22166 ;
  assign n41958 = ~n22167 ;
  assign n22168 = n154 & n41958 ;
  assign n22159 = n154 | n22158 ;
  assign n41959 = ~n22159 ;
  assign n22169 = n41959 & n22166 ;
  assign n21333 = n21324 | n21325 ;
  assign n41960 = ~n21333 ;
  assign n21976 = n41960 & n140 ;
  assign n21977 = n21110 | n21976 ;
  assign n41961 = ~n21325 ;
  assign n21331 = n21110 & n41961 ;
  assign n21332 = n41545 & n21331 ;
  assign n22188 = n21332 & n22030 ;
  assign n41962 = ~n22188 ;
  assign n22189 = n21977 & n41962 ;
  assign n22200 = n22169 | n22189 ;
  assign n41963 = ~n22168 ;
  assign n22201 = n41963 & n22200 ;
  assign n41964 = ~n22201 ;
  assign n22202 = n11067 & n41964 ;
  assign n21359 = n21328 | n21345 ;
  assign n41965 = ~n21359 ;
  assign n21885 = n41965 & n140 ;
  assign n21886 = n21124 | n21885 ;
  assign n21330 = n21124 & n41555 ;
  assign n41966 = ~n21345 ;
  assign n21358 = n21330 & n41966 ;
  assign n22146 = n21358 & n22030 ;
  assign n41967 = ~n22146 ;
  assign n22147 = n21886 & n41967 ;
  assign n22170 = n41946 & n22161 ;
  assign n22171 = n21938 | n22170 ;
  assign n41968 = ~n22163 ;
  assign n22172 = n41968 & n22171 ;
  assign n41969 = ~n22172 ;
  assign n22173 = n153 & n41969 ;
  assign n22174 = n41956 & n22171 ;
  assign n22175 = n21883 | n22174 ;
  assign n41970 = ~n22173 ;
  assign n22176 = n41970 & n22175 ;
  assign n41971 = ~n22176 ;
  assign n22177 = n154 & n41971 ;
  assign n22178 = n11067 | n22177 ;
  assign n41972 = ~n22178 ;
  assign n22219 = n41972 & n22200 ;
  assign n22220 = n22147 | n22219 ;
  assign n41973 = ~n22202 ;
  assign n22221 = n41973 & n22220 ;
  assign n41974 = ~n22221 ;
  assign n22222 = n156 & n41974 ;
  assign n21357 = n21348 | n21349 ;
  assign n41975 = ~n21357 ;
  assign n21877 = n41975 & n140 ;
  assign n21878 = n21128 | n21877 ;
  assign n41976 = ~n21349 ;
  assign n21355 = n21128 & n41976 ;
  assign n21356 = n41561 & n21355 ;
  assign n21981 = n21356 & n140 ;
  assign n41977 = ~n21981 ;
  assign n21982 = n21878 & n41977 ;
  assign n22203 = n10657 | n22202 ;
  assign n41978 = ~n22203 ;
  assign n22223 = n41978 & n22220 ;
  assign n22224 = n21982 | n22223 ;
  assign n41979 = ~n22222 ;
  assign n22225 = n41979 & n22224 ;
  assign n41980 = ~n22225 ;
  assign n22226 = n157 & n41980 ;
  assign n21383 = n21352 | n21369 ;
  assign n41981 = ~n21383 ;
  assign n21871 = n41981 & n140 ;
  assign n21872 = n21097 | n21871 ;
  assign n21354 = n21097 & n41571 ;
  assign n41982 = ~n21369 ;
  assign n21382 = n21354 & n41982 ;
  assign n21914 = n21382 & n140 ;
  assign n41983 = ~n21914 ;
  assign n21915 = n21872 & n41983 ;
  assign n22179 = n41959 & n22175 ;
  assign n22192 = n22179 | n22189 ;
  assign n41984 = ~n22177 ;
  assign n22193 = n41984 & n22192 ;
  assign n41985 = ~n22193 ;
  assign n22194 = n155 & n41985 ;
  assign n22195 = n41972 & n22192 ;
  assign n22196 = n22147 | n22195 ;
  assign n41986 = ~n22194 ;
  assign n22197 = n41986 & n22196 ;
  assign n41987 = ~n22197 ;
  assign n22198 = n10657 & n41987 ;
  assign n22199 = n157 | n22198 ;
  assign n41988 = ~n22199 ;
  assign n22239 = n41988 & n22224 ;
  assign n22240 = n21915 | n22239 ;
  assign n41989 = ~n22226 ;
  assign n22241 = n41989 & n22240 ;
  assign n41990 = ~n22241 ;
  assign n22242 = n158 & n41990 ;
  assign n41991 = ~n21373 ;
  assign n21379 = n21072 & n41991 ;
  assign n21380 = n41577 & n21379 ;
  assign n21860 = n21380 & n140 ;
  assign n21381 = n21372 | n21373 ;
  assign n41992 = ~n21381 ;
  assign n21925 = n41992 & n140 ;
  assign n21926 = n21072 | n21925 ;
  assign n41993 = ~n21860 ;
  assign n21927 = n41993 & n21926 ;
  assign n22227 = n158 | n22226 ;
  assign n41994 = ~n22227 ;
  assign n22243 = n41994 & n22240 ;
  assign n22244 = n21927 | n22243 ;
  assign n41995 = ~n22242 ;
  assign n22245 = n41995 & n22244 ;
  assign n41996 = ~n22245 ;
  assign n22246 = n8857 & n41996 ;
  assign n22204 = n22196 & n41978 ;
  assign n22205 = n21982 | n22204 ;
  assign n41997 = ~n22198 ;
  assign n22206 = n41997 & n22205 ;
  assign n41998 = ~n22206 ;
  assign n22207 = n157 & n41998 ;
  assign n22208 = n41988 & n22205 ;
  assign n22209 = n21915 | n22208 ;
  assign n41999 = ~n22207 ;
  assign n22210 = n41999 & n22209 ;
  assign n42000 = ~n22210 ;
  assign n22211 = n158 & n42000 ;
  assign n22212 = n8857 | n22211 ;
  assign n42001 = ~n22212 ;
  assign n22249 = n42001 & n22244 ;
  assign n21407 = n21376 | n21393 ;
  assign n42002 = ~n21407 ;
  assign n21833 = n42002 & n140 ;
  assign n21834 = n21108 | n21833 ;
  assign n21378 = n21108 & n41587 ;
  assign n42003 = ~n21393 ;
  assign n21406 = n21378 & n42003 ;
  assign n22252 = n21406 & n22030 ;
  assign n42004 = ~n22252 ;
  assign n22253 = n21834 & n42004 ;
  assign n22256 = n22249 | n22253 ;
  assign n42005 = ~n22246 ;
  assign n22257 = n42005 & n22256 ;
  assign n42006 = ~n22257 ;
  assign n22258 = n160 & n42006 ;
  assign n21400 = n21396 | n21397 ;
  assign n42007 = ~n21400 ;
  assign n21867 = n42007 & n140 ;
  assign n21868 = n21052 | n21867 ;
  assign n42008 = ~n21397 ;
  assign n21398 = n21052 & n42008 ;
  assign n21399 = n41593 & n21398 ;
  assign n21873 = n21399 & n140 ;
  assign n42009 = ~n21873 ;
  assign n21874 = n21868 & n42009 ;
  assign n22247 = n160 | n22246 ;
  assign n42010 = ~n22247 ;
  assign n22259 = n42010 & n22256 ;
  assign n22260 = n21874 | n22259 ;
  assign n42011 = ~n22258 ;
  assign n22261 = n42011 & n22260 ;
  assign n42012 = ~n22261 ;
  assign n22262 = n161 & n42012 ;
  assign n21431 = n21403 | n21417 ;
  assign n42013 = ~n21431 ;
  assign n21854 = n42013 & n140 ;
  assign n21855 = n21030 | n21854 ;
  assign n21405 = n21030 & n41603 ;
  assign n42014 = ~n21417 ;
  assign n21430 = n21405 & n42014 ;
  assign n21863 = n21430 & n140 ;
  assign n42015 = ~n21863 ;
  assign n21864 = n21855 & n42015 ;
  assign n22228 = n22209 & n41994 ;
  assign n22229 = n21927 | n22228 ;
  assign n42016 = ~n22211 ;
  assign n22230 = n42016 & n22229 ;
  assign n42017 = ~n22230 ;
  assign n22231 = n159 & n42017 ;
  assign n22232 = n42001 & n22229 ;
  assign n22265 = n22232 | n22253 ;
  assign n42018 = ~n22231 ;
  assign n22266 = n42018 & n22265 ;
  assign n42019 = ~n22266 ;
  assign n22267 = n8534 & n42019 ;
  assign n22268 = n161 | n22267 ;
  assign n42020 = ~n22268 ;
  assign n22269 = n22260 & n42020 ;
  assign n22270 = n21864 | n22269 ;
  assign n42021 = ~n22262 ;
  assign n22271 = n42021 & n22270 ;
  assign n42022 = ~n22271 ;
  assign n22272 = n162 & n42022 ;
  assign n21429 = n21420 | n21421 ;
  assign n42023 = ~n21429 ;
  assign n21953 = n42023 & n140 ;
  assign n21954 = n21102 | n21953 ;
  assign n42024 = ~n21421 ;
  assign n21427 = n21102 & n42024 ;
  assign n21428 = n41609 & n21427 ;
  assign n22033 = n21428 & n22030 ;
  assign n42025 = ~n22033 ;
  assign n22034 = n21954 & n42025 ;
  assign n22263 = n162 | n22262 ;
  assign n42026 = ~n22263 ;
  assign n22273 = n42026 & n22270 ;
  assign n22274 = n22034 | n22273 ;
  assign n42027 = ~n22272 ;
  assign n22275 = n42027 & n22274 ;
  assign n42028 = ~n22275 ;
  assign n22276 = n6889 & n42028 ;
  assign n21455 = n21424 | n21441 ;
  assign n42029 = ~n21455 ;
  assign n21842 = n42029 & n140 ;
  assign n21843 = n21120 | n21842 ;
  assign n21426 = n21120 & n41619 ;
  assign n42030 = ~n21441 ;
  assign n21454 = n21426 & n42030 ;
  assign n21849 = n21454 & n140 ;
  assign n42031 = ~n21849 ;
  assign n21850 = n21843 & n42031 ;
  assign n22279 = n42010 & n22265 ;
  assign n22280 = n21874 | n22279 ;
  assign n42032 = ~n22267 ;
  assign n22281 = n42032 & n22280 ;
  assign n42033 = ~n22281 ;
  assign n22282 = n161 & n42033 ;
  assign n22283 = n42020 & n22280 ;
  assign n22284 = n21864 | n22283 ;
  assign n42034 = ~n22282 ;
  assign n22285 = n42034 & n22284 ;
  assign n42035 = ~n22285 ;
  assign n22286 = n162 & n42035 ;
  assign n22287 = n6889 | n22286 ;
  assign n42036 = ~n22287 ;
  assign n22288 = n22274 & n42036 ;
  assign n22289 = n21850 | n22288 ;
  assign n42037 = ~n22276 ;
  assign n22290 = n42037 & n22289 ;
  assign n42038 = ~n22290 ;
  assign n22291 = n164 & n42038 ;
  assign n42039 = ~n21445 ;
  assign n21451 = n21039 & n42039 ;
  assign n21452 = n41625 & n21451 ;
  assign n21884 = n21452 & n140 ;
  assign n21453 = n21444 | n21445 ;
  assign n42040 = ~n21453 ;
  assign n21978 = n42040 & n140 ;
  assign n21979 = n21039 | n21978 ;
  assign n42041 = ~n21884 ;
  assign n21980 = n42041 & n21979 ;
  assign n22277 = n6600 | n22276 ;
  assign n42042 = ~n22277 ;
  assign n22292 = n42042 & n22289 ;
  assign n22293 = n21980 | n22292 ;
  assign n42043 = ~n22291 ;
  assign n22294 = n42043 & n22293 ;
  assign n42044 = ~n22294 ;
  assign n22295 = n165 & n42044 ;
  assign n21479 = n21448 | n21465 ;
  assign n42045 = ~n21479 ;
  assign n21856 = n42045 & n140 ;
  assign n21857 = n21079 | n21856 ;
  assign n21450 = n21079 & n41635 ;
  assign n42046 = ~n21465 ;
  assign n21478 = n21450 & n42046 ;
  assign n21964 = n21478 & n140 ;
  assign n42047 = ~n21964 ;
  assign n21965 = n21857 & n42047 ;
  assign n22298 = n42026 & n22284 ;
  assign n22299 = n22034 | n22298 ;
  assign n42048 = ~n22286 ;
  assign n22300 = n42048 & n22299 ;
  assign n42049 = ~n22300 ;
  assign n22301 = n163 & n42049 ;
  assign n22302 = n42036 & n22299 ;
  assign n22303 = n21850 | n22302 ;
  assign n42050 = ~n22301 ;
  assign n22304 = n42050 & n22303 ;
  assign n42051 = ~n22304 ;
  assign n22305 = n6600 & n42051 ;
  assign n22306 = n165 | n22305 ;
  assign n42052 = ~n22306 ;
  assign n22307 = n22293 & n42052 ;
  assign n22308 = n21965 | n22307 ;
  assign n42053 = ~n22295 ;
  assign n22309 = n42053 & n22308 ;
  assign n42054 = ~n22309 ;
  assign n22310 = n166 & n42054 ;
  assign n42055 = ~n21469 ;
  assign n21475 = n21013 & n42055 ;
  assign n21476 = n41641 & n21475 ;
  assign n21841 = n21476 & n140 ;
  assign n21477 = n21468 | n21469 ;
  assign n42056 = ~n21477 ;
  assign n21968 = n42056 & n140 ;
  assign n21969 = n21013 | n21968 ;
  assign n42057 = ~n21841 ;
  assign n21970 = n42057 & n21969 ;
  assign n22296 = n166 | n22295 ;
  assign n42058 = ~n22296 ;
  assign n22311 = n42058 & n22308 ;
  assign n22312 = n21970 | n22311 ;
  assign n42059 = ~n22310 ;
  assign n22313 = n42059 & n22312 ;
  assign n42060 = ~n22313 ;
  assign n22314 = n5352 & n42060 ;
  assign n21503 = n21472 | n21489 ;
  assign n42061 = ~n21503 ;
  assign n21839 = n42061 & n140 ;
  assign n21840 = n21117 | n21839 ;
  assign n21474 = n21117 & n41651 ;
  assign n42062 = ~n21489 ;
  assign n21502 = n21474 & n42062 ;
  assign n22148 = n21502 & n22030 ;
  assign n42063 = ~n22148 ;
  assign n22149 = n21840 & n42063 ;
  assign n22317 = n42042 & n22303 ;
  assign n22318 = n21980 | n22317 ;
  assign n42064 = ~n22305 ;
  assign n22319 = n42064 & n22318 ;
  assign n42065 = ~n22319 ;
  assign n22320 = n165 & n42065 ;
  assign n22321 = n42052 & n22318 ;
  assign n22324 = n21965 | n22321 ;
  assign n42066 = ~n22320 ;
  assign n22325 = n42066 & n22324 ;
  assign n42067 = ~n22325 ;
  assign n22326 = n166 & n42067 ;
  assign n22327 = n5352 | n22326 ;
  assign n42068 = ~n22327 ;
  assign n22328 = n22312 & n42068 ;
  assign n22329 = n22149 | n22328 ;
  assign n42069 = ~n22314 ;
  assign n22330 = n42069 & n22329 ;
  assign n42070 = ~n22330 ;
  assign n22331 = n168 & n42070 ;
  assign n42071 = ~n21493 ;
  assign n21499 = n21005 & n42071 ;
  assign n21500 = n41657 & n21499 ;
  assign n21827 = n21500 & n140 ;
  assign n21501 = n21492 | n21493 ;
  assign n42072 = ~n21501 ;
  assign n21830 = n42072 & n140 ;
  assign n21831 = n21005 | n21830 ;
  assign n42073 = ~n21827 ;
  assign n21832 = n42073 & n21831 ;
  assign n22315 = n4934 | n22314 ;
  assign n42074 = ~n22315 ;
  assign n22332 = n42074 & n22329 ;
  assign n22333 = n21832 | n22332 ;
  assign n42075 = ~n22331 ;
  assign n22334 = n42075 & n22333 ;
  assign n42076 = ~n22334 ;
  assign n22335 = n169 & n42076 ;
  assign n21498 = n21132 & n41667 ;
  assign n42077 = ~n21513 ;
  assign n21526 = n21498 & n42077 ;
  assign n21829 = n21526 & n140 ;
  assign n21527 = n21496 | n21513 ;
  assign n42078 = ~n21527 ;
  assign n21851 = n42078 & n140 ;
  assign n21852 = n21132 | n21851 ;
  assign n42079 = ~n21829 ;
  assign n21853 = n42079 & n21852 ;
  assign n22338 = n42058 & n22324 ;
  assign n22339 = n21970 | n22338 ;
  assign n42080 = ~n22326 ;
  assign n22340 = n42080 & n22339 ;
  assign n42081 = ~n22340 ;
  assign n22341 = n167 & n42081 ;
  assign n22342 = n42068 & n22339 ;
  assign n22343 = n22149 | n22342 ;
  assign n42082 = ~n22341 ;
  assign n22344 = n42082 & n22343 ;
  assign n42083 = ~n22344 ;
  assign n22345 = n4934 & n42083 ;
  assign n22346 = n169 | n22345 ;
  assign n42084 = ~n22346 ;
  assign n22347 = n22333 & n42084 ;
  assign n22348 = n21853 | n22347 ;
  assign n42085 = ~n22335 ;
  assign n22349 = n42085 & n22348 ;
  assign n42086 = ~n22349 ;
  assign n22350 = n170 & n42086 ;
  assign n21525 = n21516 | n21517 ;
  assign n42087 = ~n21525 ;
  assign n21825 = n42087 & n140 ;
  assign n21826 = n21037 | n21825 ;
  assign n42088 = ~n21517 ;
  assign n21523 = n21037 & n42088 ;
  assign n21524 = n41673 & n21523 ;
  assign n22250 = n21524 & n22030 ;
  assign n42089 = ~n22250 ;
  assign n22251 = n21826 & n42089 ;
  assign n22336 = n170 | n22335 ;
  assign n42090 = ~n22336 ;
  assign n22351 = n42090 & n22348 ;
  assign n22352 = n22251 | n22351 ;
  assign n42091 = ~n22350 ;
  assign n22353 = n42091 & n22352 ;
  assign n42092 = ~n22353 ;
  assign n22354 = n3940 & n42092 ;
  assign n21551 = n21520 | n21537 ;
  assign n42093 = ~n21551 ;
  assign n21861 = n42093 & n140 ;
  assign n21862 = n21047 | n21861 ;
  assign n21522 = n21047 & n41683 ;
  assign n42094 = ~n21537 ;
  assign n21550 = n21522 & n42094 ;
  assign n22035 = n21550 & n22030 ;
  assign n42095 = ~n22035 ;
  assign n22036 = n21862 & n42095 ;
  assign n22357 = n42074 & n22343 ;
  assign n22358 = n21832 | n22357 ;
  assign n42096 = ~n22345 ;
  assign n22359 = n42096 & n22358 ;
  assign n42097 = ~n22359 ;
  assign n22360 = n169 & n42097 ;
  assign n22361 = n42084 & n22358 ;
  assign n22362 = n21853 | n22361 ;
  assign n42098 = ~n22360 ;
  assign n22363 = n42098 & n22362 ;
  assign n42099 = ~n22363 ;
  assign n22364 = n170 & n42099 ;
  assign n22365 = n3940 | n22364 ;
  assign n42100 = ~n22365 ;
  assign n22366 = n22352 & n42100 ;
  assign n22367 = n22036 | n22366 ;
  assign n42101 = ~n22354 ;
  assign n22368 = n42101 & n22367 ;
  assign n42102 = ~n22368 ;
  assign n22369 = n172 & n42102 ;
  assign n42103 = ~n21541 ;
  assign n21547 = n21018 & n42103 ;
  assign n21548 = n41689 & n21547 ;
  assign n21828 = n21548 & n140 ;
  assign n21549 = n21540 | n21541 ;
  assign n42104 = ~n21549 ;
  assign n21844 = n42104 & n140 ;
  assign n21845 = n21018 | n21844 ;
  assign n42105 = ~n21828 ;
  assign n21846 = n42105 & n21845 ;
  assign n22355 = n3631 | n22354 ;
  assign n42106 = ~n22355 ;
  assign n22370 = n42106 & n22367 ;
  assign n22371 = n21846 | n22370 ;
  assign n42107 = ~n22369 ;
  assign n22372 = n42107 & n22371 ;
  assign n42108 = ~n22372 ;
  assign n22373 = n173 & n42108 ;
  assign n21575 = n21544 | n21561 ;
  assign n42109 = ~n21575 ;
  assign n21887 = n42109 & n140 ;
  assign n21888 = n21134 | n21887 ;
  assign n21546 = n21134 & n41699 ;
  assign n42110 = ~n21561 ;
  assign n21574 = n21546 & n42110 ;
  assign n21893 = n21574 & n140 ;
  assign n42111 = ~n21893 ;
  assign n21894 = n21888 & n42111 ;
  assign n22376 = n42090 & n22362 ;
  assign n22377 = n22251 | n22376 ;
  assign n42112 = ~n22364 ;
  assign n22378 = n42112 & n22377 ;
  assign n42113 = ~n22378 ;
  assign n22379 = n171 & n42113 ;
  assign n22380 = n42100 & n22377 ;
  assign n22381 = n22036 | n22380 ;
  assign n42114 = ~n22379 ;
  assign n22382 = n42114 & n22381 ;
  assign n42115 = ~n22382 ;
  assign n22383 = n3631 & n42115 ;
  assign n22384 = n173 | n22383 ;
  assign n42116 = ~n22384 ;
  assign n22385 = n22371 & n42116 ;
  assign n22386 = n21894 | n22385 ;
  assign n42117 = ~n22373 ;
  assign n22387 = n42117 & n22386 ;
  assign n42118 = ~n22387 ;
  assign n22388 = n174 & n42118 ;
  assign n42119 = ~n21565 ;
  assign n21571 = n21138 & n42119 ;
  assign n21572 = n41705 & n21571 ;
  assign n21835 = n21572 & n140 ;
  assign n21573 = n21564 | n21565 ;
  assign n42120 = ~n21573 ;
  assign n21836 = n42120 & n140 ;
  assign n21837 = n21138 | n21836 ;
  assign n42121 = ~n21835 ;
  assign n21838 = n42121 & n21837 ;
  assign n22374 = n174 | n22373 ;
  assign n42122 = ~n22374 ;
  assign n22389 = n42122 & n22386 ;
  assign n22390 = n21838 | n22389 ;
  assign n42123 = ~n22388 ;
  assign n22391 = n42123 & n22390 ;
  assign n42124 = ~n22391 ;
  assign n22392 = n2753 & n42124 ;
  assign n21570 = n21113 & n41715 ;
  assign n42125 = ~n21585 ;
  assign n21598 = n21570 & n42125 ;
  assign n21985 = n21598 & n140 ;
  assign n21599 = n21568 | n21585 ;
  assign n42126 = ~n21599 ;
  assign n21988 = n42126 & n140 ;
  assign n21989 = n21113 | n21988 ;
  assign n42127 = ~n21985 ;
  assign n21990 = n42127 & n21989 ;
  assign n22395 = n42106 & n22381 ;
  assign n22396 = n21846 | n22395 ;
  assign n42128 = ~n22383 ;
  assign n22397 = n42128 & n22396 ;
  assign n42129 = ~n22397 ;
  assign n22398 = n173 & n42129 ;
  assign n22399 = n42116 & n22396 ;
  assign n22400 = n21894 | n22399 ;
  assign n42130 = ~n22398 ;
  assign n22401 = n42130 & n22400 ;
  assign n42131 = ~n22401 ;
  assign n22402 = n174 & n42131 ;
  assign n22403 = n2753 | n22402 ;
  assign n42132 = ~n22403 ;
  assign n22404 = n22390 & n42132 ;
  assign n22405 = n21990 | n22404 ;
  assign n42133 = ~n22392 ;
  assign n22406 = n42133 & n22405 ;
  assign n42134 = ~n22406 ;
  assign n22407 = n176 & n42134 ;
  assign n42135 = ~n21589 ;
  assign n21595 = n21140 & n42135 ;
  assign n21596 = n41721 & n21595 ;
  assign n21916 = n21596 & n140 ;
  assign n21597 = n21588 | n21589 ;
  assign n42136 = ~n21597 ;
  assign n21991 = n42136 & n140 ;
  assign n21992 = n21140 | n21991 ;
  assign n42137 = ~n21916 ;
  assign n21993 = n42137 & n21992 ;
  assign n22393 = n2431 | n22392 ;
  assign n42138 = ~n22393 ;
  assign n22408 = n42138 & n22405 ;
  assign n22409 = n21993 | n22408 ;
  assign n42139 = ~n22407 ;
  assign n22410 = n42139 & n22409 ;
  assign n42140 = ~n22410 ;
  assign n22411 = n177 & n42140 ;
  assign n21594 = n21144 & n41731 ;
  assign n42141 = ~n21609 ;
  assign n21622 = n21594 & n42141 ;
  assign n21994 = n21622 & n140 ;
  assign n21623 = n21592 | n21609 ;
  assign n42142 = ~n21623 ;
  assign n21995 = n42142 & n140 ;
  assign n21996 = n21144 | n21995 ;
  assign n42143 = ~n21994 ;
  assign n21997 = n42143 & n21996 ;
  assign n22414 = n42122 & n22400 ;
  assign n22415 = n21838 | n22414 ;
  assign n42144 = ~n22402 ;
  assign n22416 = n42144 & n22415 ;
  assign n42145 = ~n22416 ;
  assign n22417 = n175 & n42145 ;
  assign n22418 = n42132 & n22415 ;
  assign n22419 = n21990 | n22418 ;
  assign n42146 = ~n22417 ;
  assign n22420 = n42146 & n22419 ;
  assign n42147 = ~n22420 ;
  assign n22421 = n2431 & n42147 ;
  assign n22422 = n177 | n22421 ;
  assign n42148 = ~n22422 ;
  assign n22423 = n22409 & n42148 ;
  assign n22424 = n21997 | n22423 ;
  assign n42149 = ~n22411 ;
  assign n22425 = n42149 & n22424 ;
  assign n42150 = ~n22425 ;
  assign n22426 = n178 & n42150 ;
  assign n21621 = n21612 | n21613 ;
  assign n42151 = ~n21621 ;
  assign n21847 = n42151 & n140 ;
  assign n21848 = n21148 | n21847 ;
  assign n42152 = ~n21613 ;
  assign n21619 = n21148 & n42152 ;
  assign n21620 = n41737 & n21619 ;
  assign n21983 = n21620 & n140 ;
  assign n42153 = ~n21983 ;
  assign n21984 = n21848 & n42153 ;
  assign n22412 = n178 | n22411 ;
  assign n42154 = ~n22412 ;
  assign n22427 = n42154 & n22424 ;
  assign n22428 = n21984 | n22427 ;
  assign n42155 = ~n22426 ;
  assign n22429 = n42155 & n22428 ;
  assign n42156 = ~n22429 ;
  assign n22430 = n1707 & n42156 ;
  assign n21647 = n21616 | n21633 ;
  assign n42157 = ~n21647 ;
  assign n21858 = n42157 & n140 ;
  assign n21859 = n21152 | n21858 ;
  assign n21618 = n21152 & n41747 ;
  assign n42158 = ~n21633 ;
  assign n21646 = n21618 & n42158 ;
  assign n22031 = n21646 & n22030 ;
  assign n42159 = ~n22031 ;
  assign n22032 = n21859 & n42159 ;
  assign n22433 = n42138 & n22419 ;
  assign n22434 = n21993 | n22433 ;
  assign n42160 = ~n22421 ;
  assign n22435 = n42160 & n22434 ;
  assign n42161 = ~n22435 ;
  assign n22436 = n177 & n42161 ;
  assign n22437 = n42148 & n22434 ;
  assign n22438 = n21997 | n22437 ;
  assign n42162 = ~n22436 ;
  assign n22439 = n42162 & n22438 ;
  assign n42163 = ~n22439 ;
  assign n22440 = n178 & n42163 ;
  assign n22441 = n1707 | n22440 ;
  assign n42164 = ~n22441 ;
  assign n22442 = n22428 & n42164 ;
  assign n22443 = n22032 | n22442 ;
  assign n42165 = ~n22430 ;
  assign n22444 = n42165 & n22443 ;
  assign n42166 = ~n22444 ;
  assign n22445 = n180 & n42166 ;
  assign n21645 = n21636 | n21637 ;
  assign n42167 = ~n21645 ;
  assign n21906 = n42167 & n140 ;
  assign n21907 = n21155 | n21906 ;
  assign n42168 = ~n21637 ;
  assign n21643 = n21155 & n42168 ;
  assign n21644 = n41753 & n21643 ;
  assign n21998 = n21644 & n140 ;
  assign n42169 = ~n21998 ;
  assign n21999 = n21907 & n42169 ;
  assign n22431 = n1487 | n22430 ;
  assign n42170 = ~n22431 ;
  assign n22446 = n42170 & n22443 ;
  assign n22447 = n21999 | n22446 ;
  assign n42171 = ~n22445 ;
  assign n22448 = n42171 & n22447 ;
  assign n42172 = ~n22448 ;
  assign n22449 = n181 & n42172 ;
  assign n21642 = n21160 & n41763 ;
  assign n42173 = ~n21657 ;
  assign n21669 = n21642 & n42173 ;
  assign n22000 = n21669 & n140 ;
  assign n21668 = n21640 | n21657 ;
  assign n42174 = ~n21668 ;
  assign n22003 = n42174 & n140 ;
  assign n22004 = n21160 | n22003 ;
  assign n42175 = ~n22000 ;
  assign n22005 = n42175 & n22004 ;
  assign n22452 = n42154 & n22438 ;
  assign n22453 = n21984 | n22452 ;
  assign n42176 = ~n22440 ;
  assign n22454 = n42176 & n22453 ;
  assign n42177 = ~n22454 ;
  assign n22455 = n179 & n42177 ;
  assign n22456 = n42164 & n22453 ;
  assign n22457 = n22032 | n22456 ;
  assign n42178 = ~n22455 ;
  assign n22458 = n42178 & n22457 ;
  assign n42179 = ~n22458 ;
  assign n22459 = n1487 & n42179 ;
  assign n22460 = n181 | n22459 ;
  assign n42180 = ~n22460 ;
  assign n22461 = n22447 & n42180 ;
  assign n22462 = n22005 | n22461 ;
  assign n42181 = ~n22449 ;
  assign n22463 = n42181 & n22462 ;
  assign n42182 = ~n22463 ;
  assign n22464 = n182 & n42182 ;
  assign n21695 = n21661 | n21677 ;
  assign n42183 = ~n21695 ;
  assign n21962 = n42183 & n140 ;
  assign n21963 = n21164 | n21962 ;
  assign n42184 = ~n21661 ;
  assign n21667 = n21164 & n42184 ;
  assign n21694 = n21667 & n41790 ;
  assign n21986 = n21694 & n140 ;
  assign n42185 = ~n21986 ;
  assign n21987 = n21963 & n42185 ;
  assign n22450 = n182 | n22449 ;
  assign n42186 = ~n22450 ;
  assign n22465 = n42186 & n22462 ;
  assign n22466 = n21987 | n22465 ;
  assign n42187 = ~n22464 ;
  assign n22467 = n42187 & n22466 ;
  assign n42188 = ~n22467 ;
  assign n22468 = n996 & n42188 ;
  assign n22470 = n42170 & n22457 ;
  assign n22471 = n21999 | n22470 ;
  assign n42189 = ~n22459 ;
  assign n22472 = n42189 & n22471 ;
  assign n42190 = ~n22472 ;
  assign n22473 = n181 & n42190 ;
  assign n22474 = n42180 & n22471 ;
  assign n22475 = n22005 | n22474 ;
  assign n42191 = ~n22473 ;
  assign n22476 = n42191 & n22475 ;
  assign n42192 = ~n22476 ;
  assign n22477 = n182 & n42192 ;
  assign n22478 = n183 | n22477 ;
  assign n42193 = ~n22478 ;
  assign n22479 = n22466 & n42193 ;
  assign n21692 = n21664 | n21679 ;
  assign n42194 = ~n21692 ;
  assign n22001 = n42194 & n140 ;
  assign n22002 = n21166 | n22001 ;
  assign n21665 = n21166 & n41779 ;
  assign n42195 = ~n21679 ;
  assign n21693 = n21665 & n42195 ;
  assign n22542 = n21693 & n22030 ;
  assign n42196 = ~n22542 ;
  assign n22543 = n22002 & n42196 ;
  assign n22546 = n22479 | n22543 ;
  assign n42197 = ~n22468 ;
  assign n22547 = n42197 & n22546 ;
  assign n42198 = ~n22547 ;
  assign n22548 = n184 & n42198 ;
  assign n42199 = ~n21683 ;
  assign n21689 = n21169 & n42199 ;
  assign n21690 = n41785 & n21689 ;
  assign n22006 = n21690 & n140 ;
  assign n21691 = n21682 | n21683 ;
  assign n42200 = ~n21691 ;
  assign n22007 = n42200 & n140 ;
  assign n22008 = n21169 | n22007 ;
  assign n42201 = ~n22006 ;
  assign n22009 = n42201 & n22008 ;
  assign n22469 = n838 | n22468 ;
  assign n42202 = ~n22469 ;
  assign n22549 = n42202 & n22546 ;
  assign n22550 = n22009 | n22549 ;
  assign n42203 = ~n22548 ;
  assign n22551 = n42203 & n22550 ;
  assign n42204 = ~n22551 ;
  assign n22552 = n185 & n42204 ;
  assign n21719 = n21686 | n21705 ;
  assign n42205 = ~n21719 ;
  assign n21928 = n42205 & n140 ;
  assign n21929 = n21174 | n21928 ;
  assign n21688 = n21174 & n41795 ;
  assign n42206 = ~n21705 ;
  assign n21718 = n21688 & n42206 ;
  assign n22010 = n21718 & n140 ;
  assign n42207 = ~n22010 ;
  assign n22011 = n21929 & n42207 ;
  assign n22480 = n42186 & n22475 ;
  assign n22481 = n21987 | n22480 ;
  assign n42208 = ~n22477 ;
  assign n22482 = n42208 & n22481 ;
  assign n42209 = ~n22482 ;
  assign n22483 = n183 & n42209 ;
  assign n22484 = n42193 & n22481 ;
  assign n22555 = n22484 | n22543 ;
  assign n42210 = ~n22483 ;
  assign n22556 = n42210 & n22555 ;
  assign n42211 = ~n22556 ;
  assign n22557 = n838 & n42211 ;
  assign n22558 = n185 | n22557 ;
  assign n42212 = ~n22558 ;
  assign n22559 = n22550 & n42212 ;
  assign n22560 = n22011 | n22559 ;
  assign n42213 = ~n22552 ;
  assign n22561 = n42213 & n22560 ;
  assign n42214 = ~n22561 ;
  assign n22562 = n186 & n42214 ;
  assign n42215 = ~n21709 ;
  assign n21715 = n21176 & n42215 ;
  assign n21716 = n41801 & n21715 ;
  assign n22014 = n21716 & n140 ;
  assign n21717 = n21708 | n21709 ;
  assign n42216 = ~n21717 ;
  assign n22015 = n42216 & n140 ;
  assign n22016 = n21176 | n22015 ;
  assign n42217 = ~n22014 ;
  assign n22017 = n42217 & n22016 ;
  assign n22553 = n186 | n22552 ;
  assign n42218 = ~n22553 ;
  assign n22563 = n42218 & n22560 ;
  assign n22564 = n22017 | n22563 ;
  assign n42219 = ~n22562 ;
  assign n22565 = n42219 & n22564 ;
  assign n42220 = ~n22565 ;
  assign n22566 = n528 & n42220 ;
  assign n21736 = n21712 | n21729 ;
  assign n42221 = ~n21736 ;
  assign n21909 = n42221 & n140 ;
  assign n21910 = n21178 | n21909 ;
  assign n21714 = n21178 & n41811 ;
  assign n42222 = ~n21729 ;
  assign n21735 = n21714 & n42222 ;
  assign n22018 = n21735 & n140 ;
  assign n42223 = ~n22018 ;
  assign n22019 = n21910 & n42223 ;
  assign n22569 = n42202 & n22555 ;
  assign n22570 = n22009 | n22569 ;
  assign n42224 = ~n22557 ;
  assign n22571 = n42224 & n22570 ;
  assign n42225 = ~n22571 ;
  assign n22572 = n185 & n42225 ;
  assign n22573 = n42212 & n22570 ;
  assign n22574 = n22011 | n22573 ;
  assign n42226 = ~n22572 ;
  assign n22575 = n42226 & n22574 ;
  assign n42227 = ~n22575 ;
  assign n22576 = n186 & n42227 ;
  assign n22577 = n528 | n22576 ;
  assign n42228 = ~n22577 ;
  assign n22578 = n22564 & n42228 ;
  assign n22579 = n22019 | n22578 ;
  assign n42229 = ~n22566 ;
  assign n22580 = n42229 & n22579 ;
  assign n42230 = ~n22580 ;
  assign n22581 = n188 & n42230 ;
  assign n22567 = n413 | n22566 ;
  assign n42231 = ~n22567 ;
  assign n22582 = n42231 & n22579 ;
  assign n42232 = ~n21733 ;
  assign n21785 = n42232 & n21766 ;
  assign n21786 = n41817 & n21785 ;
  assign n21975 = n21786 & n140 ;
  assign n21734 = n21732 | n21733 ;
  assign n42233 = ~n21734 ;
  assign n21898 = n42233 & n140 ;
  assign n22623 = n21766 | n21898 ;
  assign n42234 = ~n21975 ;
  assign n22624 = n42234 & n22623 ;
  assign n22625 = n22582 | n22624 ;
  assign n42235 = ~n22581 ;
  assign n22626 = n42235 & n22625 ;
  assign n42236 = ~n22626 ;
  assign n22627 = n189 & n42236 ;
  assign n21784 = n21769 | n21772 ;
  assign n42237 = ~n21784 ;
  assign n21899 = n42237 & n140 ;
  assign n21900 = n21182 | n21899 ;
  assign n21770 = n21182 & n41827 ;
  assign n42238 = ~n21772 ;
  assign n21783 = n21770 & n42238 ;
  assign n22020 = n21783 & n140 ;
  assign n42239 = ~n22020 ;
  assign n22021 = n21900 & n42239 ;
  assign n22583 = n42218 & n22574 ;
  assign n22584 = n22017 | n22583 ;
  assign n42240 = ~n22576 ;
  assign n22585 = n42240 & n22584 ;
  assign n42241 = ~n22585 ;
  assign n22586 = n187 & n42241 ;
  assign n22587 = n42228 & n22584 ;
  assign n22588 = n22019 | n22587 ;
  assign n42242 = ~n22586 ;
  assign n22589 = n42242 & n22588 ;
  assign n42243 = ~n22589 ;
  assign n22590 = n413 & n42243 ;
  assign n22591 = n189 | n22590 ;
  assign n42244 = ~n22591 ;
  assign n22630 = n42244 & n22625 ;
  assign n22631 = n22021 | n22630 ;
  assign n42245 = ~n22627 ;
  assign n22632 = n42245 & n22631 ;
  assign n42246 = ~n22632 ;
  assign n22633 = n190 & n42246 ;
  assign n22615 = n41832 & n21791 ;
  assign n42247 = ~n22615 ;
  assign n22616 = n21184 & n42247 ;
  assign n22617 = n41833 & n22616 ;
  assign n22618 = n140 & n22617 ;
  assign n22619 = n21775 | n22615 ;
  assign n42248 = ~n22619 ;
  assign n22620 = n140 & n42248 ;
  assign n22621 = n21184 | n22620 ;
  assign n42249 = ~n22618 ;
  assign n22622 = n42249 & n22621 ;
  assign n22628 = n190 | n22627 ;
  assign n42250 = ~n22628 ;
  assign n22634 = n42250 & n22631 ;
  assign n22635 = n22622 | n22634 ;
  assign n42251 = ~n22633 ;
  assign n22636 = n42251 & n22635 ;
  assign n42252 = ~n22636 ;
  assign n22637 = n287 & n42252 ;
  assign n21800 = n21779 | n21795 ;
  assign n42253 = ~n21800 ;
  assign n21865 = n42253 & n140 ;
  assign n21866 = n21055 | n21865 ;
  assign n21782 = n21055 & n41847 ;
  assign n42254 = ~n21795 ;
  assign n21799 = n21782 & n42254 ;
  assign n21869 = n21799 & n140 ;
  assign n42255 = ~n21869 ;
  assign n21870 = n21866 & n42255 ;
  assign n22592 = n42231 & n22588 ;
  assign n22642 = n22592 | n22624 ;
  assign n42256 = ~n22590 ;
  assign n22643 = n42256 & n22642 ;
  assign n42257 = ~n22643 ;
  assign n22644 = n189 & n42257 ;
  assign n22645 = n42244 & n22642 ;
  assign n22646 = n22021 | n22645 ;
  assign n42258 = ~n22644 ;
  assign n22647 = n42258 & n22646 ;
  assign n42259 = ~n22647 ;
  assign n22648 = n190 & n42259 ;
  assign n22653 = n287 | n22648 ;
  assign n42260 = ~n22653 ;
  assign n22654 = n22635 & n42260 ;
  assign n22655 = n21870 | n22654 ;
  assign n42261 = ~n22637 ;
  assign n22656 = n42261 & n22655 ;
  assign n22657 = n22612 | n22656 ;
  assign n22658 = n31336 & n22657 ;
  assign n21754 = n21129 | n21750 ;
  assign n42262 = ~n21754 ;
  assign n21755 = n21027 & n42262 ;
  assign n21756 = n41857 & n21755 ;
  assign n21808 = n21756 & n41858 ;
  assign n21819 = n21808 & n41859 ;
  assign n21811 = n192 & n21810 ;
  assign n42263 = ~n21130 ;
  assign n22022 = n42263 & n140 ;
  assign n42264 = ~n22022 ;
  assign n22023 = n21809 & n42264 ;
  assign n42265 = ~n22023 ;
  assign n22024 = n21811 & n42265 ;
  assign n22025 = n21819 | n22024 ;
  assign n22638 = n22611 & n42261 ;
  assign n22659 = n22638 & n22655 ;
  assign n22660 = n22025 | n22659 ;
  assign n22661 = n22658 | n22660 ;
  assign n22649 = n191 | n22648 ;
  assign n42266 = ~n22649 ;
  assign n22650 = n22635 & n42266 ;
  assign n22652 = n22637 | n22650 ;
  assign n22681 = n42250 & n22646 ;
  assign n22682 = n22622 | n22681 ;
  assign n42267 = ~n22648 ;
  assign n22683 = n42267 & n22682 ;
  assign n42268 = ~n22683 ;
  assign n22684 = n191 & n42268 ;
  assign n22685 = n42266 & n22682 ;
  assign n22686 = n21870 | n22685 ;
  assign n42269 = ~n22684 ;
  assign n22687 = n42269 & n22686 ;
  assign n22688 = n22612 | n22687 ;
  assign n22689 = n31336 & n22688 ;
  assign n22690 = n22638 & n22686 ;
  assign n22691 = n22025 | n22690 ;
  assign n139 = n22689 | n22691 ;
  assign n42270 = ~n22652 ;
  assign n23186 = n42270 & n139 ;
  assign n23187 = n21870 | n23186 ;
  assign n22639 = n21870 & n42261 ;
  assign n42271 = ~n22650 ;
  assign n22651 = n22639 & n42271 ;
  assign n23465 = n22651 & n139 ;
  assign n42272 = ~n23465 ;
  assign n23466 = n23187 & n42272 ;
  assign n22670 = n22611 | n22656 ;
  assign n42273 = ~n22670 ;
  assign n23485 = n42273 & n139 ;
  assign n23486 = n22659 | n23485 ;
  assign n23487 = n23466 | n23486 ;
  assign n42274 = ~n21819 ;
  assign n21892 = n42274 & n140 ;
  assign n42275 = ~n22024 ;
  assign n22026 = n21892 & n42275 ;
  assign n42276 = ~n22659 ;
  assign n22672 = n22026 & n42276 ;
  assign n42277 = ~n22658 ;
  assign n22673 = n42277 & n22672 ;
  assign n42278 = ~n239 ;
  assign n22732 = n42278 & n139 ;
  assign n22734 = n22673 | n22732 ;
  assign n22735 = x22 & n22734 ;
  assign n22674 = x22 | n22673 ;
  assign n22736 = n22674 | n22732 ;
  assign n42279 = ~n22735 ;
  assign n22737 = n42279 & n22736 ;
  assign n242 = x18 | x19 ;
  assign n42280 = ~x20 ;
  assign n244 = n42280 & n242 ;
  assign n42281 = ~n22661 ;
  assign n22665 = x20 & n42281 ;
  assign n22666 = n244 | n22665 ;
  assign n42282 = ~n22666 ;
  assign n22667 = n22030 & n42282 ;
  assign n22668 = n141 | n22667 ;
  assign n22727 = n42280 & n139 ;
  assign n42283 = ~n22727 ;
  assign n22728 = x21 & n42283 ;
  assign n22733 = n22728 | n22732 ;
  assign n243 = x20 | n242 ;
  assign n21757 = n243 & n41856 ;
  assign n21758 = n41857 & n21757 ;
  assign n21807 = n21758 & n41858 ;
  assign n21821 = n21807 & n41859 ;
  assign n22799 = x20 & n139 ;
  assign n42284 = ~n22799 ;
  assign n22800 = n21821 & n42284 ;
  assign n22801 = n22733 | n22800 ;
  assign n42285 = ~n22668 ;
  assign n22807 = n42285 & n22801 ;
  assign n22808 = n22737 | n22807 ;
  assign n22669 = n140 & n42282 ;
  assign n42286 = ~n22669 ;
  assign n22811 = n42286 & n22801 ;
  assign n42287 = ~n22811 ;
  assign n22812 = n141 & n42287 ;
  assign n22813 = n142 | n22812 ;
  assign n42288 = ~n22813 ;
  assign n22814 = n22808 & n42288 ;
  assign n22144 = n21902 | n22039 ;
  assign n42289 = ~n22144 ;
  assign n22778 = n42289 & n139 ;
  assign n22779 = n21941 | n22778 ;
  assign n22145 = n21941 & n42289 ;
  assign n22820 = n22145 & n139 ;
  assign n42290 = ~n22820 ;
  assign n22821 = n22779 & n42290 ;
  assign n22822 = n22814 | n22821 ;
  assign n42291 = ~n22667 ;
  assign n22802 = n42291 & n22801 ;
  assign n42292 = ~n22802 ;
  assign n22803 = n141 & n42292 ;
  assign n22824 = n243 & n42284 ;
  assign n42293 = ~n22824 ;
  assign n22825 = n140 & n42293 ;
  assign n22826 = n141 | n22825 ;
  assign n42294 = ~n22826 ;
  assign n22827 = n22801 & n42294 ;
  assign n22828 = n22737 | n22827 ;
  assign n42295 = ~n22803 ;
  assign n22829 = n42295 & n22828 ;
  assign n42296 = ~n22829 ;
  assign n22830 = n142 & n42296 ;
  assign n42297 = ~n22830 ;
  assign n22831 = n22822 & n42297 ;
  assign n42298 = ~n22831 ;
  assign n22832 = n19362 & n42298 ;
  assign n21951 = n21943 | n21947 ;
  assign n42299 = ~n21951 ;
  assign n22780 = n42299 & n139 ;
  assign n22781 = n21921 | n22780 ;
  assign n42300 = ~n21943 ;
  assign n21945 = n21921 & n42300 ;
  assign n42301 = ~n21947 ;
  assign n21950 = n21945 & n42301 ;
  assign n22784 = n21950 & n139 ;
  assign n42302 = ~n22784 ;
  assign n22785 = n22781 & n42302 ;
  assign n22836 = n19362 | n22830 ;
  assign n42303 = ~n22836 ;
  assign n22837 = n22822 & n42303 ;
  assign n22838 = n22785 | n22837 ;
  assign n42304 = ~n22832 ;
  assign n22839 = n42304 & n22838 ;
  assign n42305 = ~n22839 ;
  assign n22840 = n144 & n42305 ;
  assign n22833 = n144 | n22832 ;
  assign n42306 = ~n22833 ;
  assign n22841 = n42306 & n22838 ;
  assign n22062 = n21973 & n41876 ;
  assign n42307 = ~n21949 ;
  assign n22063 = n42307 & n22062 ;
  assign n22768 = n22063 & n139 ;
  assign n22064 = n21949 | n22061 ;
  assign n42308 = ~n22064 ;
  assign n22864 = n42308 & n139 ;
  assign n22865 = n21973 | n22864 ;
  assign n42309 = ~n22768 ;
  assign n22866 = n42309 & n22865 ;
  assign n22867 = n22841 | n22866 ;
  assign n42310 = ~n22840 ;
  assign n22868 = n42310 & n22867 ;
  assign n42311 = ~n22868 ;
  assign n22869 = n145 & n42311 ;
  assign n22060 = n22045 | n22048 ;
  assign n42312 = ~n22060 ;
  assign n22758 = n42312 & n139 ;
  assign n22759 = n21913 | n22758 ;
  assign n42313 = ~n22048 ;
  assign n22058 = n21913 & n42313 ;
  assign n22059 = n41904 & n22058 ;
  assign n22782 = n22059 & n139 ;
  assign n42314 = ~n22782 ;
  assign n22783 = n22759 & n42314 ;
  assign n22804 = n142 | n22803 ;
  assign n42315 = ~n22804 ;
  assign n22809 = n42315 & n22808 ;
  assign n22823 = n22809 | n22821 ;
  assign n22846 = n22823 & n42303 ;
  assign n22847 = n22785 | n22846 ;
  assign n22849 = n22823 & n42297 ;
  assign n42316 = ~n22849 ;
  assign n22850 = n143 & n42316 ;
  assign n42317 = ~n22850 ;
  assign n22851 = n22847 & n42317 ;
  assign n42318 = ~n22851 ;
  assign n22852 = n18797 & n42318 ;
  assign n22853 = n145 | n22852 ;
  assign n42319 = ~n22853 ;
  assign n22871 = n42319 & n22867 ;
  assign n22872 = n22783 | n22871 ;
  assign n42320 = ~n22869 ;
  assign n22873 = n42320 & n22872 ;
  assign n42321 = ~n22873 ;
  assign n22874 = n146 & n42321 ;
  assign n22870 = n146 | n22869 ;
  assign n42322 = ~n22870 ;
  assign n22875 = n42322 & n22872 ;
  assign n22057 = n22051 | n22052 ;
  assign n42323 = ~n22057 ;
  assign n22858 = n42323 & n139 ;
  assign n22859 = n21961 | n22858 ;
  assign n22088 = n21961 & n41893 ;
  assign n42324 = ~n22052 ;
  assign n22089 = n42324 & n22088 ;
  assign n22898 = n22089 & n139 ;
  assign n42325 = ~n22898 ;
  assign n22899 = n22859 & n42325 ;
  assign n22900 = n22875 | n22899 ;
  assign n42326 = ~n22874 ;
  assign n22901 = n42326 & n22900 ;
  assign n42327 = ~n22901 ;
  assign n22902 = n16322 & n42327 ;
  assign n22087 = n22055 | n22075 ;
  assign n42328 = ~n22087 ;
  assign n22707 = n42328 & n139 ;
  assign n22708 = n21890 | n22707 ;
  assign n42329 = ~n22075 ;
  assign n22085 = n21890 & n42329 ;
  assign n22086 = n41920 & n22085 ;
  assign n22862 = n22086 & n139 ;
  assign n42330 = ~n22862 ;
  assign n22863 = n22708 & n42330 ;
  assign n22848 = n42306 & n22847 ;
  assign n22882 = n22848 | n22866 ;
  assign n42331 = ~n22852 ;
  assign n22883 = n42331 & n22882 ;
  assign n42332 = ~n22883 ;
  assign n22884 = n145 & n42332 ;
  assign n22885 = n42319 & n22882 ;
  assign n22886 = n22783 | n22885 ;
  assign n42333 = ~n22884 ;
  assign n22887 = n42333 & n22886 ;
  assign n42334 = ~n22887 ;
  assign n22888 = n146 & n42334 ;
  assign n22889 = n147 | n22888 ;
  assign n42335 = ~n22889 ;
  assign n22904 = n42335 & n22900 ;
  assign n22905 = n22863 | n22904 ;
  assign n42336 = ~n22902 ;
  assign n22906 = n42336 & n22905 ;
  assign n42337 = ~n22906 ;
  assign n22907 = n148 & n42337 ;
  assign n22903 = n148 | n22902 ;
  assign n42338 = ~n22903 ;
  assign n22908 = n42338 & n22905 ;
  assign n22111 = n21935 & n41909 ;
  assign n42339 = ~n22079 ;
  assign n22112 = n42339 & n22111 ;
  assign n22893 = n22112 & n139 ;
  assign n22084 = n22078 | n22079 ;
  assign n42340 = ~n22084 ;
  assign n22929 = n42340 & n139 ;
  assign n22930 = n21935 | n22929 ;
  assign n42341 = ~n22893 ;
  assign n22931 = n42341 & n22930 ;
  assign n22932 = n22908 | n22931 ;
  assign n42342 = ~n22907 ;
  assign n22933 = n42342 & n22932 ;
  assign n42343 = ~n22933 ;
  assign n22934 = n149 & n42343 ;
  assign n42344 = ~n22099 ;
  assign n22108 = n21958 & n42344 ;
  assign n22109 = n41933 & n22108 ;
  assign n22788 = n22109 & n139 ;
  assign n22110 = n22082 | n22099 ;
  assign n42345 = ~n22110 ;
  assign n22793 = n42345 & n139 ;
  assign n22794 = n21958 | n22793 ;
  assign n42346 = ~n22788 ;
  assign n22795 = n42346 & n22794 ;
  assign n22890 = n42322 & n22886 ;
  assign n22915 = n22890 | n22899 ;
  assign n42347 = ~n22888 ;
  assign n22916 = n42347 & n22915 ;
  assign n42348 = ~n22916 ;
  assign n22917 = n147 & n42348 ;
  assign n22918 = n42335 & n22915 ;
  assign n22919 = n22863 | n22918 ;
  assign n42349 = ~n22917 ;
  assign n22920 = n42349 & n22919 ;
  assign n42350 = ~n22920 ;
  assign n22921 = n15807 & n42350 ;
  assign n22922 = n149 | n22921 ;
  assign n42351 = ~n22922 ;
  assign n22936 = n42351 & n22932 ;
  assign n22937 = n22795 | n22936 ;
  assign n42352 = ~n22934 ;
  assign n22938 = n42352 & n22937 ;
  assign n42353 = ~n22938 ;
  assign n22939 = n150 & n42353 ;
  assign n22131 = n21905 & n41925 ;
  assign n42354 = ~n22103 ;
  assign n22132 = n42354 & n22131 ;
  assign n22897 = n22132 & n139 ;
  assign n22133 = n22103 | n22120 ;
  assign n42355 = ~n22133 ;
  assign n22924 = n42355 & n139 ;
  assign n22925 = n21905 | n22924 ;
  assign n42356 = ~n22897 ;
  assign n22926 = n42356 & n22925 ;
  assign n22935 = n150 | n22934 ;
  assign n42357 = ~n22935 ;
  assign n22940 = n42357 & n22937 ;
  assign n22941 = n22926 | n22940 ;
  assign n42358 = ~n22939 ;
  assign n22942 = n42358 & n22941 ;
  assign n42359 = ~n22942 ;
  assign n22943 = n13662 & n42359 ;
  assign n22923 = n42338 & n22919 ;
  assign n22951 = n22923 | n22931 ;
  assign n42360 = ~n22921 ;
  assign n22952 = n42360 & n22951 ;
  assign n42361 = ~n22952 ;
  assign n22953 = n149 & n42361 ;
  assign n22954 = n42351 & n22951 ;
  assign n22955 = n22795 | n22954 ;
  assign n42362 = ~n22953 ;
  assign n22956 = n42362 & n22955 ;
  assign n42363 = ~n22956 ;
  assign n22957 = n150 & n42363 ;
  assign n22958 = n151 | n22957 ;
  assign n42364 = ~n22958 ;
  assign n22959 = n22941 & n42364 ;
  assign n22130 = n22106 | n22122 ;
  assign n42365 = ~n22130 ;
  assign n22891 = n42365 & n139 ;
  assign n22892 = n21967 | n22891 ;
  assign n42366 = ~n22122 ;
  assign n22128 = n21967 & n42366 ;
  assign n22129 = n41952 & n22128 ;
  assign n22968 = n22129 & n139 ;
  assign n42367 = ~n22968 ;
  assign n22969 = n22892 & n42367 ;
  assign n22987 = n22959 | n22969 ;
  assign n42368 = ~n22943 ;
  assign n22988 = n42368 & n22987 ;
  assign n42369 = ~n22988 ;
  assign n22989 = n152 & n42369 ;
  assign n22186 = n41941 & n22151 ;
  assign n42370 = ~n22126 ;
  assign n22187 = n42370 & n22186 ;
  assign n22746 = n22187 & n139 ;
  assign n22127 = n22125 | n22126 ;
  assign n42371 = ~n22127 ;
  assign n22855 = n42371 & n139 ;
  assign n22856 = n22151 | n22855 ;
  assign n42372 = ~n22746 ;
  assign n22857 = n42372 & n22856 ;
  assign n22944 = n152 | n22943 ;
  assign n42373 = ~n22944 ;
  assign n22990 = n42373 & n22987 ;
  assign n22991 = n22857 | n22990 ;
  assign n42374 = ~n22989 ;
  assign n22992 = n42374 & n22991 ;
  assign n42375 = ~n22992 ;
  assign n22993 = n153 & n42375 ;
  assign n22185 = n22163 | n22170 ;
  assign n42376 = ~n22185 ;
  assign n22740 = n42376 & n139 ;
  assign n22741 = n21938 | n22740 ;
  assign n42377 = ~n22170 ;
  assign n22183 = n21938 & n42377 ;
  assign n22184 = n41968 & n22183 ;
  assign n22791 = n22184 & n139 ;
  assign n42378 = ~n22791 ;
  assign n22792 = n22741 & n42378 ;
  assign n22963 = n42357 & n22955 ;
  assign n22964 = n22926 | n22963 ;
  assign n42379 = ~n22957 ;
  assign n22965 = n42379 & n22964 ;
  assign n42380 = ~n22965 ;
  assign n22966 = n151 & n42380 ;
  assign n22967 = n42364 & n22964 ;
  assign n22970 = n22967 | n22969 ;
  assign n42381 = ~n22966 ;
  assign n22971 = n42381 & n22970 ;
  assign n42382 = ~n22971 ;
  assign n22972 = n13079 & n42382 ;
  assign n22973 = n153 | n22972 ;
  assign n42383 = ~n22973 ;
  assign n23005 = n42383 & n22991 ;
  assign n23006 = n22792 | n23005 ;
  assign n42384 = ~n22993 ;
  assign n23007 = n42384 & n23006 ;
  assign n42385 = ~n23007 ;
  assign n23008 = n154 & n42385 ;
  assign n22182 = n22173 | n22174 ;
  assign n42386 = ~n22182 ;
  assign n22751 = n42386 & n139 ;
  assign n22752 = n21883 | n22751 ;
  assign n22160 = n21883 & n41957 ;
  assign n42387 = ~n22174 ;
  assign n22181 = n22160 & n42387 ;
  assign n22796 = n22181 & n139 ;
  assign n42388 = ~n22796 ;
  assign n22797 = n22752 & n42388 ;
  assign n22994 = n154 | n22993 ;
  assign n42389 = ~n22994 ;
  assign n23009 = n42389 & n23006 ;
  assign n23010 = n22797 | n23009 ;
  assign n42390 = ~n23008 ;
  assign n23011 = n42390 & n23010 ;
  assign n42391 = ~n23011 ;
  assign n23012 = n11067 & n42391 ;
  assign n22180 = n22177 | n22179 ;
  assign n42392 = ~n22180 ;
  assign n22742 = n42392 & n139 ;
  assign n22743 = n22189 | n22742 ;
  assign n42393 = ~n22179 ;
  assign n22190 = n42393 & n22189 ;
  assign n22191 = n41984 & n22190 ;
  assign n22744 = n22191 & n139 ;
  assign n42394 = ~n22744 ;
  assign n22745 = n22743 & n42394 ;
  assign n22975 = n42373 & n22970 ;
  assign n22976 = n22857 | n22975 ;
  assign n42395 = ~n22972 ;
  assign n22977 = n42395 & n22976 ;
  assign n42396 = ~n22977 ;
  assign n22978 = n153 & n42396 ;
  assign n22979 = n42383 & n22976 ;
  assign n22980 = n22792 | n22979 ;
  assign n42397 = ~n22978 ;
  assign n22981 = n42397 & n22980 ;
  assign n42398 = ~n22981 ;
  assign n22982 = n154 & n42398 ;
  assign n22983 = n11067 | n22982 ;
  assign n42399 = ~n22983 ;
  assign n23024 = n42399 & n23010 ;
  assign n23025 = n22745 | n23024 ;
  assign n42400 = ~n23012 ;
  assign n23026 = n42400 & n23025 ;
  assign n42401 = ~n23026 ;
  assign n23027 = n156 & n42401 ;
  assign n22218 = n22195 | n22202 ;
  assign n42402 = ~n22218 ;
  assign n22738 = n42402 & n139 ;
  assign n22739 = n22147 | n22738 ;
  assign n22216 = n22147 & n41973 ;
  assign n42403 = ~n22195 ;
  assign n22217 = n42403 & n22216 ;
  assign n22771 = n22217 & n139 ;
  assign n42404 = ~n22771 ;
  assign n22772 = n22739 & n42404 ;
  assign n23013 = n10657 | n23012 ;
  assign n42405 = ~n23013 ;
  assign n23028 = n42405 & n23025 ;
  assign n23029 = n22772 | n23028 ;
  assign n42406 = ~n23027 ;
  assign n23030 = n42406 & n23029 ;
  assign n42407 = ~n23030 ;
  assign n23031 = n157 & n42407 ;
  assign n42408 = ~n22204 ;
  assign n22213 = n21982 & n42408 ;
  assign n22214 = n41997 & n22213 ;
  assign n22726 = n22214 & n139 ;
  assign n22215 = n22198 | n22204 ;
  assign n42409 = ~n22215 ;
  assign n22775 = n42409 & n139 ;
  assign n22776 = n21982 | n22775 ;
  assign n42410 = ~n22726 ;
  assign n22777 = n42410 & n22776 ;
  assign n22995 = n22980 & n42389 ;
  assign n22996 = n22797 | n22995 ;
  assign n42411 = ~n22982 ;
  assign n22997 = n42411 & n22996 ;
  assign n42412 = ~n22997 ;
  assign n22998 = n155 & n42412 ;
  assign n22999 = n42399 & n22996 ;
  assign n23000 = n22745 | n22999 ;
  assign n42413 = ~n22998 ;
  assign n23001 = n42413 & n23000 ;
  assign n42414 = ~n23001 ;
  assign n23002 = n10657 & n42414 ;
  assign n23003 = n157 | n23002 ;
  assign n42415 = ~n23003 ;
  assign n23043 = n42415 & n23029 ;
  assign n23044 = n22777 | n23043 ;
  assign n42416 = ~n23031 ;
  assign n23045 = n42416 & n23044 ;
  assign n42417 = ~n23045 ;
  assign n23046 = n158 & n42417 ;
  assign n22238 = n22208 | n22226 ;
  assign n42418 = ~n22238 ;
  assign n22716 = n42418 & n139 ;
  assign n22717 = n21915 | n22716 ;
  assign n22236 = n21915 & n41989 ;
  assign n42419 = ~n22208 ;
  assign n22237 = n42419 & n22236 ;
  assign n22721 = n22237 & n139 ;
  assign n42420 = ~n22721 ;
  assign n22722 = n22717 & n42420 ;
  assign n23032 = n158 | n23031 ;
  assign n42421 = ~n23032 ;
  assign n23047 = n42421 & n23044 ;
  assign n23048 = n22722 | n23047 ;
  assign n42422 = ~n23046 ;
  assign n23049 = n42422 & n23048 ;
  assign n42423 = ~n23049 ;
  assign n23050 = n8857 & n42423 ;
  assign n42424 = ~n22228 ;
  assign n22233 = n21927 & n42424 ;
  assign n22234 = n42016 & n22233 ;
  assign n22715 = n22234 & n139 ;
  assign n22235 = n22211 | n22228 ;
  assign n42425 = ~n22235 ;
  assign n22753 = n42425 & n139 ;
  assign n22754 = n21927 | n22753 ;
  assign n42426 = ~n22715 ;
  assign n22755 = n42426 & n22754 ;
  assign n23014 = n23000 & n42405 ;
  assign n23015 = n22772 | n23014 ;
  assign n42427 = ~n23002 ;
  assign n23016 = n42427 & n23015 ;
  assign n42428 = ~n23016 ;
  assign n23017 = n157 & n42428 ;
  assign n23018 = n42415 & n23015 ;
  assign n23019 = n22777 | n23018 ;
  assign n42429 = ~n23017 ;
  assign n23020 = n42429 & n23019 ;
  assign n42430 = ~n23020 ;
  assign n23021 = n158 & n42430 ;
  assign n23022 = n8857 | n23021 ;
  assign n42431 = ~n23022 ;
  assign n23062 = n42431 & n23048 ;
  assign n23063 = n22755 | n23062 ;
  assign n42432 = ~n23050 ;
  assign n23064 = n42432 & n23063 ;
  assign n42433 = ~n23064 ;
  assign n23065 = n160 & n42433 ;
  assign n22248 = n22232 | n22246 ;
  assign n42434 = ~n22248 ;
  assign n22713 = n42434 & n139 ;
  assign n22714 = n22253 | n22713 ;
  assign n22254 = n42005 & n22253 ;
  assign n42435 = ~n22232 ;
  assign n22255 = n42435 & n22254 ;
  assign n22786 = n22255 & n139 ;
  assign n42436 = ~n22786 ;
  assign n22787 = n22714 & n42436 ;
  assign n23051 = n160 | n23050 ;
  assign n42437 = ~n23051 ;
  assign n23066 = n42437 & n23063 ;
  assign n23067 = n22787 | n23066 ;
  assign n42438 = ~n23065 ;
  assign n23068 = n42438 & n23067 ;
  assign n42439 = ~n23068 ;
  assign n23069 = n161 & n42439 ;
  assign n22541 = n22267 | n22279 ;
  assign n42440 = ~n22541 ;
  assign n22789 = n42440 & n139 ;
  assign n22790 = n21874 | n22789 ;
  assign n42441 = ~n22279 ;
  assign n22539 = n21874 & n42441 ;
  assign n22540 = n42032 & n22539 ;
  assign n22860 = n22540 & n139 ;
  assign n42442 = ~n22860 ;
  assign n22861 = n22790 & n42442 ;
  assign n23033 = n23019 & n42421 ;
  assign n23034 = n22722 | n23033 ;
  assign n42443 = ~n23021 ;
  assign n23035 = n42443 & n23034 ;
  assign n42444 = ~n23035 ;
  assign n23036 = n159 & n42444 ;
  assign n23037 = n42431 & n23034 ;
  assign n23038 = n22755 | n23037 ;
  assign n42445 = ~n23036 ;
  assign n23039 = n42445 & n23038 ;
  assign n42446 = ~n23039 ;
  assign n23040 = n8534 & n42446 ;
  assign n23041 = n161 | n23040 ;
  assign n42447 = ~n23041 ;
  assign n23081 = n42447 & n23067 ;
  assign n23082 = n22861 | n23081 ;
  assign n42448 = ~n23069 ;
  assign n23083 = n42448 & n23082 ;
  assign n42449 = ~n23083 ;
  assign n23084 = n162 & n42449 ;
  assign n22264 = n21864 & n42021 ;
  assign n42450 = ~n22283 ;
  assign n22537 = n22264 & n42450 ;
  assign n22710 = n22537 & n139 ;
  assign n22538 = n22282 | n22283 ;
  assign n42451 = ~n22538 ;
  assign n22723 = n42451 & n139 ;
  assign n22724 = n21864 | n22723 ;
  assign n42452 = ~n22710 ;
  assign n22725 = n42452 & n22724 ;
  assign n23070 = n162 | n23069 ;
  assign n42453 = ~n23070 ;
  assign n23085 = n42453 & n23082 ;
  assign n23086 = n22725 | n23085 ;
  assign n42454 = ~n23084 ;
  assign n23087 = n42454 & n23086 ;
  assign n42455 = ~n23087 ;
  assign n23088 = n6889 & n42455 ;
  assign n42456 = ~n22298 ;
  assign n22534 = n22034 & n42456 ;
  assign n22535 = n42048 & n22534 ;
  assign n22664 = n22535 & n22661 ;
  assign n22536 = n22286 | n22298 ;
  assign n42457 = ~n22536 ;
  assign n22748 = n42457 & n139 ;
  assign n22749 = n22034 | n22748 ;
  assign n42458 = ~n22664 ;
  assign n22750 = n42458 & n22749 ;
  assign n23052 = n23038 & n42437 ;
  assign n23053 = n22787 | n23052 ;
  assign n42459 = ~n23040 ;
  assign n23054 = n42459 & n23053 ;
  assign n42460 = ~n23054 ;
  assign n23055 = n161 & n42460 ;
  assign n23056 = n42447 & n23053 ;
  assign n23057 = n22861 | n23056 ;
  assign n42461 = ~n23055 ;
  assign n23058 = n42461 & n23057 ;
  assign n42462 = ~n23058 ;
  assign n23059 = n162 & n42462 ;
  assign n23060 = n6889 | n23059 ;
  assign n42463 = ~n23060 ;
  assign n23100 = n42463 & n23086 ;
  assign n23101 = n22750 | n23100 ;
  assign n42464 = ~n23088 ;
  assign n23102 = n42464 & n23101 ;
  assign n42465 = ~n23102 ;
  assign n23103 = n164 & n42465 ;
  assign n22278 = n21850 & n42037 ;
  assign n42466 = ~n22302 ;
  assign n22532 = n22278 & n42466 ;
  assign n22706 = n22532 & n139 ;
  assign n22533 = n22276 | n22302 ;
  assign n42467 = ~n22533 ;
  assign n22765 = n42467 & n139 ;
  assign n22766 = n21850 | n22765 ;
  assign n42468 = ~n22706 ;
  assign n22767 = n42468 & n22766 ;
  assign n23089 = n6600 | n23088 ;
  assign n42469 = ~n23089 ;
  assign n23104 = n42469 & n23101 ;
  assign n23105 = n22767 | n23104 ;
  assign n42470 = ~n23103 ;
  assign n23106 = n42470 & n23105 ;
  assign n42471 = ~n23106 ;
  assign n23107 = n165 & n42471 ;
  assign n22531 = n22305 | n22317 ;
  assign n42472 = ~n22531 ;
  assign n22701 = n42472 & n139 ;
  assign n22702 = n21980 | n22701 ;
  assign n42473 = ~n22317 ;
  assign n22529 = n21980 & n42473 ;
  assign n22530 = n42064 & n22529 ;
  assign n22769 = n22530 & n139 ;
  assign n42474 = ~n22769 ;
  assign n22770 = n22702 & n42474 ;
  assign n23071 = n23057 & n42453 ;
  assign n23072 = n22725 | n23071 ;
  assign n42475 = ~n23059 ;
  assign n23073 = n42475 & n23072 ;
  assign n42476 = ~n23073 ;
  assign n23074 = n163 & n42476 ;
  assign n23075 = n42463 & n23072 ;
  assign n23076 = n22750 | n23075 ;
  assign n42477 = ~n23074 ;
  assign n23077 = n42477 & n23076 ;
  assign n42478 = ~n23077 ;
  assign n23078 = n6600 & n42478 ;
  assign n23079 = n165 | n23078 ;
  assign n42479 = ~n23079 ;
  assign n23119 = n42479 & n23105 ;
  assign n23120 = n22770 | n23119 ;
  assign n42480 = ~n23107 ;
  assign n23121 = n42480 & n23120 ;
  assign n42481 = ~n23121 ;
  assign n23122 = n166 & n42481 ;
  assign n22297 = n21965 & n42053 ;
  assign n42482 = ~n22321 ;
  assign n22322 = n22297 & n42482 ;
  assign n22705 = n22322 & n139 ;
  assign n22323 = n22295 | n22321 ;
  assign n42483 = ~n22323 ;
  assign n22729 = n42483 & n139 ;
  assign n22730 = n21965 | n22729 ;
  assign n42484 = ~n22705 ;
  assign n22731 = n42484 & n22730 ;
  assign n23108 = n166 | n23107 ;
  assign n42485 = ~n23108 ;
  assign n23123 = n42485 & n23120 ;
  assign n23124 = n22731 | n23123 ;
  assign n42486 = ~n23122 ;
  assign n23125 = n42486 & n23124 ;
  assign n42487 = ~n23125 ;
  assign n23126 = n5352 & n42487 ;
  assign n42488 = ~n22338 ;
  assign n22526 = n21970 & n42488 ;
  assign n22527 = n42080 & n22526 ;
  assign n22698 = n22527 & n139 ;
  assign n22528 = n22326 | n22338 ;
  assign n42489 = ~n22528 ;
  assign n22760 = n42489 & n139 ;
  assign n22761 = n21970 | n22760 ;
  assign n42490 = ~n22698 ;
  assign n22762 = n42490 & n22761 ;
  assign n23090 = n23076 & n42469 ;
  assign n23091 = n22767 | n23090 ;
  assign n42491 = ~n23078 ;
  assign n23092 = n42491 & n23091 ;
  assign n42492 = ~n23092 ;
  assign n23093 = n165 & n42492 ;
  assign n23094 = n42479 & n23091 ;
  assign n23095 = n22770 | n23094 ;
  assign n42493 = ~n23093 ;
  assign n23096 = n42493 & n23095 ;
  assign n42494 = ~n23096 ;
  assign n23097 = n166 & n42494 ;
  assign n23098 = n5352 | n23097 ;
  assign n42495 = ~n23098 ;
  assign n23133 = n42495 & n23124 ;
  assign n23134 = n22762 | n23133 ;
  assign n42496 = ~n23126 ;
  assign n23135 = n42496 & n23134 ;
  assign n42497 = ~n23135 ;
  assign n23136 = n168 & n42497 ;
  assign n22525 = n22314 | n22342 ;
  assign n42498 = ~n22525 ;
  assign n22694 = n42498 & n139 ;
  assign n22695 = n22149 | n22694 ;
  assign n22316 = n22149 & n42069 ;
  assign n42499 = ~n22342 ;
  assign n22524 = n22316 & n42499 ;
  assign n22696 = n22524 & n139 ;
  assign n42500 = ~n22696 ;
  assign n22697 = n22695 & n42500 ;
  assign n23127 = n4934 | n23126 ;
  assign n42501 = ~n23127 ;
  assign n23137 = n42501 & n23134 ;
  assign n23138 = n22697 | n23137 ;
  assign n42502 = ~n23136 ;
  assign n23139 = n42502 & n23138 ;
  assign n42503 = ~n23139 ;
  assign n23140 = n169 & n42503 ;
  assign n23109 = n23095 & n42485 ;
  assign n23110 = n22731 | n23109 ;
  assign n42504 = ~n23097 ;
  assign n23111 = n42504 & n23110 ;
  assign n42505 = ~n23111 ;
  assign n23112 = n167 & n42505 ;
  assign n23113 = n42495 & n23110 ;
  assign n23114 = n22762 | n23113 ;
  assign n42506 = ~n23112 ;
  assign n23115 = n42506 & n23114 ;
  assign n42507 = ~n23115 ;
  assign n23116 = n4934 & n42507 ;
  assign n23117 = n169 | n23116 ;
  assign n42508 = ~n23117 ;
  assign n23142 = n42508 & n23138 ;
  assign n42509 = ~n22357 ;
  assign n22521 = n21832 & n42509 ;
  assign n22522 = n42096 & n22521 ;
  assign n22693 = n22522 & n139 ;
  assign n22523 = n22345 | n22357 ;
  assign n42510 = ~n22523 ;
  assign n23188 = n42510 & n139 ;
  assign n23189 = n21832 | n23188 ;
  assign n42511 = ~n22693 ;
  assign n23190 = n42511 & n23189 ;
  assign n23198 = n23142 | n23190 ;
  assign n42512 = ~n23140 ;
  assign n23199 = n42512 & n23198 ;
  assign n42513 = ~n23199 ;
  assign n23200 = n170 & n42513 ;
  assign n23141 = n170 | n23140 ;
  assign n42514 = ~n23141 ;
  assign n23201 = n42514 & n23198 ;
  assign n22337 = n21853 & n42085 ;
  assign n42515 = ~n22361 ;
  assign n22519 = n22337 & n42515 ;
  assign n22709 = n22519 & n139 ;
  assign n22520 = n22360 | n22361 ;
  assign n42516 = ~n22520 ;
  assign n23205 = n42516 & n139 ;
  assign n23206 = n21853 | n23205 ;
  assign n42517 = ~n22709 ;
  assign n23207 = n42517 & n23206 ;
  assign n23208 = n23201 | n23207 ;
  assign n42518 = ~n23200 ;
  assign n23209 = n42518 & n23208 ;
  assign n42519 = ~n23209 ;
  assign n23210 = n3940 & n42519 ;
  assign n42520 = ~n22376 ;
  assign n22517 = n22251 & n42520 ;
  assign n22518 = n42112 & n22517 ;
  assign n22747 = n22518 & n139 ;
  assign n22516 = n22364 | n22376 ;
  assign n42521 = ~n22516 ;
  assign n22894 = n42521 & n139 ;
  assign n22895 = n22251 | n22894 ;
  assign n42522 = ~n22747 ;
  assign n22896 = n42522 & n22895 ;
  assign n23128 = n23114 & n42501 ;
  assign n23129 = n22697 | n23128 ;
  assign n42523 = ~n23116 ;
  assign n23130 = n42523 & n23129 ;
  assign n42524 = ~n23130 ;
  assign n23131 = n169 & n42524 ;
  assign n23132 = n42508 & n23129 ;
  assign n23191 = n23132 | n23190 ;
  assign n42525 = ~n23131 ;
  assign n23192 = n42525 & n23191 ;
  assign n42526 = ~n23192 ;
  assign n23193 = n170 & n42526 ;
  assign n23194 = n3940 | n23193 ;
  assign n42527 = ~n23194 ;
  assign n23212 = n42527 & n23208 ;
  assign n23213 = n22896 | n23212 ;
  assign n42528 = ~n23210 ;
  assign n23214 = n42528 & n23213 ;
  assign n42529 = ~n23214 ;
  assign n23215 = n172 & n42529 ;
  assign n23211 = n3631 | n23210 ;
  assign n42530 = ~n23211 ;
  assign n23216 = n42530 & n23213 ;
  assign n22356 = n22036 & n42101 ;
  assign n42531 = ~n22380 ;
  assign n22514 = n22356 & n42531 ;
  assign n23232 = n22514 & n139 ;
  assign n22515 = n22354 | n22380 ;
  assign n42532 = ~n22515 ;
  assign n23233 = n42532 & n139 ;
  assign n23234 = n22036 | n23233 ;
  assign n42533 = ~n23232 ;
  assign n23235 = n42533 & n23234 ;
  assign n23236 = n23216 | n23235 ;
  assign n42534 = ~n23215 ;
  assign n23237 = n42534 & n23236 ;
  assign n42535 = ~n23237 ;
  assign n23238 = n173 & n42535 ;
  assign n23195 = n42514 & n23191 ;
  assign n23223 = n23195 | n23207 ;
  assign n42536 = ~n23193 ;
  assign n23224 = n42536 & n23223 ;
  assign n42537 = ~n23224 ;
  assign n23225 = n171 & n42537 ;
  assign n23226 = n42527 & n23223 ;
  assign n23227 = n22896 | n23226 ;
  assign n42538 = ~n23225 ;
  assign n23228 = n42538 & n23227 ;
  assign n42539 = ~n23228 ;
  assign n23229 = n3631 & n42539 ;
  assign n23230 = n173 | n23229 ;
  assign n42540 = ~n23230 ;
  assign n23240 = n42540 & n23236 ;
  assign n42541 = ~n22395 ;
  assign n22511 = n21846 & n42541 ;
  assign n22512 = n42128 & n22511 ;
  assign n22663 = n22512 & n22661 ;
  assign n22513 = n22383 | n22395 ;
  assign n42542 = ~n22513 ;
  assign n23248 = n42542 & n139 ;
  assign n23249 = n21846 | n23248 ;
  assign n42543 = ~n22663 ;
  assign n23250 = n42543 & n23249 ;
  assign n23253 = n23240 | n23250 ;
  assign n42544 = ~n23238 ;
  assign n23254 = n42544 & n23253 ;
  assign n42545 = ~n23254 ;
  assign n23255 = n174 & n42545 ;
  assign n23239 = n174 | n23238 ;
  assign n42546 = ~n23239 ;
  assign n23256 = n42546 & n23253 ;
  assign n22510 = n22373 | n22399 ;
  assign n42547 = ~n22510 ;
  assign n22756 = n42547 & n139 ;
  assign n22757 = n21894 | n22756 ;
  assign n22375 = n21894 & n42117 ;
  assign n42548 = ~n22399 ;
  assign n22509 = n22375 & n42548 ;
  assign n23263 = n22509 & n139 ;
  assign n42549 = ~n23263 ;
  assign n23264 = n22757 & n42549 ;
  assign n23265 = n23256 | n23264 ;
  assign n42550 = ~n23255 ;
  assign n23266 = n42550 & n23265 ;
  assign n42551 = ~n23266 ;
  assign n23267 = n2753 & n42551 ;
  assign n22508 = n22402 | n22414 ;
  assign n42552 = ~n22508 ;
  assign n22927 = n42552 & n139 ;
  assign n22928 = n21838 | n22927 ;
  assign n42553 = ~n22414 ;
  assign n22506 = n21838 & n42553 ;
  assign n22507 = n42144 & n22506 ;
  assign n23203 = n22507 & n139 ;
  assign n42554 = ~n23203 ;
  assign n23204 = n22928 & n42554 ;
  assign n23231 = n42530 & n23227 ;
  assign n23244 = n23231 | n23235 ;
  assign n42555 = ~n23229 ;
  assign n23245 = n42555 & n23244 ;
  assign n42556 = ~n23245 ;
  assign n23246 = n173 & n42556 ;
  assign n23247 = n42540 & n23244 ;
  assign n23258 = n23247 | n23250 ;
  assign n42557 = ~n23246 ;
  assign n23259 = n42557 & n23258 ;
  assign n42558 = ~n23259 ;
  assign n23260 = n174 & n42558 ;
  assign n23261 = n2753 | n23260 ;
  assign n42559 = ~n23261 ;
  assign n23269 = n42559 & n23265 ;
  assign n23270 = n23204 | n23269 ;
  assign n42560 = ~n23267 ;
  assign n23271 = n42560 & n23270 ;
  assign n42561 = ~n23271 ;
  assign n23272 = n176 & n42561 ;
  assign n23268 = n2431 | n23267 ;
  assign n42562 = ~n23268 ;
  assign n23273 = n42562 & n23270 ;
  assign n22394 = n21990 & n42133 ;
  assign n42563 = ~n22418 ;
  assign n22504 = n22394 & n42563 ;
  assign n23289 = n22504 & n139 ;
  assign n22505 = n22392 | n22418 ;
  assign n42564 = ~n22505 ;
  assign n23292 = n42564 & n139 ;
  assign n23293 = n21990 | n23292 ;
  assign n42565 = ~n23289 ;
  assign n23294 = n42565 & n23293 ;
  assign n23295 = n23273 | n23294 ;
  assign n42566 = ~n23272 ;
  assign n23296 = n42566 & n23295 ;
  assign n42567 = ~n23296 ;
  assign n23297 = n177 & n42567 ;
  assign n23262 = n42546 & n23258 ;
  assign n23280 = n23262 | n23264 ;
  assign n42568 = ~n23260 ;
  assign n23281 = n42568 & n23280 ;
  assign n42569 = ~n23281 ;
  assign n23282 = n175 & n42569 ;
  assign n23283 = n42559 & n23280 ;
  assign n23284 = n23204 | n23283 ;
  assign n42570 = ~n23282 ;
  assign n23285 = n42570 & n23284 ;
  assign n42571 = ~n23285 ;
  assign n23286 = n2431 & n42571 ;
  assign n23287 = n177 | n23286 ;
  assign n42572 = ~n23287 ;
  assign n23299 = n42572 & n23295 ;
  assign n22501 = n22421 | n22433 ;
  assign n42573 = ~n22501 ;
  assign n22763 = n42573 & n139 ;
  assign n22764 = n21993 | n22763 ;
  assign n42574 = ~n22433 ;
  assign n22502 = n21993 & n42574 ;
  assign n22503 = n42160 & n22502 ;
  assign n23307 = n22503 & n139 ;
  assign n42575 = ~n23307 ;
  assign n23308 = n22764 & n42575 ;
  assign n23316 = n23299 | n23308 ;
  assign n42576 = ~n23297 ;
  assign n23317 = n42576 & n23316 ;
  assign n42577 = ~n23317 ;
  assign n23318 = n178 & n42577 ;
  assign n23298 = n178 | n23297 ;
  assign n42578 = ~n23298 ;
  assign n23319 = n42578 & n23316 ;
  assign n22413 = n21997 & n42149 ;
  assign n42579 = ~n22437 ;
  assign n22499 = n22413 & n42579 ;
  assign n23322 = n22499 & n139 ;
  assign n22500 = n22436 | n22437 ;
  assign n42580 = ~n22500 ;
  assign n23323 = n42580 & n139 ;
  assign n23324 = n21997 | n23323 ;
  assign n42581 = ~n23322 ;
  assign n23325 = n42581 & n23324 ;
  assign n23326 = n23319 | n23325 ;
  assign n42582 = ~n23318 ;
  assign n23327 = n42582 & n23326 ;
  assign n42583 = ~n23327 ;
  assign n23328 = n1707 & n42583 ;
  assign n23288 = n42562 & n23284 ;
  assign n23303 = n23288 | n23294 ;
  assign n42584 = ~n23286 ;
  assign n23304 = n42584 & n23303 ;
  assign n42585 = ~n23304 ;
  assign n23305 = n177 & n42585 ;
  assign n23306 = n42572 & n23303 ;
  assign n23309 = n23306 | n23308 ;
  assign n42586 = ~n23305 ;
  assign n23310 = n42586 & n23309 ;
  assign n42587 = ~n23310 ;
  assign n23311 = n178 & n42587 ;
  assign n23312 = n1707 | n23311 ;
  assign n42588 = ~n23312 ;
  assign n23330 = n42588 & n23326 ;
  assign n42589 = ~n22452 ;
  assign n22496 = n21984 & n42589 ;
  assign n22497 = n42176 & n22496 ;
  assign n23338 = n22497 & n139 ;
  assign n22498 = n22440 | n22452 ;
  assign n42590 = ~n22498 ;
  assign n23339 = n42590 & n139 ;
  assign n23340 = n21984 | n23339 ;
  assign n42591 = ~n23338 ;
  assign n23341 = n42591 & n23340 ;
  assign n23349 = n23330 | n23341 ;
  assign n42592 = ~n23328 ;
  assign n23350 = n42592 & n23349 ;
  assign n42593 = ~n23350 ;
  assign n23351 = n180 & n42593 ;
  assign n23329 = n1487 | n23328 ;
  assign n42594 = ~n23329 ;
  assign n23352 = n42594 & n23349 ;
  assign n22495 = n22455 | n22456 ;
  assign n42595 = ~n22495 ;
  assign n23290 = n42595 & n139 ;
  assign n23291 = n22032 | n23290 ;
  assign n22432 = n22032 & n42165 ;
  assign n42596 = ~n22456 ;
  assign n22494 = n22432 & n42596 ;
  assign n23354 = n22494 & n139 ;
  assign n42597 = ~n23354 ;
  assign n23355 = n23291 & n42597 ;
  assign n23356 = n23352 | n23355 ;
  assign n42598 = ~n23351 ;
  assign n23357 = n42598 & n23356 ;
  assign n42599 = ~n23357 ;
  assign n23358 = n181 & n42599 ;
  assign n23313 = n42578 & n23309 ;
  assign n23334 = n23313 | n23325 ;
  assign n42600 = ~n23311 ;
  assign n23335 = n42600 & n23334 ;
  assign n42601 = ~n23335 ;
  assign n23336 = n179 & n42601 ;
  assign n23337 = n42588 & n23334 ;
  assign n23342 = n23337 | n23341 ;
  assign n42602 = ~n23336 ;
  assign n23343 = n42602 & n23342 ;
  assign n42603 = ~n23343 ;
  assign n23344 = n1487 & n42603 ;
  assign n23345 = n181 | n23344 ;
  assign n42604 = ~n23345 ;
  assign n23360 = n42604 & n23356 ;
  assign n22493 = n22459 | n22470 ;
  assign n42605 = ~n22493 ;
  assign n22699 = n42605 & n139 ;
  assign n22700 = n21999 | n22699 ;
  assign n42606 = ~n22470 ;
  assign n22491 = n21999 & n42606 ;
  assign n22492 = n42189 & n22491 ;
  assign n23368 = n22492 & n139 ;
  assign n42607 = ~n23368 ;
  assign n23369 = n22700 & n42607 ;
  assign n23377 = n23360 | n23369 ;
  assign n42608 = ~n23358 ;
  assign n23378 = n42608 & n23377 ;
  assign n42609 = ~n23378 ;
  assign n23379 = n182 & n42609 ;
  assign n23359 = n182 | n23358 ;
  assign n42610 = ~n23359 ;
  assign n23380 = n42610 & n23377 ;
  assign n22451 = n22005 & n42181 ;
  assign n42611 = ~n22474 ;
  assign n22489 = n22451 & n42611 ;
  assign n22817 = n22489 & n139 ;
  assign n22490 = n22473 | n22474 ;
  assign n42612 = ~n22490 ;
  assign n23382 = n42612 & n139 ;
  assign n23383 = n22005 | n23382 ;
  assign n42613 = ~n22817 ;
  assign n23384 = n42613 & n23383 ;
  assign n23385 = n23380 | n23384 ;
  assign n42614 = ~n23379 ;
  assign n23386 = n42614 & n23385 ;
  assign n42615 = ~n23386 ;
  assign n23387 = n996 & n42615 ;
  assign n23346 = n42594 & n23342 ;
  assign n23364 = n23346 | n23355 ;
  assign n42616 = ~n23344 ;
  assign n23365 = n42616 & n23364 ;
  assign n42617 = ~n23365 ;
  assign n23366 = n181 & n42617 ;
  assign n23367 = n42604 & n23364 ;
  assign n23370 = n23367 | n23369 ;
  assign n42618 = ~n23366 ;
  assign n23371 = n42618 & n23370 ;
  assign n42619 = ~n23371 ;
  assign n23372 = n182 & n42619 ;
  assign n23373 = n183 | n23372 ;
  assign n42620 = ~n23373 ;
  assign n23389 = n42620 & n23385 ;
  assign n22488 = n22477 | n22480 ;
  assign n42621 = ~n22488 ;
  assign n22818 = n42621 & n139 ;
  assign n22819 = n21987 | n22818 ;
  assign n42622 = ~n22480 ;
  assign n22486 = n21987 & n42622 ;
  assign n22487 = n42208 & n22486 ;
  assign n23397 = n22487 & n139 ;
  assign n42623 = ~n23397 ;
  assign n23398 = n22819 & n42623 ;
  assign n23406 = n23389 | n23398 ;
  assign n42624 = ~n23387 ;
  assign n23407 = n42624 & n23406 ;
  assign n42625 = ~n23407 ;
  assign n23408 = n184 & n42625 ;
  assign n23388 = n838 | n23387 ;
  assign n42626 = ~n23388 ;
  assign n23409 = n42626 & n23406 ;
  assign n22544 = n42197 & n22543 ;
  assign n42627 = ~n22484 ;
  assign n22545 = n42627 & n22544 ;
  assign n22798 = n22545 & n139 ;
  assign n22485 = n22468 | n22484 ;
  assign n42628 = ~n22485 ;
  assign n23411 = n42628 & n139 ;
  assign n23412 = n22543 | n23411 ;
  assign n42629 = ~n22798 ;
  assign n23413 = n42629 & n23412 ;
  assign n23414 = n23409 | n23413 ;
  assign n42630 = ~n23408 ;
  assign n23415 = n42630 & n23414 ;
  assign n42631 = ~n23415 ;
  assign n23416 = n185 & n42631 ;
  assign n23374 = n42610 & n23370 ;
  assign n23393 = n23374 | n23384 ;
  assign n42632 = ~n23372 ;
  assign n23394 = n42632 & n23393 ;
  assign n42633 = ~n23394 ;
  assign n23395 = n183 & n42633 ;
  assign n23396 = n42620 & n23393 ;
  assign n23399 = n23396 | n23398 ;
  assign n42634 = ~n23395 ;
  assign n23400 = n42634 & n23399 ;
  assign n42635 = ~n23400 ;
  assign n23401 = n838 & n42635 ;
  assign n23402 = n185 | n23401 ;
  assign n42636 = ~n23402 ;
  assign n23418 = n42636 & n23414 ;
  assign n42637 = ~n22569 ;
  assign n22601 = n22009 & n42637 ;
  assign n22602 = n42224 & n22601 ;
  assign n23321 = n22602 & n139 ;
  assign n22603 = n22557 | n22569 ;
  assign n42638 = ~n22603 ;
  assign n23426 = n42638 & n139 ;
  assign n23427 = n22009 | n23426 ;
  assign n42639 = ~n23321 ;
  assign n23428 = n42639 & n23427 ;
  assign n23445 = n23418 | n23428 ;
  assign n42640 = ~n23416 ;
  assign n23446 = n42640 & n23445 ;
  assign n42641 = ~n23446 ;
  assign n23447 = n186 & n42641 ;
  assign n22600 = n22572 | n22573 ;
  assign n42642 = ~n22600 ;
  assign n22711 = n42642 & n139 ;
  assign n22712 = n22011 | n22711 ;
  assign n22554 = n22011 & n42213 ;
  assign n42643 = ~n22573 ;
  assign n22599 = n22554 & n42643 ;
  assign n22773 = n22599 & n139 ;
  assign n42644 = ~n22773 ;
  assign n22774 = n22712 & n42644 ;
  assign n23417 = n186 | n23416 ;
  assign n42645 = ~n23417 ;
  assign n23448 = n42645 & n23445 ;
  assign n23449 = n22774 | n23448 ;
  assign n42646 = ~n23447 ;
  assign n23450 = n42646 & n23449 ;
  assign n42647 = ~n23450 ;
  assign n23451 = n528 & n42647 ;
  assign n22598 = n22576 | n22583 ;
  assign n42648 = ~n22598 ;
  assign n22703 = n42648 & n139 ;
  assign n22704 = n22017 | n22703 ;
  assign n42649 = ~n22583 ;
  assign n22596 = n22017 & n42649 ;
  assign n22597 = n42240 & n22596 ;
  assign n22718 = n22597 & n139 ;
  assign n42650 = ~n22718 ;
  assign n22719 = n22704 & n42650 ;
  assign n23403 = n42626 & n23399 ;
  assign n23422 = n23403 | n23413 ;
  assign n42651 = ~n23401 ;
  assign n23423 = n42651 & n23422 ;
  assign n42652 = ~n23423 ;
  assign n23424 = n185 & n42652 ;
  assign n23425 = n42636 & n23422 ;
  assign n23429 = n23425 | n23428 ;
  assign n42653 = ~n23424 ;
  assign n23430 = n42653 & n23429 ;
  assign n42654 = ~n23430 ;
  assign n23431 = n186 & n42654 ;
  assign n23432 = n528 | n23431 ;
  assign n42655 = ~n23432 ;
  assign n23454 = n42655 & n23449 ;
  assign n23455 = n22719 | n23454 ;
  assign n42656 = ~n23451 ;
  assign n23456 = n42656 & n23455 ;
  assign n42657 = ~n23456 ;
  assign n23457 = n188 & n42657 ;
  assign n23452 = n413 | n23451 ;
  assign n42658 = ~n23452 ;
  assign n23458 = n42658 & n23455 ;
  assign n22568 = n22019 & n42229 ;
  assign n42659 = ~n22587 ;
  assign n22594 = n22568 & n42659 ;
  assign n22720 = n22594 & n139 ;
  assign n22595 = n22586 | n22587 ;
  assign n42660 = ~n22595 ;
  assign n23469 = n42660 & n139 ;
  assign n23470 = n22019 | n23469 ;
  assign n42661 = ~n22720 ;
  assign n23471 = n42661 & n23470 ;
  assign n23472 = n23458 | n23471 ;
  assign n42662 = ~n23457 ;
  assign n23473 = n42662 & n23472 ;
  assign n42663 = ~n23473 ;
  assign n23474 = n189 & n42663 ;
  assign n23434 = n42645 & n23429 ;
  assign n23435 = n22774 | n23434 ;
  assign n42664 = ~n23431 ;
  assign n23436 = n42664 & n23435 ;
  assign n42665 = ~n23436 ;
  assign n23437 = n187 & n42665 ;
  assign n23438 = n42655 & n23435 ;
  assign n23439 = n22719 | n23438 ;
  assign n42666 = ~n23437 ;
  assign n23440 = n42666 & n23439 ;
  assign n42667 = ~n23440 ;
  assign n23441 = n413 & n42667 ;
  assign n23442 = n189 | n23441 ;
  assign n42668 = ~n23442 ;
  assign n23476 = n42668 & n23472 ;
  assign n42669 = ~n22592 ;
  assign n22640 = n42669 & n22624 ;
  assign n22641 = n42256 & n22640 ;
  assign n22662 = n22641 & n22661 ;
  assign n22593 = n22590 | n22592 ;
  assign n42670 = ~n22593 ;
  assign n23484 = n42670 & n139 ;
  assign n23508 = n22624 | n23484 ;
  assign n42671 = ~n22662 ;
  assign n23509 = n42671 & n23508 ;
  assign n23512 = n23476 | n23509 ;
  assign n42672 = ~n23474 ;
  assign n23513 = n42672 & n23512 ;
  assign n42673 = ~n23513 ;
  assign n23514 = n190 & n42673 ;
  assign n22629 = n22021 & n42245 ;
  assign n42674 = ~n22645 ;
  assign n23502 = n22629 & n42674 ;
  assign n23503 = n139 & n23502 ;
  assign n23504 = n22644 | n22645 ;
  assign n42675 = ~n23504 ;
  assign n23505 = n139 & n42675 ;
  assign n23506 = n22021 | n23505 ;
  assign n42676 = ~n23503 ;
  assign n23507 = n42676 & n23506 ;
  assign n23475 = n190 | n23474 ;
  assign n42677 = ~n23475 ;
  assign n23515 = n42677 & n23512 ;
  assign n23516 = n23507 | n23515 ;
  assign n42678 = ~n23514 ;
  assign n23517 = n42678 & n23516 ;
  assign n42679 = ~n23517 ;
  assign n23518 = n287 & n42679 ;
  assign n42680 = ~n22681 ;
  assign n23495 = n22622 & n42680 ;
  assign n23496 = n42267 & n23495 ;
  assign n23497 = n139 & n23496 ;
  assign n23498 = n22648 | n22681 ;
  assign n42681 = ~n23498 ;
  assign n23499 = n139 & n42681 ;
  assign n23500 = n22622 | n23499 ;
  assign n42682 = ~n23497 ;
  assign n23501 = n42682 & n23500 ;
  assign n23453 = n23439 & n42658 ;
  assign n23480 = n23453 | n23471 ;
  assign n42683 = ~n23441 ;
  assign n23481 = n42683 & n23480 ;
  assign n42684 = ~n23481 ;
  assign n23482 = n189 & n42684 ;
  assign n23483 = n42668 & n23480 ;
  assign n23521 = n23483 | n23509 ;
  assign n42685 = ~n23482 ;
  assign n23522 = n42685 & n23521 ;
  assign n42686 = ~n23522 ;
  assign n23523 = n190 & n42686 ;
  assign n23524 = n287 | n23523 ;
  assign n42687 = ~n23524 ;
  assign n23525 = n23516 & n42687 ;
  assign n23529 = n23501 | n23525 ;
  assign n42688 = ~n23518 ;
  assign n23530 = n42688 & n23529 ;
  assign n23531 = n23487 | n23530 ;
  assign n23532 = n31336 & n23531 ;
  assign n22607 = n21819 | n22606 ;
  assign n42689 = ~n22607 ;
  assign n22613 = n42689 & n22610 ;
  assign n22614 = n42275 & n22613 ;
  assign n22677 = n22614 & n42276 ;
  assign n22678 = n42277 & n22677 ;
  assign n22671 = n192 & n22670 ;
  assign n42690 = ~n22611 ;
  assign n23488 = n42690 & n139 ;
  assign n42691 = ~n23488 ;
  assign n23489 = n22656 & n42691 ;
  assign n42692 = ~n23489 ;
  assign n23490 = n22671 & n42692 ;
  assign n23491 = n22678 | n23490 ;
  assign n23519 = n23466 & n42688 ;
  assign n23535 = n23519 & n23529 ;
  assign n23544 = n23491 | n23535 ;
  assign n138 = n23532 | n23544 ;
  assign n248 = x14 | x15 ;
  assign n249 = x16 | n248 ;
  assign n42693 = ~n23525 ;
  assign n23526 = n23501 & n42693 ;
  assign n23527 = n42688 & n23526 ;
  assign n23753 = n23527 & n138 ;
  assign n23528 = n23518 | n23525 ;
  assign n42694 = ~n23528 ;
  assign n23755 = n42694 & n138 ;
  assign n23756 = n23501 | n23755 ;
  assign n42695 = ~n23753 ;
  assign n23757 = n42695 & n23756 ;
  assign n23533 = n23466 | n23530 ;
  assign n42696 = ~n23533 ;
  assign n23765 = n42696 & n138 ;
  assign n23766 = n23535 | n23765 ;
  assign n23767 = n23757 | n23766 ;
  assign n42697 = ~n22678 ;
  assign n22679 = n22661 & n42697 ;
  assign n42698 = ~n23490 ;
  assign n23492 = n22679 & n42698 ;
  assign n42699 = ~n23535 ;
  assign n23536 = n23492 & n42699 ;
  assign n42700 = ~n23532 ;
  assign n23537 = n42700 & n23536 ;
  assign n42701 = ~n242 ;
  assign n23613 = n42701 & n138 ;
  assign n23614 = n23537 | n23613 ;
  assign n23615 = x20 & n23614 ;
  assign n23538 = x20 | n23537 ;
  assign n23616 = n23538 | n23613 ;
  assign n42702 = ~n23615 ;
  assign n23617 = n42702 & n23616 ;
  assign n245 = x16 | x17 ;
  assign n42703 = ~x18 ;
  assign n247 = n42703 & n245 ;
  assign n42704 = ~n138 ;
  assign n23775 = x18 & n42704 ;
  assign n23776 = n247 | n23775 ;
  assign n42705 = ~n23776 ;
  assign n23777 = n22661 & n42705 ;
  assign n23778 = n22030 | n23777 ;
  assign n246 = x18 | n245 ;
  assign n21820 = n246 & n42274 ;
  assign n22027 = n21820 & n42275 ;
  assign n22675 = n22027 & n42276 ;
  assign n22676 = n42277 & n22675 ;
  assign n23645 = x18 & n138 ;
  assign n42706 = ~n23645 ;
  assign n23774 = n22676 & n42706 ;
  assign n23780 = n42703 & n138 ;
  assign n42707 = ~n23780 ;
  assign n23781 = x19 & n42707 ;
  assign n23782 = n23613 | n23781 ;
  assign n23783 = n23774 | n23782 ;
  assign n42708 = ~n23778 ;
  assign n23784 = n42708 & n23783 ;
  assign n23785 = n23617 | n23784 ;
  assign n23646 = n246 & n42706 ;
  assign n42709 = ~n23646 ;
  assign n23647 = n139 & n42709 ;
  assign n42710 = ~n23647 ;
  assign n23788 = n42710 & n23783 ;
  assign n42711 = ~n23788 ;
  assign n23789 = n22030 & n42711 ;
  assign n42712 = ~n23789 ;
  assign n23790 = n23785 & n42712 ;
  assign n42713 = ~n23790 ;
  assign n23791 = n141 & n42713 ;
  assign n22805 = n22669 | n22800 ;
  assign n42714 = ~n22805 ;
  assign n23623 = n42714 & n138 ;
  assign n23624 = n22733 | n23623 ;
  assign n22806 = n22733 & n42714 ;
  assign n23772 = n22806 & n138 ;
  assign n42715 = ~n23772 ;
  assign n23773 = n23624 & n42715 ;
  assign n23796 = n141 | n23789 ;
  assign n42716 = ~n23796 ;
  assign n23797 = n23785 & n42716 ;
  assign n23798 = n23773 | n23797 ;
  assign n42717 = ~n23791 ;
  assign n23799 = n42717 & n23798 ;
  assign n42718 = ~n23799 ;
  assign n23800 = n142 & n42718 ;
  assign n42719 = ~n22807 ;
  assign n22810 = n22737 & n42719 ;
  assign n42720 = ~n22812 ;
  assign n22815 = n22810 & n42720 ;
  assign n23596 = n22815 & n138 ;
  assign n22816 = n22807 | n22812 ;
  assign n42721 = ~n22816 ;
  assign n23605 = n42721 & n138 ;
  assign n23606 = n22737 | n23605 ;
  assign n42722 = ~n23596 ;
  assign n23607 = n42722 & n23606 ;
  assign n23792 = n142 | n23791 ;
  assign n42723 = ~n23792 ;
  assign n23801 = n42723 & n23798 ;
  assign n23802 = n23607 | n23801 ;
  assign n42724 = ~n23800 ;
  assign n23803 = n42724 & n23802 ;
  assign n42725 = ~n23803 ;
  assign n23804 = n19362 & n42725 ;
  assign n22854 = n22814 | n22830 ;
  assign n42726 = ~n22854 ;
  assign n23600 = n42726 & n138 ;
  assign n23601 = n22821 | n23600 ;
  assign n22834 = n22821 & n42297 ;
  assign n42727 = ~n22814 ;
  assign n22835 = n42727 & n22834 ;
  assign n23768 = n22835 & n138 ;
  assign n42728 = ~n23768 ;
  assign n23769 = n23601 & n42728 ;
  assign n23811 = n140 & n42711 ;
  assign n23648 = n140 | n23647 ;
  assign n42729 = ~n23648 ;
  assign n23812 = n42729 & n23783 ;
  assign n23813 = n23617 | n23812 ;
  assign n42730 = ~n23811 ;
  assign n23814 = n42730 & n23813 ;
  assign n42731 = ~n23814 ;
  assign n23815 = n141 & n42731 ;
  assign n23816 = n42716 & n23813 ;
  assign n23817 = n23773 | n23816 ;
  assign n42732 = ~n23815 ;
  assign n23818 = n42732 & n23817 ;
  assign n42733 = ~n23818 ;
  assign n23819 = n142 & n42733 ;
  assign n23820 = n143 | n23819 ;
  assign n42734 = ~n23820 ;
  assign n23821 = n23802 & n42734 ;
  assign n23822 = n23769 | n23821 ;
  assign n42735 = ~n23804 ;
  assign n23823 = n42735 & n23822 ;
  assign n42736 = ~n23823 ;
  assign n23824 = n144 & n42736 ;
  assign n42737 = ~n22837 ;
  assign n22844 = n22785 & n42737 ;
  assign n22845 = n42304 & n22844 ;
  assign n23593 = n22845 & n138 ;
  assign n22843 = n22832 | n22837 ;
  assign n42738 = ~n22843 ;
  assign n23620 = n42738 & n138 ;
  assign n23621 = n22785 | n23620 ;
  assign n42739 = ~n23593 ;
  assign n23622 = n42739 & n23621 ;
  assign n23805 = n144 | n23804 ;
  assign n42740 = ~n23805 ;
  assign n23825 = n42740 & n23822 ;
  assign n23826 = n23622 | n23825 ;
  assign n42741 = ~n23824 ;
  assign n23827 = n42741 & n23826 ;
  assign n42742 = ~n23827 ;
  assign n23828 = n145 & n42742 ;
  assign n22842 = n22840 | n22841 ;
  assign n42743 = ~n22842 ;
  assign n23603 = n42743 & n138 ;
  assign n23604 = n22866 | n23603 ;
  assign n22880 = n42331 & n22866 ;
  assign n42744 = ~n22841 ;
  assign n22881 = n42744 & n22880 ;
  assign n23618 = n22881 & n138 ;
  assign n42745 = ~n23618 ;
  assign n23619 = n23604 & n42745 ;
  assign n23836 = n42723 & n23817 ;
  assign n23837 = n23607 | n23836 ;
  assign n42746 = ~n23819 ;
  assign n23838 = n42746 & n23837 ;
  assign n42747 = ~n23838 ;
  assign n23839 = n143 & n42747 ;
  assign n23840 = n42734 & n23837 ;
  assign n23841 = n23769 | n23840 ;
  assign n42748 = ~n23839 ;
  assign n23842 = n42748 & n23841 ;
  assign n42749 = ~n23842 ;
  assign n23843 = n18797 & n42749 ;
  assign n23844 = n145 | n23843 ;
  assign n42750 = ~n23844 ;
  assign n23845 = n23826 & n42750 ;
  assign n23846 = n23619 | n23845 ;
  assign n42751 = ~n23828 ;
  assign n23847 = n42751 & n23846 ;
  assign n42752 = ~n23847 ;
  assign n23848 = n146 & n42752 ;
  assign n22879 = n22869 | n22871 ;
  assign n42753 = ~n22879 ;
  assign n23630 = n42753 & n138 ;
  assign n23631 = n22783 | n23630 ;
  assign n42754 = ~n22871 ;
  assign n22877 = n22783 & n42754 ;
  assign n22878 = n42320 & n22877 ;
  assign n23659 = n22878 & n138 ;
  assign n42755 = ~n23659 ;
  assign n23660 = n23631 & n42755 ;
  assign n23829 = n146 | n23828 ;
  assign n42756 = ~n23829 ;
  assign n23849 = n42756 & n23846 ;
  assign n23850 = n23660 | n23849 ;
  assign n42757 = ~n23848 ;
  assign n23851 = n42757 & n23850 ;
  assign n42758 = ~n23851 ;
  assign n23852 = n16322 & n42758 ;
  assign n22913 = n42347 & n22899 ;
  assign n42759 = ~n22875 ;
  assign n22914 = n42759 & n22913 ;
  assign n23571 = n22914 & n138 ;
  assign n22876 = n22874 | n22875 ;
  assign n42760 = ~n22876 ;
  assign n23632 = n42760 & n138 ;
  assign n23633 = n22899 | n23632 ;
  assign n42761 = ~n23571 ;
  assign n23634 = n42761 & n23633 ;
  assign n23860 = n42740 & n23841 ;
  assign n23861 = n23622 | n23860 ;
  assign n42762 = ~n23843 ;
  assign n23862 = n42762 & n23861 ;
  assign n42763 = ~n23862 ;
  assign n23863 = n145 & n42763 ;
  assign n23864 = n42750 & n23861 ;
  assign n23865 = n23619 | n23864 ;
  assign n42764 = ~n23863 ;
  assign n23866 = n42764 & n23865 ;
  assign n42765 = ~n23866 ;
  assign n23867 = n146 & n42765 ;
  assign n23868 = n147 | n23867 ;
  assign n42766 = ~n23868 ;
  assign n23869 = n23850 & n42766 ;
  assign n23870 = n23634 | n23869 ;
  assign n42767 = ~n23852 ;
  assign n23871 = n42767 & n23870 ;
  assign n42768 = ~n23871 ;
  assign n23872 = n148 & n42768 ;
  assign n22910 = n22902 | n22904 ;
  assign n42769 = ~n22910 ;
  assign n23650 = n42769 & n138 ;
  assign n23651 = n22863 | n23650 ;
  assign n42770 = ~n22904 ;
  assign n22911 = n22863 & n42770 ;
  assign n22912 = n42336 & n22911 ;
  assign n23670 = n22912 & n138 ;
  assign n42771 = ~n23670 ;
  assign n23671 = n23651 & n42771 ;
  assign n23853 = n148 | n23852 ;
  assign n42772 = ~n23853 ;
  assign n23873 = n42772 & n23870 ;
  assign n23876 = n23671 | n23873 ;
  assign n42773 = ~n23872 ;
  assign n23877 = n42773 & n23876 ;
  assign n42774 = ~n23877 ;
  assign n23878 = n149 & n42774 ;
  assign n22909 = n22907 | n22908 ;
  assign n42775 = ~n22909 ;
  assign n23678 = n42775 & n138 ;
  assign n23679 = n22931 | n23678 ;
  assign n22949 = n42360 & n22931 ;
  assign n42776 = ~n22908 ;
  assign n22950 = n42776 & n22949 ;
  assign n23689 = n22950 & n138 ;
  assign n42777 = ~n23689 ;
  assign n23690 = n23679 & n42777 ;
  assign n23884 = n42756 & n23865 ;
  assign n23885 = n23660 | n23884 ;
  assign n42778 = ~n23867 ;
  assign n23886 = n42778 & n23885 ;
  assign n42779 = ~n23886 ;
  assign n23887 = n147 & n42779 ;
  assign n23888 = n42766 & n23885 ;
  assign n23889 = n23634 | n23888 ;
  assign n42780 = ~n23887 ;
  assign n23890 = n42780 & n23889 ;
  assign n42781 = ~n23890 ;
  assign n23891 = n15807 & n42781 ;
  assign n23892 = n149 | n23891 ;
  assign n42782 = ~n23892 ;
  assign n23893 = n23876 & n42782 ;
  assign n23894 = n23690 | n23893 ;
  assign n42783 = ~n23878 ;
  assign n23895 = n42783 & n23894 ;
  assign n42784 = ~n23895 ;
  assign n23896 = n150 & n42784 ;
  assign n22948 = n22934 | n22936 ;
  assign n42785 = ~n22948 ;
  assign n23549 = n42785 & n138 ;
  assign n23550 = n22795 | n23549 ;
  assign n42786 = ~n22936 ;
  assign n22946 = n22795 & n42786 ;
  assign n22947 = n42352 & n22946 ;
  assign n23676 = n22947 & n138 ;
  assign n42787 = ~n23676 ;
  assign n23677 = n23550 & n42787 ;
  assign n23879 = n150 | n23878 ;
  assign n42788 = ~n23879 ;
  assign n23897 = n42788 & n23894 ;
  assign n23898 = n23677 | n23897 ;
  assign n42789 = ~n23896 ;
  assign n23899 = n42789 & n23898 ;
  assign n42790 = ~n23899 ;
  assign n23900 = n13662 & n42790 ;
  assign n22945 = n22939 | n22940 ;
  assign n42791 = ~n22945 ;
  assign n23663 = n42791 & n138 ;
  assign n23664 = n22926 | n23663 ;
  assign n22961 = n22926 & n42379 ;
  assign n42792 = ~n22940 ;
  assign n22962 = n42792 & n22961 ;
  assign n23687 = n22962 & n138 ;
  assign n42793 = ~n23687 ;
  assign n23688 = n23664 & n42793 ;
  assign n23908 = n42772 & n23889 ;
  assign n23909 = n23671 | n23908 ;
  assign n42794 = ~n23891 ;
  assign n23910 = n42794 & n23909 ;
  assign n42795 = ~n23910 ;
  assign n23911 = n149 & n42795 ;
  assign n23912 = n42782 & n23909 ;
  assign n23913 = n23690 | n23912 ;
  assign n42796 = ~n23911 ;
  assign n23914 = n42796 & n23913 ;
  assign n42797 = ~n23914 ;
  assign n23915 = n150 & n42797 ;
  assign n23916 = n151 | n23915 ;
  assign n42798 = ~n23916 ;
  assign n23917 = n23898 & n42798 ;
  assign n23918 = n23688 | n23917 ;
  assign n42799 = ~n23900 ;
  assign n23919 = n42799 & n23918 ;
  assign n42800 = ~n23919 ;
  assign n23920 = n152 & n42800 ;
  assign n42801 = ~n22959 ;
  assign n22985 = n42801 & n22969 ;
  assign n22986 = n42368 & n22985 ;
  assign n23639 = n22986 & n138 ;
  assign n22960 = n22943 | n22959 ;
  assign n42802 = ~n22960 ;
  assign n23667 = n42802 & n138 ;
  assign n23668 = n22969 | n23667 ;
  assign n42803 = ~n23639 ;
  assign n23669 = n42803 & n23668 ;
  assign n23901 = n152 | n23900 ;
  assign n42804 = ~n23901 ;
  assign n23921 = n42804 & n23918 ;
  assign n23922 = n23669 | n23921 ;
  assign n42805 = ~n23920 ;
  assign n23923 = n42805 & n23922 ;
  assign n42806 = ~n23923 ;
  assign n23924 = n153 & n42806 ;
  assign n22974 = n22857 & n42395 ;
  assign n42807 = ~n22990 ;
  assign n23184 = n22974 & n42807 ;
  assign n23653 = n23184 & n138 ;
  assign n23185 = n22989 | n22990 ;
  assign n42808 = ~n23185 ;
  assign n23693 = n42808 & n138 ;
  assign n23694 = n22857 | n23693 ;
  assign n42809 = ~n23653 ;
  assign n23695 = n42809 & n23694 ;
  assign n23932 = n42788 & n23913 ;
  assign n23933 = n23677 | n23932 ;
  assign n42810 = ~n23915 ;
  assign n23934 = n42810 & n23933 ;
  assign n42811 = ~n23934 ;
  assign n23935 = n151 & n42811 ;
  assign n23936 = n42798 & n23933 ;
  assign n23937 = n23688 | n23936 ;
  assign n42812 = ~n23935 ;
  assign n23938 = n42812 & n23937 ;
  assign n42813 = ~n23938 ;
  assign n23939 = n13079 & n42813 ;
  assign n23940 = n153 | n23939 ;
  assign n42814 = ~n23940 ;
  assign n23941 = n23922 & n42814 ;
  assign n23942 = n23695 | n23941 ;
  assign n42815 = ~n23924 ;
  assign n23943 = n42815 & n23942 ;
  assign n42816 = ~n23943 ;
  assign n23944 = n154 & n42816 ;
  assign n42817 = ~n23005 ;
  assign n23181 = n22792 & n42817 ;
  assign n23182 = n42384 & n23181 ;
  assign n23590 = n23182 & n138 ;
  assign n23183 = n22993 | n23005 ;
  assign n42818 = ~n23183 ;
  assign n23684 = n42818 & n138 ;
  assign n23685 = n22792 | n23684 ;
  assign n42819 = ~n23590 ;
  assign n23686 = n42819 & n23685 ;
  assign n23925 = n154 | n23924 ;
  assign n42820 = ~n23925 ;
  assign n23945 = n42820 & n23942 ;
  assign n23946 = n23686 | n23945 ;
  assign n42821 = ~n23944 ;
  assign n23947 = n42821 & n23946 ;
  assign n42822 = ~n23947 ;
  assign n23948 = n11067 & n42822 ;
  assign n22984 = n22797 & n42411 ;
  assign n42823 = ~n23009 ;
  assign n23179 = n22984 & n42823 ;
  assign n23589 = n23179 & n138 ;
  assign n23180 = n23008 | n23009 ;
  assign n42824 = ~n23180 ;
  assign n23635 = n42824 & n138 ;
  assign n23636 = n22797 | n23635 ;
  assign n42825 = ~n23589 ;
  assign n23637 = n42825 & n23636 ;
  assign n23956 = n42804 & n23937 ;
  assign n23957 = n23669 | n23956 ;
  assign n42826 = ~n23939 ;
  assign n23958 = n42826 & n23957 ;
  assign n42827 = ~n23958 ;
  assign n23959 = n153 & n42827 ;
  assign n23960 = n42814 & n23957 ;
  assign n23961 = n23695 | n23960 ;
  assign n42828 = ~n23959 ;
  assign n23962 = n42828 & n23961 ;
  assign n42829 = ~n23962 ;
  assign n23963 = n154 & n42829 ;
  assign n23964 = n11067 | n23963 ;
  assign n42830 = ~n23964 ;
  assign n23965 = n23946 & n42830 ;
  assign n23966 = n23637 | n23965 ;
  assign n42831 = ~n23948 ;
  assign n23967 = n42831 & n23966 ;
  assign n42832 = ~n23967 ;
  assign n23968 = n156 & n42832 ;
  assign n23178 = n23012 | n23024 ;
  assign n42833 = ~n23178 ;
  assign n23587 = n42833 & n138 ;
  assign n23588 = n22745 | n23587 ;
  assign n42834 = ~n23024 ;
  assign n23176 = n22745 & n42834 ;
  assign n23177 = n42400 & n23176 ;
  assign n23665 = n23177 & n138 ;
  assign n42835 = ~n23665 ;
  assign n23666 = n23588 & n42835 ;
  assign n23949 = n10657 | n23948 ;
  assign n42836 = ~n23949 ;
  assign n23969 = n42836 & n23966 ;
  assign n23970 = n23666 | n23969 ;
  assign n42837 = ~n23968 ;
  assign n23971 = n42837 & n23970 ;
  assign n42838 = ~n23971 ;
  assign n23972 = n157 & n42838 ;
  assign n23004 = n22772 & n42427 ;
  assign n42839 = ~n23028 ;
  assign n23174 = n23004 & n42839 ;
  assign n23578 = n23174 & n138 ;
  assign n23175 = n23027 | n23028 ;
  assign n42840 = ~n23175 ;
  assign n23579 = n42840 & n138 ;
  assign n23580 = n22772 | n23579 ;
  assign n42841 = ~n23578 ;
  assign n23581 = n42841 & n23580 ;
  assign n23980 = n42820 & n23961 ;
  assign n23981 = n23686 | n23980 ;
  assign n42842 = ~n23963 ;
  assign n23982 = n42842 & n23981 ;
  assign n42843 = ~n23982 ;
  assign n23983 = n155 & n42843 ;
  assign n23984 = n42830 & n23981 ;
  assign n23985 = n23637 | n23984 ;
  assign n42844 = ~n23983 ;
  assign n23986 = n42844 & n23985 ;
  assign n42845 = ~n23986 ;
  assign n23987 = n10657 & n42845 ;
  assign n23988 = n157 | n23987 ;
  assign n42846 = ~n23988 ;
  assign n23989 = n23970 & n42846 ;
  assign n23990 = n23581 | n23989 ;
  assign n42847 = ~n23972 ;
  assign n23991 = n42847 & n23990 ;
  assign n42848 = ~n23991 ;
  assign n23992 = n158 & n42848 ;
  assign n23173 = n23031 | n23043 ;
  assign n42849 = ~n23173 ;
  assign n23572 = n42849 & n138 ;
  assign n23573 = n22777 | n23572 ;
  assign n42850 = ~n23043 ;
  assign n23171 = n22777 & n42850 ;
  assign n23172 = n42416 & n23171 ;
  assign n23661 = n23172 & n138 ;
  assign n42851 = ~n23661 ;
  assign n23662 = n23573 & n42851 ;
  assign n23974 = n158 | n23972 ;
  assign n42852 = ~n23974 ;
  assign n23993 = n42852 & n23990 ;
  assign n23994 = n23662 | n23993 ;
  assign n42853 = ~n23992 ;
  assign n23995 = n42853 & n23994 ;
  assign n42854 = ~n23995 ;
  assign n23996 = n8857 & n42854 ;
  assign n23023 = n22722 & n42443 ;
  assign n42855 = ~n23047 ;
  assign n23169 = n23023 & n42855 ;
  assign n23564 = n23169 & n138 ;
  assign n23170 = n23046 | n23047 ;
  assign n42856 = ~n23170 ;
  assign n23565 = n42856 & n138 ;
  assign n23566 = n22722 | n23565 ;
  assign n42857 = ~n23564 ;
  assign n23567 = n42857 & n23566 ;
  assign n24004 = n42836 & n23985 ;
  assign n24005 = n23666 | n24004 ;
  assign n42858 = ~n23987 ;
  assign n24006 = n42858 & n24005 ;
  assign n42859 = ~n24006 ;
  assign n24007 = n157 & n42859 ;
  assign n24008 = n42846 & n24005 ;
  assign n24009 = n23581 | n24008 ;
  assign n42860 = ~n24007 ;
  assign n24010 = n42860 & n24009 ;
  assign n42861 = ~n24010 ;
  assign n24011 = n158 & n42861 ;
  assign n24012 = n8857 | n24011 ;
  assign n42862 = ~n24012 ;
  assign n24013 = n23994 & n42862 ;
  assign n24014 = n23567 | n24013 ;
  assign n42863 = ~n23996 ;
  assign n24015 = n42863 & n24014 ;
  assign n42864 = ~n24015 ;
  assign n24016 = n160 & n42864 ;
  assign n42865 = ~n23062 ;
  assign n23166 = n22755 & n42865 ;
  assign n23167 = n42432 & n23166 ;
  assign n23559 = n23167 & n138 ;
  assign n23168 = n23050 | n23062 ;
  assign n42866 = ~n23168 ;
  assign n23560 = n42866 & n138 ;
  assign n23561 = n22755 | n23560 ;
  assign n42867 = ~n23559 ;
  assign n23562 = n42867 & n23561 ;
  assign n23997 = n160 | n23996 ;
  assign n42868 = ~n23997 ;
  assign n24017 = n42868 & n24014 ;
  assign n24018 = n23562 | n24017 ;
  assign n42869 = ~n24016 ;
  assign n24019 = n42869 & n24018 ;
  assign n42870 = ~n24019 ;
  assign n24020 = n161 & n42870 ;
  assign n23042 = n22787 & n42459 ;
  assign n42871 = ~n23066 ;
  assign n23164 = n23042 & n42871 ;
  assign n23558 = n23164 & n138 ;
  assign n23165 = n23065 | n23066 ;
  assign n42872 = ~n23165 ;
  assign n23584 = n42872 & n138 ;
  assign n23585 = n22787 | n23584 ;
  assign n42873 = ~n23558 ;
  assign n23586 = n42873 & n23585 ;
  assign n24028 = n42852 & n24009 ;
  assign n24029 = n23662 | n24028 ;
  assign n42874 = ~n24011 ;
  assign n24030 = n42874 & n24029 ;
  assign n42875 = ~n24030 ;
  assign n24031 = n159 & n42875 ;
  assign n24032 = n42862 & n24029 ;
  assign n24033 = n23567 | n24032 ;
  assign n42876 = ~n24031 ;
  assign n24034 = n42876 & n24033 ;
  assign n42877 = ~n24034 ;
  assign n24035 = n8534 & n42877 ;
  assign n24036 = n161 | n24035 ;
  assign n42878 = ~n24036 ;
  assign n24037 = n24018 & n42878 ;
  assign n24038 = n23586 | n24037 ;
  assign n42879 = ~n24020 ;
  assign n24039 = n42879 & n24038 ;
  assign n42880 = ~n24039 ;
  assign n24040 = n162 & n42880 ;
  assign n23163 = n23069 | n23081 ;
  assign n42881 = ~n23163 ;
  assign n23657 = n42881 & n138 ;
  assign n23658 = n22861 | n23657 ;
  assign n42882 = ~n23081 ;
  assign n23161 = n22861 & n42882 ;
  assign n23162 = n42448 & n23161 ;
  assign n23674 = n23162 & n138 ;
  assign n42883 = ~n23674 ;
  assign n23675 = n23658 & n42883 ;
  assign n24021 = n162 | n24020 ;
  assign n42884 = ~n24021 ;
  assign n24041 = n42884 & n24038 ;
  assign n24042 = n23675 | n24041 ;
  assign n42885 = ~n24040 ;
  assign n24043 = n42885 & n24042 ;
  assign n42886 = ~n24043 ;
  assign n24044 = n6889 & n42886 ;
  assign n23061 = n22725 & n42475 ;
  assign n42887 = ~n23085 ;
  assign n23159 = n23061 & n42887 ;
  assign n23557 = n23159 & n138 ;
  assign n23160 = n23084 | n23085 ;
  assign n42888 = ~n23160 ;
  assign n23568 = n42888 & n138 ;
  assign n23569 = n22725 | n23568 ;
  assign n42889 = ~n23557 ;
  assign n23570 = n42889 & n23569 ;
  assign n24052 = n42868 & n24033 ;
  assign n24053 = n23562 | n24052 ;
  assign n42890 = ~n24035 ;
  assign n24054 = n42890 & n24053 ;
  assign n42891 = ~n24054 ;
  assign n24055 = n161 & n42891 ;
  assign n24056 = n42878 & n24053 ;
  assign n24057 = n23586 | n24056 ;
  assign n42892 = ~n24055 ;
  assign n24058 = n42892 & n24057 ;
  assign n42893 = ~n24058 ;
  assign n24059 = n162 & n42893 ;
  assign n24060 = n6889 | n24059 ;
  assign n42894 = ~n24060 ;
  assign n24061 = n24042 & n42894 ;
  assign n24062 = n23570 | n24061 ;
  assign n42895 = ~n24044 ;
  assign n24063 = n42895 & n24062 ;
  assign n42896 = ~n24063 ;
  assign n24064 = n164 & n42896 ;
  assign n42897 = ~n23100 ;
  assign n23156 = n22750 & n42897 ;
  assign n23157 = n42464 & n23156 ;
  assign n23553 = n23157 & n138 ;
  assign n23158 = n23088 | n23100 ;
  assign n42898 = ~n23158 ;
  assign n23554 = n42898 & n138 ;
  assign n23555 = n22750 | n23554 ;
  assign n42899 = ~n23553 ;
  assign n23556 = n42899 & n23555 ;
  assign n24046 = n6600 | n24044 ;
  assign n42900 = ~n24046 ;
  assign n24065 = n42900 & n24062 ;
  assign n24066 = n23556 | n24065 ;
  assign n42901 = ~n24064 ;
  assign n24067 = n42901 & n24066 ;
  assign n42902 = ~n24067 ;
  assign n24068 = n165 & n42902 ;
  assign n23155 = n23103 | n23104 ;
  assign n42903 = ~n23155 ;
  assign n23547 = n42903 & n138 ;
  assign n23548 = n22767 | n23547 ;
  assign n23080 = n22767 & n42491 ;
  assign n42904 = ~n23104 ;
  assign n23154 = n23080 & n42904 ;
  assign n23608 = n23154 & n138 ;
  assign n42905 = ~n23608 ;
  assign n23609 = n23548 & n42905 ;
  assign n24076 = n42884 & n24057 ;
  assign n24077 = n23675 | n24076 ;
  assign n42906 = ~n24059 ;
  assign n24078 = n42906 & n24077 ;
  assign n42907 = ~n24078 ;
  assign n24079 = n163 & n42907 ;
  assign n24080 = n42894 & n24077 ;
  assign n24081 = n23570 | n24080 ;
  assign n42908 = ~n24079 ;
  assign n24082 = n42908 & n24081 ;
  assign n42909 = ~n24082 ;
  assign n24083 = n6600 & n42909 ;
  assign n24084 = n165 | n24083 ;
  assign n42910 = ~n24084 ;
  assign n24085 = n24066 & n42910 ;
  assign n24086 = n23609 | n24085 ;
  assign n42911 = ~n24068 ;
  assign n24087 = n42911 & n24086 ;
  assign n42912 = ~n24087 ;
  assign n24088 = n166 & n42912 ;
  assign n42913 = ~n23119 ;
  assign n23151 = n22770 & n42913 ;
  assign n23152 = n42480 & n23151 ;
  assign n23546 = n23152 & n138 ;
  assign n23153 = n23107 | n23119 ;
  assign n42914 = ~n23153 ;
  assign n23597 = n42914 & n138 ;
  assign n23598 = n22770 | n23597 ;
  assign n42915 = ~n23546 ;
  assign n23599 = n42915 & n23598 ;
  assign n24069 = n166 | n24068 ;
  assign n42916 = ~n24069 ;
  assign n24089 = n42916 & n24086 ;
  assign n24090 = n23599 | n24089 ;
  assign n42917 = ~n24088 ;
  assign n24091 = n42917 & n24090 ;
  assign n42918 = ~n24091 ;
  assign n24092 = n5352 & n42918 ;
  assign n23150 = n23122 | n23123 ;
  assign n42919 = ~n23150 ;
  assign n23582 = n42919 & n138 ;
  assign n23583 = n22731 | n23582 ;
  assign n23099 = n22731 & n42504 ;
  assign n42920 = ~n23123 ;
  assign n23149 = n23099 & n42920 ;
  assign n23594 = n23149 & n138 ;
  assign n42921 = ~n23594 ;
  assign n23595 = n23583 & n42921 ;
  assign n24100 = n42900 & n24081 ;
  assign n24101 = n23556 | n24100 ;
  assign n42922 = ~n24083 ;
  assign n24102 = n42922 & n24101 ;
  assign n42923 = ~n24102 ;
  assign n24103 = n165 & n42923 ;
  assign n24104 = n42910 & n24101 ;
  assign n24105 = n23609 | n24104 ;
  assign n42924 = ~n24103 ;
  assign n24106 = n42924 & n24105 ;
  assign n42925 = ~n24106 ;
  assign n24107 = n166 & n42925 ;
  assign n24108 = n5352 | n24107 ;
  assign n42926 = ~n24108 ;
  assign n24109 = n24090 & n42926 ;
  assign n24110 = n23595 | n24109 ;
  assign n42927 = ~n24092 ;
  assign n24111 = n42927 & n24110 ;
  assign n42928 = ~n24111 ;
  assign n24112 = n168 & n42928 ;
  assign n42929 = ~n23133 ;
  assign n23146 = n22762 & n42929 ;
  assign n23147 = n42496 & n23146 ;
  assign n23652 = n23147 & n138 ;
  assign n23148 = n23126 | n23133 ;
  assign n42930 = ~n23148 ;
  assign n23680 = n42930 & n138 ;
  assign n23681 = n22762 | n23680 ;
  assign n42931 = ~n23652 ;
  assign n23682 = n42931 & n23681 ;
  assign n24093 = n4934 | n24092 ;
  assign n42932 = ~n24093 ;
  assign n24113 = n42932 & n24110 ;
  assign n24114 = n23682 | n24113 ;
  assign n42933 = ~n24112 ;
  assign n24115 = n42933 & n24114 ;
  assign n42934 = ~n24115 ;
  assign n24116 = n169 & n42934 ;
  assign n23145 = n23136 | n23137 ;
  assign n42935 = ~n23145 ;
  assign n23574 = n42935 & n138 ;
  assign n23575 = n22697 | n23574 ;
  assign n23118 = n22697 & n42523 ;
  assign n42936 = ~n23137 ;
  assign n23144 = n23118 & n42936 ;
  assign n23696 = n23144 & n138 ;
  assign n42937 = ~n23696 ;
  assign n23697 = n23575 & n42937 ;
  assign n24124 = n42916 & n24105 ;
  assign n24125 = n23599 | n24124 ;
  assign n42938 = ~n24107 ;
  assign n24126 = n42938 & n24125 ;
  assign n42939 = ~n24126 ;
  assign n24127 = n167 & n42939 ;
  assign n24128 = n42926 & n24125 ;
  assign n24129 = n23595 | n24128 ;
  assign n42940 = ~n24127 ;
  assign n24130 = n42940 & n24129 ;
  assign n42941 = ~n24130 ;
  assign n24131 = n4934 & n42941 ;
  assign n24132 = n169 | n24131 ;
  assign n42942 = ~n24132 ;
  assign n24133 = n24114 & n42942 ;
  assign n24134 = n23697 | n24133 ;
  assign n42943 = ~n24116 ;
  assign n24135 = n42943 & n24134 ;
  assign n42944 = ~n24135 ;
  assign n24136 = n170 & n42944 ;
  assign n23143 = n23140 | n23142 ;
  assign n42945 = ~n23143 ;
  assign n23698 = n42945 & n138 ;
  assign n23699 = n23190 | n23698 ;
  assign n42946 = ~n23142 ;
  assign n23196 = n42946 & n23190 ;
  assign n23197 = n42512 & n23196 ;
  assign n23701 = n23197 & n138 ;
  assign n42947 = ~n23701 ;
  assign n23702 = n23699 & n42947 ;
  assign n24117 = n170 | n24116 ;
  assign n42948 = ~n24117 ;
  assign n24137 = n42948 & n24134 ;
  assign n24138 = n23702 | n24137 ;
  assign n42949 = ~n24136 ;
  assign n24139 = n42949 & n24138 ;
  assign n42950 = ~n24139 ;
  assign n24140 = n3940 & n42950 ;
  assign n23202 = n23200 | n23201 ;
  assign n42951 = ~n23202 ;
  assign n23703 = n42951 & n138 ;
  assign n23704 = n23207 | n23703 ;
  assign n23221 = n42536 & n23207 ;
  assign n42952 = ~n23201 ;
  assign n23222 = n42952 & n23221 ;
  assign n23705 = n23222 & n138 ;
  assign n42953 = ~n23705 ;
  assign n23706 = n23704 & n42953 ;
  assign n24148 = n42932 & n24129 ;
  assign n24149 = n23682 | n24148 ;
  assign n42954 = ~n24131 ;
  assign n24150 = n42954 & n24149 ;
  assign n42955 = ~n24150 ;
  assign n24151 = n169 & n42955 ;
  assign n24152 = n42942 & n24149 ;
  assign n24153 = n23697 | n24152 ;
  assign n42956 = ~n24151 ;
  assign n24154 = n42956 & n24153 ;
  assign n42957 = ~n24154 ;
  assign n24155 = n170 & n42957 ;
  assign n24156 = n3940 | n24155 ;
  assign n42958 = ~n24156 ;
  assign n24157 = n24138 & n42958 ;
  assign n24158 = n23706 | n24157 ;
  assign n42959 = ~n24140 ;
  assign n24159 = n42959 & n24158 ;
  assign n42960 = ~n24159 ;
  assign n24160 = n172 & n42960 ;
  assign n23220 = n23210 | n23212 ;
  assign n42961 = ~n23220 ;
  assign n23707 = n42961 & n138 ;
  assign n23708 = n22896 | n23707 ;
  assign n42962 = ~n23212 ;
  assign n23218 = n22896 & n42962 ;
  assign n23219 = n42528 & n23218 ;
  assign n23711 = n23219 & n138 ;
  assign n42963 = ~n23711 ;
  assign n23712 = n23708 & n42963 ;
  assign n24141 = n3631 | n24140 ;
  assign n42964 = ~n24141 ;
  assign n24161 = n42964 & n24158 ;
  assign n24162 = n23712 | n24161 ;
  assign n42965 = ~n24160 ;
  assign n24163 = n42965 & n24162 ;
  assign n42966 = ~n24163 ;
  assign n24164 = n173 & n42966 ;
  assign n23217 = n23215 | n23216 ;
  assign n42967 = ~n23217 ;
  assign n23640 = n42967 & n138 ;
  assign n23641 = n23235 | n23640 ;
  assign n23242 = n42555 & n23235 ;
  assign n42968 = ~n23216 ;
  assign n23243 = n42968 & n23242 ;
  assign n23691 = n23243 & n138 ;
  assign n42969 = ~n23691 ;
  assign n23692 = n23641 & n42969 ;
  assign n24172 = n42948 & n24153 ;
  assign n24173 = n23702 | n24172 ;
  assign n42970 = ~n24155 ;
  assign n24174 = n42970 & n24173 ;
  assign n42971 = ~n24174 ;
  assign n24175 = n171 & n42971 ;
  assign n24176 = n42958 & n24173 ;
  assign n24177 = n23706 | n24176 ;
  assign n42972 = ~n24175 ;
  assign n24178 = n42972 & n24177 ;
  assign n42973 = ~n24178 ;
  assign n24179 = n3631 & n42973 ;
  assign n24180 = n173 | n24179 ;
  assign n42974 = ~n24180 ;
  assign n24181 = n24162 & n42974 ;
  assign n24182 = n23692 | n24181 ;
  assign n42975 = ~n24164 ;
  assign n24183 = n42975 & n24182 ;
  assign n42976 = ~n24183 ;
  assign n24184 = n174 & n42976 ;
  assign n42977 = ~n23240 ;
  assign n23251 = n42977 & n23250 ;
  assign n23252 = n42544 & n23251 ;
  assign n23700 = n23252 & n138 ;
  assign n23241 = n23238 | n23240 ;
  assign n42978 = ~n23241 ;
  assign n23713 = n42978 & n138 ;
  assign n23714 = n23250 | n23713 ;
  assign n42979 = ~n23700 ;
  assign n23715 = n42979 & n23714 ;
  assign n24165 = n174 | n24164 ;
  assign n42980 = ~n24165 ;
  assign n24185 = n42980 & n24182 ;
  assign n24186 = n23715 | n24185 ;
  assign n42981 = ~n24184 ;
  assign n24187 = n42981 & n24186 ;
  assign n42982 = ~n24187 ;
  assign n24188 = n2753 & n42982 ;
  assign n23278 = n42568 & n23264 ;
  assign n42983 = ~n23256 ;
  assign n23279 = n42983 & n23278 ;
  assign n23610 = n23279 & n138 ;
  assign n23257 = n23255 | n23256 ;
  assign n42984 = ~n23257 ;
  assign n23654 = n42984 & n138 ;
  assign n23655 = n23264 | n23654 ;
  assign n42985 = ~n23610 ;
  assign n23656 = n42985 & n23655 ;
  assign n24196 = n42964 & n24177 ;
  assign n24197 = n23712 | n24196 ;
  assign n42986 = ~n24179 ;
  assign n24198 = n42986 & n24197 ;
  assign n42987 = ~n24198 ;
  assign n24199 = n173 & n42987 ;
  assign n24200 = n42974 & n24197 ;
  assign n24201 = n23692 | n24200 ;
  assign n42988 = ~n24199 ;
  assign n24202 = n42988 & n24201 ;
  assign n42989 = ~n24202 ;
  assign n24203 = n174 & n42989 ;
  assign n24204 = n2753 | n24203 ;
  assign n42990 = ~n24204 ;
  assign n24205 = n24186 & n42990 ;
  assign n24206 = n23656 | n24205 ;
  assign n42991 = ~n24188 ;
  assign n24207 = n42991 & n24206 ;
  assign n42992 = ~n24207 ;
  assign n24208 = n176 & n42992 ;
  assign n42993 = ~n23269 ;
  assign n23275 = n23204 & n42993 ;
  assign n23276 = n42560 & n23275 ;
  assign n23642 = n23276 & n138 ;
  assign n23277 = n23267 | n23269 ;
  assign n42994 = ~n23277 ;
  assign n23716 = n42994 & n138 ;
  assign n23717 = n23204 | n23716 ;
  assign n42995 = ~n23642 ;
  assign n23718 = n42995 & n23717 ;
  assign n24189 = n2431 | n24188 ;
  assign n42996 = ~n24189 ;
  assign n24209 = n42996 & n24206 ;
  assign n24210 = n23718 | n24209 ;
  assign n42997 = ~n24208 ;
  assign n24211 = n42997 & n24210 ;
  assign n42998 = ~n24211 ;
  assign n24212 = n177 & n42998 ;
  assign n23274 = n23272 | n23273 ;
  assign n42999 = ~n23274 ;
  assign n23672 = n42999 & n138 ;
  assign n23673 = n23294 | n23672 ;
  assign n23301 = n42584 & n23294 ;
  assign n43000 = ~n23273 ;
  assign n23302 = n43000 & n23301 ;
  assign n23709 = n23302 & n138 ;
  assign n43001 = ~n23709 ;
  assign n23710 = n23673 & n43001 ;
  assign n24220 = n42980 & n24201 ;
  assign n24221 = n23715 | n24220 ;
  assign n43002 = ~n24203 ;
  assign n24222 = n43002 & n24221 ;
  assign n43003 = ~n24222 ;
  assign n24223 = n175 & n43003 ;
  assign n24224 = n42990 & n24221 ;
  assign n24225 = n23656 | n24224 ;
  assign n43004 = ~n24223 ;
  assign n24226 = n43004 & n24225 ;
  assign n43005 = ~n24226 ;
  assign n24227 = n2431 & n43005 ;
  assign n24228 = n177 | n24227 ;
  assign n43006 = ~n24228 ;
  assign n24229 = n24210 & n43006 ;
  assign n24230 = n23710 | n24229 ;
  assign n43007 = ~n24212 ;
  assign n24231 = n43007 & n24230 ;
  assign n43008 = ~n24231 ;
  assign n24232 = n178 & n43008 ;
  assign n23300 = n23297 | n23299 ;
  assign n43009 = ~n23300 ;
  assign n23721 = n43009 & n138 ;
  assign n23722 = n23308 | n23721 ;
  assign n43010 = ~n23299 ;
  assign n23314 = n43010 & n23308 ;
  assign n23315 = n42576 & n23314 ;
  assign n23724 = n23315 & n138 ;
  assign n43011 = ~n23724 ;
  assign n23725 = n23722 & n43011 ;
  assign n24213 = n178 | n24212 ;
  assign n43012 = ~n24213 ;
  assign n24233 = n43012 & n24230 ;
  assign n24234 = n23725 | n24233 ;
  assign n43013 = ~n24232 ;
  assign n24235 = n43013 & n24234 ;
  assign n43014 = ~n24235 ;
  assign n24236 = n1707 & n43014 ;
  assign n23332 = n42600 & n23325 ;
  assign n43015 = ~n23319 ;
  assign n23333 = n43015 & n23332 ;
  assign n23649 = n23333 & n138 ;
  assign n23320 = n23318 | n23319 ;
  assign n43016 = ~n23320 ;
  assign n23726 = n43016 & n138 ;
  assign n23727 = n23325 | n23726 ;
  assign n43017 = ~n23649 ;
  assign n23728 = n43017 & n23727 ;
  assign n24244 = n42996 & n24225 ;
  assign n24245 = n23718 | n24244 ;
  assign n43018 = ~n24227 ;
  assign n24246 = n43018 & n24245 ;
  assign n43019 = ~n24246 ;
  assign n24247 = n177 & n43019 ;
  assign n24248 = n43006 & n24245 ;
  assign n24249 = n23710 | n24248 ;
  assign n43020 = ~n24247 ;
  assign n24250 = n43020 & n24249 ;
  assign n43021 = ~n24250 ;
  assign n24251 = n178 & n43021 ;
  assign n24252 = n1707 | n24251 ;
  assign n43022 = ~n24252 ;
  assign n24253 = n24234 & n43022 ;
  assign n24254 = n23728 | n24253 ;
  assign n43023 = ~n24236 ;
  assign n24255 = n43023 & n24254 ;
  assign n43024 = ~n24255 ;
  assign n24256 = n180 & n43024 ;
  assign n23331 = n23328 | n23330 ;
  assign n43025 = ~n23331 ;
  assign n23643 = n43025 & n138 ;
  assign n23644 = n23341 | n23643 ;
  assign n43026 = ~n23330 ;
  assign n23347 = n43026 & n23341 ;
  assign n23348 = n42592 & n23347 ;
  assign n23729 = n23348 & n138 ;
  assign n43027 = ~n23729 ;
  assign n23730 = n23644 & n43027 ;
  assign n24237 = n1487 | n24236 ;
  assign n43028 = ~n24237 ;
  assign n24257 = n43028 & n24254 ;
  assign n24258 = n23730 | n24257 ;
  assign n43029 = ~n24256 ;
  assign n24259 = n43029 & n24258 ;
  assign n43030 = ~n24259 ;
  assign n24260 = n181 & n43030 ;
  assign n23362 = n42616 & n23355 ;
  assign n43031 = ~n23352 ;
  assign n23363 = n43031 & n23362 ;
  assign n23683 = n23363 & n138 ;
  assign n23353 = n23351 | n23352 ;
  assign n43032 = ~n23353 ;
  assign n23731 = n43032 & n138 ;
  assign n23732 = n23355 | n23731 ;
  assign n43033 = ~n23683 ;
  assign n23733 = n43033 & n23732 ;
  assign n24268 = n43012 & n24249 ;
  assign n24269 = n23725 | n24268 ;
  assign n43034 = ~n24251 ;
  assign n24270 = n43034 & n24269 ;
  assign n43035 = ~n24270 ;
  assign n24271 = n179 & n43035 ;
  assign n24272 = n43022 & n24269 ;
  assign n24273 = n23728 | n24272 ;
  assign n43036 = ~n24271 ;
  assign n24274 = n43036 & n24273 ;
  assign n43037 = ~n24274 ;
  assign n24275 = n1487 & n43037 ;
  assign n24276 = n181 | n24275 ;
  assign n43038 = ~n24276 ;
  assign n24277 = n24258 & n43038 ;
  assign n24278 = n23733 | n24277 ;
  assign n43039 = ~n24260 ;
  assign n24279 = n43039 & n24278 ;
  assign n43040 = ~n24279 ;
  assign n24280 = n182 & n43040 ;
  assign n43041 = ~n23360 ;
  assign n23375 = n43041 & n23369 ;
  assign n23376 = n42608 & n23375 ;
  assign n23563 = n23376 & n138 ;
  assign n23361 = n23358 | n23360 ;
  assign n43042 = ~n23361 ;
  assign n23734 = n43042 & n138 ;
  assign n23735 = n23369 | n23734 ;
  assign n43043 = ~n23563 ;
  assign n23736 = n43043 & n23735 ;
  assign n24261 = n182 | n24260 ;
  assign n43044 = ~n24261 ;
  assign n24281 = n43044 & n24278 ;
  assign n24282 = n23736 | n24281 ;
  assign n43045 = ~n24280 ;
  assign n24283 = n43045 & n24282 ;
  assign n43046 = ~n24283 ;
  assign n24284 = n996 & n43046 ;
  assign n23381 = n23379 | n23380 ;
  assign n43047 = ~n23381 ;
  assign n23576 = n43047 & n138 ;
  assign n23577 = n23384 | n23576 ;
  assign n23391 = n42632 & n23384 ;
  assign n43048 = ~n23380 ;
  assign n23392 = n43048 & n23391 ;
  assign n23737 = n23392 & n138 ;
  assign n43049 = ~n23737 ;
  assign n23738 = n23577 & n43049 ;
  assign n24292 = n43028 & n24273 ;
  assign n24293 = n23730 | n24292 ;
  assign n43050 = ~n24275 ;
  assign n24294 = n43050 & n24293 ;
  assign n43051 = ~n24294 ;
  assign n24295 = n181 & n43051 ;
  assign n24296 = n43038 & n24293 ;
  assign n24297 = n23733 | n24296 ;
  assign n43052 = ~n24295 ;
  assign n24298 = n43052 & n24297 ;
  assign n43053 = ~n24298 ;
  assign n24299 = n182 & n43053 ;
  assign n24300 = n183 | n24299 ;
  assign n43054 = ~n24300 ;
  assign n24301 = n24282 & n43054 ;
  assign n24302 = n23738 | n24301 ;
  assign n43055 = ~n24284 ;
  assign n24303 = n43055 & n24302 ;
  assign n43056 = ~n24303 ;
  assign n24304 = n184 & n43056 ;
  assign n23390 = n23387 | n23389 ;
  assign n43057 = ~n23390 ;
  assign n23739 = n43057 & n138 ;
  assign n23740 = n23398 | n23739 ;
  assign n43058 = ~n23389 ;
  assign n23404 = n43058 & n23398 ;
  assign n23405 = n42624 & n23404 ;
  assign n23741 = n23405 & n138 ;
  assign n43059 = ~n23741 ;
  assign n23742 = n23740 & n43059 ;
  assign n24285 = n838 | n24284 ;
  assign n43060 = ~n24285 ;
  assign n24305 = n43060 & n24302 ;
  assign n24306 = n23742 | n24305 ;
  assign n43061 = ~n24304 ;
  assign n24307 = n43061 & n24306 ;
  assign n43062 = ~n24307 ;
  assign n24308 = n185 & n43062 ;
  assign n23420 = n42651 & n23413 ;
  assign n43063 = ~n23409 ;
  assign n23421 = n43063 & n23420 ;
  assign n23638 = n23421 & n138 ;
  assign n23410 = n23408 | n23409 ;
  assign n43064 = ~n23410 ;
  assign n23743 = n43064 & n138 ;
  assign n23744 = n23413 | n23743 ;
  assign n43065 = ~n23638 ;
  assign n23745 = n43065 & n23744 ;
  assign n24316 = n43044 & n24297 ;
  assign n24317 = n23736 | n24316 ;
  assign n43066 = ~n24299 ;
  assign n24318 = n43066 & n24317 ;
  assign n43067 = ~n24318 ;
  assign n24319 = n183 & n43067 ;
  assign n24320 = n43054 & n24317 ;
  assign n24321 = n23738 | n24320 ;
  assign n43068 = ~n24319 ;
  assign n24322 = n43068 & n24321 ;
  assign n43069 = ~n24322 ;
  assign n24323 = n838 & n43069 ;
  assign n24324 = n185 | n24323 ;
  assign n43070 = ~n24324 ;
  assign n24325 = n24306 & n43070 ;
  assign n24326 = n23745 | n24325 ;
  assign n43071 = ~n24308 ;
  assign n24327 = n43071 & n24326 ;
  assign n43072 = ~n24327 ;
  assign n24328 = n186 & n43072 ;
  assign n43073 = ~n23418 ;
  assign n23443 = n43073 & n23428 ;
  assign n23444 = n42640 & n23443 ;
  assign n23602 = n23444 & n138 ;
  assign n23419 = n23416 | n23418 ;
  assign n43074 = ~n23419 ;
  assign n23625 = n43074 & n138 ;
  assign n23626 = n23428 | n23625 ;
  assign n43075 = ~n23602 ;
  assign n23627 = n43075 & n23626 ;
  assign n24309 = n186 | n24308 ;
  assign n43076 = ~n24309 ;
  assign n24329 = n43076 & n24326 ;
  assign n24330 = n23627 | n24329 ;
  assign n43077 = ~n24328 ;
  assign n24331 = n43077 & n24330 ;
  assign n43078 = ~n24331 ;
  assign n24332 = n528 & n43078 ;
  assign n23464 = n23447 | n23448 ;
  assign n43079 = ~n23464 ;
  assign n23746 = n43079 & n138 ;
  assign n23747 = n22774 | n23746 ;
  assign n23433 = n22774 & n42664 ;
  assign n43080 = ~n23448 ;
  assign n23463 = n23433 & n43080 ;
  assign n23748 = n23463 & n138 ;
  assign n43081 = ~n23748 ;
  assign n23749 = n23747 & n43081 ;
  assign n24340 = n43060 & n24321 ;
  assign n24341 = n23742 | n24340 ;
  assign n43082 = ~n24323 ;
  assign n24342 = n43082 & n24341 ;
  assign n43083 = ~n24342 ;
  assign n24343 = n185 & n43083 ;
  assign n24344 = n43070 & n24341 ;
  assign n24345 = n23745 | n24344 ;
  assign n43084 = ~n24343 ;
  assign n24346 = n43084 & n24345 ;
  assign n43085 = ~n24346 ;
  assign n24347 = n186 & n43085 ;
  assign n24348 = n528 | n24347 ;
  assign n43086 = ~n24348 ;
  assign n24349 = n24330 & n43086 ;
  assign n24350 = n23749 | n24349 ;
  assign n43087 = ~n24332 ;
  assign n24351 = n43087 & n24350 ;
  assign n43088 = ~n24351 ;
  assign n24352 = n188 & n43088 ;
  assign n23462 = n23451 | n23454 ;
  assign n43089 = ~n23462 ;
  assign n23591 = n43089 & n138 ;
  assign n23592 = n22719 | n23591 ;
  assign n43090 = ~n23454 ;
  assign n23460 = n22719 & n43090 ;
  assign n23461 = n42656 & n23460 ;
  assign n23611 = n23461 & n138 ;
  assign n43091 = ~n23611 ;
  assign n23612 = n23592 & n43091 ;
  assign n24334 = n413 | n24332 ;
  assign n43092 = ~n24334 ;
  assign n24353 = n43092 & n24350 ;
  assign n24354 = n23612 | n24353 ;
  assign n43093 = ~n24352 ;
  assign n24355 = n43093 & n24354 ;
  assign n43094 = ~n24355 ;
  assign n24356 = n189 & n43094 ;
  assign n23459 = n23457 | n23458 ;
  assign n43095 = ~n23459 ;
  assign n23628 = n43095 & n138 ;
  assign n23629 = n23471 | n23628 ;
  assign n23478 = n42683 & n23471 ;
  assign n43096 = ~n23458 ;
  assign n23479 = n43096 & n23478 ;
  assign n23719 = n23479 & n138 ;
  assign n43097 = ~n23719 ;
  assign n23720 = n23629 & n43097 ;
  assign n24364 = n43076 & n24345 ;
  assign n24365 = n23627 | n24364 ;
  assign n43098 = ~n24347 ;
  assign n24366 = n43098 & n24365 ;
  assign n43099 = ~n24366 ;
  assign n24367 = n187 & n43099 ;
  assign n24368 = n43086 & n24365 ;
  assign n24369 = n23749 | n24368 ;
  assign n43100 = ~n24367 ;
  assign n24370 = n43100 & n24369 ;
  assign n43101 = ~n24370 ;
  assign n24371 = n413 & n43101 ;
  assign n24372 = n189 | n24371 ;
  assign n43102 = ~n24372 ;
  assign n24373 = n24354 & n43102 ;
  assign n24374 = n23720 | n24373 ;
  assign n43103 = ~n24356 ;
  assign n24375 = n43103 & n24374 ;
  assign n43104 = ~n24375 ;
  assign n24376 = n190 & n43104 ;
  assign n43105 = ~n23476 ;
  assign n23510 = n43105 & n23509 ;
  assign n23511 = n42672 & n23510 ;
  assign n23723 = n23511 & n138 ;
  assign n23477 = n23474 | n23476 ;
  assign n43106 = ~n23477 ;
  assign n23750 = n43106 & n138 ;
  assign n23751 = n23509 | n23750 ;
  assign n43107 = ~n23723 ;
  assign n23752 = n43107 & n23751 ;
  assign n24357 = n190 | n24356 ;
  assign n43108 = ~n24357 ;
  assign n24377 = n43108 & n24374 ;
  assign n24378 = n23752 | n24377 ;
  assign n43109 = ~n24376 ;
  assign n24379 = n43109 & n24378 ;
  assign n43110 = ~n24379 ;
  assign n24380 = n287 & n43110 ;
  assign n24387 = n43092 & n24369 ;
  assign n24388 = n23612 | n24387 ;
  assign n43111 = ~n24371 ;
  assign n24389 = n43111 & n24388 ;
  assign n43112 = ~n24389 ;
  assign n24390 = n189 & n43112 ;
  assign n24391 = n43102 & n24388 ;
  assign n24392 = n23720 | n24391 ;
  assign n43113 = ~n24390 ;
  assign n24393 = n43113 & n24392 ;
  assign n43114 = ~n24393 ;
  assign n24394 = n190 & n43114 ;
  assign n24395 = n287 | n24394 ;
  assign n43115 = ~n24395 ;
  assign n24396 = n24378 & n43115 ;
  assign n23520 = n23514 | n23515 ;
  assign n43116 = ~n23520 ;
  assign n23551 = n43116 & n138 ;
  assign n23552 = n23507 | n23551 ;
  assign n43117 = ~n23523 ;
  assign n24399 = n23507 & n43117 ;
  assign n43118 = ~n23515 ;
  assign n24400 = n43118 & n24399 ;
  assign n24401 = n138 & n24400 ;
  assign n43119 = ~n24401 ;
  assign n24402 = n23552 & n43119 ;
  assign n24405 = n24396 | n24402 ;
  assign n43120 = ~n24380 ;
  assign n24406 = n43120 & n24405 ;
  assign n24409 = n23767 | n24406 ;
  assign n24410 = n31336 & n24409 ;
  assign n23467 = n22678 | n23465 ;
  assign n43121 = ~n23467 ;
  assign n23468 = n23187 & n43121 ;
  assign n23493 = n23468 & n42698 ;
  assign n23539 = n23493 & n42699 ;
  assign n23540 = n42700 & n23539 ;
  assign n23534 = n192 & n23533 ;
  assign n43122 = ~n23466 ;
  assign n23759 = n43122 & n138 ;
  assign n43123 = ~n23759 ;
  assign n23760 = n23530 & n43123 ;
  assign n43124 = ~n23760 ;
  assign n23761 = n23534 & n43124 ;
  assign n23763 = n23540 | n23761 ;
  assign n24381 = n23757 & n43120 ;
  assign n24411 = n24381 & n24405 ;
  assign n24412 = n23763 | n24411 ;
  assign n137 = n24410 | n24412 ;
  assign n24491 = x16 & n137 ;
  assign n43125 = ~n24491 ;
  assign n24492 = n249 & n43125 ;
  assign n43126 = ~n24492 ;
  assign n24493 = n138 & n43126 ;
  assign n22680 = n249 & n42697 ;
  assign n23494 = n22680 & n42698 ;
  assign n23542 = n23494 & n42699 ;
  assign n23543 = n42700 & n23542 ;
  assign n24631 = n23543 & n43125 ;
  assign n43127 = ~n245 ;
  assign n24495 = n43127 & n137 ;
  assign n43128 = ~x16 ;
  assign n24639 = n43128 & n137 ;
  assign n43129 = ~n24639 ;
  assign n24640 = x17 & n43129 ;
  assign n24641 = n24495 | n24640 ;
  assign n24642 = n24631 | n24641 ;
  assign n43130 = ~n24493 ;
  assign n24644 = n43130 & n24642 ;
  assign n43131 = ~n24644 ;
  assign n24645 = n22661 & n43131 ;
  assign n250 = n43128 & n248 ;
  assign n43132 = ~n137 ;
  assign n24634 = x16 & n43132 ;
  assign n24635 = n250 | n24634 ;
  assign n43133 = ~n24635 ;
  assign n24636 = n138 & n43133 ;
  assign n24637 = n22661 | n24636 ;
  assign n43134 = ~n24637 ;
  assign n24643 = n43134 & n24642 ;
  assign n43135 = ~n23540 ;
  assign n23770 = n43135 & n138 ;
  assign n43136 = ~n23761 ;
  assign n23771 = n43136 & n23770 ;
  assign n43137 = ~n24411 ;
  assign n24651 = n23771 & n43137 ;
  assign n43138 = ~n24410 ;
  assign n24652 = n43138 & n24651 ;
  assign n24653 = n24495 | n24652 ;
  assign n24654 = x18 & n24653 ;
  assign n24655 = x18 | n24652 ;
  assign n24656 = n24495 | n24655 ;
  assign n43139 = ~n24654 ;
  assign n24657 = n43139 & n24656 ;
  assign n24658 = n24643 | n24657 ;
  assign n43140 = ~n24645 ;
  assign n24659 = n43140 & n24658 ;
  assign n43141 = ~n24659 ;
  assign n24660 = n22030 & n43141 ;
  assign n23779 = n23774 | n23777 ;
  assign n43142 = ~n23779 ;
  assign n24538 = n43142 & n137 ;
  assign n24539 = n23782 | n24538 ;
  assign n23787 = n43142 & n23782 ;
  assign n24546 = n23787 & n137 ;
  assign n43143 = ~n24546 ;
  assign n24547 = n24539 & n43143 ;
  assign n24646 = n22030 | n24645 ;
  assign n43144 = ~n24646 ;
  assign n24663 = n43144 & n24658 ;
  assign n24664 = n24547 | n24663 ;
  assign n43145 = ~n24660 ;
  assign n24665 = n43145 & n24664 ;
  assign n43146 = ~n24665 ;
  assign n24666 = n141 & n43146 ;
  assign n43147 = ~n23784 ;
  assign n23786 = n23617 & n43147 ;
  assign n23794 = n23786 & n42712 ;
  assign n24455 = n23794 & n137 ;
  assign n23795 = n23784 | n23789 ;
  assign n43148 = ~n23795 ;
  assign n24483 = n43148 & n137 ;
  assign n24484 = n23617 | n24483 ;
  assign n43149 = ~n24455 ;
  assign n24485 = n43149 & n24484 ;
  assign n24661 = n141 | n24660 ;
  assign n43150 = ~n24661 ;
  assign n24667 = n43150 & n24664 ;
  assign n24671 = n24485 | n24667 ;
  assign n43151 = ~n24666 ;
  assign n24672 = n43151 & n24671 ;
  assign n43152 = ~n24672 ;
  assign n24673 = n142 & n43152 ;
  assign n23809 = n23791 | n23797 ;
  assign n43153 = ~n23809 ;
  assign n24481 = n43153 & n137 ;
  assign n24482 = n23773 | n24481 ;
  assign n23793 = n23773 & n42717 ;
  assign n43154 = ~n23797 ;
  assign n23810 = n23793 & n43154 ;
  assign n24632 = n23810 & n137 ;
  assign n43155 = ~n24632 ;
  assign n24633 = n24482 & n43155 ;
  assign n24647 = n139 & n43131 ;
  assign n24494 = n139 | n24493 ;
  assign n43156 = ~n24494 ;
  assign n24649 = n43156 & n24642 ;
  assign n24680 = n24649 | n24657 ;
  assign n43157 = ~n24647 ;
  assign n24681 = n43157 & n24680 ;
  assign n43158 = ~n24681 ;
  assign n24682 = n140 & n43158 ;
  assign n24683 = n43144 & n24680 ;
  assign n24684 = n24547 | n24683 ;
  assign n43159 = ~n24682 ;
  assign n24685 = n43159 & n24684 ;
  assign n43160 = ~n24685 ;
  assign n24686 = n141 & n43160 ;
  assign n24687 = n142 | n24686 ;
  assign n43161 = ~n24687 ;
  assign n24688 = n24671 & n43161 ;
  assign n24689 = n24633 | n24688 ;
  assign n43162 = ~n24673 ;
  assign n24690 = n43162 & n24689 ;
  assign n43163 = ~n24690 ;
  assign n24691 = n143 & n43163 ;
  assign n23835 = n23801 | n23819 ;
  assign n43164 = ~n23835 ;
  assign n24466 = n43164 & n137 ;
  assign n24467 = n23607 | n24466 ;
  assign n43165 = ~n23801 ;
  assign n23807 = n23607 & n43165 ;
  assign n23808 = n42724 & n23807 ;
  assign n24468 = n23808 & n137 ;
  assign n43166 = ~n24468 ;
  assign n24469 = n24467 & n43166 ;
  assign n24674 = n143 | n24673 ;
  assign n43167 = ~n24674 ;
  assign n24692 = n43167 & n24689 ;
  assign n43168 = ~n24692 ;
  assign n24693 = n24469 & n43168 ;
  assign n43169 = ~n24691 ;
  assign n24694 = n43169 & n24693 ;
  assign n24696 = n24469 | n24692 ;
  assign n24697 = n43169 & n24696 ;
  assign n43170 = ~n24697 ;
  assign n24698 = n18797 & n43170 ;
  assign n23806 = n23769 & n42735 ;
  assign n43171 = ~n23821 ;
  assign n23833 = n23806 & n43171 ;
  assign n24496 = n23833 & n137 ;
  assign n23834 = n23804 | n23821 ;
  assign n43172 = ~n23834 ;
  assign n24510 = n43172 & n137 ;
  assign n24511 = n23769 | n24510 ;
  assign n43173 = ~n24496 ;
  assign n24512 = n43173 & n24511 ;
  assign n24703 = n43150 & n24684 ;
  assign n24704 = n24485 | n24703 ;
  assign n43174 = ~n24686 ;
  assign n24705 = n43174 & n24704 ;
  assign n43175 = ~n24705 ;
  assign n24706 = n142 & n43175 ;
  assign n24707 = n43161 & n24704 ;
  assign n24708 = n24633 | n24707 ;
  assign n43176 = ~n24706 ;
  assign n24709 = n43176 & n24708 ;
  assign n43177 = ~n24709 ;
  assign n24710 = n19362 & n43177 ;
  assign n24711 = n144 | n24710 ;
  assign n43178 = ~n24711 ;
  assign n24712 = n24696 & n43178 ;
  assign n24713 = n24512 | n24712 ;
  assign n43179 = ~n24698 ;
  assign n24714 = n43179 & n24713 ;
  assign n43180 = ~n24714 ;
  assign n24715 = n145 & n43180 ;
  assign n23859 = n23825 | n23843 ;
  assign n43181 = ~n23859 ;
  assign n24460 = n43181 & n137 ;
  assign n24461 = n23622 | n24460 ;
  assign n43182 = ~n23825 ;
  assign n23831 = n23622 & n43182 ;
  assign n23832 = n42741 & n23831 ;
  assign n24515 = n23832 & n137 ;
  assign n43183 = ~n24515 ;
  assign n24516 = n24461 & n43183 ;
  assign n24699 = n145 | n24698 ;
  assign n43184 = ~n24699 ;
  assign n24716 = n43184 & n24713 ;
  assign n24717 = n24516 | n24716 ;
  assign n43185 = ~n24715 ;
  assign n24718 = n43185 & n24717 ;
  assign n43186 = ~n24718 ;
  assign n24719 = n146 & n43186 ;
  assign n23858 = n23828 | n23845 ;
  assign n43187 = ~n23858 ;
  assign n24450 = n43187 & n137 ;
  assign n24451 = n23619 | n24450 ;
  assign n23830 = n23619 & n42751 ;
  assign n43188 = ~n23845 ;
  assign n23857 = n23830 & n43188 ;
  assign n24526 = n23857 & n137 ;
  assign n43189 = ~n24526 ;
  assign n24527 = n24451 & n43189 ;
  assign n24725 = n43167 & n24708 ;
  assign n24726 = n24469 | n24725 ;
  assign n43190 = ~n24710 ;
  assign n24727 = n43190 & n24726 ;
  assign n43191 = ~n24727 ;
  assign n24728 = n144 & n43191 ;
  assign n24729 = n43178 & n24726 ;
  assign n24730 = n24512 | n24729 ;
  assign n43192 = ~n24728 ;
  assign n24731 = n43192 & n24730 ;
  assign n43193 = ~n24731 ;
  assign n24732 = n145 & n43193 ;
  assign n24733 = n146 | n24732 ;
  assign n43194 = ~n24733 ;
  assign n24734 = n24717 & n43194 ;
  assign n24735 = n24527 | n24734 ;
  assign n43195 = ~n24719 ;
  assign n24736 = n43195 & n24735 ;
  assign n43196 = ~n24736 ;
  assign n24737 = n147 & n43196 ;
  assign n43197 = ~n23849 ;
  assign n23855 = n23660 & n43197 ;
  assign n23856 = n42757 & n23855 ;
  assign n24472 = n23856 & n137 ;
  assign n23883 = n23849 | n23867 ;
  assign n43198 = ~n23883 ;
  assign n24543 = n43198 & n137 ;
  assign n24544 = n23660 | n24543 ;
  assign n43199 = ~n24472 ;
  assign n24545 = n43199 & n24544 ;
  assign n24720 = n147 | n24719 ;
  assign n43200 = ~n24720 ;
  assign n24738 = n43200 & n24735 ;
  assign n24739 = n24545 | n24738 ;
  assign n43201 = ~n24737 ;
  assign n24740 = n43201 & n24739 ;
  assign n43202 = ~n24740 ;
  assign n24741 = n15807 & n43202 ;
  assign n23854 = n23634 & n42767 ;
  assign n43203 = ~n23869 ;
  assign n23881 = n23854 & n43203 ;
  assign n24477 = n23881 & n137 ;
  assign n23882 = n23852 | n23869 ;
  assign n43204 = ~n23882 ;
  assign n24498 = n43204 & n137 ;
  assign n24499 = n23634 | n24498 ;
  assign n43205 = ~n24477 ;
  assign n24500 = n43205 & n24499 ;
  assign n24751 = n43184 & n24730 ;
  assign n24752 = n24516 | n24751 ;
  assign n43206 = ~n24732 ;
  assign n24753 = n43206 & n24752 ;
  assign n43207 = ~n24753 ;
  assign n24754 = n146 & n43207 ;
  assign n24755 = n43194 & n24752 ;
  assign n24756 = n24527 | n24755 ;
  assign n43208 = ~n24754 ;
  assign n24757 = n43208 & n24756 ;
  assign n43209 = ~n24757 ;
  assign n24758 = n16322 & n43209 ;
  assign n24759 = n148 | n24758 ;
  assign n43210 = ~n24759 ;
  assign n24760 = n24739 & n43210 ;
  assign n24761 = n24500 | n24760 ;
  assign n43211 = ~n24741 ;
  assign n24762 = n43211 & n24761 ;
  assign n43212 = ~n24762 ;
  assign n24763 = n149 & n43212 ;
  assign n23907 = n23873 | n23891 ;
  assign n43213 = ~n23907 ;
  assign n24552 = n43213 & n137 ;
  assign n24553 = n23671 | n24552 ;
  assign n43214 = ~n23873 ;
  assign n23874 = n23671 & n43214 ;
  assign n23875 = n42773 & n23874 ;
  assign n24554 = n23875 & n137 ;
  assign n43215 = ~n24554 ;
  assign n24555 = n24553 & n43215 ;
  assign n24742 = n149 | n24741 ;
  assign n43216 = ~n24742 ;
  assign n24764 = n43216 & n24761 ;
  assign n24765 = n24555 | n24764 ;
  assign n43217 = ~n24763 ;
  assign n24766 = n43217 & n24765 ;
  assign n43218 = ~n24766 ;
  assign n24767 = n150 & n43218 ;
  assign n23880 = n23690 & n42783 ;
  assign n43219 = ~n23893 ;
  assign n23905 = n23880 & n43219 ;
  assign n24551 = n23905 & n137 ;
  assign n23906 = n23878 | n23893 ;
  assign n43220 = ~n23906 ;
  assign n24556 = n43220 & n137 ;
  assign n24557 = n23690 | n24556 ;
  assign n43221 = ~n24551 ;
  assign n24558 = n43221 & n24557 ;
  assign n24775 = n43200 & n24756 ;
  assign n24776 = n24545 | n24775 ;
  assign n43222 = ~n24758 ;
  assign n24777 = n43222 & n24776 ;
  assign n43223 = ~n24777 ;
  assign n24778 = n148 & n43223 ;
  assign n24779 = n43210 & n24776 ;
  assign n24780 = n24500 | n24779 ;
  assign n43224 = ~n24778 ;
  assign n24781 = n43224 & n24780 ;
  assign n43225 = ~n24781 ;
  assign n24782 = n149 & n43225 ;
  assign n24783 = n150 | n24782 ;
  assign n43226 = ~n24783 ;
  assign n24784 = n24765 & n43226 ;
  assign n24785 = n24558 | n24784 ;
  assign n43227 = ~n24767 ;
  assign n24786 = n43227 & n24785 ;
  assign n43228 = ~n24786 ;
  assign n24787 = n151 & n43228 ;
  assign n43229 = ~n23897 ;
  assign n23903 = n23677 & n43229 ;
  assign n23904 = n42789 & n23903 ;
  assign n24505 = n23904 & n137 ;
  assign n23931 = n23897 | n23915 ;
  assign n43230 = ~n23931 ;
  assign n24517 = n43230 & n137 ;
  assign n24518 = n23677 | n24517 ;
  assign n43231 = ~n24505 ;
  assign n24519 = n43231 & n24518 ;
  assign n24768 = n151 | n24767 ;
  assign n43232 = ~n24768 ;
  assign n24788 = n43232 & n24785 ;
  assign n24789 = n24519 | n24788 ;
  assign n43233 = ~n24787 ;
  assign n24790 = n43233 & n24789 ;
  assign n43234 = ~n24790 ;
  assign n24791 = n13079 & n43234 ;
  assign n23930 = n23900 | n23917 ;
  assign n43235 = ~n23930 ;
  assign n24524 = n43235 & n137 ;
  assign n24525 = n23688 | n24524 ;
  assign n23902 = n23688 & n42799 ;
  assign n43236 = ~n23917 ;
  assign n23929 = n23902 & n43236 ;
  assign n24561 = n23929 & n137 ;
  assign n43237 = ~n24561 ;
  assign n24562 = n24525 & n43237 ;
  assign n24799 = n43216 & n24780 ;
  assign n24800 = n24555 | n24799 ;
  assign n43238 = ~n24782 ;
  assign n24801 = n43238 & n24800 ;
  assign n43239 = ~n24801 ;
  assign n24802 = n150 & n43239 ;
  assign n24803 = n43226 & n24800 ;
  assign n24804 = n24558 | n24803 ;
  assign n43240 = ~n24802 ;
  assign n24805 = n43240 & n24804 ;
  assign n43241 = ~n24805 ;
  assign n24806 = n13662 & n43241 ;
  assign n24807 = n152 | n24806 ;
  assign n43242 = ~n24807 ;
  assign n24808 = n24789 & n43242 ;
  assign n24809 = n24562 | n24808 ;
  assign n43243 = ~n24791 ;
  assign n24810 = n43243 & n24809 ;
  assign n43244 = ~n24810 ;
  assign n24811 = n153 & n43244 ;
  assign n23955 = n23921 | n23939 ;
  assign n43245 = ~n23955 ;
  assign n24488 = n43245 & n137 ;
  assign n24489 = n23669 | n24488 ;
  assign n43246 = ~n23921 ;
  assign n23927 = n23669 & n43246 ;
  assign n23928 = n42805 & n23927 ;
  assign n24508 = n23928 & n137 ;
  assign n43247 = ~n24508 ;
  assign n24509 = n24489 & n43247 ;
  assign n24792 = n153 | n24791 ;
  assign n43248 = ~n24792 ;
  assign n24812 = n43248 & n24809 ;
  assign n24813 = n24509 | n24812 ;
  assign n43249 = ~n24811 ;
  assign n24814 = n43249 & n24813 ;
  assign n43250 = ~n24814 ;
  assign n24815 = n154 & n43250 ;
  assign n23954 = n23924 | n23941 ;
  assign n43251 = ~n23954 ;
  assign n24456 = n43251 & n137 ;
  assign n24457 = n23695 | n24456 ;
  assign n23926 = n23695 & n42815 ;
  assign n43252 = ~n23941 ;
  assign n23953 = n23926 & n43252 ;
  assign n24506 = n23953 & n137 ;
  assign n43253 = ~n24506 ;
  assign n24507 = n24457 & n43253 ;
  assign n24823 = n43232 & n24804 ;
  assign n24824 = n24519 | n24823 ;
  assign n43254 = ~n24806 ;
  assign n24825 = n43254 & n24824 ;
  assign n43255 = ~n24825 ;
  assign n24826 = n152 & n43255 ;
  assign n24827 = n43242 & n24824 ;
  assign n24828 = n24562 | n24827 ;
  assign n43256 = ~n24826 ;
  assign n24829 = n43256 & n24828 ;
  assign n43257 = ~n24829 ;
  assign n24830 = n153 & n43257 ;
  assign n24831 = n154 | n24830 ;
  assign n43258 = ~n24831 ;
  assign n24832 = n24813 & n43258 ;
  assign n24833 = n24507 | n24832 ;
  assign n43259 = ~n24815 ;
  assign n24834 = n43259 & n24833 ;
  assign n43260 = ~n24834 ;
  assign n24835 = n155 & n43260 ;
  assign n43261 = ~n23945 ;
  assign n23951 = n23686 & n43261 ;
  assign n23952 = n42821 & n23951 ;
  assign n24490 = n23952 & n137 ;
  assign n23979 = n23945 | n23963 ;
  assign n43262 = ~n23979 ;
  assign n24535 = n43262 & n137 ;
  assign n24536 = n23686 | n24535 ;
  assign n43263 = ~n24490 ;
  assign n24537 = n43263 & n24536 ;
  assign n24816 = n11067 | n24815 ;
  assign n43264 = ~n24816 ;
  assign n24836 = n43264 & n24833 ;
  assign n24837 = n24537 | n24836 ;
  assign n43265 = ~n24835 ;
  assign n24838 = n43265 & n24837 ;
  assign n43266 = ~n24838 ;
  assign n24839 = n10657 & n43266 ;
  assign n23950 = n23637 & n42831 ;
  assign n43267 = ~n23965 ;
  assign n23977 = n23950 & n43267 ;
  assign n24454 = n23977 & n137 ;
  assign n23978 = n23948 | n23965 ;
  assign n43268 = ~n23978 ;
  assign n24478 = n43268 & n137 ;
  assign n24479 = n23637 | n24478 ;
  assign n43269 = ~n24454 ;
  assign n24480 = n43269 & n24479 ;
  assign n24847 = n43248 & n24828 ;
  assign n24848 = n24509 | n24847 ;
  assign n43270 = ~n24830 ;
  assign n24849 = n43270 & n24848 ;
  assign n43271 = ~n24849 ;
  assign n24850 = n154 & n43271 ;
  assign n24851 = n43258 & n24848 ;
  assign n24852 = n24507 | n24851 ;
  assign n43272 = ~n24850 ;
  assign n24853 = n43272 & n24852 ;
  assign n43273 = ~n24853 ;
  assign n24854 = n11067 & n43273 ;
  assign n24855 = n10657 | n24854 ;
  assign n43274 = ~n24855 ;
  assign n24856 = n24837 & n43274 ;
  assign n24857 = n24480 | n24856 ;
  assign n43275 = ~n24839 ;
  assign n24858 = n43275 & n24857 ;
  assign n43276 = ~n24858 ;
  assign n24859 = n157 & n43276 ;
  assign n24003 = n23969 | n23987 ;
  assign n43277 = ~n24003 ;
  assign n24452 = n43277 & n137 ;
  assign n24453 = n23666 | n24452 ;
  assign n43278 = ~n23969 ;
  assign n23975 = n23666 & n43278 ;
  assign n23976 = n42837 & n23975 ;
  assign n24475 = n23976 & n137 ;
  assign n43279 = ~n24475 ;
  assign n24476 = n24453 & n43279 ;
  assign n24841 = n157 | n24839 ;
  assign n43280 = ~n24841 ;
  assign n24860 = n43280 & n24857 ;
  assign n24861 = n24476 | n24860 ;
  assign n43281 = ~n24859 ;
  assign n24862 = n43281 & n24861 ;
  assign n43282 = ~n24862 ;
  assign n24863 = n158 & n43282 ;
  assign n23973 = n23581 & n42847 ;
  assign n43283 = ~n23989 ;
  assign n24001 = n23973 & n43283 ;
  assign n24449 = n24001 & n137 ;
  assign n24002 = n23972 | n23989 ;
  assign n43284 = ~n24002 ;
  assign n24540 = n43284 & n137 ;
  assign n24541 = n23581 | n24540 ;
  assign n43285 = ~n24449 ;
  assign n24542 = n43285 & n24541 ;
  assign n24871 = n43264 & n24852 ;
  assign n24872 = n24537 | n24871 ;
  assign n43286 = ~n24854 ;
  assign n24873 = n43286 & n24872 ;
  assign n43287 = ~n24873 ;
  assign n24874 = n156 & n43287 ;
  assign n24875 = n43274 & n24872 ;
  assign n24876 = n24480 | n24875 ;
  assign n43288 = ~n24874 ;
  assign n24877 = n43288 & n24876 ;
  assign n43289 = ~n24877 ;
  assign n24878 = n157 & n43289 ;
  assign n24879 = n158 | n24878 ;
  assign n43290 = ~n24879 ;
  assign n24880 = n24861 & n43290 ;
  assign n24881 = n24542 | n24880 ;
  assign n43291 = ~n24863 ;
  assign n24882 = n43291 & n24881 ;
  assign n43292 = ~n24882 ;
  assign n24883 = n159 & n43292 ;
  assign n43293 = ~n23993 ;
  assign n23999 = n23662 & n43293 ;
  assign n24000 = n42853 & n23999 ;
  assign n24448 = n24000 & n137 ;
  assign n24027 = n23993 | n24011 ;
  assign n43294 = ~n24027 ;
  assign n24528 = n43294 & n137 ;
  assign n24529 = n23662 | n24528 ;
  assign n43295 = ~n24448 ;
  assign n24530 = n43295 & n24529 ;
  assign n24864 = n8857 | n24863 ;
  assign n43296 = ~n24864 ;
  assign n24884 = n43296 & n24881 ;
  assign n24885 = n24530 | n24884 ;
  assign n43297 = ~n24883 ;
  assign n24886 = n43297 & n24885 ;
  assign n43298 = ~n24886 ;
  assign n24887 = n8534 & n43298 ;
  assign n23998 = n23567 & n42863 ;
  assign n43299 = ~n24013 ;
  assign n24025 = n23998 & n43299 ;
  assign n24444 = n24025 & n137 ;
  assign n24026 = n23996 | n24013 ;
  assign n43300 = ~n24026 ;
  assign n24445 = n43300 & n137 ;
  assign n24446 = n23567 | n24445 ;
  assign n43301 = ~n24444 ;
  assign n24447 = n43301 & n24446 ;
  assign n24895 = n43280 & n24876 ;
  assign n24896 = n24476 | n24895 ;
  assign n43302 = ~n24878 ;
  assign n24897 = n43302 & n24896 ;
  assign n43303 = ~n24897 ;
  assign n24898 = n158 & n43303 ;
  assign n24899 = n43290 & n24896 ;
  assign n24900 = n24542 | n24899 ;
  assign n43304 = ~n24898 ;
  assign n24901 = n43304 & n24900 ;
  assign n43305 = ~n24901 ;
  assign n24902 = n8857 & n43305 ;
  assign n24903 = n160 | n24902 ;
  assign n43306 = ~n24903 ;
  assign n24904 = n24885 & n43306 ;
  assign n24905 = n24447 | n24904 ;
  assign n43307 = ~n24887 ;
  assign n24906 = n43307 & n24905 ;
  assign n43308 = ~n24906 ;
  assign n24907 = n161 & n43308 ;
  assign n43309 = ~n24017 ;
  assign n24023 = n23562 & n43309 ;
  assign n24024 = n42869 & n24023 ;
  assign n24436 = n24024 & n137 ;
  assign n24051 = n24017 | n24035 ;
  assign n43310 = ~n24051 ;
  assign n24439 = n43310 & n137 ;
  assign n24440 = n23562 | n24439 ;
  assign n43311 = ~n24436 ;
  assign n24441 = n43311 & n24440 ;
  assign n24888 = n161 | n24887 ;
  assign n43312 = ~n24888 ;
  assign n24908 = n43312 & n24905 ;
  assign n24909 = n24441 | n24908 ;
  assign n43313 = ~n24907 ;
  assign n24910 = n43313 & n24909 ;
  assign n43314 = ~n24910 ;
  assign n24911 = n162 & n43314 ;
  assign n24050 = n24020 | n24037 ;
  assign n43315 = ~n24050 ;
  assign n24437 = n43315 & n137 ;
  assign n24438 = n23586 | n24437 ;
  assign n24022 = n23586 & n42879 ;
  assign n43316 = ~n24037 ;
  assign n24049 = n24022 & n43316 ;
  assign n24522 = n24049 & n137 ;
  assign n43317 = ~n24522 ;
  assign n24523 = n24438 & n43317 ;
  assign n24919 = n43296 & n24900 ;
  assign n24920 = n24530 | n24919 ;
  assign n43318 = ~n24902 ;
  assign n24921 = n43318 & n24920 ;
  assign n43319 = ~n24921 ;
  assign n24922 = n160 & n43319 ;
  assign n24923 = n43306 & n24920 ;
  assign n24924 = n24447 | n24923 ;
  assign n43320 = ~n24922 ;
  assign n24925 = n43320 & n24924 ;
  assign n43321 = ~n24925 ;
  assign n24926 = n161 & n43321 ;
  assign n24927 = n162 | n24926 ;
  assign n43322 = ~n24927 ;
  assign n24928 = n24909 & n43322 ;
  assign n24929 = n24523 | n24928 ;
  assign n43323 = ~n24911 ;
  assign n24930 = n43323 & n24929 ;
  assign n43324 = ~n24930 ;
  assign n24931 = n163 & n43324 ;
  assign n43325 = ~n24041 ;
  assign n24047 = n23675 & n43325 ;
  assign n24048 = n42885 & n24047 ;
  assign n24427 = n24048 & n137 ;
  assign n24075 = n24041 | n24059 ;
  assign n43326 = ~n24075 ;
  assign n24433 = n43326 & n137 ;
  assign n24434 = n23675 | n24433 ;
  assign n43327 = ~n24427 ;
  assign n24435 = n43327 & n24434 ;
  assign n24912 = n6889 | n24911 ;
  assign n43328 = ~n24912 ;
  assign n24932 = n43328 & n24929 ;
  assign n24933 = n24435 | n24932 ;
  assign n43329 = ~n24931 ;
  assign n24934 = n43329 & n24933 ;
  assign n43330 = ~n24934 ;
  assign n24935 = n6600 & n43330 ;
  assign n24045 = n23570 & n42895 ;
  assign n43331 = ~n24061 ;
  assign n24073 = n24045 & n43331 ;
  assign n24420 = n24073 & n137 ;
  assign n24074 = n24044 | n24061 ;
  assign n43332 = ~n24074 ;
  assign n24424 = n43332 & n137 ;
  assign n24425 = n23570 | n24424 ;
  assign n43333 = ~n24420 ;
  assign n24426 = n43333 & n24425 ;
  assign n24941 = n43312 & n24924 ;
  assign n24942 = n24441 | n24941 ;
  assign n43334 = ~n24926 ;
  assign n24943 = n43334 & n24942 ;
  assign n43335 = ~n24943 ;
  assign n24944 = n162 & n43335 ;
  assign n24945 = n43322 & n24942 ;
  assign n24946 = n24523 | n24945 ;
  assign n43336 = ~n24944 ;
  assign n24947 = n43336 & n24946 ;
  assign n43337 = ~n24947 ;
  assign n24948 = n6889 & n43337 ;
  assign n24949 = n6600 | n24948 ;
  assign n43338 = ~n24949 ;
  assign n24950 = n24933 & n43338 ;
  assign n24951 = n24426 | n24950 ;
  assign n43339 = ~n24935 ;
  assign n24952 = n43339 & n24951 ;
  assign n43340 = ~n24952 ;
  assign n24953 = n165 & n43340 ;
  assign n24099 = n24065 | n24083 ;
  assign n43341 = ~n24099 ;
  assign n24415 = n43341 & n137 ;
  assign n24416 = n23556 | n24415 ;
  assign n43342 = ~n24065 ;
  assign n24071 = n23556 & n43342 ;
  assign n24072 = n42901 & n24071 ;
  assign n24417 = n24072 & n137 ;
  assign n43343 = ~n24417 ;
  assign n24418 = n24416 & n43343 ;
  assign n24936 = n165 | n24935 ;
  assign n43344 = ~n24936 ;
  assign n24954 = n43344 & n24951 ;
  assign n24955 = n24418 | n24954 ;
  assign n43345 = ~n24953 ;
  assign n24956 = n43345 & n24955 ;
  assign n43346 = ~n24956 ;
  assign n24957 = n166 & n43346 ;
  assign n24098 = n24068 | n24085 ;
  assign n43347 = ~n24098 ;
  assign n24531 = n43347 & n137 ;
  assign n24532 = n23609 | n24531 ;
  assign n24070 = n23609 & n42911 ;
  assign n43348 = ~n24085 ;
  assign n24097 = n24070 & n43348 ;
  assign n24533 = n24097 & n137 ;
  assign n43349 = ~n24533 ;
  assign n24534 = n24532 & n43349 ;
  assign n24967 = n43328 & n24946 ;
  assign n24968 = n24435 | n24967 ;
  assign n43350 = ~n24948 ;
  assign n24969 = n43350 & n24968 ;
  assign n43351 = ~n24969 ;
  assign n24970 = n164 & n43351 ;
  assign n24971 = n43338 & n24968 ;
  assign n24972 = n24426 | n24971 ;
  assign n43352 = ~n24970 ;
  assign n24973 = n43352 & n24972 ;
  assign n43353 = ~n24973 ;
  assign n24974 = n165 & n43353 ;
  assign n24975 = n166 | n24974 ;
  assign n43354 = ~n24975 ;
  assign n24976 = n24955 & n43354 ;
  assign n24977 = n24534 | n24976 ;
  assign n43355 = ~n24957 ;
  assign n24978 = n43355 & n24977 ;
  assign n43356 = ~n24978 ;
  assign n24979 = n167 & n43356 ;
  assign n43357 = ~n24089 ;
  assign n24095 = n23599 & n43357 ;
  assign n24096 = n42917 & n24095 ;
  assign n24414 = n24096 & n137 ;
  assign n24123 = n24089 | n24107 ;
  assign n43358 = ~n24123 ;
  assign n24502 = n43358 & n137 ;
  assign n24503 = n23599 | n24502 ;
  assign n43359 = ~n24414 ;
  assign n24504 = n43359 & n24503 ;
  assign n24958 = n5352 | n24957 ;
  assign n43360 = ~n24958 ;
  assign n24980 = n43360 & n24977 ;
  assign n24981 = n24504 | n24980 ;
  assign n43361 = ~n24979 ;
  assign n24982 = n43361 & n24981 ;
  assign n43362 = ~n24982 ;
  assign n24983 = n4934 & n43362 ;
  assign n24122 = n24092 | n24109 ;
  assign n43363 = ~n24122 ;
  assign n24473 = n43363 & n137 ;
  assign n24474 = n23595 | n24473 ;
  assign n24094 = n23595 & n42927 ;
  assign n43364 = ~n24109 ;
  assign n24121 = n24094 & n43364 ;
  assign n24564 = n24121 & n137 ;
  assign n43365 = ~n24564 ;
  assign n24565 = n24474 & n43365 ;
  assign n24991 = n43344 & n24972 ;
  assign n24992 = n24418 | n24991 ;
  assign n43366 = ~n24974 ;
  assign n24993 = n43366 & n24992 ;
  assign n43367 = ~n24993 ;
  assign n24994 = n166 & n43367 ;
  assign n24995 = n43354 & n24992 ;
  assign n24996 = n24534 | n24995 ;
  assign n43368 = ~n24994 ;
  assign n24997 = n43368 & n24996 ;
  assign n43369 = ~n24997 ;
  assign n24998 = n5352 & n43369 ;
  assign n24999 = n4934 | n24998 ;
  assign n43370 = ~n24999 ;
  assign n25000 = n24981 & n43370 ;
  assign n25001 = n24565 | n25000 ;
  assign n43371 = ~n24983 ;
  assign n25002 = n43371 & n25001 ;
  assign n43372 = ~n25002 ;
  assign n25003 = n169 & n43372 ;
  assign n43373 = ~n24113 ;
  assign n24119 = n23682 & n43373 ;
  assign n24120 = n42933 & n24119 ;
  assign n24566 = n24120 & n137 ;
  assign n24147 = n24113 | n24131 ;
  assign n43374 = ~n24147 ;
  assign n24567 = n43374 & n137 ;
  assign n24568 = n23682 | n24567 ;
  assign n43375 = ~n24566 ;
  assign n24569 = n43375 & n24568 ;
  assign n24984 = n169 | n24983 ;
  assign n43376 = ~n24984 ;
  assign n25004 = n43376 & n25001 ;
  assign n25005 = n24569 | n25004 ;
  assign n43377 = ~n25003 ;
  assign n25006 = n43377 & n25005 ;
  assign n43378 = ~n25006 ;
  assign n25007 = n170 & n43378 ;
  assign n24146 = n24116 | n24133 ;
  assign n43379 = ~n24146 ;
  assign n24559 = n43379 & n137 ;
  assign n24560 = n23697 | n24559 ;
  assign n24118 = n23697 & n42943 ;
  assign n43380 = ~n24133 ;
  assign n24145 = n24118 & n43380 ;
  assign n24570 = n24145 & n137 ;
  assign n43381 = ~n24570 ;
  assign n24571 = n24560 & n43381 ;
  assign n25015 = n43360 & n24996 ;
  assign n25016 = n24504 | n25015 ;
  assign n43382 = ~n24998 ;
  assign n25017 = n43382 & n25016 ;
  assign n43383 = ~n25017 ;
  assign n25018 = n168 & n43383 ;
  assign n25019 = n43370 & n25016 ;
  assign n25020 = n24565 | n25019 ;
  assign n43384 = ~n25018 ;
  assign n25021 = n43384 & n25020 ;
  assign n43385 = ~n25021 ;
  assign n25022 = n169 & n43385 ;
  assign n25023 = n170 | n25022 ;
  assign n43386 = ~n25023 ;
  assign n25024 = n25005 & n43386 ;
  assign n25025 = n24571 | n25024 ;
  assign n43387 = ~n25007 ;
  assign n25026 = n43387 & n25025 ;
  assign n43388 = ~n25026 ;
  assign n25027 = n171 & n43388 ;
  assign n24171 = n24137 | n24155 ;
  assign n43389 = ~n24171 ;
  assign n24421 = n43389 & n137 ;
  assign n24422 = n23702 | n24421 ;
  assign n43390 = ~n24137 ;
  assign n24143 = n23702 & n43390 ;
  assign n24144 = n42949 & n24143 ;
  assign n24428 = n24144 & n137 ;
  assign n43391 = ~n24428 ;
  assign n24429 = n24422 & n43391 ;
  assign n25008 = n3940 | n25007 ;
  assign n43392 = ~n25008 ;
  assign n25028 = n43392 & n25025 ;
  assign n25029 = n24429 | n25028 ;
  assign n43393 = ~n25027 ;
  assign n25030 = n43393 & n25029 ;
  assign n43394 = ~n25030 ;
  assign n25031 = n3631 & n43394 ;
  assign n24142 = n23706 & n42959 ;
  assign n43395 = ~n24157 ;
  assign n24169 = n24142 & n43395 ;
  assign n24419 = n24169 & n137 ;
  assign n24170 = n24140 | n24157 ;
  assign n43396 = ~n24170 ;
  assign n24430 = n43396 & n137 ;
  assign n24431 = n23706 | n24430 ;
  assign n43397 = ~n24419 ;
  assign n24432 = n43397 & n24431 ;
  assign n25037 = n43376 & n25020 ;
  assign n25038 = n24569 | n25037 ;
  assign n43398 = ~n25022 ;
  assign n25039 = n43398 & n25038 ;
  assign n43399 = ~n25039 ;
  assign n25040 = n170 & n43399 ;
  assign n25041 = n43386 & n25038 ;
  assign n25042 = n24571 | n25041 ;
  assign n43400 = ~n25040 ;
  assign n25043 = n43400 & n25042 ;
  assign n43401 = ~n25043 ;
  assign n25044 = n3940 & n43401 ;
  assign n25045 = n3631 | n25044 ;
  assign n43402 = ~n25045 ;
  assign n25046 = n25029 & n43402 ;
  assign n25047 = n24432 | n25046 ;
  assign n43403 = ~n25031 ;
  assign n25048 = n43403 & n25047 ;
  assign n43404 = ~n25048 ;
  assign n25049 = n173 & n43404 ;
  assign n24195 = n24161 | n24179 ;
  assign n43405 = ~n24195 ;
  assign n24442 = n43405 & n137 ;
  assign n24443 = n23712 | n24442 ;
  assign n43406 = ~n24161 ;
  assign n24167 = n23712 & n43406 ;
  assign n24168 = n42965 & n24167 ;
  assign n24572 = n24168 & n137 ;
  assign n43407 = ~n24572 ;
  assign n24573 = n24443 & n43407 ;
  assign n25032 = n173 | n25031 ;
  assign n43408 = ~n25032 ;
  assign n25050 = n43408 & n25047 ;
  assign n25051 = n24573 | n25050 ;
  assign n43409 = ~n25049 ;
  assign n25052 = n43409 & n25051 ;
  assign n43410 = ~n25052 ;
  assign n25053 = n174 & n43410 ;
  assign n24194 = n24164 | n24181 ;
  assign n43411 = ~n24194 ;
  assign n24462 = n43411 & n137 ;
  assign n24463 = n23692 | n24462 ;
  assign n24166 = n23692 & n42975 ;
  assign n43412 = ~n24181 ;
  assign n24193 = n24166 & n43412 ;
  assign n24574 = n24193 & n137 ;
  assign n43413 = ~n24574 ;
  assign n24575 = n24463 & n43413 ;
  assign n25063 = n43392 & n25042 ;
  assign n25064 = n24429 | n25063 ;
  assign n43414 = ~n25044 ;
  assign n25065 = n43414 & n25064 ;
  assign n43415 = ~n25065 ;
  assign n25066 = n172 & n43415 ;
  assign n25067 = n43402 & n25064 ;
  assign n25068 = n24432 | n25067 ;
  assign n43416 = ~n25066 ;
  assign n25069 = n43416 & n25068 ;
  assign n43417 = ~n25069 ;
  assign n25070 = n173 & n43417 ;
  assign n25071 = n174 | n25070 ;
  assign n43418 = ~n25071 ;
  assign n25072 = n25051 & n43418 ;
  assign n25073 = n24575 | n25072 ;
  assign n43419 = ~n25053 ;
  assign n25074 = n43419 & n25073 ;
  assign n43420 = ~n25074 ;
  assign n25075 = n175 & n43420 ;
  assign n43421 = ~n24185 ;
  assign n24191 = n23715 & n43421 ;
  assign n24192 = n42981 & n24191 ;
  assign n24423 = n24192 & n137 ;
  assign n24219 = n24185 | n24203 ;
  assign n43422 = ~n24219 ;
  assign n24578 = n43422 & n137 ;
  assign n24579 = n23715 | n24578 ;
  assign n43423 = ~n24423 ;
  assign n24580 = n43423 & n24579 ;
  assign n25054 = n2753 | n25053 ;
  assign n43424 = ~n25054 ;
  assign n25076 = n43424 & n25073 ;
  assign n25077 = n24580 | n25076 ;
  assign n43425 = ~n25075 ;
  assign n25078 = n43425 & n25077 ;
  assign n43426 = ~n25078 ;
  assign n25079 = n2431 & n43426 ;
  assign n24218 = n24188 | n24205 ;
  assign n43427 = ~n24218 ;
  assign n24581 = n43427 & n137 ;
  assign n24582 = n23656 | n24581 ;
  assign n24190 = n23656 & n42991 ;
  assign n43428 = ~n24205 ;
  assign n24217 = n24190 & n43428 ;
  assign n24583 = n24217 & n137 ;
  assign n43429 = ~n24583 ;
  assign n24584 = n24582 & n43429 ;
  assign n25087 = n43408 & n25068 ;
  assign n25088 = n24573 | n25087 ;
  assign n43430 = ~n25070 ;
  assign n25089 = n43430 & n25088 ;
  assign n43431 = ~n25089 ;
  assign n25090 = n174 & n43431 ;
  assign n25091 = n43418 & n25088 ;
  assign n25092 = n24575 | n25091 ;
  assign n43432 = ~n25090 ;
  assign n25093 = n43432 & n25092 ;
  assign n43433 = ~n25093 ;
  assign n25094 = n2753 & n43433 ;
  assign n25095 = n2431 | n25094 ;
  assign n43434 = ~n25095 ;
  assign n25096 = n25077 & n43434 ;
  assign n25097 = n24584 | n25096 ;
  assign n43435 = ~n25079 ;
  assign n25098 = n43435 & n25097 ;
  assign n43436 = ~n25098 ;
  assign n25099 = n177 & n43436 ;
  assign n24243 = n24209 | n24227 ;
  assign n43437 = ~n24243 ;
  assign n24513 = n43437 & n137 ;
  assign n24514 = n23718 | n24513 ;
  assign n43438 = ~n24209 ;
  assign n24215 = n23718 & n43438 ;
  assign n24216 = n42997 & n24215 ;
  assign n24585 = n24216 & n137 ;
  assign n43439 = ~n24585 ;
  assign n24586 = n24514 & n43439 ;
  assign n25080 = n177 | n25079 ;
  assign n43440 = ~n25080 ;
  assign n25100 = n43440 & n25097 ;
  assign n25101 = n24586 | n25100 ;
  assign n43441 = ~n25099 ;
  assign n25102 = n43441 & n25101 ;
  assign n43442 = ~n25102 ;
  assign n25103 = n178 & n43442 ;
  assign n24242 = n24212 | n24229 ;
  assign n43443 = ~n24242 ;
  assign n24589 = n43443 & n137 ;
  assign n24590 = n23710 | n24589 ;
  assign n24214 = n23710 & n43007 ;
  assign n43444 = ~n24229 ;
  assign n24241 = n24214 & n43444 ;
  assign n24591 = n24241 & n137 ;
  assign n43445 = ~n24591 ;
  assign n24592 = n24590 & n43445 ;
  assign n25111 = n43424 & n25092 ;
  assign n25112 = n24580 | n25111 ;
  assign n43446 = ~n25094 ;
  assign n25113 = n43446 & n25112 ;
  assign n43447 = ~n25113 ;
  assign n25114 = n176 & n43447 ;
  assign n25115 = n43434 & n25112 ;
  assign n25116 = n24584 | n25115 ;
  assign n43448 = ~n25114 ;
  assign n25117 = n43448 & n25116 ;
  assign n43449 = ~n25117 ;
  assign n25118 = n177 & n43449 ;
  assign n25119 = n178 | n25118 ;
  assign n43450 = ~n25119 ;
  assign n25120 = n25101 & n43450 ;
  assign n25121 = n24592 | n25120 ;
  assign n43451 = ~n25103 ;
  assign n25122 = n43451 & n25121 ;
  assign n43452 = ~n25122 ;
  assign n25123 = n179 & n43452 ;
  assign n43453 = ~n24233 ;
  assign n24239 = n23725 & n43453 ;
  assign n24240 = n43013 & n24239 ;
  assign n24501 = n24240 & n137 ;
  assign n24267 = n24233 | n24251 ;
  assign n43454 = ~n24267 ;
  assign n24548 = n43454 & n137 ;
  assign n24549 = n23725 | n24548 ;
  assign n43455 = ~n24501 ;
  assign n24550 = n43455 & n24549 ;
  assign n25104 = n1707 | n25103 ;
  assign n43456 = ~n25104 ;
  assign n25124 = n43456 & n25121 ;
  assign n25125 = n24550 | n25124 ;
  assign n43457 = ~n25123 ;
  assign n25126 = n43457 & n25125 ;
  assign n43458 = ~n25126 ;
  assign n25127 = n1487 & n43458 ;
  assign n24266 = n24236 | n24253 ;
  assign n43459 = ~n24266 ;
  assign n24593 = n43459 & n137 ;
  assign n24594 = n23728 | n24593 ;
  assign n24238 = n23728 & n43023 ;
  assign n43460 = ~n24253 ;
  assign n24265 = n24238 & n43460 ;
  assign n24595 = n24265 & n137 ;
  assign n43461 = ~n24595 ;
  assign n24596 = n24594 & n43461 ;
  assign n25133 = n43440 & n25116 ;
  assign n25134 = n24586 | n25133 ;
  assign n43462 = ~n25118 ;
  assign n25135 = n43462 & n25134 ;
  assign n43463 = ~n25135 ;
  assign n25136 = n178 & n43463 ;
  assign n25137 = n43450 & n25134 ;
  assign n25138 = n24592 | n25137 ;
  assign n43464 = ~n25136 ;
  assign n25139 = n43464 & n25138 ;
  assign n43465 = ~n25139 ;
  assign n25140 = n1707 & n43465 ;
  assign n25141 = n1487 | n25140 ;
  assign n43466 = ~n25141 ;
  assign n25142 = n25125 & n43466 ;
  assign n25143 = n24596 | n25142 ;
  assign n43467 = ~n25127 ;
  assign n25144 = n43467 & n25143 ;
  assign n43468 = ~n25144 ;
  assign n25145 = n181 & n43468 ;
  assign n24291 = n24257 | n24275 ;
  assign n43469 = ~n24291 ;
  assign n24597 = n43469 & n137 ;
  assign n24598 = n23730 | n24597 ;
  assign n43470 = ~n24257 ;
  assign n24263 = n23730 & n43470 ;
  assign n24264 = n43029 & n24263 ;
  assign n24599 = n24264 & n137 ;
  assign n43471 = ~n24599 ;
  assign n24600 = n24598 & n43471 ;
  assign n25128 = n181 | n25127 ;
  assign n43472 = ~n25128 ;
  assign n25146 = n43472 & n25143 ;
  assign n25147 = n24600 | n25146 ;
  assign n43473 = ~n25145 ;
  assign n25148 = n43473 & n25147 ;
  assign n43474 = ~n25148 ;
  assign n25149 = n182 & n43474 ;
  assign n24290 = n24260 | n24277 ;
  assign n43475 = ~n24290 ;
  assign n24486 = n43475 & n137 ;
  assign n24487 = n23733 | n24486 ;
  assign n24262 = n23733 & n43039 ;
  assign n43476 = ~n24277 ;
  assign n24289 = n24262 & n43476 ;
  assign n24520 = n24289 & n137 ;
  assign n43477 = ~n24520 ;
  assign n24521 = n24487 & n43477 ;
  assign n25159 = n43456 & n25138 ;
  assign n25160 = n24550 | n25159 ;
  assign n43478 = ~n25140 ;
  assign n25161 = n43478 & n25160 ;
  assign n43479 = ~n25161 ;
  assign n25162 = n180 & n43479 ;
  assign n25163 = n43466 & n25160 ;
  assign n25164 = n24596 | n25163 ;
  assign n43480 = ~n25162 ;
  assign n25165 = n43480 & n25164 ;
  assign n43481 = ~n25165 ;
  assign n25166 = n181 & n43481 ;
  assign n25167 = n182 | n25166 ;
  assign n43482 = ~n25167 ;
  assign n25168 = n25147 & n43482 ;
  assign n25169 = n24521 | n25168 ;
  assign n43483 = ~n25149 ;
  assign n25170 = n43483 & n25169 ;
  assign n43484 = ~n25170 ;
  assign n25171 = n183 & n43484 ;
  assign n24315 = n24281 | n24299 ;
  assign n43485 = ~n24315 ;
  assign n24458 = n43485 & n137 ;
  assign n24459 = n23736 | n24458 ;
  assign n43486 = ~n24281 ;
  assign n24287 = n23736 & n43486 ;
  assign n24288 = n43045 & n24287 ;
  assign n24601 = n24288 & n137 ;
  assign n43487 = ~n24601 ;
  assign n24602 = n24459 & n43487 ;
  assign n25150 = n183 | n25149 ;
  assign n43488 = ~n25150 ;
  assign n25172 = n43488 & n25169 ;
  assign n25173 = n24602 | n25172 ;
  assign n43489 = ~n25171 ;
  assign n25174 = n43489 & n25173 ;
  assign n43490 = ~n25174 ;
  assign n25175 = n838 & n43490 ;
  assign n24314 = n24284 | n24301 ;
  assign n43491 = ~n24314 ;
  assign n24603 = n43491 & n137 ;
  assign n24604 = n23738 | n24603 ;
  assign n24286 = n23738 & n43055 ;
  assign n43492 = ~n24301 ;
  assign n24313 = n24286 & n43492 ;
  assign n24605 = n24313 & n137 ;
  assign n43493 = ~n24605 ;
  assign n24606 = n24604 & n43493 ;
  assign n25183 = n43472 & n25164 ;
  assign n25184 = n24600 | n25183 ;
  assign n43494 = ~n25166 ;
  assign n25185 = n43494 & n25184 ;
  assign n43495 = ~n25185 ;
  assign n25186 = n182 & n43495 ;
  assign n25187 = n43482 & n25184 ;
  assign n25188 = n24521 | n25187 ;
  assign n43496 = ~n25186 ;
  assign n25189 = n43496 & n25188 ;
  assign n43497 = ~n25189 ;
  assign n25190 = n996 & n43497 ;
  assign n25191 = n838 | n25190 ;
  assign n43498 = ~n25191 ;
  assign n25192 = n25173 & n43498 ;
  assign n25193 = n24606 | n25192 ;
  assign n43499 = ~n25175 ;
  assign n25194 = n43499 & n25193 ;
  assign n43500 = ~n25194 ;
  assign n25195 = n185 & n43500 ;
  assign n24339 = n24305 | n24323 ;
  assign n43501 = ~n24339 ;
  assign n24607 = n43501 & n137 ;
  assign n24608 = n23742 | n24607 ;
  assign n43502 = ~n24305 ;
  assign n24311 = n23742 & n43502 ;
  assign n24312 = n43061 & n24311 ;
  assign n24610 = n24312 & n137 ;
  assign n43503 = ~n24610 ;
  assign n24611 = n24608 & n43503 ;
  assign n25176 = n185 | n25175 ;
  assign n43504 = ~n25176 ;
  assign n25196 = n43504 & n25193 ;
  assign n25197 = n24611 | n25196 ;
  assign n43505 = ~n25195 ;
  assign n25198 = n43505 & n25197 ;
  assign n43506 = ~n25198 ;
  assign n25199 = n186 & n43506 ;
  assign n24310 = n23745 & n43071 ;
  assign n43507 = ~n24325 ;
  assign n24337 = n24310 & n43507 ;
  assign n24563 = n24337 & n137 ;
  assign n24338 = n24308 | n24325 ;
  assign n43508 = ~n24338 ;
  assign n24612 = n43508 & n137 ;
  assign n24613 = n23745 | n24612 ;
  assign n43509 = ~n24563 ;
  assign n24614 = n43509 & n24613 ;
  assign n25207 = n43488 & n25188 ;
  assign n25208 = n24602 | n25207 ;
  assign n43510 = ~n25190 ;
  assign n25209 = n43510 & n25208 ;
  assign n43511 = ~n25209 ;
  assign n25210 = n184 & n43511 ;
  assign n25211 = n43498 & n25208 ;
  assign n25212 = n24606 | n25211 ;
  assign n43512 = ~n25210 ;
  assign n25213 = n43512 & n25212 ;
  assign n43513 = ~n25213 ;
  assign n25214 = n185 & n43513 ;
  assign n25215 = n186 | n25214 ;
  assign n43514 = ~n25215 ;
  assign n25216 = n25197 & n43514 ;
  assign n25217 = n24614 | n25216 ;
  assign n43515 = ~n25199 ;
  assign n25218 = n43515 & n25217 ;
  assign n43516 = ~n25218 ;
  assign n25219 = n187 & n43516 ;
  assign n43517 = ~n24329 ;
  assign n24335 = n23627 & n43517 ;
  assign n24336 = n43077 & n24335 ;
  assign n24497 = n24336 & n137 ;
  assign n24363 = n24329 | n24347 ;
  assign n43518 = ~n24363 ;
  assign n24615 = n43518 & n137 ;
  assign n24616 = n23627 | n24615 ;
  assign n43519 = ~n24497 ;
  assign n24617 = n43519 & n24616 ;
  assign n25200 = n528 | n25199 ;
  assign n43520 = ~n25200 ;
  assign n25220 = n43520 & n25217 ;
  assign n25221 = n24617 | n25220 ;
  assign n43521 = ~n25219 ;
  assign n25222 = n43521 & n25221 ;
  assign n43522 = ~n25222 ;
  assign n25223 = n413 & n43522 ;
  assign n24362 = n24332 | n24349 ;
  assign n43523 = ~n24362 ;
  assign n24464 = n43523 & n137 ;
  assign n24465 = n23749 | n24464 ;
  assign n24333 = n23749 & n43087 ;
  assign n43524 = ~n24349 ;
  assign n24361 = n24333 & n43524 ;
  assign n24576 = n24361 & n137 ;
  assign n43525 = ~n24576 ;
  assign n24577 = n24465 & n43525 ;
  assign n25229 = n43504 & n25212 ;
  assign n25230 = n24611 | n25229 ;
  assign n43526 = ~n25214 ;
  assign n25231 = n43526 & n25230 ;
  assign n43527 = ~n25231 ;
  assign n25232 = n186 & n43527 ;
  assign n25233 = n43514 & n25230 ;
  assign n25234 = n24614 | n25233 ;
  assign n43528 = ~n25232 ;
  assign n25235 = n43528 & n25234 ;
  assign n43529 = ~n25235 ;
  assign n25236 = n528 & n43529 ;
  assign n25237 = n413 | n25236 ;
  assign n43530 = ~n25237 ;
  assign n25238 = n25221 & n43530 ;
  assign n25239 = n24577 | n25238 ;
  assign n43531 = ~n25223 ;
  assign n25240 = n43531 & n25239 ;
  assign n43532 = ~n25240 ;
  assign n25241 = n189 & n43532 ;
  assign n24386 = n24353 | n24371 ;
  assign n43533 = ~n24386 ;
  assign n24618 = n43533 & n137 ;
  assign n24619 = n23612 | n24618 ;
  assign n43534 = ~n24353 ;
  assign n24359 = n23612 & n43534 ;
  assign n24360 = n43093 & n24359 ;
  assign n24621 = n24360 & n137 ;
  assign n43535 = ~n24621 ;
  assign n24622 = n24619 & n43535 ;
  assign n25224 = n189 | n25223 ;
  assign n43536 = ~n25224 ;
  assign n25242 = n43536 & n25239 ;
  assign n25243 = n24622 | n25242 ;
  assign n43537 = ~n25241 ;
  assign n25244 = n43537 & n25243 ;
  assign n43538 = ~n25244 ;
  assign n25245 = n190 & n43538 ;
  assign n24385 = n24356 | n24373 ;
  assign n43539 = ~n24385 ;
  assign n24470 = n43539 & n137 ;
  assign n24471 = n23720 | n24470 ;
  assign n24358 = n23720 & n43103 ;
  assign n43540 = ~n24373 ;
  assign n24384 = n24358 & n43540 ;
  assign n24587 = n24384 & n137 ;
  assign n43541 = ~n24587 ;
  assign n24588 = n24471 & n43541 ;
  assign n25253 = n43520 & n25234 ;
  assign n25254 = n24617 | n25253 ;
  assign n43542 = ~n25236 ;
  assign n25255 = n43542 & n25254 ;
  assign n43543 = ~n25255 ;
  assign n25256 = n188 & n43543 ;
  assign n25257 = n43530 & n25254 ;
  assign n25258 = n24577 | n25257 ;
  assign n43544 = ~n25256 ;
  assign n25259 = n43544 & n25258 ;
  assign n43545 = ~n25259 ;
  assign n25260 = n189 & n43545 ;
  assign n25261 = n190 | n25260 ;
  assign n43546 = ~n25261 ;
  assign n25262 = n25243 & n43546 ;
  assign n25263 = n24588 | n25262 ;
  assign n43547 = ~n25245 ;
  assign n25268 = n43547 & n25263 ;
  assign n43548 = ~n25268 ;
  assign n25269 = n191 & n43548 ;
  assign n24398 = n24377 | n24394 ;
  assign n43549 = ~n24398 ;
  assign n24623 = n43549 & n137 ;
  assign n24624 = n23752 | n24623 ;
  assign n43550 = ~n24377 ;
  assign n24382 = n23752 & n43550 ;
  assign n24383 = n43109 & n24382 ;
  assign n24625 = n24383 & n137 ;
  assign n43551 = ~n24625 ;
  assign n24626 = n24624 & n43551 ;
  assign n25246 = n191 | n25245 ;
  assign n43552 = ~n25246 ;
  assign n25271 = n43552 & n25263 ;
  assign n25272 = n24626 | n25271 ;
  assign n43553 = ~n25269 ;
  assign n25273 = n43553 & n25272 ;
  assign n24407 = n23757 | n24406 ;
  assign n43554 = ~n24407 ;
  assign n24627 = n43554 & n137 ;
  assign n25281 = n24411 | n24627 ;
  assign n24403 = n43120 & n24402 ;
  assign n43555 = ~n24396 ;
  assign n24404 = n43555 & n24403 ;
  assign n24620 = n24404 & n137 ;
  assign n24397 = n24380 | n24396 ;
  assign n43556 = ~n24397 ;
  assign n24609 = n43556 & n137 ;
  assign n25292 = n24402 | n24609 ;
  assign n43557 = ~n24620 ;
  assign n25293 = n43557 & n25292 ;
  assign n25294 = n25281 | n25293 ;
  assign n25295 = n25273 | n25294 ;
  assign n25296 = n31336 & n25295 ;
  assign n24408 = n192 & n24407 ;
  assign n43558 = ~n23757 ;
  assign n24628 = n43558 & n137 ;
  assign n43559 = ~n24628 ;
  assign n24629 = n24406 & n43559 ;
  assign n43560 = ~n24629 ;
  assign n24630 = n24408 & n43560 ;
  assign n23754 = n23540 | n23753 ;
  assign n43561 = ~n23754 ;
  assign n23758 = n43561 & n23756 ;
  assign n23764 = n23758 & n43136 ;
  assign n25282 = n23764 & n43137 ;
  assign n25283 = n43138 & n25282 ;
  assign n25284 = n24630 | n25283 ;
  assign n25301 = n43553 & n25293 ;
  assign n25302 = n25272 & n25301 ;
  assign n25303 = n25284 | n25302 ;
  assign n136 = n25296 | n25303 ;
  assign n25435 = n24694 & n136 ;
  assign n24695 = n24691 | n24692 ;
  assign n43562 = ~n24695 ;
  assign n25438 = n43562 & n136 ;
  assign n25439 = n24469 | n25438 ;
  assign n43563 = ~n25435 ;
  assign n25440 = n43563 & n25439 ;
  assign n251 = x12 | x13 ;
  assign n252 = x14 | n251 ;
  assign n23541 = n252 & n43135 ;
  assign n23762 = n23541 & n43136 ;
  assign n25290 = n23762 & n43137 ;
  assign n25291 = n43138 & n25290 ;
  assign n25400 = x14 & n136 ;
  assign n43564 = ~n25400 ;
  assign n25401 = n25291 & n43564 ;
  assign n43565 = ~n248 ;
  assign n25379 = n43565 & n136 ;
  assign n43566 = ~x14 ;
  assign n25405 = n43566 & n136 ;
  assign n43567 = ~n25405 ;
  assign n25406 = x15 & n43567 ;
  assign n25407 = n25379 | n25406 ;
  assign n25408 = n25401 | n25407 ;
  assign n253 = n43566 & n251 ;
  assign n25247 = n287 | n25245 ;
  assign n43568 = ~n25247 ;
  assign n25264 = n43568 & n25263 ;
  assign n25265 = n24626 | n25264 ;
  assign n25270 = n25265 & n43553 ;
  assign n25297 = n25270 | n25294 ;
  assign n25298 = n31336 & n25297 ;
  assign n25515 = n25265 & n25301 ;
  assign n25516 = n25284 | n25515 ;
  assign n25517 = n25298 | n25516 ;
  assign n43569 = ~n25517 ;
  assign n25536 = x14 & n43569 ;
  assign n25537 = n253 | n25536 ;
  assign n43570 = ~n25537 ;
  assign n25538 = n137 & n43570 ;
  assign n43571 = ~n25538 ;
  assign n25539 = n25408 & n43571 ;
  assign n43572 = ~n25539 ;
  assign n25540 = n138 & n43572 ;
  assign n25413 = n252 & n43564 ;
  assign n43573 = ~n25413 ;
  assign n25414 = n137 & n43573 ;
  assign n25415 = n138 | n25414 ;
  assign n43574 = ~n25415 ;
  assign n25416 = n25408 & n43574 ;
  assign n43575 = ~n25283 ;
  assign n25287 = n137 & n43575 ;
  assign n43576 = ~n24630 ;
  assign n25288 = n43576 & n25287 ;
  assign n43577 = ~n25515 ;
  assign n25553 = n25288 & n43577 ;
  assign n43578 = ~n25296 ;
  assign n25554 = n43578 & n25553 ;
  assign n25555 = n25379 | n25554 ;
  assign n25556 = x16 & n25555 ;
  assign n25557 = x16 | n25554 ;
  assign n25558 = n25379 | n25557 ;
  assign n43579 = ~n25556 ;
  assign n25559 = n43579 & n25558 ;
  assign n25560 = n25416 | n25559 ;
  assign n43580 = ~n25540 ;
  assign n25561 = n43580 & n25560 ;
  assign n43581 = ~n25561 ;
  assign n25562 = n22661 & n43581 ;
  assign n24638 = n24631 | n24636 ;
  assign n43582 = ~n24638 ;
  assign n24650 = n43582 & n24641 ;
  assign n25309 = n24650 & n136 ;
  assign n25384 = n43582 & n136 ;
  assign n25385 = n24641 | n25384 ;
  assign n43583 = ~n25309 ;
  assign n25386 = n43583 & n25385 ;
  assign n43584 = ~n25414 ;
  assign n25417 = n25408 & n43584 ;
  assign n43585 = ~n25417 ;
  assign n25418 = n138 & n43585 ;
  assign n25419 = n22661 | n25418 ;
  assign n25544 = n138 | n25538 ;
  assign n43586 = ~n25544 ;
  assign n25545 = n25408 & n43586 ;
  assign n25568 = n25545 | n25559 ;
  assign n43587 = ~n25419 ;
  assign n25569 = n43587 & n25568 ;
  assign n25570 = n25386 | n25569 ;
  assign n43588 = ~n25562 ;
  assign n25571 = n43588 & n25570 ;
  assign n43589 = ~n25571 ;
  assign n25572 = n22030 & n43589 ;
  assign n43590 = ~n24643 ;
  assign n24678 = n43590 & n24657 ;
  assign n24679 = n43157 & n24678 ;
  assign n25376 = n24679 & n136 ;
  assign n24648 = n24643 | n24647 ;
  assign n43591 = ~n24648 ;
  assign n25389 = n43591 & n136 ;
  assign n25390 = n24657 | n25389 ;
  assign n43592 = ~n25376 ;
  assign n25391 = n43592 & n25390 ;
  assign n25563 = n22030 | n25562 ;
  assign n43593 = ~n25563 ;
  assign n25574 = n43593 & n25570 ;
  assign n25575 = n25391 | n25574 ;
  assign n43594 = ~n25572 ;
  assign n25576 = n43594 & n25575 ;
  assign n43595 = ~n25576 ;
  assign n25577 = n141 & n43595 ;
  assign n24662 = n24547 & n43145 ;
  assign n43596 = ~n24663 ;
  assign n24676 = n24662 & n43596 ;
  assign n25372 = n24676 & n136 ;
  assign n24677 = n24660 | n24663 ;
  assign n43597 = ~n24677 ;
  assign n25443 = n43597 & n136 ;
  assign n25444 = n24547 | n25443 ;
  assign n43598 = ~n25372 ;
  assign n25445 = n43598 & n25444 ;
  assign n25573 = n141 | n25572 ;
  assign n43599 = ~n25573 ;
  assign n25578 = n43599 & n25575 ;
  assign n25579 = n25445 | n25578 ;
  assign n43600 = ~n25577 ;
  assign n25580 = n43600 & n25579 ;
  assign n43601 = ~n25580 ;
  assign n25581 = n142 & n43601 ;
  assign n24670 = n24666 | n24667 ;
  assign n43602 = ~n24670 ;
  assign n25343 = n43602 & n136 ;
  assign n25344 = n24485 | n25343 ;
  assign n43603 = ~n24667 ;
  assign n24668 = n24485 & n43603 ;
  assign n24669 = n43151 & n24668 ;
  assign n25526 = n24669 & n25517 ;
  assign n43604 = ~n25526 ;
  assign n25527 = n25344 & n43604 ;
  assign n25564 = n139 & n43581 ;
  assign n25541 = n139 | n25540 ;
  assign n43605 = ~n25541 ;
  assign n25587 = n43605 & n25568 ;
  assign n25588 = n25386 | n25587 ;
  assign n43606 = ~n25564 ;
  assign n25589 = n43606 & n25588 ;
  assign n43607 = ~n25589 ;
  assign n25590 = n140 & n43607 ;
  assign n25591 = n43593 & n25588 ;
  assign n25592 = n25391 | n25591 ;
  assign n43608 = ~n25590 ;
  assign n25593 = n43608 & n25592 ;
  assign n43609 = ~n25593 ;
  assign n25594 = n141 & n43609 ;
  assign n25595 = n142 | n25594 ;
  assign n43610 = ~n25595 ;
  assign n25596 = n25579 & n43610 ;
  assign n25597 = n25527 | n25596 ;
  assign n43611 = ~n25581 ;
  assign n25598 = n43611 & n25597 ;
  assign n43612 = ~n25598 ;
  assign n25599 = n143 & n43612 ;
  assign n24675 = n24633 & n43162 ;
  assign n43613 = ~n24688 ;
  assign n24701 = n24675 & n43613 ;
  assign n25425 = n24701 & n136 ;
  assign n24702 = n24673 | n24688 ;
  assign n43614 = ~n24702 ;
  assign n25429 = n43614 & n136 ;
  assign n25430 = n24633 | n25429 ;
  assign n43615 = ~n25425 ;
  assign n25431 = n43615 & n25430 ;
  assign n25582 = n143 | n25581 ;
  assign n43616 = ~n25582 ;
  assign n25600 = n43616 & n25597 ;
  assign n25601 = n25431 | n25600 ;
  assign n43617 = ~n25599 ;
  assign n25602 = n43617 & n25601 ;
  assign n43618 = ~n25602 ;
  assign n25603 = n18797 & n43618 ;
  assign n25611 = n43599 & n25592 ;
  assign n25612 = n25445 | n25611 ;
  assign n43619 = ~n25594 ;
  assign n25613 = n43619 & n25612 ;
  assign n43620 = ~n25613 ;
  assign n25614 = n142 & n43620 ;
  assign n25615 = n43610 & n25612 ;
  assign n25616 = n25527 | n25615 ;
  assign n43621 = ~n25614 ;
  assign n25617 = n43621 & n25616 ;
  assign n43622 = ~n25617 ;
  assign n25618 = n19362 & n43622 ;
  assign n25619 = n144 | n25618 ;
  assign n43623 = ~n25619 ;
  assign n25620 = n25601 & n43623 ;
  assign n25632 = n25603 | n25620 ;
  assign n25621 = n25440 | n25620 ;
  assign n43624 = ~n25603 ;
  assign n25622 = n43624 & n25621 ;
  assign n43625 = ~n25622 ;
  assign n25623 = n145 & n43625 ;
  assign n24700 = n24512 & n43179 ;
  assign n43626 = ~n24712 ;
  assign n24723 = n24700 & n43626 ;
  assign n25412 = n24723 & n136 ;
  assign n24724 = n24698 | n24712 ;
  assign n43627 = ~n24724 ;
  assign n25426 = n43627 & n136 ;
  assign n25427 = n24512 | n25426 ;
  assign n43628 = ~n25412 ;
  assign n25428 = n43628 & n25427 ;
  assign n25604 = n145 | n25603 ;
  assign n43629 = ~n25604 ;
  assign n25624 = n43629 & n25621 ;
  assign n25625 = n25428 | n25624 ;
  assign n43630 = ~n25623 ;
  assign n25626 = n43630 & n25625 ;
  assign n43631 = ~n25626 ;
  assign n25627 = n146 & n43631 ;
  assign n24750 = n24716 | n24732 ;
  assign n43632 = ~n24750 ;
  assign n25340 = n43632 & n136 ;
  assign n25341 = n24516 | n25340 ;
  assign n43633 = ~n24716 ;
  assign n24722 = n24516 & n43633 ;
  assign n24749 = n24722 & n43206 ;
  assign n25452 = n24749 & n136 ;
  assign n43634 = ~n25452 ;
  assign n25453 = n25341 & n43634 ;
  assign n25635 = n43616 & n25616 ;
  assign n25636 = n25431 | n25635 ;
  assign n43635 = ~n25618 ;
  assign n25637 = n43635 & n25636 ;
  assign n43636 = ~n25637 ;
  assign n25638 = n144 & n43636 ;
  assign n25639 = n43623 & n25636 ;
  assign n25640 = n25440 | n25639 ;
  assign n43637 = ~n25638 ;
  assign n25641 = n43637 & n25640 ;
  assign n43638 = ~n25641 ;
  assign n25642 = n145 & n43638 ;
  assign n25643 = n146 | n25642 ;
  assign n43639 = ~n25643 ;
  assign n25644 = n25625 & n43639 ;
  assign n25645 = n25453 | n25644 ;
  assign n43640 = ~n25627 ;
  assign n25646 = n43640 & n25645 ;
  assign n43641 = ~n25646 ;
  assign n25647 = n147 & n43641 ;
  assign n24748 = n24719 | n24734 ;
  assign n43642 = ~n24748 ;
  assign n25370 = n43642 & n136 ;
  assign n25371 = n24527 | n25370 ;
  assign n24721 = n24527 & n43195 ;
  assign n43643 = ~n24734 ;
  assign n24747 = n24721 & n43643 ;
  assign n25387 = n24747 & n136 ;
  assign n43644 = ~n25387 ;
  assign n25388 = n25371 & n43644 ;
  assign n25628 = n147 | n25627 ;
  assign n43645 = ~n25628 ;
  assign n25648 = n43645 & n25645 ;
  assign n25649 = n25388 | n25648 ;
  assign n43646 = ~n25647 ;
  assign n25650 = n43646 & n25649 ;
  assign n43647 = ~n25650 ;
  assign n25651 = n15807 & n43647 ;
  assign n43648 = ~n24738 ;
  assign n24744 = n24545 & n43648 ;
  assign n24745 = n43201 & n24744 ;
  assign n25411 = n24745 & n136 ;
  assign n24746 = n24737 | n24738 ;
  assign n43649 = ~n24746 ;
  assign n25420 = n43649 & n136 ;
  assign n25421 = n24545 | n25420 ;
  assign n43650 = ~n25411 ;
  assign n25422 = n43650 & n25421 ;
  assign n25659 = n43629 & n25640 ;
  assign n25660 = n25428 | n25659 ;
  assign n43651 = ~n25642 ;
  assign n25661 = n43651 & n25660 ;
  assign n43652 = ~n25661 ;
  assign n25662 = n146 & n43652 ;
  assign n25663 = n43639 & n25660 ;
  assign n25664 = n25453 | n25663 ;
  assign n43653 = ~n25662 ;
  assign n25665 = n43653 & n25664 ;
  assign n43654 = ~n25665 ;
  assign n25666 = n16322 & n43654 ;
  assign n25667 = n148 | n25666 ;
  assign n43655 = ~n25667 ;
  assign n25668 = n25649 & n43655 ;
  assign n25669 = n25422 | n25668 ;
  assign n43656 = ~n25651 ;
  assign n25670 = n43656 & n25669 ;
  assign n43657 = ~n25670 ;
  assign n25671 = n149 & n43657 ;
  assign n24773 = n24741 | n24760 ;
  assign n43658 = ~n24773 ;
  assign n25432 = n43658 & n136 ;
  assign n25433 = n24500 | n25432 ;
  assign n24743 = n24500 & n43211 ;
  assign n43659 = ~n24760 ;
  assign n24774 = n24743 & n43659 ;
  assign n25532 = n24774 & n25517 ;
  assign n43660 = ~n25532 ;
  assign n25533 = n25433 & n43660 ;
  assign n25652 = n149 | n25651 ;
  assign n43661 = ~n25652 ;
  assign n25672 = n43661 & n25669 ;
  assign n25673 = n25533 | n25672 ;
  assign n43662 = ~n25671 ;
  assign n25674 = n43662 & n25673 ;
  assign n43663 = ~n25674 ;
  assign n25675 = n150 & n43663 ;
  assign n43664 = ~n24764 ;
  assign n24770 = n24555 & n43664 ;
  assign n24771 = n43217 & n24770 ;
  assign n25434 = n24771 & n136 ;
  assign n24772 = n24763 | n24764 ;
  assign n43665 = ~n24772 ;
  assign n25446 = n43665 & n136 ;
  assign n25447 = n24555 | n25446 ;
  assign n43666 = ~n25434 ;
  assign n25448 = n43666 & n25447 ;
  assign n25683 = n43645 & n25664 ;
  assign n25684 = n25388 | n25683 ;
  assign n43667 = ~n25666 ;
  assign n25685 = n43667 & n25684 ;
  assign n43668 = ~n25685 ;
  assign n25686 = n148 & n43668 ;
  assign n25687 = n43655 & n25684 ;
  assign n25688 = n25422 | n25687 ;
  assign n43669 = ~n25686 ;
  assign n25689 = n43669 & n25688 ;
  assign n43670 = ~n25689 ;
  assign n25690 = n149 & n43670 ;
  assign n25691 = n150 | n25690 ;
  assign n43671 = ~n25691 ;
  assign n25692 = n25673 & n43671 ;
  assign n25693 = n25448 | n25692 ;
  assign n43672 = ~n25675 ;
  assign n25694 = n43672 & n25693 ;
  assign n43673 = ~n25694 ;
  assign n25695 = n151 & n43673 ;
  assign n24769 = n24558 & n43227 ;
  assign n43674 = ~n24784 ;
  assign n24797 = n24769 & n43674 ;
  assign n25455 = n24797 & n136 ;
  assign n24798 = n24767 | n24784 ;
  assign n43675 = ~n24798 ;
  assign n25456 = n43675 & n136 ;
  assign n25457 = n24558 | n25456 ;
  assign n43676 = ~n25455 ;
  assign n25458 = n43676 & n25457 ;
  assign n25676 = n151 | n25675 ;
  assign n43677 = ~n25676 ;
  assign n25696 = n43677 & n25693 ;
  assign n25697 = n25458 | n25696 ;
  assign n43678 = ~n25695 ;
  assign n25698 = n43678 & n25697 ;
  assign n43679 = ~n25698 ;
  assign n25699 = n13079 & n43679 ;
  assign n43680 = ~n24788 ;
  assign n24794 = n24519 & n43680 ;
  assign n24795 = n43233 & n24794 ;
  assign n25358 = n24795 & n136 ;
  assign n24796 = n24787 | n24788 ;
  assign n43681 = ~n24796 ;
  assign n25367 = n43681 & n136 ;
  assign n25368 = n24519 | n25367 ;
  assign n43682 = ~n25358 ;
  assign n25369 = n43682 & n25368 ;
  assign n25706 = n43661 & n25688 ;
  assign n25707 = n25533 | n25706 ;
  assign n43683 = ~n25690 ;
  assign n25708 = n43683 & n25707 ;
  assign n43684 = ~n25708 ;
  assign n25709 = n150 & n43684 ;
  assign n25710 = n43671 & n25707 ;
  assign n25711 = n25448 | n25710 ;
  assign n43685 = ~n25709 ;
  assign n25712 = n43685 & n25711 ;
  assign n43686 = ~n25712 ;
  assign n25713 = n13662 & n43686 ;
  assign n25714 = n152 | n25713 ;
  assign n43687 = ~n25714 ;
  assign n25715 = n25697 & n43687 ;
  assign n25716 = n25369 | n25715 ;
  assign n43688 = ~n25699 ;
  assign n25717 = n43688 & n25716 ;
  assign n43689 = ~n25717 ;
  assign n25718 = n153 & n43689 ;
  assign n24822 = n24791 | n24808 ;
  assign n43690 = ~n24822 ;
  assign n25352 = n43690 & n136 ;
  assign n25353 = n24562 | n25352 ;
  assign n24793 = n24562 & n43243 ;
  assign n43691 = ~n24808 ;
  assign n24821 = n24793 & n43691 ;
  assign n25356 = n24821 & n136 ;
  assign n43692 = ~n25356 ;
  assign n25357 = n25353 & n43692 ;
  assign n25700 = n153 | n25699 ;
  assign n43693 = ~n25700 ;
  assign n25719 = n43693 & n25716 ;
  assign n25720 = n25357 | n25719 ;
  assign n43694 = ~n25718 ;
  assign n25721 = n43694 & n25720 ;
  assign n43695 = ~n25721 ;
  assign n25722 = n154 & n43695 ;
  assign n43696 = ~n24812 ;
  assign n24818 = n24509 & n43696 ;
  assign n24819 = n43249 & n24818 ;
  assign n25351 = n24819 & n136 ;
  assign n24820 = n24811 | n24812 ;
  assign n43697 = ~n24820 ;
  assign n25359 = n43697 & n136 ;
  assign n25360 = n24509 | n25359 ;
  assign n43698 = ~n25351 ;
  assign n25361 = n43698 & n25360 ;
  assign n25730 = n43677 & n25711 ;
  assign n25731 = n25458 | n25730 ;
  assign n43699 = ~n25713 ;
  assign n25732 = n43699 & n25731 ;
  assign n43700 = ~n25732 ;
  assign n25733 = n152 & n43700 ;
  assign n25734 = n43687 & n25731 ;
  assign n25735 = n25369 | n25734 ;
  assign n43701 = ~n25733 ;
  assign n25736 = n43701 & n25735 ;
  assign n43702 = ~n25736 ;
  assign n25737 = n153 & n43702 ;
  assign n25738 = n154 | n25737 ;
  assign n43703 = ~n25738 ;
  assign n25739 = n25720 & n43703 ;
  assign n25740 = n25361 | n25739 ;
  assign n43704 = ~n25722 ;
  assign n25741 = n43704 & n25740 ;
  assign n43705 = ~n25741 ;
  assign n25742 = n155 & n43705 ;
  assign n24846 = n24815 | n24832 ;
  assign n43706 = ~n24846 ;
  assign n25436 = n43706 & n136 ;
  assign n25437 = n24507 | n25436 ;
  assign n24817 = n24507 & n43259 ;
  assign n43707 = ~n24832 ;
  assign n24845 = n24817 & n43707 ;
  assign n25520 = n24845 & n25517 ;
  assign n43708 = ~n25520 ;
  assign n25521 = n25437 & n43708 ;
  assign n25723 = n11067 | n25722 ;
  assign n43709 = ~n25723 ;
  assign n25743 = n43709 & n25740 ;
  assign n25744 = n25521 | n25743 ;
  assign n43710 = ~n25742 ;
  assign n25745 = n43710 & n25744 ;
  assign n43711 = ~n25745 ;
  assign n25746 = n10657 & n43711 ;
  assign n24844 = n24835 | n24836 ;
  assign n43712 = ~n24844 ;
  assign n25345 = n43712 & n136 ;
  assign n25346 = n24537 | n25345 ;
  assign n43713 = ~n24836 ;
  assign n24842 = n24537 & n43713 ;
  assign n24843 = n43265 & n24842 ;
  assign n25349 = n24843 & n136 ;
  assign n43714 = ~n25349 ;
  assign n25350 = n25346 & n43714 ;
  assign n25754 = n43693 & n25735 ;
  assign n25755 = n25357 | n25754 ;
  assign n43715 = ~n25737 ;
  assign n25756 = n43715 & n25755 ;
  assign n43716 = ~n25756 ;
  assign n25757 = n154 & n43716 ;
  assign n25758 = n43703 & n25755 ;
  assign n25759 = n25361 | n25758 ;
  assign n43717 = ~n25757 ;
  assign n25760 = n43717 & n25759 ;
  assign n43718 = ~n25760 ;
  assign n25761 = n11067 & n43718 ;
  assign n25762 = n10657 | n25761 ;
  assign n43719 = ~n25762 ;
  assign n25763 = n25744 & n43719 ;
  assign n25764 = n25350 | n25763 ;
  assign n43720 = ~n25746 ;
  assign n25765 = n43720 & n25764 ;
  assign n43721 = ~n25765 ;
  assign n25766 = n157 & n43721 ;
  assign n24869 = n24839 | n24856 ;
  assign n43722 = ~n24869 ;
  assign n25335 = n43722 & n136 ;
  assign n25336 = n24480 | n25335 ;
  assign n24840 = n24480 & n43275 ;
  assign n43723 = ~n24856 ;
  assign n24870 = n24840 & n43723 ;
  assign n25338 = n24870 & n136 ;
  assign n43724 = ~n25338 ;
  assign n25339 = n25336 & n43724 ;
  assign n25747 = n157 | n25746 ;
  assign n43725 = ~n25747 ;
  assign n25767 = n43725 & n25764 ;
  assign n25768 = n25339 | n25767 ;
  assign n43726 = ~n25766 ;
  assign n25769 = n43726 & n25768 ;
  assign n43727 = ~n25769 ;
  assign n25770 = n158 & n43727 ;
  assign n24868 = n24859 | n24860 ;
  assign n43728 = ~n24868 ;
  assign n25330 = n43728 & n136 ;
  assign n25331 = n24476 | n25330 ;
  assign n43729 = ~n24860 ;
  assign n24866 = n24476 & n43729 ;
  assign n24867 = n43281 & n24866 ;
  assign n25333 = n24867 & n136 ;
  assign n43730 = ~n25333 ;
  assign n25334 = n25331 & n43730 ;
  assign n25779 = n43709 & n25759 ;
  assign n25780 = n25521 | n25779 ;
  assign n43731 = ~n25761 ;
  assign n25781 = n43731 & n25780 ;
  assign n43732 = ~n25781 ;
  assign n25782 = n156 & n43732 ;
  assign n25783 = n43719 & n25780 ;
  assign n25784 = n25350 | n25783 ;
  assign n43733 = ~n25782 ;
  assign n25785 = n43733 & n25784 ;
  assign n43734 = ~n25785 ;
  assign n25786 = n157 & n43734 ;
  assign n25787 = n158 | n25786 ;
  assign n43735 = ~n25787 ;
  assign n25788 = n25768 & n43735 ;
  assign n25789 = n25334 | n25788 ;
  assign n43736 = ~n25770 ;
  assign n25790 = n43736 & n25789 ;
  assign n43737 = ~n25790 ;
  assign n25791 = n159 & n43737 ;
  assign n24894 = n24863 | n24880 ;
  assign n43738 = ~n24894 ;
  assign n25326 = n43738 & n136 ;
  assign n25327 = n24542 | n25326 ;
  assign n24865 = n24542 & n43291 ;
  assign n43739 = ~n24880 ;
  assign n24893 = n24865 & n43739 ;
  assign n25524 = n24893 & n25517 ;
  assign n43740 = ~n25524 ;
  assign n25525 = n25327 & n43740 ;
  assign n25771 = n8857 | n25770 ;
  assign n43741 = ~n25771 ;
  assign n25792 = n43741 & n25789 ;
  assign n25793 = n25525 | n25792 ;
  assign n43742 = ~n25791 ;
  assign n25794 = n43742 & n25793 ;
  assign n43743 = ~n25794 ;
  assign n25795 = n8534 & n43743 ;
  assign n43744 = ~n24884 ;
  assign n24890 = n24530 & n43744 ;
  assign n24891 = n43297 & n24890 ;
  assign n25322 = n24891 & n136 ;
  assign n24892 = n24883 | n24884 ;
  assign n43745 = ~n24892 ;
  assign n25395 = n43745 & n136 ;
  assign n25396 = n24530 | n25395 ;
  assign n43746 = ~n25322 ;
  assign n25397 = n43746 & n25396 ;
  assign n25802 = n43725 & n25784 ;
  assign n25803 = n25339 | n25802 ;
  assign n43747 = ~n25786 ;
  assign n25804 = n43747 & n25803 ;
  assign n43748 = ~n25804 ;
  assign n25805 = n158 & n43748 ;
  assign n25806 = n43735 & n25803 ;
  assign n25807 = n25334 | n25806 ;
  assign n43749 = ~n25805 ;
  assign n25808 = n43749 & n25807 ;
  assign n43750 = ~n25808 ;
  assign n25809 = n8857 & n43750 ;
  assign n25810 = n160 | n25809 ;
  assign n43751 = ~n25810 ;
  assign n25811 = n25793 & n43751 ;
  assign n25812 = n25397 | n25811 ;
  assign n43752 = ~n25795 ;
  assign n25813 = n43752 & n25812 ;
  assign n43753 = ~n25813 ;
  assign n25814 = n161 & n43753 ;
  assign n24918 = n24887 | n24904 ;
  assign n43754 = ~n24918 ;
  assign n25441 = n43754 & n136 ;
  assign n25442 = n24447 | n25441 ;
  assign n24889 = n24447 & n43307 ;
  assign n43755 = ~n24904 ;
  assign n24917 = n24889 & n43755 ;
  assign n25522 = n24917 & n25517 ;
  assign n43756 = ~n25522 ;
  assign n25523 = n25442 & n43756 ;
  assign n25796 = n161 | n25795 ;
  assign n43757 = ~n25796 ;
  assign n25815 = n43757 & n25812 ;
  assign n25816 = n25523 | n25815 ;
  assign n43758 = ~n25814 ;
  assign n25817 = n43758 & n25816 ;
  assign n43759 = ~n25817 ;
  assign n25818 = n162 & n43759 ;
  assign n24916 = n24907 | n24908 ;
  assign n43760 = ~n24916 ;
  assign n25320 = n43760 & n136 ;
  assign n25321 = n24441 | n25320 ;
  assign n43761 = ~n24908 ;
  assign n24914 = n24441 & n43761 ;
  assign n24915 = n43313 & n24914 ;
  assign n25328 = n24915 & n136 ;
  assign n43762 = ~n25328 ;
  assign n25329 = n25321 & n43762 ;
  assign n25826 = n43741 & n25807 ;
  assign n25827 = n25525 | n25826 ;
  assign n43763 = ~n25809 ;
  assign n25828 = n43763 & n25827 ;
  assign n43764 = ~n25828 ;
  assign n25829 = n160 & n43764 ;
  assign n25830 = n43751 & n25827 ;
  assign n25831 = n25397 | n25830 ;
  assign n43765 = ~n25829 ;
  assign n25832 = n43765 & n25831 ;
  assign n43766 = ~n25832 ;
  assign n25833 = n161 & n43766 ;
  assign n25834 = n162 | n25833 ;
  assign n43767 = ~n25834 ;
  assign n25835 = n25816 & n43767 ;
  assign n25836 = n25329 | n25835 ;
  assign n43768 = ~n25818 ;
  assign n25837 = n43768 & n25836 ;
  assign n43769 = ~n25837 ;
  assign n25838 = n163 & n43769 ;
  assign n24913 = n24523 & n43323 ;
  assign n43770 = ~n24928 ;
  assign n24939 = n24913 & n43770 ;
  assign n25316 = n24939 & n136 ;
  assign n24940 = n24911 | n24928 ;
  assign n43771 = ~n24940 ;
  assign n25317 = n43771 & n136 ;
  assign n25318 = n24523 | n25317 ;
  assign n43772 = ~n25316 ;
  assign n25319 = n43772 & n25318 ;
  assign n25819 = n6889 | n25818 ;
  assign n43773 = ~n25819 ;
  assign n25839 = n43773 & n25836 ;
  assign n25840 = n25319 | n25839 ;
  assign n43774 = ~n25838 ;
  assign n25841 = n43774 & n25840 ;
  assign n43775 = ~n25841 ;
  assign n25842 = n6600 & n43775 ;
  assign n43776 = ~n24932 ;
  assign n24938 = n24435 & n43776 ;
  assign n24965 = n24938 & n43350 ;
  assign n25342 = n24965 & n136 ;
  assign n24966 = n24932 | n24948 ;
  assign n43777 = ~n24966 ;
  assign n25373 = n43777 & n136 ;
  assign n25374 = n24435 | n25373 ;
  assign n43778 = ~n25342 ;
  assign n25375 = n43778 & n25374 ;
  assign n25850 = n43757 & n25831 ;
  assign n25851 = n25523 | n25850 ;
  assign n43779 = ~n25833 ;
  assign n25852 = n43779 & n25851 ;
  assign n43780 = ~n25852 ;
  assign n25853 = n162 & n43780 ;
  assign n25854 = n43767 & n25851 ;
  assign n25855 = n25329 | n25854 ;
  assign n43781 = ~n25853 ;
  assign n25856 = n43781 & n25855 ;
  assign n43782 = ~n25856 ;
  assign n25857 = n6889 & n43782 ;
  assign n25858 = n6600 | n25857 ;
  assign n43783 = ~n25858 ;
  assign n25859 = n25840 & n43783 ;
  assign n25860 = n25375 | n25859 ;
  assign n43784 = ~n25842 ;
  assign n25861 = n43784 & n25860 ;
  assign n43785 = ~n25861 ;
  assign n25862 = n165 & n43785 ;
  assign n24964 = n24935 | n24950 ;
  assign n43786 = ~n24964 ;
  assign n25314 = n43786 & n136 ;
  assign n25315 = n24426 | n25314 ;
  assign n24937 = n24426 & n43339 ;
  assign n43787 = ~n24950 ;
  assign n24963 = n24937 & n43787 ;
  assign n25530 = n24963 & n25517 ;
  assign n43788 = ~n25530 ;
  assign n25531 = n25315 & n43788 ;
  assign n25843 = n165 | n25842 ;
  assign n43789 = ~n25843 ;
  assign n25863 = n43789 & n25860 ;
  assign n25864 = n25531 | n25863 ;
  assign n43790 = ~n25862 ;
  assign n25865 = n43790 & n25864 ;
  assign n43791 = ~n25865 ;
  assign n25866 = n166 & n43791 ;
  assign n24962 = n24953 | n24954 ;
  assign n43792 = ~n24962 ;
  assign n25310 = n43792 & n136 ;
  assign n25311 = n24418 | n25310 ;
  assign n43793 = ~n24954 ;
  assign n24960 = n24418 & n43793 ;
  assign n24961 = n43345 & n24960 ;
  assign n25382 = n24961 & n136 ;
  assign n43794 = ~n25382 ;
  assign n25383 = n25311 & n43794 ;
  assign n25875 = n43773 & n25855 ;
  assign n25876 = n25319 | n25875 ;
  assign n43795 = ~n25857 ;
  assign n25877 = n43795 & n25876 ;
  assign n43796 = ~n25877 ;
  assign n25878 = n164 & n43796 ;
  assign n25879 = n43783 & n25876 ;
  assign n25880 = n25375 | n25879 ;
  assign n43797 = ~n25878 ;
  assign n25881 = n43797 & n25880 ;
  assign n43798 = ~n25881 ;
  assign n25882 = n165 & n43798 ;
  assign n25883 = n166 | n25882 ;
  assign n43799 = ~n25883 ;
  assign n25884 = n25864 & n43799 ;
  assign n25885 = n25383 | n25884 ;
  assign n43800 = ~n25866 ;
  assign n25886 = n43800 & n25885 ;
  assign n43801 = ~n25886 ;
  assign n25887 = n167 & n43801 ;
  assign n24990 = n24957 | n24976 ;
  assign n43802 = ~n24990 ;
  assign n25347 = n43802 & n136 ;
  assign n25348 = n24534 | n25347 ;
  assign n24959 = n24534 & n43355 ;
  assign n43803 = ~n24976 ;
  assign n24989 = n24959 & n43803 ;
  assign n25534 = n24989 & n25517 ;
  assign n43804 = ~n25534 ;
  assign n25535 = n25348 & n43804 ;
  assign n25867 = n5352 | n25866 ;
  assign n43805 = ~n25867 ;
  assign n25888 = n43805 & n25885 ;
  assign n25889 = n25535 | n25888 ;
  assign n43806 = ~n25887 ;
  assign n25890 = n43806 & n25889 ;
  assign n43807 = ~n25890 ;
  assign n25891 = n4934 & n43807 ;
  assign n24988 = n24979 | n24980 ;
  assign n43808 = ~n24988 ;
  assign n25307 = n43808 & n136 ;
  assign n25308 = n24504 | n25307 ;
  assign n43809 = ~n24980 ;
  assign n24986 = n24504 & n43809 ;
  assign n24987 = n43361 & n24986 ;
  assign n25380 = n24987 & n136 ;
  assign n43810 = ~n25380 ;
  assign n25381 = n25308 & n43810 ;
  assign n25899 = n43789 & n25880 ;
  assign n25900 = n25531 | n25899 ;
  assign n43811 = ~n25882 ;
  assign n25901 = n43811 & n25900 ;
  assign n43812 = ~n25901 ;
  assign n25902 = n166 & n43812 ;
  assign n25903 = n43799 & n25900 ;
  assign n25904 = n25383 | n25903 ;
  assign n43813 = ~n25902 ;
  assign n25905 = n43813 & n25904 ;
  assign n43814 = ~n25905 ;
  assign n25906 = n5352 & n43814 ;
  assign n25907 = n4934 | n25906 ;
  assign n43815 = ~n25907 ;
  assign n25908 = n25889 & n43815 ;
  assign n25909 = n25381 | n25908 ;
  assign n43816 = ~n25891 ;
  assign n25910 = n43816 & n25909 ;
  assign n43817 = ~n25910 ;
  assign n25911 = n169 & n43817 ;
  assign n25014 = n24983 | n25000 ;
  assign n43818 = ~n25014 ;
  assign n25305 = n43818 & n136 ;
  assign n25306 = n24565 | n25305 ;
  assign n24985 = n24565 & n43371 ;
  assign n43819 = ~n25000 ;
  assign n25013 = n24985 & n43819 ;
  assign n25518 = n25013 & n25517 ;
  assign n43820 = ~n25518 ;
  assign n25519 = n25306 & n43820 ;
  assign n25892 = n169 | n25891 ;
  assign n43821 = ~n25892 ;
  assign n25912 = n43821 & n25909 ;
  assign n25913 = n25519 | n25912 ;
  assign n43822 = ~n25911 ;
  assign n25914 = n43822 & n25913 ;
  assign n43823 = ~n25914 ;
  assign n25915 = n170 & n43823 ;
  assign n43824 = ~n25004 ;
  assign n25010 = n24569 & n43824 ;
  assign n25011 = n43377 & n25010 ;
  assign n25337 = n25011 & n136 ;
  assign n25012 = n25003 | n25004 ;
  assign n43825 = ~n25012 ;
  assign n25459 = n43825 & n136 ;
  assign n25460 = n24569 | n25459 ;
  assign n43826 = ~n25337 ;
  assign n25461 = n43826 & n25460 ;
  assign n25923 = n43805 & n25904 ;
  assign n25924 = n25535 | n25923 ;
  assign n43827 = ~n25906 ;
  assign n25925 = n43827 & n25924 ;
  assign n43828 = ~n25925 ;
  assign n25926 = n168 & n43828 ;
  assign n25927 = n43815 & n25924 ;
  assign n25928 = n25381 | n25927 ;
  assign n43829 = ~n25926 ;
  assign n25929 = n43829 & n25928 ;
  assign n43830 = ~n25929 ;
  assign n25930 = n169 & n43830 ;
  assign n25931 = n170 | n25930 ;
  assign n43831 = ~n25931 ;
  assign n25932 = n25913 & n43831 ;
  assign n25933 = n25461 | n25932 ;
  assign n43832 = ~n25915 ;
  assign n25934 = n43832 & n25933 ;
  assign n43833 = ~n25934 ;
  assign n25935 = n171 & n43833 ;
  assign n25009 = n24571 & n43387 ;
  assign n43834 = ~n25024 ;
  assign n25035 = n25009 & n43834 ;
  assign n25463 = n25035 & n136 ;
  assign n25036 = n25007 | n25024 ;
  assign n43835 = ~n25036 ;
  assign n25464 = n43835 & n136 ;
  assign n25465 = n24571 | n25464 ;
  assign n43836 = ~n25463 ;
  assign n25466 = n43836 & n25465 ;
  assign n25916 = n3940 | n25915 ;
  assign n43837 = ~n25916 ;
  assign n25936 = n43837 & n25933 ;
  assign n25938 = n25466 | n25936 ;
  assign n43838 = ~n25935 ;
  assign n25939 = n43838 & n25938 ;
  assign n43839 = ~n25939 ;
  assign n25940 = n3631 & n43839 ;
  assign n43840 = ~n25028 ;
  assign n25034 = n24429 & n43840 ;
  assign n25061 = n25034 & n43414 ;
  assign n25462 = n25061 & n136 ;
  assign n25062 = n25028 | n25044 ;
  assign n43841 = ~n25062 ;
  assign n25467 = n43841 & n136 ;
  assign n25468 = n24429 | n25467 ;
  assign n43842 = ~n25462 ;
  assign n25469 = n43842 & n25468 ;
  assign n25947 = n43821 & n25928 ;
  assign n25948 = n25519 | n25947 ;
  assign n43843 = ~n25930 ;
  assign n25949 = n43843 & n25948 ;
  assign n43844 = ~n25949 ;
  assign n25950 = n170 & n43844 ;
  assign n25951 = n43831 & n25948 ;
  assign n25952 = n25461 | n25951 ;
  assign n43845 = ~n25950 ;
  assign n25953 = n43845 & n25952 ;
  assign n43846 = ~n25953 ;
  assign n25954 = n3940 & n43846 ;
  assign n25955 = n3631 | n25954 ;
  assign n43847 = ~n25955 ;
  assign n25956 = n25938 & n43847 ;
  assign n25957 = n25469 | n25956 ;
  assign n43848 = ~n25940 ;
  assign n25958 = n43848 & n25957 ;
  assign n43849 = ~n25958 ;
  assign n25959 = n173 & n43849 ;
  assign n25060 = n25031 | n25046 ;
  assign n43850 = ~n25060 ;
  assign n25354 = n43850 & n136 ;
  assign n25355 = n24432 | n25354 ;
  assign n25033 = n24432 & n43403 ;
  assign n43851 = ~n25046 ;
  assign n25059 = n25033 & n43851 ;
  assign n25470 = n25059 & n136 ;
  assign n43852 = ~n25470 ;
  assign n25471 = n25355 & n43852 ;
  assign n25941 = n173 | n25940 ;
  assign n43853 = ~n25941 ;
  assign n25960 = n43853 & n25957 ;
  assign n25961 = n25471 | n25960 ;
  assign n43854 = ~n25959 ;
  assign n25962 = n43854 & n25961 ;
  assign n43855 = ~n25962 ;
  assign n25963 = n174 & n43855 ;
  assign n43856 = ~n25050 ;
  assign n25056 = n24573 & n43856 ;
  assign n25057 = n43409 & n25056 ;
  assign n25472 = n25057 & n136 ;
  assign n25058 = n25049 | n25050 ;
  assign n43857 = ~n25058 ;
  assign n25473 = n43857 & n136 ;
  assign n25474 = n24573 | n25473 ;
  assign n43858 = ~n25472 ;
  assign n25475 = n43858 & n25474 ;
  assign n25971 = n43837 & n25952 ;
  assign n25972 = n25466 | n25971 ;
  assign n43859 = ~n25954 ;
  assign n25973 = n43859 & n25972 ;
  assign n43860 = ~n25973 ;
  assign n25974 = n172 & n43860 ;
  assign n25975 = n43847 & n25972 ;
  assign n25976 = n25469 | n25975 ;
  assign n43861 = ~n25974 ;
  assign n25977 = n43861 & n25976 ;
  assign n43862 = ~n25977 ;
  assign n25978 = n173 & n43862 ;
  assign n25979 = n174 | n25978 ;
  assign n43863 = ~n25979 ;
  assign n25980 = n25961 & n43863 ;
  assign n25981 = n25475 | n25980 ;
  assign n43864 = ~n25963 ;
  assign n25982 = n43864 & n25981 ;
  assign n43865 = ~n25982 ;
  assign n25983 = n175 & n43865 ;
  assign n25086 = n25053 | n25072 ;
  assign n43866 = ~n25086 ;
  assign n25476 = n43866 & n136 ;
  assign n25477 = n24575 | n25476 ;
  assign n25055 = n24575 & n43419 ;
  assign n43867 = ~n25072 ;
  assign n25085 = n25055 & n43867 ;
  assign n25528 = n25085 & n25517 ;
  assign n43868 = ~n25528 ;
  assign n25529 = n25477 & n43868 ;
  assign n25964 = n2753 | n25963 ;
  assign n43869 = ~n25964 ;
  assign n25984 = n43869 & n25981 ;
  assign n25985 = n25529 | n25984 ;
  assign n43870 = ~n25983 ;
  assign n25986 = n43870 & n25985 ;
  assign n43871 = ~n25986 ;
  assign n25987 = n2431 & n43871 ;
  assign n25084 = n25075 | n25076 ;
  assign n43872 = ~n25084 ;
  assign n25312 = n43872 & n136 ;
  assign n25313 = n24580 | n25312 ;
  assign n43873 = ~n25076 ;
  assign n25082 = n24580 & n43873 ;
  assign n25083 = n43425 & n25082 ;
  assign n25409 = n25083 & n136 ;
  assign n43874 = ~n25409 ;
  assign n25410 = n25313 & n43874 ;
  assign n25995 = n43853 & n25976 ;
  assign n25996 = n25471 | n25995 ;
  assign n43875 = ~n25978 ;
  assign n25997 = n43875 & n25996 ;
  assign n43876 = ~n25997 ;
  assign n25998 = n174 & n43876 ;
  assign n25999 = n43863 & n25996 ;
  assign n26000 = n25475 | n25999 ;
  assign n43877 = ~n25998 ;
  assign n26001 = n43877 & n26000 ;
  assign n43878 = ~n26001 ;
  assign n26002 = n2753 & n43878 ;
  assign n26003 = n2431 | n26002 ;
  assign n43879 = ~n26003 ;
  assign n26004 = n25985 & n43879 ;
  assign n26005 = n25410 | n26004 ;
  assign n43880 = ~n25987 ;
  assign n26006 = n43880 & n26005 ;
  assign n43881 = ~n26006 ;
  assign n26007 = n177 & n43881 ;
  assign n25110 = n25079 | n25096 ;
  assign n43882 = ~n25110 ;
  assign n25478 = n43882 & n136 ;
  assign n25479 = n24584 | n25478 ;
  assign n25081 = n24584 & n43435 ;
  assign n43883 = ~n25096 ;
  assign n25109 = n25081 & n43883 ;
  assign n25547 = n25109 & n25517 ;
  assign n43884 = ~n25547 ;
  assign n25548 = n25479 & n43884 ;
  assign n25988 = n177 | n25987 ;
  assign n43885 = ~n25988 ;
  assign n26008 = n43885 & n26005 ;
  assign n26009 = n25548 | n26008 ;
  assign n43886 = ~n26007 ;
  assign n26010 = n43886 & n26009 ;
  assign n43887 = ~n26010 ;
  assign n26011 = n178 & n43887 ;
  assign n25108 = n25099 | n25100 ;
  assign n43888 = ~n25108 ;
  assign n25323 = n43888 & n136 ;
  assign n25324 = n24586 | n25323 ;
  assign n43889 = ~n25100 ;
  assign n25106 = n24586 & n43889 ;
  assign n25107 = n43441 & n25106 ;
  assign n25480 = n25107 & n136 ;
  assign n43890 = ~n25480 ;
  assign n25481 = n25324 & n43890 ;
  assign n26019 = n43869 & n26000 ;
  assign n26020 = n25529 | n26019 ;
  assign n43891 = ~n26002 ;
  assign n26021 = n43891 & n26020 ;
  assign n43892 = ~n26021 ;
  assign n26022 = n176 & n43892 ;
  assign n26023 = n43879 & n26020 ;
  assign n26024 = n25410 | n26023 ;
  assign n43893 = ~n26022 ;
  assign n26025 = n43893 & n26024 ;
  assign n43894 = ~n26025 ;
  assign n26026 = n177 & n43894 ;
  assign n26027 = n178 | n26026 ;
  assign n43895 = ~n26027 ;
  assign n26028 = n26009 & n43895 ;
  assign n26029 = n25481 | n26028 ;
  assign n43896 = ~n26011 ;
  assign n26030 = n43896 & n26029 ;
  assign n43897 = ~n26030 ;
  assign n26031 = n179 & n43897 ;
  assign n25132 = n25103 | n25120 ;
  assign n43898 = ~n25132 ;
  assign n25486 = n43898 & n136 ;
  assign n25487 = n24592 | n25486 ;
  assign n25105 = n24592 & n43451 ;
  assign n43899 = ~n25120 ;
  assign n25131 = n25105 & n43899 ;
  assign n25549 = n25131 & n25517 ;
  assign n43900 = ~n25549 ;
  assign n25550 = n25487 & n43900 ;
  assign n26012 = n1707 | n26011 ;
  assign n43901 = ~n26012 ;
  assign n26032 = n43901 & n26029 ;
  assign n26033 = n25550 | n26032 ;
  assign n43902 = ~n26031 ;
  assign n26034 = n43902 & n26033 ;
  assign n43903 = ~n26034 ;
  assign n26035 = n1487 & n43903 ;
  assign n25158 = n25124 | n25140 ;
  assign n43904 = ~n25158 ;
  assign n25423 = n43904 & n136 ;
  assign n25424 = n24550 | n25423 ;
  assign n43905 = ~n25124 ;
  assign n25130 = n24550 & n43905 ;
  assign n25157 = n25130 & n43478 ;
  assign n25490 = n25157 & n136 ;
  assign n43906 = ~n25490 ;
  assign n25491 = n25424 & n43906 ;
  assign n26043 = n43885 & n26024 ;
  assign n26044 = n25548 | n26043 ;
  assign n43907 = ~n26026 ;
  assign n26045 = n43907 & n26044 ;
  assign n43908 = ~n26045 ;
  assign n26046 = n178 & n43908 ;
  assign n26047 = n43895 & n26044 ;
  assign n26048 = n25481 | n26047 ;
  assign n43909 = ~n26046 ;
  assign n26049 = n43909 & n26048 ;
  assign n43910 = ~n26049 ;
  assign n26050 = n1707 & n43910 ;
  assign n26051 = n1487 | n26050 ;
  assign n43911 = ~n26051 ;
  assign n26052 = n26033 & n43911 ;
  assign n26053 = n25491 | n26052 ;
  assign n43912 = ~n26035 ;
  assign n26054 = n43912 & n26053 ;
  assign n43913 = ~n26054 ;
  assign n26055 = n181 & n43913 ;
  assign n25129 = n24596 & n43467 ;
  assign n43914 = ~n25142 ;
  assign n25155 = n25129 & n43914 ;
  assign n25482 = n25155 & n136 ;
  assign n25156 = n25127 | n25142 ;
  assign n43915 = ~n25156 ;
  assign n25492 = n43915 & n136 ;
  assign n25493 = n24596 | n25492 ;
  assign n43916 = ~n25482 ;
  assign n25494 = n43916 & n25493 ;
  assign n26036 = n181 | n26035 ;
  assign n43917 = ~n26036 ;
  assign n26056 = n43917 & n26053 ;
  assign n26057 = n25494 | n26056 ;
  assign n43918 = ~n26055 ;
  assign n26058 = n43918 & n26057 ;
  assign n43919 = ~n26058 ;
  assign n26059 = n182 & n43919 ;
  assign n43920 = ~n25146 ;
  assign n25152 = n24600 & n43920 ;
  assign n25153 = n43473 & n25152 ;
  assign n25495 = n25153 & n136 ;
  assign n25154 = n25145 | n25146 ;
  assign n43921 = ~n25154 ;
  assign n25496 = n43921 & n136 ;
  assign n25497 = n24600 | n25496 ;
  assign n43922 = ~n25495 ;
  assign n25498 = n43922 & n25497 ;
  assign n26067 = n43901 & n26048 ;
  assign n26068 = n25550 | n26067 ;
  assign n43923 = ~n26050 ;
  assign n26069 = n43923 & n26068 ;
  assign n43924 = ~n26069 ;
  assign n26070 = n180 & n43924 ;
  assign n26071 = n43911 & n26068 ;
  assign n26072 = n25491 | n26071 ;
  assign n43925 = ~n26070 ;
  assign n26073 = n43925 & n26072 ;
  assign n43926 = ~n26073 ;
  assign n26074 = n181 & n43926 ;
  assign n26075 = n182 | n26074 ;
  assign n43927 = ~n26075 ;
  assign n26076 = n26057 & n43927 ;
  assign n26077 = n25498 | n26076 ;
  assign n43928 = ~n26059 ;
  assign n26078 = n43928 & n26077 ;
  assign n43929 = ~n26078 ;
  assign n26079 = n183 & n43929 ;
  assign n25151 = n24521 & n43483 ;
  assign n43930 = ~n25168 ;
  assign n25181 = n25151 & n43930 ;
  assign n25325 = n25181 & n136 ;
  assign n25182 = n25149 | n25168 ;
  assign n43931 = ~n25182 ;
  assign n25501 = n43931 & n136 ;
  assign n25502 = n24521 | n25501 ;
  assign n43932 = ~n25325 ;
  assign n25503 = n43932 & n25502 ;
  assign n26060 = n183 | n26059 ;
  assign n43933 = ~n26060 ;
  assign n26080 = n43933 & n26077 ;
  assign n26081 = n25503 | n26080 ;
  assign n43934 = ~n26079 ;
  assign n26082 = n43934 & n26081 ;
  assign n43935 = ~n26082 ;
  assign n26083 = n838 & n43935 ;
  assign n25180 = n25171 | n25172 ;
  assign n43936 = ~n25180 ;
  assign n25488 = n43936 & n136 ;
  assign n25489 = n24602 | n25488 ;
  assign n43937 = ~n25172 ;
  assign n25178 = n24602 & n43937 ;
  assign n25179 = n43489 & n25178 ;
  assign n25504 = n25179 & n136 ;
  assign n43938 = ~n25504 ;
  assign n25505 = n25489 & n43938 ;
  assign n26091 = n43917 & n26072 ;
  assign n26092 = n25494 | n26091 ;
  assign n43939 = ~n26074 ;
  assign n26093 = n43939 & n26092 ;
  assign n43940 = ~n26093 ;
  assign n26094 = n182 & n43940 ;
  assign n26095 = n43927 & n26092 ;
  assign n26096 = n25498 | n26095 ;
  assign n43941 = ~n26094 ;
  assign n26097 = n43941 & n26096 ;
  assign n43942 = ~n26097 ;
  assign n26098 = n996 & n43942 ;
  assign n26099 = n838 | n26098 ;
  assign n43943 = ~n26099 ;
  assign n26100 = n26081 & n43943 ;
  assign n26101 = n25505 | n26100 ;
  assign n43944 = ~n26083 ;
  assign n26102 = n43944 & n26101 ;
  assign n43945 = ~n26102 ;
  assign n26103 = n185 & n43945 ;
  assign n25206 = n25175 | n25192 ;
  assign n43946 = ~n25206 ;
  assign n25398 = n43946 & n136 ;
  assign n25399 = n24606 | n25398 ;
  assign n25177 = n24606 & n43499 ;
  assign n43947 = ~n25192 ;
  assign n25205 = n25177 & n43947 ;
  assign n25551 = n25205 & n25517 ;
  assign n43948 = ~n25551 ;
  assign n25552 = n25399 & n43948 ;
  assign n26084 = n185 | n26083 ;
  assign n43949 = ~n26084 ;
  assign n26104 = n43949 & n26101 ;
  assign n26105 = n25552 | n26104 ;
  assign n43950 = ~n26103 ;
  assign n26106 = n43950 & n26105 ;
  assign n43951 = ~n26106 ;
  assign n26107 = n186 & n43951 ;
  assign n43952 = ~n25196 ;
  assign n25202 = n24611 & n43952 ;
  assign n25203 = n43505 & n25202 ;
  assign n25332 = n25203 & n136 ;
  assign n25204 = n25195 | n25196 ;
  assign n43953 = ~n25204 ;
  assign n25506 = n43953 & n136 ;
  assign n25507 = n24611 | n25506 ;
  assign n43954 = ~n25332 ;
  assign n25508 = n43954 & n25507 ;
  assign n26115 = n43933 & n26096 ;
  assign n26116 = n25503 | n26115 ;
  assign n43955 = ~n26098 ;
  assign n26117 = n43955 & n26116 ;
  assign n43956 = ~n26117 ;
  assign n26118 = n184 & n43956 ;
  assign n26119 = n43943 & n26116 ;
  assign n26120 = n25505 | n26119 ;
  assign n43957 = ~n26118 ;
  assign n26121 = n43957 & n26120 ;
  assign n43958 = ~n26121 ;
  assign n26122 = n185 & n43958 ;
  assign n26123 = n186 | n26122 ;
  assign n43959 = ~n26123 ;
  assign n26124 = n26105 & n43959 ;
  assign n26125 = n25508 | n26124 ;
  assign n43960 = ~n26107 ;
  assign n26126 = n43960 & n26125 ;
  assign n43961 = ~n26126 ;
  assign n26127 = n187 & n43961 ;
  assign n25201 = n24614 & n43515 ;
  assign n43962 = ~n25216 ;
  assign n25227 = n25201 & n43962 ;
  assign n25402 = n25227 & n136 ;
  assign n25228 = n25199 | n25216 ;
  assign n43963 = ~n25228 ;
  assign n25449 = n43963 & n136 ;
  assign n25450 = n24614 | n25449 ;
  assign n43964 = ~n25402 ;
  assign n25451 = n43964 & n25450 ;
  assign n26108 = n528 | n26107 ;
  assign n43965 = ~n26108 ;
  assign n26128 = n43965 & n26125 ;
  assign n26129 = n25451 | n26128 ;
  assign n43966 = ~n26127 ;
  assign n26130 = n43966 & n26129 ;
  assign n43967 = ~n26130 ;
  assign n26131 = n413 & n43967 ;
  assign n43968 = ~n25220 ;
  assign n25226 = n24617 & n43968 ;
  assign n25251 = n25226 & n43542 ;
  assign n25362 = n25251 & n136 ;
  assign n25252 = n25220 | n25236 ;
  assign n43969 = ~n25252 ;
  assign n25509 = n43969 & n136 ;
  assign n25510 = n24617 | n25509 ;
  assign n43970 = ~n25362 ;
  assign n25511 = n43970 & n25510 ;
  assign n26139 = n43949 & n26120 ;
  assign n26140 = n25552 | n26139 ;
  assign n43971 = ~n26122 ;
  assign n26141 = n43971 & n26140 ;
  assign n43972 = ~n26141 ;
  assign n26142 = n186 & n43972 ;
  assign n26143 = n43959 & n26140 ;
  assign n26144 = n25508 | n26143 ;
  assign n43973 = ~n26142 ;
  assign n26145 = n43973 & n26144 ;
  assign n43974 = ~n26145 ;
  assign n26146 = n528 & n43974 ;
  assign n26147 = n413 | n26146 ;
  assign n43975 = ~n26147 ;
  assign n26148 = n26129 & n43975 ;
  assign n26149 = n25511 | n26148 ;
  assign n43976 = ~n26131 ;
  assign n26150 = n43976 & n26149 ;
  assign n43977 = ~n26150 ;
  assign n26151 = n189 & n43977 ;
  assign n25225 = n24577 & n43531 ;
  assign n43978 = ~n25238 ;
  assign n25249 = n25225 & n43978 ;
  assign n25454 = n25249 & n136 ;
  assign n25250 = n25223 | n25238 ;
  assign n43979 = ~n25250 ;
  assign n25483 = n43979 & n136 ;
  assign n25484 = n24577 | n25483 ;
  assign n43980 = ~n25454 ;
  assign n25485 = n43980 & n25484 ;
  assign n26132 = n189 | n26131 ;
  assign n43981 = ~n26132 ;
  assign n26152 = n43981 & n26149 ;
  assign n26153 = n25485 | n26152 ;
  assign n43982 = ~n26151 ;
  assign n26154 = n43982 & n26153 ;
  assign n43983 = ~n26154 ;
  assign n26155 = n190 & n43983 ;
  assign n25277 = n43536 & n25258 ;
  assign n25280 = n25241 | n25277 ;
  assign n43984 = ~n25280 ;
  assign n25363 = n43984 & n136 ;
  assign n25364 = n24622 | n25363 ;
  assign n43985 = ~n25277 ;
  assign n25278 = n24622 & n43985 ;
  assign n25279 = n43537 & n25278 ;
  assign n25499 = n25279 & n136 ;
  assign n43986 = ~n25499 ;
  assign n25500 = n25364 & n43986 ;
  assign n26163 = n43965 & n26144 ;
  assign n26164 = n25451 | n26163 ;
  assign n43987 = ~n26146 ;
  assign n26165 = n43987 & n26164 ;
  assign n43988 = ~n26165 ;
  assign n26166 = n188 & n43988 ;
  assign n26167 = n43975 & n26164 ;
  assign n26168 = n25511 | n26167 ;
  assign n43989 = ~n26166 ;
  assign n26169 = n43989 & n26168 ;
  assign n43990 = ~n26169 ;
  assign n26170 = n189 & n43990 ;
  assign n26171 = n190 | n26170 ;
  assign n43991 = ~n26171 ;
  assign n26172 = n26153 & n43991 ;
  assign n26173 = n25500 | n26172 ;
  assign n43992 = ~n26155 ;
  assign n26174 = n43992 & n26173 ;
  assign n43993 = ~n26174 ;
  assign n26175 = n191 & n43993 ;
  assign n25267 = n25245 | n25262 ;
  assign n43994 = ~n25267 ;
  assign n25365 = n43994 & n136 ;
  assign n25366 = n24588 | n25365 ;
  assign n25248 = n24588 & n43547 ;
  assign n43995 = ~n25262 ;
  assign n25266 = n25248 & n43995 ;
  assign n25512 = n25266 & n136 ;
  assign n43996 = ~n25512 ;
  assign n25513 = n25366 & n43996 ;
  assign n26156 = n191 | n26155 ;
  assign n43997 = ~n26156 ;
  assign n26176 = n43997 & n26173 ;
  assign n26177 = n25513 | n26176 ;
  assign n43998 = ~n26175 ;
  assign n26178 = n43998 & n26177 ;
  assign n25276 = n25269 | n25271 ;
  assign n43999 = ~n25276 ;
  assign n25377 = n43999 & n136 ;
  assign n25378 = n24626 | n25377 ;
  assign n44000 = ~n25271 ;
  assign n25274 = n24626 & n44000 ;
  assign n25275 = n43553 & n25274 ;
  assign n25403 = n25275 & n136 ;
  assign n44001 = ~n25403 ;
  assign n25404 = n25378 & n44001 ;
  assign n25299 = n25270 | n25293 ;
  assign n44002 = ~n25299 ;
  assign n25514 = n44002 & n136 ;
  assign n26207 = n25514 | n25515 ;
  assign n26208 = n25404 | n26207 ;
  assign n26209 = n26178 | n26208 ;
  assign n26210 = n31336 & n26209 ;
  assign n26185 = n43981 & n26168 ;
  assign n26186 = n25485 | n26185 ;
  assign n44003 = ~n26170 ;
  assign n26187 = n44003 & n26186 ;
  assign n44004 = ~n26187 ;
  assign n26188 = n190 & n44004 ;
  assign n26189 = n43991 & n26186 ;
  assign n26190 = n25500 | n26189 ;
  assign n44005 = ~n26188 ;
  assign n26191 = n44005 & n26190 ;
  assign n44006 = ~n26191 ;
  assign n26192 = n287 & n44006 ;
  assign n44007 = ~n26192 ;
  assign n26193 = n25404 & n44007 ;
  assign n26194 = n26177 & n26193 ;
  assign n25300 = n192 & n25299 ;
  assign n44008 = ~n25293 ;
  assign n25392 = n44008 & n136 ;
  assign n44009 = ~n25392 ;
  assign n25393 = n25270 & n44009 ;
  assign n44010 = ~n25393 ;
  assign n25394 = n25300 & n44010 ;
  assign n25289 = n24620 | n25283 ;
  assign n44011 = ~n25289 ;
  assign n26215 = n44011 & n25292 ;
  assign n26216 = n43576 & n26215 ;
  assign n26217 = n43577 & n26216 ;
  assign n26218 = n43578 & n26217 ;
  assign n26219 = n25394 | n26218 ;
  assign n26220 = n26194 | n26219 ;
  assign n135 = n26210 | n26220 ;
  assign n44012 = ~n25632 ;
  assign n26269 = n44012 & n135 ;
  assign n26270 = n25440 | n26269 ;
  assign n44013 = ~n25620 ;
  assign n25630 = n25440 & n44013 ;
  assign n25631 = n43624 & n25630 ;
  assign n26350 = n25631 & n135 ;
  assign n44014 = ~n26350 ;
  assign n26351 = n26270 & n44014 ;
  assign n25608 = n25581 | n25596 ;
  assign n44015 = ~n25608 ;
  assign n26236 = n44015 & n135 ;
  assign n26237 = n25527 | n26236 ;
  assign n44016 = ~n25596 ;
  assign n25606 = n25527 & n44016 ;
  assign n25607 = n43611 & n25606 ;
  assign n26346 = n25607 & n135 ;
  assign n44017 = ~n26346 ;
  assign n26347 = n26237 & n44017 ;
  assign n254 = x10 | x11 ;
  assign n255 = x12 | n254 ;
  assign n25285 = n255 & n43575 ;
  assign n25286 = n43576 & n25285 ;
  assign n26213 = n25286 & n43577 ;
  assign n26214 = n43578 & n26213 ;
  assign n26309 = x12 & n135 ;
  assign n44018 = ~n26309 ;
  assign n26330 = n26214 & n44018 ;
  assign n44019 = ~x12 ;
  assign n26232 = n44019 & n135 ;
  assign n44020 = ~n26232 ;
  assign n26233 = x13 & n44020 ;
  assign n44021 = ~n251 ;
  assign n26313 = n44021 & n135 ;
  assign n26335 = n26233 | n26313 ;
  assign n26336 = n26330 | n26335 ;
  assign n256 = n44019 & n254 ;
  assign n26157 = n287 | n26155 ;
  assign n44022 = ~n26157 ;
  assign n26196 = n44022 & n26190 ;
  assign n26197 = n25513 | n26196 ;
  assign n26198 = n44007 & n26197 ;
  assign n26211 = n26198 | n26208 ;
  assign n26212 = n31336 & n26211 ;
  assign n26199 = n26193 & n26197 ;
  assign n26441 = n26199 | n26219 ;
  assign n26442 = n26212 | n26441 ;
  assign n44023 = ~n26442 ;
  assign n26449 = x12 & n44023 ;
  assign n26450 = n256 | n26449 ;
  assign n44024 = ~n26450 ;
  assign n26451 = n25517 & n44024 ;
  assign n44025 = ~n26451 ;
  assign n26452 = n26336 & n44025 ;
  assign n44026 = ~n26452 ;
  assign n26453 = n137 & n44026 ;
  assign n26310 = n255 & n44018 ;
  assign n44027 = ~n26310 ;
  assign n26311 = n136 & n44027 ;
  assign n26312 = n137 | n26311 ;
  assign n44028 = ~n26312 ;
  assign n26337 = n44028 & n26336 ;
  assign n44029 = ~n26218 ;
  assign n26478 = n25517 & n44029 ;
  assign n44030 = ~n25394 ;
  assign n26479 = n44030 & n26478 ;
  assign n44031 = ~n26199 ;
  assign n26480 = n44031 & n26479 ;
  assign n44032 = ~n26212 ;
  assign n26481 = n44032 & n26480 ;
  assign n26482 = n26313 | n26481 ;
  assign n26483 = x14 & n26482 ;
  assign n26484 = x14 | n26481 ;
  assign n26485 = n26313 | n26484 ;
  assign n44033 = ~n26483 ;
  assign n26486 = n44033 & n26485 ;
  assign n26487 = n26337 | n26486 ;
  assign n44034 = ~n26453 ;
  assign n26488 = n44034 & n26487 ;
  assign n44035 = ~n26488 ;
  assign n26489 = n138 & n44035 ;
  assign n25542 = n25401 | n25538 ;
  assign n44036 = ~n25542 ;
  assign n26271 = n44036 & n135 ;
  assign n26272 = n25407 | n26271 ;
  assign n25543 = n25407 & n44036 ;
  assign n26315 = n25543 & n135 ;
  assign n44037 = ~n26315 ;
  assign n26316 = n26272 & n44037 ;
  assign n26454 = n138 | n26453 ;
  assign n26455 = n137 | n26451 ;
  assign n44038 = ~n26455 ;
  assign n26456 = n26336 & n44038 ;
  assign n26494 = n26456 | n26486 ;
  assign n44039 = ~n26454 ;
  assign n26495 = n44039 & n26494 ;
  assign n26496 = n26316 | n26495 ;
  assign n44040 = ~n26489 ;
  assign n26497 = n44040 & n26496 ;
  assign n44041 = ~n26497 ;
  assign n26498 = n139 & n44041 ;
  assign n44042 = ~n25545 ;
  assign n25566 = n44042 & n25559 ;
  assign n44043 = ~n25418 ;
  assign n25567 = n44043 & n25566 ;
  assign n26317 = n25567 & n135 ;
  assign n25546 = n25418 | n25545 ;
  assign n44044 = ~n25546 ;
  assign n26318 = n44044 & n135 ;
  assign n26319 = n25559 | n26318 ;
  assign n44045 = ~n26317 ;
  assign n26320 = n44045 & n26319 ;
  assign n26491 = n22661 | n26489 ;
  assign n44046 = ~n26491 ;
  assign n26499 = n44046 & n26496 ;
  assign n26500 = n26320 | n26499 ;
  assign n44047 = ~n26498 ;
  assign n26501 = n44047 & n26500 ;
  assign n44048 = ~n26501 ;
  assign n26502 = n22030 & n44048 ;
  assign n26206 = n25564 | n25569 ;
  assign n44049 = ~n26206 ;
  assign n26305 = n44049 & n135 ;
  assign n26306 = n25386 | n26305 ;
  assign n25565 = n25386 & n43606 ;
  assign n44050 = ~n25569 ;
  assign n26205 = n25565 & n44050 ;
  assign n26307 = n26205 & n135 ;
  assign n44051 = ~n26307 ;
  assign n26308 = n26306 & n44051 ;
  assign n26457 = n136 & n44024 ;
  assign n44052 = ~n26457 ;
  assign n26458 = n26336 & n44052 ;
  assign n44053 = ~n26458 ;
  assign n26459 = n137 & n44053 ;
  assign n26460 = n138 | n26459 ;
  assign n44054 = ~n26460 ;
  assign n26505 = n44054 & n26494 ;
  assign n26508 = n26316 | n26505 ;
  assign n26509 = n44040 & n26508 ;
  assign n44055 = ~n26509 ;
  assign n26510 = n22661 & n44055 ;
  assign n26511 = n140 | n26510 ;
  assign n44056 = ~n26511 ;
  assign n26512 = n26500 & n44056 ;
  assign n26513 = n26308 | n26512 ;
  assign n44057 = ~n26502 ;
  assign n26514 = n44057 & n26513 ;
  assign n44058 = ~n26514 ;
  assign n26515 = n141 & n44058 ;
  assign n25586 = n25572 | n25574 ;
  assign n44059 = ~n25586 ;
  assign n26295 = n44059 & n135 ;
  assign n26296 = n25391 | n26295 ;
  assign n44060 = ~n25574 ;
  assign n25584 = n25391 & n44060 ;
  assign n25585 = n43594 & n25584 ;
  assign n26322 = n25585 & n135 ;
  assign n44061 = ~n26322 ;
  assign n26323 = n26296 & n44061 ;
  assign n26503 = n141 | n26502 ;
  assign n44062 = ~n26503 ;
  assign n26516 = n44062 & n26513 ;
  assign n26517 = n26323 | n26516 ;
  assign n44063 = ~n26515 ;
  assign n26518 = n44063 & n26517 ;
  assign n44064 = ~n26518 ;
  assign n26519 = n142 & n44064 ;
  assign n26520 = n143 | n26519 ;
  assign n25609 = n25445 & n43619 ;
  assign n44065 = ~n25578 ;
  assign n25610 = n44065 & n25609 ;
  assign n26326 = n25610 & n135 ;
  assign n25583 = n25577 | n25578 ;
  assign n44066 = ~n25583 ;
  assign n26327 = n44066 & n135 ;
  assign n26328 = n25445 | n26327 ;
  assign n44067 = ~n26326 ;
  assign n26329 = n44067 & n26328 ;
  assign n26522 = n44046 & n26508 ;
  assign n26523 = n26320 | n26522 ;
  assign n44068 = ~n26510 ;
  assign n26524 = n44068 & n26523 ;
  assign n44069 = ~n26524 ;
  assign n26525 = n140 & n44069 ;
  assign n26526 = n44056 & n26523 ;
  assign n26529 = n26308 | n26526 ;
  assign n44070 = ~n26525 ;
  assign n26530 = n44070 & n26529 ;
  assign n44071 = ~n26530 ;
  assign n26531 = n141 & n44071 ;
  assign n26532 = n142 | n26531 ;
  assign n44072 = ~n26532 ;
  assign n26533 = n26517 & n44072 ;
  assign n26534 = n26329 | n26533 ;
  assign n44073 = ~n26520 ;
  assign n26535 = n44073 & n26534 ;
  assign n26536 = n26347 | n26535 ;
  assign n44074 = ~n26519 ;
  assign n26537 = n44074 & n26534 ;
  assign n44075 = ~n26537 ;
  assign n26538 = n143 & n44075 ;
  assign n44076 = ~n26538 ;
  assign n26539 = n26536 & n44076 ;
  assign n44077 = ~n26539 ;
  assign n26540 = n18797 & n44077 ;
  assign n26541 = n145 | n26540 ;
  assign n25633 = n25431 & n43635 ;
  assign n44078 = ~n25600 ;
  assign n25634 = n44078 & n25633 ;
  assign n26284 = n25634 & n135 ;
  assign n25605 = n25599 | n25600 ;
  assign n44079 = ~n25605 ;
  assign n26341 = n44079 & n135 ;
  assign n26342 = n25431 | n26341 ;
  assign n44080 = ~n26284 ;
  assign n26343 = n44080 & n26342 ;
  assign n26543 = n44062 & n26529 ;
  assign n26544 = n26323 | n26543 ;
  assign n44081 = ~n26531 ;
  assign n26545 = n44081 & n26544 ;
  assign n44082 = ~n26545 ;
  assign n26546 = n142 & n44082 ;
  assign n26547 = n44072 & n26544 ;
  assign n26550 = n26329 | n26547 ;
  assign n44083 = ~n26546 ;
  assign n26551 = n44083 & n26550 ;
  assign n44084 = ~n26551 ;
  assign n26552 = n19362 & n44084 ;
  assign n26553 = n144 | n26552 ;
  assign n44085 = ~n26553 ;
  assign n26554 = n26536 & n44085 ;
  assign n26555 = n26343 | n26554 ;
  assign n44086 = ~n26541 ;
  assign n26556 = n44086 & n26555 ;
  assign n26557 = n26351 | n26556 ;
  assign n26565 = n44073 & n26550 ;
  assign n26566 = n26347 | n26565 ;
  assign n44087 = ~n26552 ;
  assign n26567 = n44087 & n26566 ;
  assign n44088 = ~n26567 ;
  assign n26568 = n144 & n44088 ;
  assign n26569 = n44085 & n26566 ;
  assign n26570 = n26343 | n26569 ;
  assign n44089 = ~n26568 ;
  assign n26571 = n44089 & n26570 ;
  assign n44090 = ~n26571 ;
  assign n26572 = n145 & n44090 ;
  assign n44091 = ~n26572 ;
  assign n26573 = n26557 & n44091 ;
  assign n44092 = ~n26573 ;
  assign n26574 = n146 & n44092 ;
  assign n25629 = n25623 | n25624 ;
  assign n44093 = ~n25629 ;
  assign n26223 = n44093 & n135 ;
  assign n26224 = n25428 | n26223 ;
  assign n25657 = n25428 & n43651 ;
  assign n44094 = ~n25624 ;
  assign n25658 = n44094 & n25657 ;
  assign n26470 = n25658 & n26442 ;
  assign n44095 = ~n26470 ;
  assign n26471 = n26224 & n44095 ;
  assign n26575 = n146 | n26572 ;
  assign n44096 = ~n26575 ;
  assign n26576 = n26557 & n44096 ;
  assign n26577 = n26471 | n26576 ;
  assign n44097 = ~n26574 ;
  assign n26578 = n44097 & n26577 ;
  assign n44098 = ~n26578 ;
  assign n26579 = n16322 & n44098 ;
  assign n44099 = ~n25644 ;
  assign n25654 = n25453 & n44099 ;
  assign n25655 = n43640 & n25654 ;
  assign n26299 = n25655 & n135 ;
  assign n25656 = n25627 | n25644 ;
  assign n44100 = ~n25656 ;
  assign n26357 = n44100 & n135 ;
  assign n26358 = n25453 | n26357 ;
  assign n44101 = ~n26299 ;
  assign n26359 = n44101 & n26358 ;
  assign n44102 = ~n26540 ;
  assign n26559 = n44102 & n26555 ;
  assign n44103 = ~n26559 ;
  assign n26560 = n145 & n44103 ;
  assign n44104 = ~n26560 ;
  assign n26561 = n26557 & n44104 ;
  assign n44105 = ~n26561 ;
  assign n26562 = n146 & n44105 ;
  assign n26563 = n147 | n26562 ;
  assign n44106 = ~n26563 ;
  assign n26581 = n44106 & n26577 ;
  assign n26582 = n26359 | n26581 ;
  assign n44107 = ~n26579 ;
  assign n26583 = n44107 & n26582 ;
  assign n44108 = ~n26583 ;
  assign n26584 = n148 & n44108 ;
  assign n25681 = n25388 & n43667 ;
  assign n44109 = ~n25648 ;
  assign n25682 = n44109 & n25681 ;
  assign n26264 = n25682 & n135 ;
  assign n25653 = n25647 | n25648 ;
  assign n44110 = ~n25653 ;
  assign n26332 = n44110 & n135 ;
  assign n26333 = n25388 | n26332 ;
  assign n44111 = ~n26264 ;
  assign n26334 = n44111 & n26333 ;
  assign n26580 = n148 | n26579 ;
  assign n44112 = ~n26580 ;
  assign n26585 = n44112 & n26582 ;
  assign n26586 = n26334 | n26585 ;
  assign n44113 = ~n26584 ;
  assign n26587 = n44113 & n26586 ;
  assign n44114 = ~n26587 ;
  assign n26588 = n149 & n44114 ;
  assign n44115 = ~n25668 ;
  assign n25678 = n25422 & n44115 ;
  assign n25679 = n43656 & n25678 ;
  assign n26314 = n25679 & n135 ;
  assign n25680 = n25651 | n25668 ;
  assign n44116 = ~n25680 ;
  assign n26364 = n44116 & n135 ;
  assign n26365 = n25422 | n26364 ;
  assign n44117 = ~n26314 ;
  assign n26366 = n44117 & n26365 ;
  assign n44118 = ~n26562 ;
  assign n26596 = n44118 & n26577 ;
  assign n44119 = ~n26596 ;
  assign n26597 = n147 & n44119 ;
  assign n44120 = ~n26597 ;
  assign n26598 = n26582 & n44120 ;
  assign n44121 = ~n26598 ;
  assign n26599 = n15807 & n44121 ;
  assign n26600 = n149 | n26599 ;
  assign n44122 = ~n26600 ;
  assign n26601 = n26586 & n44122 ;
  assign n26602 = n26366 | n26601 ;
  assign n44123 = ~n26588 ;
  assign n26603 = n44123 & n26602 ;
  assign n44124 = ~n26603 ;
  assign n26604 = n150 & n44124 ;
  assign n25677 = n25671 | n25672 ;
  assign n44125 = ~n25677 ;
  assign n26293 = n44125 & n135 ;
  assign n26294 = n25533 | n26293 ;
  assign n25704 = n25533 & n43683 ;
  assign n44126 = ~n25672 ;
  assign n25705 = n44126 & n25704 ;
  assign n26368 = n25705 & n135 ;
  assign n44127 = ~n26368 ;
  assign n26369 = n26294 & n44127 ;
  assign n26589 = n150 | n26588 ;
  assign n44128 = ~n26589 ;
  assign n26605 = n44128 & n26602 ;
  assign n26606 = n26369 | n26605 ;
  assign n44129 = ~n26604 ;
  assign n26607 = n44129 & n26606 ;
  assign n44130 = ~n26607 ;
  assign n26608 = n13662 & n44130 ;
  assign n25701 = n25675 | n25692 ;
  assign n44131 = ~n25701 ;
  assign n26287 = n44131 & n135 ;
  assign n26288 = n25448 | n26287 ;
  assign n44132 = ~n25692 ;
  assign n25702 = n25448 & n44132 ;
  assign n25703 = n43672 & n25702 ;
  assign n26291 = n25703 & n135 ;
  assign n44133 = ~n26291 ;
  assign n26292 = n26288 & n44133 ;
  assign n44134 = ~n26599 ;
  assign n26616 = n26586 & n44134 ;
  assign n44135 = ~n26616 ;
  assign n26617 = n149 & n44135 ;
  assign n44136 = ~n26617 ;
  assign n26618 = n26602 & n44136 ;
  assign n44137 = ~n26618 ;
  assign n26619 = n150 & n44137 ;
  assign n26620 = n151 | n26619 ;
  assign n44138 = ~n26620 ;
  assign n26621 = n26606 & n44138 ;
  assign n26622 = n26292 | n26621 ;
  assign n44139 = ~n26608 ;
  assign n26623 = n44139 & n26622 ;
  assign n44140 = ~n26623 ;
  assign n26624 = n152 & n44140 ;
  assign n25728 = n25458 & n43699 ;
  assign n44141 = ~n25696 ;
  assign n25729 = n44141 & n25728 ;
  assign n26283 = n25729 & n135 ;
  assign n25727 = n25696 | n25713 ;
  assign n44142 = ~n25727 ;
  assign n26302 = n44142 & n135 ;
  assign n26303 = n25458 | n26302 ;
  assign n44143 = ~n26283 ;
  assign n26304 = n44143 & n26303 ;
  assign n26609 = n152 | n26608 ;
  assign n44144 = ~n26609 ;
  assign n26625 = n44144 & n26622 ;
  assign n26626 = n26304 | n26625 ;
  assign n44145 = ~n26624 ;
  assign n26627 = n44145 & n26626 ;
  assign n44146 = ~n26627 ;
  assign n26628 = n153 & n44146 ;
  assign n25726 = n25699 | n25715 ;
  assign n44147 = ~n25726 ;
  assign n26279 = n44147 & n135 ;
  assign n26280 = n25369 | n26279 ;
  assign n44148 = ~n25715 ;
  assign n25724 = n25369 & n44148 ;
  assign n25725 = n43688 & n25724 ;
  assign n26281 = n25725 & n135 ;
  assign n44149 = ~n26281 ;
  assign n26282 = n26280 & n44149 ;
  assign n44150 = ~n26619 ;
  assign n26636 = n26606 & n44150 ;
  assign n44151 = ~n26636 ;
  assign n26637 = n151 & n44151 ;
  assign n44152 = ~n26637 ;
  assign n26638 = n26622 & n44152 ;
  assign n44153 = ~n26638 ;
  assign n26639 = n13079 & n44153 ;
  assign n26640 = n153 | n26639 ;
  assign n44154 = ~n26640 ;
  assign n26641 = n26626 & n44154 ;
  assign n26642 = n26282 | n26641 ;
  assign n44155 = ~n26628 ;
  assign n26643 = n44155 & n26642 ;
  assign n44156 = ~n26643 ;
  assign n26644 = n154 & n44156 ;
  assign n25751 = n25719 | n25737 ;
  assign n44157 = ~n25751 ;
  assign n26267 = n44157 & n135 ;
  assign n26268 = n25357 | n26267 ;
  assign n25752 = n25357 & n43715 ;
  assign n44158 = ~n25719 ;
  assign n25753 = n44158 & n25752 ;
  assign n26275 = n25753 & n135 ;
  assign n44159 = ~n26275 ;
  assign n26276 = n26268 & n44159 ;
  assign n26629 = n154 | n26628 ;
  assign n44160 = ~n26629 ;
  assign n26645 = n44160 & n26642 ;
  assign n26646 = n26276 | n26645 ;
  assign n44161 = ~n26644 ;
  assign n26647 = n44161 & n26646 ;
  assign n44162 = ~n26647 ;
  assign n26648 = n11067 & n44162 ;
  assign n44163 = ~n25739 ;
  assign n25748 = n25361 & n44163 ;
  assign n25749 = n43704 & n25748 ;
  assign n26244 = n25749 & n135 ;
  assign n25750 = n25722 | n25739 ;
  assign n44164 = ~n25750 ;
  assign n26256 = n44164 & n135 ;
  assign n26257 = n25361 | n26256 ;
  assign n44165 = ~n26244 ;
  assign n26258 = n44165 & n26257 ;
  assign n44166 = ~n26639 ;
  assign n26656 = n26626 & n44166 ;
  assign n44167 = ~n26656 ;
  assign n26657 = n153 & n44167 ;
  assign n44168 = ~n26657 ;
  assign n26658 = n26642 & n44168 ;
  assign n44169 = ~n26658 ;
  assign n26659 = n154 & n44169 ;
  assign n26660 = n11067 | n26659 ;
  assign n44170 = ~n26660 ;
  assign n26661 = n26646 & n44170 ;
  assign n26662 = n26258 | n26661 ;
  assign n44171 = ~n26648 ;
  assign n26663 = n44171 & n26662 ;
  assign n44172 = ~n26663 ;
  assign n26664 = n156 & n44172 ;
  assign n25778 = n25743 | n25761 ;
  assign n44173 = ~n25778 ;
  assign n26252 = n44173 & n135 ;
  assign n26253 = n25521 | n26252 ;
  assign n25776 = n25521 & n43731 ;
  assign n44174 = ~n25743 ;
  assign n25777 = n44174 & n25776 ;
  assign n26254 = n25777 & n135 ;
  assign n44175 = ~n26254 ;
  assign n26255 = n26253 & n44175 ;
  assign n26649 = n10657 | n26648 ;
  assign n44176 = ~n26649 ;
  assign n26665 = n44176 & n26662 ;
  assign n26666 = n26255 | n26665 ;
  assign n44177 = ~n26664 ;
  assign n26667 = n44177 & n26666 ;
  assign n44178 = ~n26667 ;
  assign n26668 = n157 & n44178 ;
  assign n25775 = n25746 | n25763 ;
  assign n44179 = ~n25775 ;
  assign n26242 = n44179 & n135 ;
  assign n26243 = n25350 | n26242 ;
  assign n44180 = ~n25763 ;
  assign n25773 = n25350 & n44180 ;
  assign n25774 = n43720 & n25773 ;
  assign n26247 = n25774 & n135 ;
  assign n44181 = ~n26247 ;
  assign n26248 = n26243 & n44181 ;
  assign n44182 = ~n26659 ;
  assign n26676 = n26646 & n44182 ;
  assign n44183 = ~n26676 ;
  assign n26677 = n155 & n44183 ;
  assign n44184 = ~n26677 ;
  assign n26678 = n26662 & n44184 ;
  assign n44185 = ~n26678 ;
  assign n26679 = n10657 & n44185 ;
  assign n26680 = n157 | n26679 ;
  assign n44186 = ~n26680 ;
  assign n26681 = n26666 & n44186 ;
  assign n26682 = n26248 | n26681 ;
  assign n44187 = ~n26668 ;
  assign n26683 = n44187 & n26682 ;
  assign n44188 = ~n26683 ;
  assign n26684 = n158 & n44188 ;
  assign n25800 = n25339 & n43747 ;
  assign n44189 = ~n25767 ;
  assign n25801 = n44189 & n25800 ;
  assign n26225 = n25801 & n135 ;
  assign n25772 = n25766 | n25767 ;
  assign n44190 = ~n25772 ;
  assign n26352 = n44190 & n135 ;
  assign n26353 = n25339 | n26352 ;
  assign n44191 = ~n26225 ;
  assign n26354 = n44191 & n26353 ;
  assign n26669 = n158 | n26668 ;
  assign n44192 = ~n26669 ;
  assign n26685 = n44192 & n26682 ;
  assign n26686 = n26354 | n26685 ;
  assign n44193 = ~n26684 ;
  assign n26687 = n44193 & n26686 ;
  assign n44194 = ~n26687 ;
  assign n26688 = n8857 & n44194 ;
  assign n25799 = n25770 | n25788 ;
  assign n44195 = ~n25799 ;
  assign n26339 = n44195 & n135 ;
  assign n26340 = n25334 | n26339 ;
  assign n44196 = ~n25788 ;
  assign n25797 = n25334 & n44196 ;
  assign n25798 = n43736 & n25797 ;
  assign n26348 = n25798 & n135 ;
  assign n44197 = ~n26348 ;
  assign n26349 = n26340 & n44197 ;
  assign n44198 = ~n26679 ;
  assign n26696 = n26666 & n44198 ;
  assign n44199 = ~n26696 ;
  assign n26697 = n157 & n44199 ;
  assign n44200 = ~n26697 ;
  assign n26698 = n26682 & n44200 ;
  assign n44201 = ~n26698 ;
  assign n26699 = n158 & n44201 ;
  assign n26700 = n8857 | n26699 ;
  assign n44202 = ~n26700 ;
  assign n26701 = n26686 & n44202 ;
  assign n26702 = n26349 | n26701 ;
  assign n44203 = ~n26688 ;
  assign n26703 = n44203 & n26702 ;
  assign n44204 = ~n26703 ;
  assign n26704 = n160 & n44204 ;
  assign n25823 = n25525 & n43763 ;
  assign n44205 = ~n25792 ;
  assign n25824 = n44205 & n25823 ;
  assign n26241 = n25824 & n135 ;
  assign n25825 = n25792 | n25809 ;
  assign n44206 = ~n25825 ;
  assign n26249 = n44206 & n135 ;
  assign n26250 = n25525 | n26249 ;
  assign n44207 = ~n26241 ;
  assign n26251 = n44207 & n26250 ;
  assign n26689 = n160 | n26688 ;
  assign n44208 = ~n26689 ;
  assign n26705 = n44208 & n26702 ;
  assign n26706 = n26251 | n26705 ;
  assign n44209 = ~n26704 ;
  assign n26707 = n44209 & n26706 ;
  assign n44210 = ~n26707 ;
  assign n26708 = n161 & n44210 ;
  assign n25822 = n25795 | n25811 ;
  assign n44211 = ~n25822 ;
  assign n26239 = n44211 & n135 ;
  assign n26240 = n25397 | n26239 ;
  assign n44212 = ~n25811 ;
  assign n25820 = n25397 & n44212 ;
  assign n25821 = n43752 & n25820 ;
  assign n26360 = n25821 & n135 ;
  assign n44213 = ~n26360 ;
  assign n26361 = n26240 & n44213 ;
  assign n44214 = ~n26699 ;
  assign n26716 = n26686 & n44214 ;
  assign n44215 = ~n26716 ;
  assign n26717 = n159 & n44215 ;
  assign n44216 = ~n26717 ;
  assign n26718 = n26702 & n44216 ;
  assign n44217 = ~n26718 ;
  assign n26719 = n8534 & n44217 ;
  assign n26720 = n161 | n26719 ;
  assign n44218 = ~n26720 ;
  assign n26721 = n26706 & n44218 ;
  assign n26722 = n26361 | n26721 ;
  assign n44219 = ~n26708 ;
  assign n26723 = n44219 & n26722 ;
  assign n44220 = ~n26723 ;
  assign n26724 = n162 & n44220 ;
  assign n25847 = n25523 & n43779 ;
  assign n44221 = ~n25815 ;
  assign n25848 = n44221 & n25847 ;
  assign n26238 = n25848 & n135 ;
  assign n25849 = n25815 | n25833 ;
  assign n44222 = ~n25849 ;
  assign n26261 = n44222 & n135 ;
  assign n26262 = n25523 | n26261 ;
  assign n44223 = ~n26238 ;
  assign n26263 = n44223 & n26262 ;
  assign n26709 = n162 | n26708 ;
  assign n44224 = ~n26709 ;
  assign n26725 = n44224 & n26722 ;
  assign n26727 = n26263 | n26725 ;
  assign n44225 = ~n26724 ;
  assign n26728 = n44225 & n26727 ;
  assign n44226 = ~n26728 ;
  assign n26729 = n6889 & n44226 ;
  assign n25846 = n25818 | n25835 ;
  assign n44227 = ~n25846 ;
  assign n26230 = n44227 & n135 ;
  assign n26231 = n25329 | n26230 ;
  assign n44228 = ~n25835 ;
  assign n25844 = n25329 & n44228 ;
  assign n25845 = n43768 & n25844 ;
  assign n26234 = n25845 & n135 ;
  assign n44229 = ~n26234 ;
  assign n26235 = n26231 & n44229 ;
  assign n44230 = ~n26719 ;
  assign n26736 = n26706 & n44230 ;
  assign n44231 = ~n26736 ;
  assign n26737 = n161 & n44231 ;
  assign n44232 = ~n26737 ;
  assign n26738 = n26722 & n44232 ;
  assign n44233 = ~n26738 ;
  assign n26739 = n162 & n44233 ;
  assign n26740 = n6889 | n26739 ;
  assign n44234 = ~n26740 ;
  assign n26741 = n26727 & n44234 ;
  assign n26742 = n26235 | n26741 ;
  assign n44235 = ~n26729 ;
  assign n26743 = n44235 & n26742 ;
  assign n44236 = ~n26743 ;
  assign n26744 = n164 & n44236 ;
  assign n25874 = n25839 | n25857 ;
  assign n44237 = ~n25874 ;
  assign n26226 = n44237 & n135 ;
  assign n26227 = n25319 | n26226 ;
  assign n25872 = n25319 & n43795 ;
  assign n44238 = ~n25839 ;
  assign n25873 = n44238 & n25872 ;
  assign n26228 = n25873 & n135 ;
  assign n44239 = ~n26228 ;
  assign n26229 = n26227 & n44239 ;
  assign n26730 = n6600 | n26729 ;
  assign n44240 = ~n26730 ;
  assign n26745 = n44240 & n26742 ;
  assign n26746 = n26229 | n26745 ;
  assign n44241 = ~n26744 ;
  assign n26747 = n44241 & n26746 ;
  assign n44242 = ~n26747 ;
  assign n26748 = n165 & n44242 ;
  assign n44243 = ~n25859 ;
  assign n25869 = n25375 & n44243 ;
  assign n25870 = n43784 & n25869 ;
  assign n26222 = n25870 & n135 ;
  assign n25871 = n25842 | n25859 ;
  assign n44244 = ~n25871 ;
  assign n26371 = n44244 & n135 ;
  assign n26372 = n25375 | n26371 ;
  assign n44245 = ~n26222 ;
  assign n26373 = n44245 & n26372 ;
  assign n44246 = ~n26739 ;
  assign n26756 = n26727 & n44246 ;
  assign n44247 = ~n26756 ;
  assign n26757 = n163 & n44247 ;
  assign n44248 = ~n26757 ;
  assign n26758 = n26742 & n44248 ;
  assign n44249 = ~n26758 ;
  assign n26759 = n6600 & n44249 ;
  assign n26760 = n165 | n26759 ;
  assign n44250 = ~n26760 ;
  assign n26761 = n26746 & n44250 ;
  assign n26762 = n26373 | n26761 ;
  assign n44251 = ~n26748 ;
  assign n26763 = n44251 & n26762 ;
  assign n44252 = ~n26763 ;
  assign n26764 = n166 & n44252 ;
  assign n25868 = n25862 | n25863 ;
  assign n44253 = ~n25868 ;
  assign n26344 = n44253 & n135 ;
  assign n26345 = n25531 | n26344 ;
  assign n25897 = n25531 & n43811 ;
  assign n44254 = ~n25863 ;
  assign n25898 = n44254 & n25897 ;
  assign n26472 = n25898 & n26442 ;
  assign n44255 = ~n26472 ;
  assign n26473 = n26345 & n44255 ;
  assign n26749 = n166 | n26748 ;
  assign n44256 = ~n26749 ;
  assign n26765 = n44256 & n26762 ;
  assign n26766 = n26473 | n26765 ;
  assign n44257 = ~n26764 ;
  assign n26767 = n44257 & n26766 ;
  assign n44258 = ~n26767 ;
  assign n26768 = n5352 & n44258 ;
  assign n44259 = ~n25884 ;
  assign n25894 = n25383 & n44259 ;
  assign n25895 = n43800 & n25894 ;
  assign n26374 = n25895 & n135 ;
  assign n25896 = n25866 | n25884 ;
  assign n44260 = ~n25896 ;
  assign n26377 = n44260 & n135 ;
  assign n26378 = n25383 | n26377 ;
  assign n44261 = ~n26374 ;
  assign n26379 = n44261 & n26378 ;
  assign n44262 = ~n26759 ;
  assign n26776 = n26746 & n44262 ;
  assign n44263 = ~n26776 ;
  assign n26777 = n165 & n44263 ;
  assign n44264 = ~n26777 ;
  assign n26778 = n26762 & n44264 ;
  assign n44265 = ~n26778 ;
  assign n26779 = n166 & n44265 ;
  assign n26780 = n5352 | n26779 ;
  assign n44266 = ~n26780 ;
  assign n26781 = n26766 & n44266 ;
  assign n26782 = n26379 | n26781 ;
  assign n44267 = ~n26768 ;
  assign n26783 = n44267 & n26782 ;
  assign n44268 = ~n26783 ;
  assign n26784 = n168 & n44268 ;
  assign n25921 = n25535 & n43827 ;
  assign n44269 = ~n25888 ;
  assign n25922 = n44269 & n25921 ;
  assign n26380 = n25922 & n135 ;
  assign n25893 = n25887 | n25888 ;
  assign n44270 = ~n25893 ;
  assign n26381 = n44270 & n135 ;
  assign n26382 = n25535 | n26381 ;
  assign n44271 = ~n26380 ;
  assign n26383 = n44271 & n26382 ;
  assign n26769 = n4934 | n26768 ;
  assign n44272 = ~n26769 ;
  assign n26785 = n44272 & n26782 ;
  assign n26786 = n26383 | n26785 ;
  assign n44273 = ~n26784 ;
  assign n26787 = n44273 & n26786 ;
  assign n44274 = ~n26787 ;
  assign n26788 = n169 & n44274 ;
  assign n44275 = ~n25908 ;
  assign n25918 = n25381 & n44275 ;
  assign n25919 = n43816 & n25918 ;
  assign n26289 = n25919 & n135 ;
  assign n25920 = n25891 | n25908 ;
  assign n44276 = ~n25920 ;
  assign n26384 = n44276 & n135 ;
  assign n26385 = n25381 | n26384 ;
  assign n44277 = ~n26289 ;
  assign n26386 = n44277 & n26385 ;
  assign n44278 = ~n26779 ;
  assign n26796 = n26766 & n44278 ;
  assign n44279 = ~n26796 ;
  assign n26797 = n167 & n44279 ;
  assign n44280 = ~n26797 ;
  assign n26798 = n26782 & n44280 ;
  assign n44281 = ~n26798 ;
  assign n26799 = n4934 & n44281 ;
  assign n26800 = n169 | n26799 ;
  assign n44282 = ~n26800 ;
  assign n26801 = n26786 & n44282 ;
  assign n26802 = n26386 | n26801 ;
  assign n44283 = ~n26788 ;
  assign n26803 = n44283 & n26802 ;
  assign n44284 = ~n26803 ;
  assign n26804 = n170 & n44284 ;
  assign n25945 = n25519 & n43843 ;
  assign n44285 = ~n25912 ;
  assign n25946 = n44285 & n25945 ;
  assign n26387 = n25946 & n135 ;
  assign n25917 = n25911 | n25912 ;
  assign n44286 = ~n25917 ;
  assign n26388 = n44286 & n135 ;
  assign n26389 = n25519 | n26388 ;
  assign n44287 = ~n26387 ;
  assign n26390 = n44287 & n26389 ;
  assign n26789 = n170 | n26788 ;
  assign n44288 = ~n26789 ;
  assign n26805 = n44288 & n26802 ;
  assign n26806 = n26390 | n26805 ;
  assign n44289 = ~n26804 ;
  assign n26807 = n44289 & n26806 ;
  assign n44290 = ~n26807 ;
  assign n26808 = n3940 & n44290 ;
  assign n25944 = n25915 | n25932 ;
  assign n44291 = ~n25944 ;
  assign n26297 = n44291 & n135 ;
  assign n26298 = n25461 | n26297 ;
  assign n44292 = ~n25932 ;
  assign n25942 = n25461 & n44292 ;
  assign n25943 = n43832 & n25942 ;
  assign n26468 = n25943 & n26442 ;
  assign n44293 = ~n26468 ;
  assign n26469 = n26298 & n44293 ;
  assign n44294 = ~n26799 ;
  assign n26816 = n26786 & n44294 ;
  assign n44295 = ~n26816 ;
  assign n26817 = n169 & n44295 ;
  assign n44296 = ~n26817 ;
  assign n26818 = n26802 & n44296 ;
  assign n44297 = ~n26818 ;
  assign n26819 = n170 & n44297 ;
  assign n26820 = n3940 | n26819 ;
  assign n44298 = ~n26820 ;
  assign n26821 = n26806 & n44298 ;
  assign n26822 = n26469 | n26821 ;
  assign n44299 = ~n26808 ;
  assign n26823 = n44299 & n26822 ;
  assign n44300 = ~n26823 ;
  assign n26824 = n172 & n44300 ;
  assign n25969 = n25466 & n43859 ;
  assign n44301 = ~n25936 ;
  assign n25970 = n44301 & n25969 ;
  assign n26321 = n25970 & n135 ;
  assign n25937 = n25935 | n25936 ;
  assign n44302 = ~n25937 ;
  assign n26391 = n44302 & n135 ;
  assign n26392 = n25466 | n26391 ;
  assign n44303 = ~n26321 ;
  assign n26393 = n44303 & n26392 ;
  assign n26809 = n3631 | n26808 ;
  assign n44304 = ~n26809 ;
  assign n26825 = n44304 & n26822 ;
  assign n26826 = n26393 | n26825 ;
  assign n44305 = ~n26824 ;
  assign n26827 = n44305 & n26826 ;
  assign n44306 = ~n26827 ;
  assign n26828 = n173 & n44306 ;
  assign n25968 = n25940 | n25956 ;
  assign n44307 = ~n25968 ;
  assign n26324 = n44307 & n135 ;
  assign n26325 = n25469 | n26324 ;
  assign n44308 = ~n25956 ;
  assign n25966 = n25469 & n44308 ;
  assign n25967 = n43848 & n25966 ;
  assign n26397 = n25967 & n135 ;
  assign n44309 = ~n26397 ;
  assign n26398 = n26325 & n44309 ;
  assign n44310 = ~n26819 ;
  assign n26836 = n26806 & n44310 ;
  assign n44311 = ~n26836 ;
  assign n26837 = n171 & n44311 ;
  assign n44312 = ~n26837 ;
  assign n26838 = n26822 & n44312 ;
  assign n44313 = ~n26838 ;
  assign n26839 = n3631 & n44313 ;
  assign n26840 = n173 | n26839 ;
  assign n44314 = ~n26840 ;
  assign n26841 = n26826 & n44314 ;
  assign n26842 = n26398 | n26841 ;
  assign n44315 = ~n26828 ;
  assign n26843 = n44315 & n26842 ;
  assign n44316 = ~n26843 ;
  assign n26844 = n174 & n44316 ;
  assign n25965 = n25959 | n25960 ;
  assign n44317 = ~n25965 ;
  assign n26401 = n44317 & n135 ;
  assign n26402 = n25471 | n26401 ;
  assign n25993 = n25471 & n43875 ;
  assign n44318 = ~n25960 ;
  assign n25994 = n44318 & n25993 ;
  assign n26464 = n25994 & n26442 ;
  assign n44319 = ~n26464 ;
  assign n26465 = n26402 & n44319 ;
  assign n26829 = n174 | n26828 ;
  assign n44320 = ~n26829 ;
  assign n26845 = n44320 & n26842 ;
  assign n26846 = n26465 | n26845 ;
  assign n44321 = ~n26844 ;
  assign n26847 = n44321 & n26846 ;
  assign n44322 = ~n26847 ;
  assign n26848 = n2753 & n44322 ;
  assign n25992 = n25963 | n25980 ;
  assign n44323 = ~n25992 ;
  assign n26375 = n44323 & n135 ;
  assign n26376 = n25475 | n26375 ;
  assign n44324 = ~n25980 ;
  assign n25990 = n25475 & n44324 ;
  assign n25991 = n43864 & n25990 ;
  assign n26403 = n25991 & n135 ;
  assign n44325 = ~n26403 ;
  assign n26404 = n26376 & n44325 ;
  assign n44326 = ~n26839 ;
  assign n26856 = n26826 & n44326 ;
  assign n44327 = ~n26856 ;
  assign n26857 = n173 & n44327 ;
  assign n44328 = ~n26857 ;
  assign n26858 = n26842 & n44328 ;
  assign n44329 = ~n26858 ;
  assign n26859 = n174 & n44329 ;
  assign n26860 = n2753 | n26859 ;
  assign n44330 = ~n26860 ;
  assign n26861 = n26846 & n44330 ;
  assign n26862 = n26404 | n26861 ;
  assign n44331 = ~n26848 ;
  assign n26863 = n44331 & n26862 ;
  assign n44332 = ~n26863 ;
  assign n26864 = n176 & n44332 ;
  assign n26017 = n25529 & n43891 ;
  assign n44333 = ~n25984 ;
  assign n26018 = n44333 & n26017 ;
  assign n26331 = n26018 & n135 ;
  assign n25989 = n25983 | n25984 ;
  assign n44334 = ~n25989 ;
  assign n26405 = n44334 & n135 ;
  assign n26406 = n25529 | n26405 ;
  assign n44335 = ~n26331 ;
  assign n26407 = n44335 & n26406 ;
  assign n26849 = n2431 | n26848 ;
  assign n44336 = ~n26849 ;
  assign n26865 = n44336 & n26862 ;
  assign n26867 = n26407 | n26865 ;
  assign n44337 = ~n26864 ;
  assign n26868 = n44337 & n26867 ;
  assign n44338 = ~n26868 ;
  assign n26869 = n177 & n44338 ;
  assign n26016 = n25987 | n26004 ;
  assign n44339 = ~n26016 ;
  assign n26355 = n44339 & n135 ;
  assign n26356 = n25410 | n26355 ;
  assign n44340 = ~n26004 ;
  assign n26014 = n25410 & n44340 ;
  assign n26015 = n43880 & n26014 ;
  assign n26408 = n26015 & n135 ;
  assign n44341 = ~n26408 ;
  assign n26409 = n26356 & n44341 ;
  assign n44342 = ~n26859 ;
  assign n26876 = n26846 & n44342 ;
  assign n44343 = ~n26876 ;
  assign n26877 = n175 & n44343 ;
  assign n44344 = ~n26877 ;
  assign n26878 = n26862 & n44344 ;
  assign n44345 = ~n26878 ;
  assign n26879 = n2431 & n44345 ;
  assign n26880 = n177 | n26879 ;
  assign n44346 = ~n26880 ;
  assign n26881 = n26867 & n44346 ;
  assign n26882 = n26409 | n26881 ;
  assign n44347 = ~n26869 ;
  assign n26883 = n44347 & n26882 ;
  assign n44348 = ~n26883 ;
  assign n26884 = n178 & n44348 ;
  assign n26041 = n25548 & n43907 ;
  assign n44349 = ~n26008 ;
  assign n26042 = n44349 & n26041 ;
  assign n26410 = n26042 & n135 ;
  assign n26013 = n26007 | n26008 ;
  assign n44350 = ~n26013 ;
  assign n26411 = n44350 & n135 ;
  assign n26412 = n25548 | n26411 ;
  assign n44351 = ~n26410 ;
  assign n26413 = n44351 & n26412 ;
  assign n26870 = n178 | n26869 ;
  assign n44352 = ~n26870 ;
  assign n26885 = n44352 & n26882 ;
  assign n26887 = n26413 | n26885 ;
  assign n44353 = ~n26884 ;
  assign n26888 = n44353 & n26887 ;
  assign n44354 = ~n26888 ;
  assign n26889 = n1707 & n44354 ;
  assign n26040 = n26011 | n26028 ;
  assign n44355 = ~n26040 ;
  assign n26277 = n44355 & n135 ;
  assign n26278 = n25481 | n26277 ;
  assign n44356 = ~n26028 ;
  assign n26038 = n25481 & n44356 ;
  assign n26039 = n43896 & n26038 ;
  assign n26285 = n26039 & n135 ;
  assign n44357 = ~n26285 ;
  assign n26286 = n26278 & n44357 ;
  assign n44358 = ~n26879 ;
  assign n26896 = n26867 & n44358 ;
  assign n44359 = ~n26896 ;
  assign n26897 = n177 & n44359 ;
  assign n44360 = ~n26897 ;
  assign n26898 = n26882 & n44360 ;
  assign n44361 = ~n26898 ;
  assign n26899 = n178 & n44361 ;
  assign n26900 = n1707 | n26899 ;
  assign n44362 = ~n26900 ;
  assign n26901 = n26887 & n44362 ;
  assign n26902 = n26286 | n26901 ;
  assign n44363 = ~n26889 ;
  assign n26903 = n44363 & n26902 ;
  assign n44364 = ~n26903 ;
  assign n26904 = n180 & n44364 ;
  assign n26037 = n26031 | n26032 ;
  assign n44365 = ~n26037 ;
  assign n26265 = n44365 & n135 ;
  assign n26266 = n25550 | n26265 ;
  assign n26065 = n25550 & n43923 ;
  assign n44366 = ~n26032 ;
  assign n26066 = n44366 & n26065 ;
  assign n26466 = n26066 & n26442 ;
  assign n44367 = ~n26466 ;
  assign n26467 = n26266 & n44367 ;
  assign n26890 = n1487 | n26889 ;
  assign n44368 = ~n26890 ;
  assign n26905 = n44368 & n26902 ;
  assign n26906 = n26467 | n26905 ;
  assign n44369 = ~n26904 ;
  assign n26907 = n44369 & n26906 ;
  assign n44370 = ~n26907 ;
  assign n26908 = n181 & n44370 ;
  assign n44371 = ~n26052 ;
  assign n26062 = n25491 & n44371 ;
  assign n26063 = n43912 & n26062 ;
  assign n26414 = n26063 & n135 ;
  assign n26064 = n26035 | n26052 ;
  assign n44372 = ~n26064 ;
  assign n26415 = n44372 & n135 ;
  assign n26416 = n25491 | n26415 ;
  assign n44373 = ~n26414 ;
  assign n26417 = n44373 & n26416 ;
  assign n44374 = ~n26899 ;
  assign n26916 = n26887 & n44374 ;
  assign n44375 = ~n26916 ;
  assign n26917 = n179 & n44375 ;
  assign n44376 = ~n26917 ;
  assign n26918 = n26902 & n44376 ;
  assign n44377 = ~n26918 ;
  assign n26919 = n1487 & n44377 ;
  assign n26920 = n181 | n26919 ;
  assign n44378 = ~n26920 ;
  assign n26921 = n26906 & n44378 ;
  assign n26922 = n26417 | n26921 ;
  assign n44379 = ~n26908 ;
  assign n26923 = n44379 & n26922 ;
  assign n44380 = ~n26923 ;
  assign n26924 = n182 & n44380 ;
  assign n26061 = n26055 | n26056 ;
  assign n44381 = ~n26061 ;
  assign n26362 = n44381 & n135 ;
  assign n26363 = n25494 | n26362 ;
  assign n26089 = n25494 & n43939 ;
  assign n44382 = ~n26056 ;
  assign n26090 = n44382 & n26089 ;
  assign n26418 = n26090 & n135 ;
  assign n44383 = ~n26418 ;
  assign n26419 = n26363 & n44383 ;
  assign n26909 = n182 | n26908 ;
  assign n44384 = ~n26909 ;
  assign n26925 = n44384 & n26922 ;
  assign n26926 = n26419 | n26925 ;
  assign n44385 = ~n26924 ;
  assign n26927 = n44385 & n26926 ;
  assign n44386 = ~n26927 ;
  assign n26928 = n996 & n44386 ;
  assign n44387 = ~n26076 ;
  assign n26086 = n25498 & n44387 ;
  assign n26087 = n43928 & n26086 ;
  assign n26338 = n26087 & n135 ;
  assign n26088 = n26059 | n26076 ;
  assign n44388 = ~n26088 ;
  assign n26394 = n44388 & n135 ;
  assign n26395 = n25498 | n26394 ;
  assign n44389 = ~n26338 ;
  assign n26396 = n44389 & n26395 ;
  assign n44390 = ~n26919 ;
  assign n26936 = n26906 & n44390 ;
  assign n44391 = ~n26936 ;
  assign n26937 = n181 & n44391 ;
  assign n44392 = ~n26937 ;
  assign n26938 = n26922 & n44392 ;
  assign n44393 = ~n26938 ;
  assign n26939 = n182 & n44393 ;
  assign n26940 = n183 | n26939 ;
  assign n44394 = ~n26940 ;
  assign n26941 = n26926 & n44394 ;
  assign n26942 = n26396 | n26941 ;
  assign n44395 = ~n26928 ;
  assign n26943 = n44395 & n26942 ;
  assign n44396 = ~n26943 ;
  assign n26944 = n184 & n44396 ;
  assign n26113 = n25503 & n43955 ;
  assign n44397 = ~n26080 ;
  assign n26114 = n44397 & n26113 ;
  assign n26420 = n26114 & n135 ;
  assign n26085 = n26079 | n26080 ;
  assign n44398 = ~n26085 ;
  assign n26421 = n44398 & n135 ;
  assign n26422 = n25503 | n26421 ;
  assign n44399 = ~n26420 ;
  assign n26423 = n44399 & n26422 ;
  assign n26929 = n838 | n26928 ;
  assign n44400 = ~n26929 ;
  assign n26945 = n44400 & n26942 ;
  assign n26946 = n26423 | n26945 ;
  assign n44401 = ~n26944 ;
  assign n26947 = n44401 & n26946 ;
  assign n44402 = ~n26947 ;
  assign n26948 = n185 & n44402 ;
  assign n26112 = n26083 | n26100 ;
  assign n44403 = ~n26112 ;
  assign n26245 = n44403 & n135 ;
  assign n26246 = n25505 | n26245 ;
  assign n44404 = ~n26100 ;
  assign n26110 = n25505 & n44404 ;
  assign n26111 = n43944 & n26110 ;
  assign n26424 = n26111 & n135 ;
  assign n44405 = ~n26424 ;
  assign n26425 = n26246 & n44405 ;
  assign n44406 = ~n26939 ;
  assign n26956 = n26926 & n44406 ;
  assign n44407 = ~n26956 ;
  assign n26957 = n183 & n44407 ;
  assign n44408 = ~n26957 ;
  assign n26958 = n26942 & n44408 ;
  assign n44409 = ~n26958 ;
  assign n26959 = n838 & n44409 ;
  assign n26960 = n185 | n26959 ;
  assign n44410 = ~n26960 ;
  assign n26961 = n26946 & n44410 ;
  assign n26962 = n26425 | n26961 ;
  assign n44411 = ~n26948 ;
  assign n26963 = n44411 & n26962 ;
  assign n44412 = ~n26963 ;
  assign n26964 = n186 & n44412 ;
  assign n26109 = n26103 | n26104 ;
  assign n44413 = ~n26109 ;
  assign n26300 = n44413 & n135 ;
  assign n26301 = n25552 | n26300 ;
  assign n26137 = n25552 & n43971 ;
  assign n44414 = ~n26104 ;
  assign n26138 = n44414 & n26137 ;
  assign n26426 = n26138 & n135 ;
  assign n44415 = ~n26426 ;
  assign n26427 = n26301 & n44415 ;
  assign n26949 = n186 | n26948 ;
  assign n44416 = ~n26949 ;
  assign n26965 = n44416 & n26962 ;
  assign n26966 = n26427 | n26965 ;
  assign n44417 = ~n26964 ;
  assign n26967 = n44417 & n26966 ;
  assign n44418 = ~n26967 ;
  assign n26968 = n528 & n44418 ;
  assign n26969 = n413 | n26968 ;
  assign n44419 = ~n26124 ;
  assign n26134 = n25508 & n44419 ;
  assign n26135 = n43960 & n26134 ;
  assign n26290 = n26135 & n135 ;
  assign n26136 = n26107 | n26124 ;
  assign n44420 = ~n26136 ;
  assign n26428 = n44420 & n135 ;
  assign n26429 = n25508 | n26428 ;
  assign n44421 = ~n26290 ;
  assign n26430 = n44421 & n26429 ;
  assign n44422 = ~n26959 ;
  assign n26976 = n26946 & n44422 ;
  assign n44423 = ~n26976 ;
  assign n26977 = n185 & n44423 ;
  assign n44424 = ~n26977 ;
  assign n26978 = n26962 & n44424 ;
  assign n44425 = ~n26978 ;
  assign n26979 = n186 & n44425 ;
  assign n26980 = n528 | n26979 ;
  assign n44426 = ~n26980 ;
  assign n26981 = n26966 & n44426 ;
  assign n26982 = n26430 | n26981 ;
  assign n44427 = ~n26969 ;
  assign n26985 = n44427 & n26982 ;
  assign n26133 = n26127 | n26128 ;
  assign n44428 = ~n26133 ;
  assign n26273 = n44428 & n135 ;
  assign n26274 = n25451 | n26273 ;
  assign n26161 = n25451 & n43987 ;
  assign n44429 = ~n26128 ;
  assign n26162 = n44429 & n26161 ;
  assign n26431 = n26162 & n135 ;
  assign n44430 = ~n26431 ;
  assign n26432 = n26274 & n44430 ;
  assign n44431 = ~n26979 ;
  assign n26996 = n26966 & n44431 ;
  assign n44432 = ~n26996 ;
  assign n26997 = n187 & n44432 ;
  assign n44433 = ~n26997 ;
  assign n26998 = n26982 & n44433 ;
  assign n44434 = ~n26998 ;
  assign n26999 = n413 & n44434 ;
  assign n44435 = ~n26999 ;
  assign n27014 = n26432 & n44435 ;
  assign n44436 = ~n26985 ;
  assign n27015 = n44436 & n27014 ;
  assign n26200 = n25404 | n26198 ;
  assign n26201 = n192 & n26200 ;
  assign n44437 = ~n25404 ;
  assign n26443 = n44437 & n26442 ;
  assign n44438 = ~n26443 ;
  assign n26444 = n26198 & n44438 ;
  assign n44439 = ~n26444 ;
  assign n26445 = n26201 & n44439 ;
  assign n26195 = n25513 & n44007 ;
  assign n26202 = n43997 & n26190 ;
  assign n44440 = ~n26202 ;
  assign n26203 = n26195 & n44440 ;
  assign n26448 = n26203 & n26442 ;
  assign n26204 = n26192 | n26202 ;
  assign n44441 = ~n26204 ;
  assign n26474 = n44441 & n26442 ;
  assign n26475 = n25513 | n26474 ;
  assign n44442 = ~n26448 ;
  assign n26476 = n44442 & n26475 ;
  assign n44443 = ~n26968 ;
  assign n26983 = n44443 & n26982 ;
  assign n44444 = ~n26983 ;
  assign n26984 = n188 & n44444 ;
  assign n26986 = n26432 | n26985 ;
  assign n44445 = ~n26984 ;
  assign n26987 = n44445 & n26986 ;
  assign n44446 = ~n26987 ;
  assign n26988 = n189 & n44446 ;
  assign n26160 = n26131 | n26148 ;
  assign n44447 = ~n26160 ;
  assign n26399 = n44447 & n135 ;
  assign n26400 = n25511 | n26399 ;
  assign n44448 = ~n26148 ;
  assign n26158 = n25511 & n44448 ;
  assign n26159 = n43976 & n26158 ;
  assign n26433 = n26159 & n135 ;
  assign n44449 = ~n26433 ;
  assign n26434 = n26400 & n44449 ;
  assign n27000 = n189 | n26999 ;
  assign n44450 = ~n27000 ;
  assign n27001 = n26986 & n44450 ;
  assign n27002 = n26434 | n27001 ;
  assign n44451 = ~n26988 ;
  assign n27003 = n44451 & n27002 ;
  assign n44452 = ~n27003 ;
  assign n27004 = n190 & n44452 ;
  assign n26182 = n25485 & n44003 ;
  assign n44453 = ~n26152 ;
  assign n26183 = n44453 & n26182 ;
  assign n26370 = n26183 & n135 ;
  assign n26184 = n26152 | n26170 ;
  assign n44454 = ~n26184 ;
  assign n26435 = n44454 & n135 ;
  assign n26436 = n25485 | n26435 ;
  assign n44455 = ~n26370 ;
  assign n26437 = n44455 & n26436 ;
  assign n26989 = n190 | n26988 ;
  assign n44456 = ~n26989 ;
  assign n27005 = n44456 & n27002 ;
  assign n27006 = n26437 | n27005 ;
  assign n44457 = ~n27004 ;
  assign n27007 = n44457 & n27006 ;
  assign n44458 = ~n27007 ;
  assign n27008 = n287 & n44458 ;
  assign n44459 = ~n27008 ;
  assign n27009 = n26476 & n44459 ;
  assign n44460 = ~n26172 ;
  assign n26179 = n25500 & n44460 ;
  assign n26180 = n43992 & n26179 ;
  assign n26367 = n26180 & n135 ;
  assign n26181 = n26155 | n26172 ;
  assign n44461 = ~n26181 ;
  assign n26438 = n44461 & n135 ;
  assign n26439 = n25500 | n26438 ;
  assign n44462 = ~n26367 ;
  assign n26440 = n44462 & n26439 ;
  assign n27016 = n26986 & n44435 ;
  assign n44463 = ~n27016 ;
  assign n27017 = n189 & n44463 ;
  assign n44464 = ~n27017 ;
  assign n27018 = n27002 & n44464 ;
  assign n44465 = ~n27018 ;
  assign n27019 = n190 & n44465 ;
  assign n27020 = n287 | n27019 ;
  assign n44466 = ~n27020 ;
  assign n27021 = n27006 & n44466 ;
  assign n27022 = n26440 | n27021 ;
  assign n27023 = n27009 & n27022 ;
  assign n27024 = n26445 | n27023 ;
  assign n44467 = ~n26200 ;
  assign n26259 = n44467 & n135 ;
  assign n26260 = n26199 | n26259 ;
  assign n26477 = n26260 | n26476 ;
  assign n27028 = n44459 & n27022 ;
  assign n27029 = n26477 | n27028 ;
  assign n27030 = n31336 & n27029 ;
  assign n134 = n27024 | n27030 ;
  assign n27126 = n27015 & n134 ;
  assign n26990 = n26984 | n26985 ;
  assign n44468 = ~n26990 ;
  assign n27225 = n44468 & n134 ;
  assign n27226 = n26432 | n27225 ;
  assign n44469 = ~n27126 ;
  assign n27227 = n44469 & n27226 ;
  assign n257 = x8 | x9 ;
  assign n258 = x10 | n257 ;
  assign n27130 = x10 & n134 ;
  assign n44470 = ~n27130 ;
  assign n27131 = n258 & n44470 ;
  assign n44471 = ~n27131 ;
  assign n27132 = n135 & n44471 ;
  assign n44472 = ~n254 ;
  assign n27055 = n44472 & n134 ;
  assign n44473 = ~x10 ;
  assign n27233 = n44473 & n134 ;
  assign n44474 = ~n27233 ;
  assign n27234 = x11 & n44474 ;
  assign n27235 = n27055 | n27234 ;
  assign n27302 = n258 & n44029 ;
  assign n27303 = n44030 & n27302 ;
  assign n27304 = n44031 & n27303 ;
  assign n27305 = n44032 & n27304 ;
  assign n27306 = n44470 & n27305 ;
  assign n27307 = n27235 | n27306 ;
  assign n44475 = ~n27132 ;
  assign n27308 = n44475 & n27307 ;
  assign n44476 = ~n27308 ;
  assign n27309 = n25517 & n44476 ;
  assign n44477 = ~n26445 ;
  assign n26446 = n135 & n44477 ;
  assign n44478 = ~n27023 ;
  assign n27254 = n26446 & n44478 ;
  assign n44479 = ~n27030 ;
  assign n27255 = n44479 & n27254 ;
  assign n27256 = n27055 | n27255 ;
  assign n27257 = x12 & n27256 ;
  assign n27258 = x12 | n27255 ;
  assign n27259 = n27055 | n27258 ;
  assign n44480 = ~n27257 ;
  assign n27260 = n44480 & n27259 ;
  assign n259 = n44473 & n257 ;
  assign n44481 = ~n134 ;
  assign n27244 = x10 & n44481 ;
  assign n27245 = n259 | n27244 ;
  assign n44482 = ~n27245 ;
  assign n27246 = n26442 & n44482 ;
  assign n27247 = n25517 | n27246 ;
  assign n44483 = ~n27247 ;
  assign n27312 = n44483 & n27307 ;
  assign n27313 = n27260 | n27312 ;
  assign n44484 = ~n27309 ;
  assign n27314 = n44484 & n27313 ;
  assign n44485 = ~n27314 ;
  assign n27315 = n137 & n44485 ;
  assign n26462 = n26330 | n26457 ;
  assign n44486 = ~n26462 ;
  assign n27109 = n44486 & n134 ;
  assign n27110 = n26335 | n27109 ;
  assign n26463 = n26335 & n44486 ;
  assign n27238 = n26463 & n134 ;
  assign n44487 = ~n27238 ;
  assign n27239 = n27110 & n44487 ;
  assign n27310 = n137 | n27309 ;
  assign n44488 = ~n27310 ;
  assign n27318 = n44488 & n27313 ;
  assign n27319 = n27239 | n27318 ;
  assign n44489 = ~n27315 ;
  assign n27320 = n44489 & n27319 ;
  assign n44490 = ~n27320 ;
  assign n27321 = n138 & n44490 ;
  assign n26461 = n26456 | n26459 ;
  assign n44491 = ~n26461 ;
  assign n27053 = n44491 & n134 ;
  assign n27054 = n26486 | n27053 ;
  assign n44492 = ~n26456 ;
  assign n26492 = n44492 & n26486 ;
  assign n44493 = ~n26459 ;
  assign n26493 = n44493 & n26492 ;
  assign n27103 = n26493 & n134 ;
  assign n44494 = ~n27103 ;
  assign n27104 = n27054 & n44494 ;
  assign n27316 = n138 | n27315 ;
  assign n44495 = ~n27316 ;
  assign n27322 = n44495 & n27319 ;
  assign n27323 = n27104 | n27322 ;
  assign n44496 = ~n27321 ;
  assign n27324 = n44496 & n27323 ;
  assign n44497 = ~n27324 ;
  assign n27325 = n22661 & n44497 ;
  assign n26507 = n26489 | n26505 ;
  assign n44498 = ~n26507 ;
  assign n27119 = n44498 & n134 ;
  assign n27120 = n26316 | n27119 ;
  assign n26490 = n26316 & n44040 ;
  assign n44499 = ~n26505 ;
  assign n26506 = n26490 & n44499 ;
  assign n27242 = n26506 & n134 ;
  assign n44500 = ~n27242 ;
  assign n27243 = n27120 & n44500 ;
  assign n27311 = n136 & n44476 ;
  assign n27133 = n136 | n27132 ;
  assign n44501 = ~n27133 ;
  assign n27335 = n44501 & n27307 ;
  assign n27336 = n27260 | n27335 ;
  assign n44502 = ~n27311 ;
  assign n27337 = n44502 & n27336 ;
  assign n44503 = ~n27337 ;
  assign n27338 = n137 & n44503 ;
  assign n27339 = n44488 & n27336 ;
  assign n27340 = n27239 | n27339 ;
  assign n44504 = ~n27338 ;
  assign n27341 = n44504 & n27340 ;
  assign n44505 = ~n27341 ;
  assign n27342 = n138 & n44505 ;
  assign n27343 = n139 | n27342 ;
  assign n44506 = ~n27343 ;
  assign n27344 = n27323 & n44506 ;
  assign n27345 = n27243 | n27344 ;
  assign n44507 = ~n27325 ;
  assign n27346 = n44507 & n27345 ;
  assign n44508 = ~n27346 ;
  assign n27347 = n140 & n44508 ;
  assign n44509 = ~n26522 ;
  assign n27295 = n26320 & n44509 ;
  assign n27296 = n44068 & n27295 ;
  assign n27297 = n134 & n27296 ;
  assign n27298 = n26510 | n26522 ;
  assign n44510 = ~n27298 ;
  assign n27299 = n134 & n44510 ;
  assign n27300 = n26320 | n27299 ;
  assign n44511 = ~n27297 ;
  assign n27301 = n44511 & n27300 ;
  assign n27327 = n140 | n27325 ;
  assign n44512 = ~n27327 ;
  assign n27348 = n44512 & n27345 ;
  assign n27349 = n27301 | n27348 ;
  assign n44513 = ~n27347 ;
  assign n27350 = n44513 & n27349 ;
  assign n44514 = ~n27350 ;
  assign n27351 = n141 & n44514 ;
  assign n26528 = n26525 | n26526 ;
  assign n44515 = ~n26528 ;
  assign n27046 = n44515 & n134 ;
  assign n27047 = n26308 | n27046 ;
  assign n26504 = n26308 & n44057 ;
  assign n44516 = ~n26526 ;
  assign n26527 = n26504 & n44516 ;
  assign n27092 = n26527 & n134 ;
  assign n44517 = ~n27092 ;
  assign n27093 = n27047 & n44517 ;
  assign n27359 = n44495 & n27340 ;
  assign n27360 = n27104 | n27359 ;
  assign n44518 = ~n27342 ;
  assign n27361 = n44518 & n27360 ;
  assign n44519 = ~n27361 ;
  assign n27362 = n139 & n44519 ;
  assign n27363 = n44506 & n27360 ;
  assign n27364 = n27243 | n27363 ;
  assign n44520 = ~n27362 ;
  assign n27365 = n44520 & n27364 ;
  assign n44521 = ~n27365 ;
  assign n27366 = n22030 & n44521 ;
  assign n27367 = n141 | n27366 ;
  assign n44522 = ~n27367 ;
  assign n27368 = n27349 & n44522 ;
  assign n27369 = n27093 | n27368 ;
  assign n44523 = ~n27351 ;
  assign n27370 = n44523 & n27369 ;
  assign n44524 = ~n27370 ;
  assign n27371 = n142 & n44524 ;
  assign n44525 = ~n26543 ;
  assign n27288 = n26323 & n44525 ;
  assign n27289 = n44081 & n27288 ;
  assign n27290 = n134 & n27289 ;
  assign n27291 = n26531 | n26543 ;
  assign n44526 = ~n27291 ;
  assign n27292 = n134 & n44526 ;
  assign n27293 = n26323 | n27292 ;
  assign n44527 = ~n27290 ;
  assign n27294 = n44527 & n27293 ;
  assign n27352 = n142 | n27351 ;
  assign n44528 = ~n27352 ;
  assign n27372 = n44528 & n27369 ;
  assign n27373 = n27294 | n27372 ;
  assign n44529 = ~n27371 ;
  assign n27374 = n44529 & n27373 ;
  assign n44530 = ~n27374 ;
  assign n27375 = n19362 & n44530 ;
  assign n26521 = n26329 & n44074 ;
  assign n44531 = ~n26547 ;
  assign n26548 = n26521 & n44531 ;
  assign n27094 = n26548 & n134 ;
  assign n26549 = n26546 | n26547 ;
  assign n44532 = ~n26549 ;
  assign n27113 = n44532 & n134 ;
  assign n27114 = n26329 | n27113 ;
  assign n44533 = ~n27094 ;
  assign n27115 = n44533 & n27114 ;
  assign n27383 = n44512 & n27364 ;
  assign n27384 = n27301 | n27383 ;
  assign n44534 = ~n27366 ;
  assign n27385 = n44534 & n27384 ;
  assign n44535 = ~n27385 ;
  assign n27386 = n141 & n44535 ;
  assign n27387 = n44522 & n27384 ;
  assign n27388 = n27093 | n27387 ;
  assign n44536 = ~n27386 ;
  assign n27389 = n44536 & n27388 ;
  assign n44537 = ~n27389 ;
  assign n27390 = n142 & n44537 ;
  assign n27391 = n143 | n27390 ;
  assign n44538 = ~n27391 ;
  assign n27392 = n27373 & n44538 ;
  assign n27393 = n27115 | n27392 ;
  assign n44539 = ~n27375 ;
  assign n27394 = n44539 & n27393 ;
  assign n44540 = ~n27394 ;
  assign n27395 = n144 & n44540 ;
  assign n44541 = ~n26565 ;
  assign n27281 = n26347 & n44541 ;
  assign n27282 = n44087 & n27281 ;
  assign n27283 = n134 & n27282 ;
  assign n27284 = n26552 | n26565 ;
  assign n44542 = ~n27284 ;
  assign n27285 = n134 & n44542 ;
  assign n27286 = n26347 | n27285 ;
  assign n44543 = ~n27283 ;
  assign n27287 = n44543 & n27286 ;
  assign n27376 = n144 | n27375 ;
  assign n44544 = ~n27376 ;
  assign n27396 = n44544 & n27393 ;
  assign n27397 = n27287 | n27396 ;
  assign n44545 = ~n27395 ;
  assign n27398 = n44545 & n27397 ;
  assign n44546 = ~n27398 ;
  assign n27399 = n145 & n44546 ;
  assign n26542 = n26343 & n44102 ;
  assign n44547 = ~n26569 ;
  assign n27275 = n26542 & n44547 ;
  assign n27276 = n134 & n27275 ;
  assign n27277 = n26540 | n26569 ;
  assign n44548 = ~n27277 ;
  assign n27278 = n134 & n44548 ;
  assign n27279 = n26343 | n27278 ;
  assign n44549 = ~n27276 ;
  assign n27280 = n44549 & n27279 ;
  assign n27407 = n44528 & n27388 ;
  assign n27408 = n27294 | n27407 ;
  assign n44550 = ~n27390 ;
  assign n27409 = n44550 & n27408 ;
  assign n44551 = ~n27409 ;
  assign n27410 = n143 & n44551 ;
  assign n27411 = n44538 & n27408 ;
  assign n27412 = n27115 | n27411 ;
  assign n44552 = ~n27410 ;
  assign n27413 = n44552 & n27412 ;
  assign n44553 = ~n27413 ;
  assign n27414 = n18797 & n44553 ;
  assign n27415 = n145 | n27414 ;
  assign n44554 = ~n27415 ;
  assign n27416 = n27397 & n44554 ;
  assign n27417 = n27280 | n27416 ;
  assign n44555 = ~n27399 ;
  assign n27418 = n44555 & n27417 ;
  assign n44556 = ~n27418 ;
  assign n27419 = n146 & n44556 ;
  assign n44557 = ~n26556 ;
  assign n26558 = n26351 & n44557 ;
  assign n27269 = n26558 & n44091 ;
  assign n27270 = n134 & n27269 ;
  assign n27271 = n26556 | n26572 ;
  assign n44558 = ~n27271 ;
  assign n27272 = n134 & n44558 ;
  assign n27273 = n26351 | n27272 ;
  assign n44559 = ~n27270 ;
  assign n27274 = n44559 & n27273 ;
  assign n27400 = n146 | n27399 ;
  assign n44560 = ~n27400 ;
  assign n27420 = n44560 & n27417 ;
  assign n27421 = n27274 | n27420 ;
  assign n44561 = ~n27419 ;
  assign n27422 = n44561 & n27421 ;
  assign n44562 = ~n27422 ;
  assign n27423 = n16322 & n44562 ;
  assign n26564 = n26471 & n44118 ;
  assign n44563 = ~n26576 ;
  assign n26594 = n26564 & n44563 ;
  assign n27137 = n26594 & n134 ;
  assign n26595 = n26574 | n26576 ;
  assign n44564 = ~n26595 ;
  assign n27143 = n44564 & n134 ;
  assign n27144 = n26471 | n27143 ;
  assign n44565 = ~n27137 ;
  assign n27145 = n44565 & n27144 ;
  assign n27431 = n44544 & n27412 ;
  assign n27432 = n27287 | n27431 ;
  assign n44566 = ~n27414 ;
  assign n27433 = n44566 & n27432 ;
  assign n44567 = ~n27433 ;
  assign n27434 = n145 & n44567 ;
  assign n27435 = n44554 & n27432 ;
  assign n27436 = n27280 | n27435 ;
  assign n44568 = ~n27434 ;
  assign n27437 = n44568 & n27436 ;
  assign n44569 = ~n27437 ;
  assign n27438 = n146 & n44569 ;
  assign n27439 = n147 | n27438 ;
  assign n44570 = ~n27439 ;
  assign n27440 = n27421 & n44570 ;
  assign n27441 = n27145 | n27440 ;
  assign n44571 = ~n27423 ;
  assign n27442 = n44571 & n27441 ;
  assign n44572 = ~n27442 ;
  assign n27443 = n148 & n44572 ;
  assign n26593 = n26579 | n26581 ;
  assign n44573 = ~n26593 ;
  assign n27117 = n44573 & n134 ;
  assign n27118 = n26359 | n27117 ;
  assign n44574 = ~n26581 ;
  assign n26591 = n26359 & n44574 ;
  assign n26592 = n44107 & n26591 ;
  assign n27154 = n26592 & n134 ;
  assign n44575 = ~n27154 ;
  assign n27155 = n27118 & n44575 ;
  assign n27425 = n148 | n27423 ;
  assign n44576 = ~n27425 ;
  assign n27444 = n44576 & n27441 ;
  assign n27445 = n27155 | n27444 ;
  assign n44577 = ~n27443 ;
  assign n27446 = n44577 & n27445 ;
  assign n44578 = ~n27446 ;
  assign n27447 = n149 & n44578 ;
  assign n26590 = n26584 | n26585 ;
  assign n44579 = ~n26590 ;
  assign n27146 = n44579 & n134 ;
  assign n27147 = n26334 | n27146 ;
  assign n26614 = n26334 & n44134 ;
  assign n44580 = ~n26585 ;
  assign n26615 = n44580 & n26614 ;
  assign n27156 = n26615 & n134 ;
  assign n44581 = ~n27156 ;
  assign n27157 = n27147 & n44581 ;
  assign n27455 = n44560 & n27436 ;
  assign n27456 = n27274 | n27455 ;
  assign n44582 = ~n27438 ;
  assign n27457 = n44582 & n27456 ;
  assign n44583 = ~n27457 ;
  assign n27458 = n147 & n44583 ;
  assign n27459 = n44570 & n27456 ;
  assign n27460 = n27145 | n27459 ;
  assign n44584 = ~n27458 ;
  assign n27461 = n44584 & n27460 ;
  assign n44585 = ~n27461 ;
  assign n27462 = n15807 & n44585 ;
  assign n27463 = n149 | n27462 ;
  assign n44586 = ~n27463 ;
  assign n27464 = n27445 & n44586 ;
  assign n27465 = n27157 | n27464 ;
  assign n44587 = ~n27447 ;
  assign n27466 = n44587 & n27465 ;
  assign n44588 = ~n27466 ;
  assign n27467 = n150 & n44588 ;
  assign n44589 = ~n26601 ;
  assign n26611 = n26366 & n44589 ;
  assign n26612 = n44123 & n26611 ;
  assign n27083 = n26612 & n134 ;
  assign n26613 = n26588 | n26601 ;
  assign n44590 = ~n26613 ;
  assign n27086 = n44590 & n134 ;
  assign n27087 = n26366 | n27086 ;
  assign n44591 = ~n27083 ;
  assign n27088 = n44591 & n27087 ;
  assign n27448 = n150 | n27447 ;
  assign n44592 = ~n27448 ;
  assign n27468 = n44592 & n27465 ;
  assign n27469 = n27088 | n27468 ;
  assign n44593 = ~n27467 ;
  assign n27470 = n44593 & n27469 ;
  assign n44594 = ~n27470 ;
  assign n27471 = n13662 & n44594 ;
  assign n26610 = n26604 | n26605 ;
  assign n44595 = ~n26610 ;
  assign n27068 = n44595 & n134 ;
  assign n27069 = n26369 | n27068 ;
  assign n26634 = n26369 & n44150 ;
  assign n44596 = ~n26605 ;
  assign n26635 = n44596 & n26634 ;
  assign n27081 = n26635 & n134 ;
  assign n44597 = ~n27081 ;
  assign n27082 = n27069 & n44597 ;
  assign n27479 = n44576 & n27460 ;
  assign n27480 = n27155 | n27479 ;
  assign n44598 = ~n27462 ;
  assign n27481 = n44598 & n27480 ;
  assign n44599 = ~n27481 ;
  assign n27482 = n149 & n44599 ;
  assign n27483 = n44586 & n27480 ;
  assign n27484 = n27157 | n27483 ;
  assign n44600 = ~n27482 ;
  assign n27485 = n44600 & n27484 ;
  assign n44601 = ~n27485 ;
  assign n27486 = n150 & n44601 ;
  assign n27487 = n151 | n27486 ;
  assign n44602 = ~n27487 ;
  assign n27488 = n27469 & n44602 ;
  assign n27489 = n27082 | n27488 ;
  assign n44603 = ~n27471 ;
  assign n27490 = n44603 & n27489 ;
  assign n44604 = ~n27490 ;
  assign n27491 = n152 & n44604 ;
  assign n44605 = ~n26621 ;
  assign n26631 = n26292 & n44605 ;
  assign n26632 = n44139 & n26631 ;
  assign n27076 = n26632 & n134 ;
  assign n26633 = n26608 | n26621 ;
  assign n44606 = ~n26633 ;
  assign n27078 = n44606 & n134 ;
  assign n27079 = n26292 | n27078 ;
  assign n44607 = ~n27076 ;
  assign n27080 = n44607 & n27079 ;
  assign n27472 = n152 | n27471 ;
  assign n44608 = ~n27472 ;
  assign n27492 = n44608 & n27489 ;
  assign n27493 = n27080 | n27492 ;
  assign n44609 = ~n27491 ;
  assign n27494 = n44609 & n27493 ;
  assign n44610 = ~n27494 ;
  assign n27495 = n153 & n44610 ;
  assign n26654 = n26304 & n44166 ;
  assign n44611 = ~n26625 ;
  assign n26655 = n44611 & n26654 ;
  assign n27072 = n26655 & n134 ;
  assign n26630 = n26624 | n26625 ;
  assign n44612 = ~n26630 ;
  assign n27073 = n44612 & n134 ;
  assign n27074 = n26304 | n27073 ;
  assign n44613 = ~n27072 ;
  assign n27075 = n44613 & n27074 ;
  assign n27503 = n44592 & n27484 ;
  assign n27504 = n27088 | n27503 ;
  assign n44614 = ~n27486 ;
  assign n27505 = n44614 & n27504 ;
  assign n44615 = ~n27505 ;
  assign n27506 = n151 & n44615 ;
  assign n27507 = n44602 & n27504 ;
  assign n27508 = n27082 | n27507 ;
  assign n44616 = ~n27506 ;
  assign n27509 = n44616 & n27508 ;
  assign n44617 = ~n27509 ;
  assign n27510 = n13079 & n44617 ;
  assign n27511 = n153 | n27510 ;
  assign n44618 = ~n27511 ;
  assign n27512 = n27493 & n44618 ;
  assign n27513 = n27075 | n27512 ;
  assign n44619 = ~n27495 ;
  assign n27514 = n44619 & n27513 ;
  assign n44620 = ~n27514 ;
  assign n27515 = n154 & n44620 ;
  assign n26653 = n26628 | n26641 ;
  assign n44621 = ~n26653 ;
  assign n27066 = n44621 & n134 ;
  assign n27067 = n26282 | n27066 ;
  assign n44622 = ~n26641 ;
  assign n26651 = n26282 & n44622 ;
  assign n26652 = n44155 & n26651 ;
  assign n27111 = n26652 & n134 ;
  assign n44623 = ~n27111 ;
  assign n27112 = n27067 & n44623 ;
  assign n27496 = n154 | n27495 ;
  assign n44624 = ~n27496 ;
  assign n27516 = n44624 & n27513 ;
  assign n27517 = n27112 | n27516 ;
  assign n44625 = ~n27515 ;
  assign n27518 = n44625 & n27517 ;
  assign n44626 = ~n27518 ;
  assign n27519 = n11067 & n44626 ;
  assign n26674 = n26276 & n44182 ;
  assign n44627 = ~n26645 ;
  assign n26675 = n44627 & n26674 ;
  assign n27045 = n26675 & n134 ;
  assign n26650 = n26644 | n26645 ;
  assign n44628 = ~n26650 ;
  assign n27127 = n44628 & n134 ;
  assign n27128 = n26276 | n27127 ;
  assign n44629 = ~n27045 ;
  assign n27129 = n44629 & n27128 ;
  assign n27527 = n44608 & n27508 ;
  assign n27528 = n27080 | n27527 ;
  assign n44630 = ~n27510 ;
  assign n27529 = n44630 & n27528 ;
  assign n44631 = ~n27529 ;
  assign n27530 = n153 & n44631 ;
  assign n27531 = n44618 & n27528 ;
  assign n27532 = n27075 | n27531 ;
  assign n44632 = ~n27530 ;
  assign n27533 = n44632 & n27532 ;
  assign n44633 = ~n27533 ;
  assign n27534 = n154 & n44633 ;
  assign n27535 = n11067 | n27534 ;
  assign n44634 = ~n27535 ;
  assign n27536 = n27517 & n44634 ;
  assign n27537 = n27129 | n27536 ;
  assign n44635 = ~n27519 ;
  assign n27538 = n44635 & n27537 ;
  assign n44636 = ~n27538 ;
  assign n27539 = n156 & n44636 ;
  assign n44637 = ~n26661 ;
  assign n26671 = n26258 & n44637 ;
  assign n26672 = n44171 & n26671 ;
  assign n27056 = n26672 & n134 ;
  assign n26673 = n26648 | n26661 ;
  assign n44638 = ~n26673 ;
  assign n27062 = n44638 & n134 ;
  assign n27063 = n26258 | n27062 ;
  assign n44639 = ~n27056 ;
  assign n27064 = n44639 & n27063 ;
  assign n27521 = n10657 | n27519 ;
  assign n44640 = ~n27521 ;
  assign n27540 = n44640 & n27537 ;
  assign n27541 = n27064 | n27540 ;
  assign n44641 = ~n27539 ;
  assign n27542 = n44641 & n27541 ;
  assign n44642 = ~n27542 ;
  assign n27543 = n157 & n44642 ;
  assign n26670 = n26664 | n26665 ;
  assign n44643 = ~n26670 ;
  assign n27051 = n44643 & n134 ;
  assign n27052 = n26255 | n27051 ;
  assign n26694 = n26255 & n44198 ;
  assign n44644 = ~n26665 ;
  assign n26695 = n44644 & n26694 ;
  assign n27138 = n26695 & n134 ;
  assign n44645 = ~n27138 ;
  assign n27139 = n27052 & n44645 ;
  assign n27551 = n44624 & n27532 ;
  assign n27552 = n27112 | n27551 ;
  assign n44646 = ~n27534 ;
  assign n27553 = n44646 & n27552 ;
  assign n44647 = ~n27553 ;
  assign n27554 = n155 & n44647 ;
  assign n27555 = n44634 & n27552 ;
  assign n27556 = n27129 | n27555 ;
  assign n44648 = ~n27554 ;
  assign n27557 = n44648 & n27556 ;
  assign n44649 = ~n27557 ;
  assign n27558 = n10657 & n44649 ;
  assign n27559 = n157 | n27558 ;
  assign n44650 = ~n27559 ;
  assign n27560 = n27541 & n44650 ;
  assign n27561 = n27139 | n27560 ;
  assign n44651 = ~n27543 ;
  assign n27562 = n44651 & n27561 ;
  assign n44652 = ~n27562 ;
  assign n27563 = n158 & n44652 ;
  assign n26693 = n26668 | n26681 ;
  assign n44653 = ~n26693 ;
  assign n27049 = n44653 & n134 ;
  assign n27050 = n26248 | n27049 ;
  assign n44654 = ~n26681 ;
  assign n26691 = n26248 & n44654 ;
  assign n26692 = n44187 & n26691 ;
  assign n27070 = n26692 & n134 ;
  assign n44655 = ~n27070 ;
  assign n27071 = n27050 & n44655 ;
  assign n27544 = n158 | n27543 ;
  assign n44656 = ~n27544 ;
  assign n27564 = n44656 & n27561 ;
  assign n27565 = n27071 | n27564 ;
  assign n44657 = ~n27563 ;
  assign n27566 = n44657 & n27565 ;
  assign n44658 = ~n27566 ;
  assign n27567 = n8857 & n44658 ;
  assign n26690 = n26684 | n26685 ;
  assign n44659 = ~n26690 ;
  assign n27058 = n44659 & n134 ;
  assign n27059 = n26354 | n27058 ;
  assign n26714 = n26354 & n44214 ;
  assign n44660 = ~n26685 ;
  assign n26715 = n44660 & n26714 ;
  assign n27099 = n26715 & n134 ;
  assign n44661 = ~n27099 ;
  assign n27100 = n27059 & n44661 ;
  assign n27575 = n44640 & n27556 ;
  assign n27576 = n27064 | n27575 ;
  assign n44662 = ~n27558 ;
  assign n27577 = n44662 & n27576 ;
  assign n44663 = ~n27577 ;
  assign n27578 = n157 & n44663 ;
  assign n27579 = n44650 & n27576 ;
  assign n27580 = n27139 | n27579 ;
  assign n44664 = ~n27578 ;
  assign n27581 = n44664 & n27580 ;
  assign n44665 = ~n27581 ;
  assign n27582 = n158 & n44665 ;
  assign n27583 = n8857 | n27582 ;
  assign n44666 = ~n27583 ;
  assign n27584 = n27565 & n44666 ;
  assign n27585 = n27100 | n27584 ;
  assign n44667 = ~n27567 ;
  assign n27586 = n44667 & n27585 ;
  assign n44668 = ~n27586 ;
  assign n27587 = n160 & n44668 ;
  assign n44669 = ~n26701 ;
  assign n26711 = n26349 & n44669 ;
  assign n26712 = n44203 & n26711 ;
  assign n27048 = n26712 & n134 ;
  assign n26713 = n26688 | n26701 ;
  assign n44670 = ~n26713 ;
  assign n27140 = n44670 & n134 ;
  assign n27141 = n26349 | n27140 ;
  assign n44671 = ~n27048 ;
  assign n27142 = n44671 & n27141 ;
  assign n27568 = n160 | n27567 ;
  assign n44672 = ~n27568 ;
  assign n27588 = n44672 & n27585 ;
  assign n27591 = n27142 | n27588 ;
  assign n44673 = ~n27587 ;
  assign n27592 = n44673 & n27591 ;
  assign n44674 = ~n27592 ;
  assign n27593 = n161 & n44674 ;
  assign n26710 = n26704 | n26705 ;
  assign n44675 = ~n26710 ;
  assign n27037 = n44675 & n134 ;
  assign n27038 = n26251 | n27037 ;
  assign n26734 = n26251 & n44230 ;
  assign n44676 = ~n26705 ;
  assign n26735 = n44676 & n26734 ;
  assign n27150 = n26735 & n134 ;
  assign n44677 = ~n27150 ;
  assign n27151 = n27038 & n44677 ;
  assign n27599 = n44656 & n27580 ;
  assign n27600 = n27071 | n27599 ;
  assign n44678 = ~n27582 ;
  assign n27601 = n44678 & n27600 ;
  assign n44679 = ~n27601 ;
  assign n27602 = n159 & n44679 ;
  assign n27603 = n44666 & n27600 ;
  assign n27604 = n27100 | n27603 ;
  assign n44680 = ~n27602 ;
  assign n27605 = n44680 & n27604 ;
  assign n44681 = ~n27605 ;
  assign n27606 = n8534 & n44681 ;
  assign n27607 = n161 | n27606 ;
  assign n44682 = ~n27607 ;
  assign n27608 = n27591 & n44682 ;
  assign n27609 = n27151 | n27608 ;
  assign n44683 = ~n27593 ;
  assign n27610 = n44683 & n27609 ;
  assign n44684 = ~n27610 ;
  assign n27611 = n162 & n44684 ;
  assign n26733 = n26708 | n26721 ;
  assign n44685 = ~n26733 ;
  assign n27043 = n44685 & n134 ;
  assign n27044 = n26361 | n27043 ;
  assign n44686 = ~n26721 ;
  assign n26731 = n26361 & n44686 ;
  assign n26732 = n44219 & n26731 ;
  assign n27105 = n26732 & n134 ;
  assign n44687 = ~n27105 ;
  assign n27106 = n27044 & n44687 ;
  assign n27594 = n162 | n27593 ;
  assign n44688 = ~n27594 ;
  assign n27612 = n44688 & n27609 ;
  assign n27613 = n27106 | n27612 ;
  assign n44689 = ~n27611 ;
  assign n27614 = n44689 & n27613 ;
  assign n44690 = ~n27614 ;
  assign n27615 = n6889 & n44690 ;
  assign n26754 = n26263 & n44246 ;
  assign n44691 = ~n26725 ;
  assign n26755 = n44691 & n26754 ;
  assign n27032 = n26755 & n134 ;
  assign n26726 = n26724 | n26725 ;
  assign n44692 = ~n26726 ;
  assign n27033 = n44692 & n134 ;
  assign n27034 = n26263 | n27033 ;
  assign n44693 = ~n27032 ;
  assign n27035 = n44693 & n27034 ;
  assign n27623 = n44672 & n27604 ;
  assign n27624 = n27142 | n27623 ;
  assign n44694 = ~n27606 ;
  assign n27625 = n44694 & n27624 ;
  assign n44695 = ~n27625 ;
  assign n27626 = n161 & n44695 ;
  assign n27627 = n44682 & n27624 ;
  assign n27628 = n27151 | n27627 ;
  assign n44696 = ~n27626 ;
  assign n27629 = n44696 & n27628 ;
  assign n44697 = ~n27629 ;
  assign n27630 = n162 & n44697 ;
  assign n27631 = n6889 | n27630 ;
  assign n44698 = ~n27631 ;
  assign n27632 = n27613 & n44698 ;
  assign n27633 = n27035 | n27632 ;
  assign n44699 = ~n27615 ;
  assign n27634 = n44699 & n27633 ;
  assign n44700 = ~n27634 ;
  assign n27635 = n164 & n44700 ;
  assign n26753 = n26729 | n26741 ;
  assign n44701 = ~n26753 ;
  assign n27041 = n44701 & n134 ;
  assign n27042 = n26235 | n27041 ;
  assign n44702 = ~n26741 ;
  assign n26751 = n26235 & n44702 ;
  assign n26752 = n44235 & n26751 ;
  assign n27148 = n26752 & n134 ;
  assign n44703 = ~n27148 ;
  assign n27149 = n27042 & n44703 ;
  assign n27616 = n6600 | n27615 ;
  assign n44704 = ~n27616 ;
  assign n27636 = n44704 & n27633 ;
  assign n27637 = n27149 | n27636 ;
  assign n44705 = ~n27635 ;
  assign n27638 = n44705 & n27637 ;
  assign n44706 = ~n27638 ;
  assign n27639 = n165 & n44706 ;
  assign n26774 = n26229 & n44262 ;
  assign n44707 = ~n26745 ;
  assign n26775 = n44707 & n26774 ;
  assign n27101 = n26775 & n134 ;
  assign n26750 = n26744 | n26745 ;
  assign n44708 = ~n26750 ;
  assign n27158 = n44708 & n134 ;
  assign n27159 = n26229 | n27158 ;
  assign n44709 = ~n27101 ;
  assign n27160 = n44709 & n27159 ;
  assign n27647 = n44688 & n27628 ;
  assign n27648 = n27106 | n27647 ;
  assign n44710 = ~n27630 ;
  assign n27649 = n44710 & n27648 ;
  assign n44711 = ~n27649 ;
  assign n27650 = n163 & n44711 ;
  assign n27651 = n44698 & n27648 ;
  assign n27652 = n27035 | n27651 ;
  assign n44712 = ~n27650 ;
  assign n27653 = n44712 & n27652 ;
  assign n44713 = ~n27653 ;
  assign n27654 = n6600 & n44713 ;
  assign n27655 = n165 | n27654 ;
  assign n44714 = ~n27655 ;
  assign n27656 = n27637 & n44714 ;
  assign n27657 = n27160 | n27656 ;
  assign n44715 = ~n27639 ;
  assign n27658 = n44715 & n27657 ;
  assign n44716 = ~n27658 ;
  assign n27659 = n166 & n44716 ;
  assign n26771 = n26748 | n26761 ;
  assign n44717 = ~n26771 ;
  assign n27161 = n44717 & n134 ;
  assign n27162 = n26373 | n27161 ;
  assign n44718 = ~n26761 ;
  assign n26772 = n26373 & n44718 ;
  assign n26773 = n44251 & n26772 ;
  assign n27164 = n26773 & n134 ;
  assign n44719 = ~n27164 ;
  assign n27165 = n27162 & n44719 ;
  assign n27640 = n166 | n27639 ;
  assign n44720 = ~n27640 ;
  assign n27660 = n44720 & n27657 ;
  assign n27663 = n27165 | n27660 ;
  assign n44721 = ~n27659 ;
  assign n27664 = n44721 & n27663 ;
  assign n44722 = ~n27664 ;
  assign n27665 = n5352 & n44722 ;
  assign n26794 = n26473 & n44278 ;
  assign n44723 = ~n26765 ;
  assign n26795 = n44723 & n26794 ;
  assign n27077 = n26795 & n134 ;
  assign n26770 = n26764 | n26765 ;
  assign n44724 = ~n26770 ;
  assign n27168 = n44724 & n134 ;
  assign n27169 = n26473 | n27168 ;
  assign n44725 = ~n27077 ;
  assign n27170 = n44725 & n27169 ;
  assign n27671 = n44704 & n27652 ;
  assign n27672 = n27149 | n27671 ;
  assign n44726 = ~n27654 ;
  assign n27673 = n44726 & n27672 ;
  assign n44727 = ~n27673 ;
  assign n27674 = n165 & n44727 ;
  assign n27675 = n44714 & n27672 ;
  assign n27676 = n27160 | n27675 ;
  assign n44728 = ~n27674 ;
  assign n27677 = n44728 & n27676 ;
  assign n44729 = ~n27677 ;
  assign n27678 = n166 & n44729 ;
  assign n27679 = n5352 | n27678 ;
  assign n44730 = ~n27679 ;
  assign n27680 = n27663 & n44730 ;
  assign n27681 = n27170 | n27680 ;
  assign n44731 = ~n27665 ;
  assign n27682 = n44731 & n27681 ;
  assign n44732 = ~n27682 ;
  assign n27683 = n168 & n44732 ;
  assign n26793 = n26768 | n26781 ;
  assign n44733 = ~n26793 ;
  assign n27171 = n44733 & n134 ;
  assign n27172 = n26379 | n27171 ;
  assign n44734 = ~n26781 ;
  assign n26791 = n26379 & n44734 ;
  assign n26792 = n44267 & n26791 ;
  assign n27173 = n26792 & n134 ;
  assign n44735 = ~n27173 ;
  assign n27174 = n27172 & n44735 ;
  assign n27666 = n4934 | n27665 ;
  assign n44736 = ~n27666 ;
  assign n27684 = n44736 & n27681 ;
  assign n27685 = n27174 | n27684 ;
  assign n44737 = ~n27683 ;
  assign n27686 = n44737 & n27685 ;
  assign n44738 = ~n27686 ;
  assign n27687 = n169 & n44738 ;
  assign n26814 = n26383 & n44294 ;
  assign n44739 = ~n26785 ;
  assign n26815 = n44739 & n26814 ;
  assign n27163 = n26815 & n134 ;
  assign n26790 = n26784 | n26785 ;
  assign n44740 = ~n26790 ;
  assign n27175 = n44740 & n134 ;
  assign n27176 = n26383 | n27175 ;
  assign n44741 = ~n27163 ;
  assign n27177 = n44741 & n27176 ;
  assign n27695 = n44720 & n27676 ;
  assign n27696 = n27165 | n27695 ;
  assign n44742 = ~n27678 ;
  assign n27697 = n44742 & n27696 ;
  assign n44743 = ~n27697 ;
  assign n27698 = n167 & n44743 ;
  assign n27699 = n44730 & n27696 ;
  assign n27700 = n27170 | n27699 ;
  assign n44744 = ~n27698 ;
  assign n27701 = n44744 & n27700 ;
  assign n44745 = ~n27701 ;
  assign n27702 = n4934 & n44745 ;
  assign n27703 = n169 | n27702 ;
  assign n44746 = ~n27703 ;
  assign n27704 = n27685 & n44746 ;
  assign n27705 = n27177 | n27704 ;
  assign n44747 = ~n27687 ;
  assign n27706 = n44747 & n27705 ;
  assign n44748 = ~n27706 ;
  assign n27707 = n170 & n44748 ;
  assign n26813 = n26788 | n26801 ;
  assign n44749 = ~n26813 ;
  assign n27095 = n44749 & n134 ;
  assign n27096 = n26386 | n27095 ;
  assign n44750 = ~n26801 ;
  assign n26811 = n26386 & n44750 ;
  assign n26812 = n44283 & n26811 ;
  assign n27179 = n26812 & n134 ;
  assign n44751 = ~n27179 ;
  assign n27180 = n27096 & n44751 ;
  assign n27689 = n170 | n27687 ;
  assign n44752 = ~n27689 ;
  assign n27708 = n44752 & n27705 ;
  assign n27709 = n27180 | n27708 ;
  assign n44753 = ~n27707 ;
  assign n27710 = n44753 & n27709 ;
  assign n44754 = ~n27710 ;
  assign n27711 = n3940 & n44754 ;
  assign n26834 = n26390 & n44310 ;
  assign n44755 = ~n26805 ;
  assign n26835 = n44755 & n26834 ;
  assign n27102 = n26835 & n134 ;
  assign n26810 = n26804 | n26805 ;
  assign n44756 = ~n26810 ;
  assign n27121 = n44756 & n134 ;
  assign n27122 = n26390 | n27121 ;
  assign n44757 = ~n27102 ;
  assign n27123 = n44757 & n27122 ;
  assign n27719 = n44736 & n27700 ;
  assign n27720 = n27174 | n27719 ;
  assign n44758 = ~n27702 ;
  assign n27721 = n44758 & n27720 ;
  assign n44759 = ~n27721 ;
  assign n27722 = n169 & n44759 ;
  assign n27723 = n44746 & n27720 ;
  assign n27724 = n27177 | n27723 ;
  assign n44760 = ~n27722 ;
  assign n27725 = n44760 & n27724 ;
  assign n44761 = ~n27725 ;
  assign n27726 = n170 & n44761 ;
  assign n27727 = n3940 | n27726 ;
  assign n44762 = ~n27727 ;
  assign n27728 = n27709 & n44762 ;
  assign n27729 = n27123 | n27728 ;
  assign n44763 = ~n27711 ;
  assign n27730 = n44763 & n27729 ;
  assign n44764 = ~n27730 ;
  assign n27731 = n172 & n44764 ;
  assign n26833 = n26808 | n26821 ;
  assign n44765 = ~n26833 ;
  assign n27181 = n44765 & n134 ;
  assign n27182 = n26469 | n27181 ;
  assign n44766 = ~n26821 ;
  assign n26831 = n26469 & n44766 ;
  assign n26832 = n44299 & n26831 ;
  assign n27185 = n26832 & n134 ;
  assign n44767 = ~n27185 ;
  assign n27186 = n27182 & n44767 ;
  assign n27712 = n3631 | n27711 ;
  assign n44768 = ~n27712 ;
  assign n27732 = n44768 & n27729 ;
  assign n27733 = n27186 | n27732 ;
  assign n44769 = ~n27731 ;
  assign n27734 = n44769 & n27733 ;
  assign n44770 = ~n27734 ;
  assign n27735 = n173 & n44770 ;
  assign n26830 = n26824 | n26825 ;
  assign n44771 = ~n26830 ;
  assign n27060 = n44771 & n134 ;
  assign n27061 = n26393 | n27060 ;
  assign n26854 = n26393 & n44326 ;
  assign n44772 = ~n26825 ;
  assign n26855 = n44772 & n26854 ;
  assign n27187 = n26855 & n134 ;
  assign n44773 = ~n27187 ;
  assign n27188 = n27061 & n44773 ;
  assign n27743 = n44752 & n27724 ;
  assign n27744 = n27180 | n27743 ;
  assign n44774 = ~n27726 ;
  assign n27745 = n44774 & n27744 ;
  assign n44775 = ~n27745 ;
  assign n27746 = n171 & n44775 ;
  assign n27747 = n44762 & n27744 ;
  assign n27748 = n27123 | n27747 ;
  assign n44776 = ~n27746 ;
  assign n27749 = n44776 & n27748 ;
  assign n44777 = ~n27749 ;
  assign n27750 = n3631 & n44777 ;
  assign n27751 = n173 | n27750 ;
  assign n44778 = ~n27751 ;
  assign n27752 = n27733 & n44778 ;
  assign n27753 = n27188 | n27752 ;
  assign n44779 = ~n27735 ;
  assign n27754 = n44779 & n27753 ;
  assign n44780 = ~n27754 ;
  assign n27755 = n174 & n44780 ;
  assign n26851 = n26828 | n26841 ;
  assign n44781 = ~n26851 ;
  assign n27189 = n44781 & n134 ;
  assign n27190 = n26398 | n27189 ;
  assign n44782 = ~n26841 ;
  assign n26852 = n26398 & n44782 ;
  assign n26853 = n44315 & n26852 ;
  assign n27193 = n26853 & n134 ;
  assign n44783 = ~n27193 ;
  assign n27194 = n27190 & n44783 ;
  assign n27736 = n174 | n27735 ;
  assign n44784 = ~n27736 ;
  assign n27756 = n44784 & n27753 ;
  assign n27757 = n27194 | n27756 ;
  assign n44785 = ~n27755 ;
  assign n27758 = n44785 & n27757 ;
  assign n44786 = ~n27758 ;
  assign n27759 = n2753 & n44786 ;
  assign n26874 = n26465 & n44342 ;
  assign n44787 = ~n26845 ;
  assign n26875 = n44787 & n26874 ;
  assign n27178 = n26875 & n134 ;
  assign n26850 = n26844 | n26845 ;
  assign n44788 = ~n26850 ;
  assign n27195 = n44788 & n134 ;
  assign n27196 = n26465 | n27195 ;
  assign n44789 = ~n27178 ;
  assign n27197 = n44789 & n27196 ;
  assign n27767 = n44768 & n27748 ;
  assign n27768 = n27186 | n27767 ;
  assign n44790 = ~n27750 ;
  assign n27769 = n44790 & n27768 ;
  assign n44791 = ~n27769 ;
  assign n27770 = n173 & n44791 ;
  assign n27771 = n44778 & n27768 ;
  assign n27772 = n27188 | n27771 ;
  assign n44792 = ~n27770 ;
  assign n27773 = n44792 & n27772 ;
  assign n44793 = ~n27773 ;
  assign n27774 = n174 & n44793 ;
  assign n27775 = n2753 | n27774 ;
  assign n44794 = ~n27775 ;
  assign n27776 = n27757 & n44794 ;
  assign n27777 = n27197 | n27776 ;
  assign n44795 = ~n27759 ;
  assign n27778 = n44795 & n27777 ;
  assign n44796 = ~n27778 ;
  assign n27779 = n176 & n44796 ;
  assign n44797 = ~n26861 ;
  assign n26871 = n26404 & n44797 ;
  assign n26872 = n44331 & n26871 ;
  assign n27057 = n26872 & n134 ;
  assign n26873 = n26848 | n26861 ;
  assign n44798 = ~n26873 ;
  assign n27089 = n44798 & n134 ;
  assign n27090 = n26404 | n27089 ;
  assign n44799 = ~n27057 ;
  assign n27091 = n44799 & n27090 ;
  assign n27760 = n2431 | n27759 ;
  assign n44800 = ~n27760 ;
  assign n27780 = n44800 & n27777 ;
  assign n27781 = n27091 | n27780 ;
  assign n44801 = ~n27779 ;
  assign n27782 = n44801 & n27781 ;
  assign n44802 = ~n27782 ;
  assign n27783 = n177 & n44802 ;
  assign n26866 = n26864 | n26865 ;
  assign n44803 = ~n26866 ;
  assign n27198 = n44803 & n134 ;
  assign n27199 = n26407 | n27198 ;
  assign n26894 = n26407 & n44358 ;
  assign n44804 = ~n26865 ;
  assign n26895 = n44804 & n26894 ;
  assign n27200 = n26895 & n134 ;
  assign n44805 = ~n27200 ;
  assign n27201 = n27199 & n44805 ;
  assign n27791 = n44784 & n27772 ;
  assign n27792 = n27194 | n27791 ;
  assign n44806 = ~n27774 ;
  assign n27793 = n44806 & n27792 ;
  assign n44807 = ~n27793 ;
  assign n27794 = n175 & n44807 ;
  assign n27795 = n44794 & n27792 ;
  assign n27796 = n27197 | n27795 ;
  assign n44808 = ~n27794 ;
  assign n27797 = n44808 & n27796 ;
  assign n44809 = ~n27797 ;
  assign n27798 = n2431 & n44809 ;
  assign n27799 = n177 | n27798 ;
  assign n44810 = ~n27799 ;
  assign n27800 = n27781 & n44810 ;
  assign n27801 = n27201 | n27800 ;
  assign n44811 = ~n27783 ;
  assign n27802 = n44811 & n27801 ;
  assign n44812 = ~n27802 ;
  assign n27803 = n178 & n44812 ;
  assign n44813 = ~n26881 ;
  assign n26891 = n26409 & n44813 ;
  assign n26892 = n44347 & n26891 ;
  assign n27065 = n26892 & n134 ;
  assign n26893 = n26869 | n26881 ;
  assign n44814 = ~n26893 ;
  assign n27202 = n44814 & n134 ;
  assign n27203 = n26409 | n27202 ;
  assign n44815 = ~n27065 ;
  assign n27204 = n44815 & n27203 ;
  assign n27784 = n178 | n27783 ;
  assign n44816 = ~n27784 ;
  assign n27804 = n44816 & n27801 ;
  assign n27805 = n27204 | n27804 ;
  assign n44817 = ~n27803 ;
  assign n27806 = n44817 & n27805 ;
  assign n44818 = ~n27806 ;
  assign n27807 = n1707 & n44818 ;
  assign n26886 = n26884 | n26885 ;
  assign n44819 = ~n26886 ;
  assign n27205 = n44819 & n134 ;
  assign n27206 = n26413 | n27205 ;
  assign n26914 = n26413 & n44374 ;
  assign n44820 = ~n26885 ;
  assign n26915 = n44820 & n26914 ;
  assign n27207 = n26915 & n134 ;
  assign n44821 = ~n27207 ;
  assign n27208 = n27206 & n44821 ;
  assign n27815 = n44800 & n27796 ;
  assign n27816 = n27091 | n27815 ;
  assign n44822 = ~n27798 ;
  assign n27817 = n44822 & n27816 ;
  assign n44823 = ~n27817 ;
  assign n27818 = n177 & n44823 ;
  assign n27819 = n44810 & n27816 ;
  assign n27820 = n27201 | n27819 ;
  assign n44824 = ~n27818 ;
  assign n27821 = n44824 & n27820 ;
  assign n44825 = ~n27821 ;
  assign n27822 = n178 & n44825 ;
  assign n27823 = n1707 | n27822 ;
  assign n44826 = ~n27823 ;
  assign n27824 = n27805 & n44826 ;
  assign n27825 = n27208 | n27824 ;
  assign n44827 = ~n27807 ;
  assign n27826 = n44827 & n27825 ;
  assign n44828 = ~n27826 ;
  assign n27827 = n180 & n44828 ;
  assign n26913 = n26889 | n26901 ;
  assign n44829 = ~n26913 ;
  assign n27039 = n44829 & n134 ;
  assign n27040 = n26286 | n27039 ;
  assign n44830 = ~n26901 ;
  assign n26911 = n26286 & n44830 ;
  assign n26912 = n44363 & n26911 ;
  assign n27124 = n26912 & n134 ;
  assign n44831 = ~n27124 ;
  assign n27125 = n27040 & n44831 ;
  assign n27808 = n1487 | n27807 ;
  assign n44832 = ~n27808 ;
  assign n27828 = n44832 & n27825 ;
  assign n27829 = n27125 | n27828 ;
  assign n44833 = ~n27827 ;
  assign n27830 = n44833 & n27829 ;
  assign n44834 = ~n27830 ;
  assign n27831 = n181 & n44834 ;
  assign n26910 = n26904 | n26905 ;
  assign n44835 = ~n26910 ;
  assign n27183 = n44835 & n134 ;
  assign n27184 = n26467 | n27183 ;
  assign n26934 = n26467 & n44390 ;
  assign n44836 = ~n26905 ;
  assign n26935 = n44836 & n26934 ;
  assign n27191 = n26935 & n134 ;
  assign n44837 = ~n27191 ;
  assign n27192 = n27184 & n44837 ;
  assign n27839 = n44816 & n27820 ;
  assign n27840 = n27204 | n27839 ;
  assign n44838 = ~n27822 ;
  assign n27841 = n44838 & n27840 ;
  assign n44839 = ~n27841 ;
  assign n27842 = n179 & n44839 ;
  assign n27843 = n44826 & n27840 ;
  assign n27844 = n27208 | n27843 ;
  assign n44840 = ~n27842 ;
  assign n27845 = n44840 & n27844 ;
  assign n44841 = ~n27845 ;
  assign n27846 = n1487 & n44841 ;
  assign n27847 = n181 | n27846 ;
  assign n44842 = ~n27847 ;
  assign n27848 = n27829 & n44842 ;
  assign n27849 = n27192 | n27848 ;
  assign n44843 = ~n27831 ;
  assign n27850 = n44843 & n27849 ;
  assign n44844 = ~n27850 ;
  assign n27851 = n182 & n44844 ;
  assign n26933 = n26908 | n26921 ;
  assign n44845 = ~n26933 ;
  assign n27084 = n44845 & n134 ;
  assign n27085 = n26417 | n27084 ;
  assign n44846 = ~n26921 ;
  assign n26931 = n26417 & n44846 ;
  assign n26932 = n44379 & n26931 ;
  assign n27152 = n26932 & n134 ;
  assign n44847 = ~n27152 ;
  assign n27153 = n27085 & n44847 ;
  assign n27832 = n182 | n27831 ;
  assign n44848 = ~n27832 ;
  assign n27852 = n44848 & n27849 ;
  assign n27855 = n27153 | n27852 ;
  assign n44849 = ~n27851 ;
  assign n27856 = n44849 & n27855 ;
  assign n44850 = ~n27856 ;
  assign n27857 = n996 & n44850 ;
  assign n26930 = n26924 | n26925 ;
  assign n44851 = ~n26930 ;
  assign n27209 = n44851 & n134 ;
  assign n27210 = n26419 | n27209 ;
  assign n26954 = n26419 & n44406 ;
  assign n44852 = ~n26925 ;
  assign n26955 = n44852 & n26954 ;
  assign n27211 = n26955 & n134 ;
  assign n44853 = ~n27211 ;
  assign n27212 = n27210 & n44853 ;
  assign n27863 = n44832 & n27844 ;
  assign n27864 = n27125 | n27863 ;
  assign n44854 = ~n27846 ;
  assign n27865 = n44854 & n27864 ;
  assign n44855 = ~n27865 ;
  assign n27866 = n181 & n44855 ;
  assign n27867 = n44842 & n27864 ;
  assign n27868 = n27192 | n27867 ;
  assign n44856 = ~n27866 ;
  assign n27869 = n44856 & n27868 ;
  assign n44857 = ~n27869 ;
  assign n27870 = n182 & n44857 ;
  assign n27871 = n183 | n27870 ;
  assign n44858 = ~n27871 ;
  assign n27872 = n27855 & n44858 ;
  assign n27873 = n27212 | n27872 ;
  assign n44859 = ~n27857 ;
  assign n27874 = n44859 & n27873 ;
  assign n44860 = ~n27874 ;
  assign n27875 = n184 & n44860 ;
  assign n26953 = n26928 | n26941 ;
  assign n44861 = ~n26953 ;
  assign n27097 = n44861 & n134 ;
  assign n27098 = n26396 | n27097 ;
  assign n44862 = ~n26941 ;
  assign n26951 = n26396 & n44862 ;
  assign n26952 = n44395 & n26951 ;
  assign n27213 = n26952 & n134 ;
  assign n44863 = ~n27213 ;
  assign n27214 = n27098 & n44863 ;
  assign n27858 = n838 | n27857 ;
  assign n44864 = ~n27858 ;
  assign n27876 = n44864 & n27873 ;
  assign n27877 = n27214 | n27876 ;
  assign n44865 = ~n27875 ;
  assign n27878 = n44865 & n27877 ;
  assign n44866 = ~n27878 ;
  assign n27879 = n185 & n44866 ;
  assign n26950 = n26944 | n26945 ;
  assign n44867 = ~n26950 ;
  assign n27215 = n44867 & n134 ;
  assign n27216 = n26423 | n27215 ;
  assign n26974 = n26423 & n44422 ;
  assign n44868 = ~n26945 ;
  assign n26975 = n44868 & n26974 ;
  assign n27217 = n26975 & n134 ;
  assign n44869 = ~n27217 ;
  assign n27218 = n27216 & n44869 ;
  assign n27887 = n44848 & n27868 ;
  assign n27888 = n27153 | n27887 ;
  assign n44870 = ~n27870 ;
  assign n27889 = n44870 & n27888 ;
  assign n44871 = ~n27889 ;
  assign n27890 = n183 & n44871 ;
  assign n27891 = n44858 & n27888 ;
  assign n27892 = n27212 | n27891 ;
  assign n44872 = ~n27890 ;
  assign n27893 = n44872 & n27892 ;
  assign n44873 = ~n27893 ;
  assign n27894 = n838 & n44873 ;
  assign n27895 = n185 | n27894 ;
  assign n44874 = ~n27895 ;
  assign n27896 = n27877 & n44874 ;
  assign n27897 = n27218 | n27896 ;
  assign n44875 = ~n27879 ;
  assign n27898 = n44875 & n27897 ;
  assign n44876 = ~n27898 ;
  assign n27899 = n186 & n44876 ;
  assign n26973 = n26948 | n26961 ;
  assign n44877 = ~n26973 ;
  assign n27107 = n44877 & n134 ;
  assign n27108 = n26425 | n27107 ;
  assign n44878 = ~n26961 ;
  assign n26971 = n26425 & n44878 ;
  assign n26972 = n44411 & n26971 ;
  assign n27219 = n26972 & n134 ;
  assign n44879 = ~n27219 ;
  assign n27220 = n27108 & n44879 ;
  assign n27880 = n186 | n27879 ;
  assign n44880 = ~n27880 ;
  assign n27900 = n44880 & n27897 ;
  assign n27903 = n27220 | n27900 ;
  assign n44881 = ~n27899 ;
  assign n27904 = n44881 & n27903 ;
  assign n44882 = ~n27904 ;
  assign n27905 = n528 & n44882 ;
  assign n26994 = n26427 & n44431 ;
  assign n44883 = ~n26965 ;
  assign n26995 = n44883 & n26994 ;
  assign n27036 = n26995 & n134 ;
  assign n26970 = n26964 | n26965 ;
  assign n44884 = ~n26970 ;
  assign n27134 = n44884 & n134 ;
  assign n27135 = n26427 | n27134 ;
  assign n44885 = ~n27036 ;
  assign n27136 = n44885 & n27135 ;
  assign n27911 = n44864 & n27892 ;
  assign n27912 = n27214 | n27911 ;
  assign n44886 = ~n27894 ;
  assign n27913 = n44886 & n27912 ;
  assign n44887 = ~n27913 ;
  assign n27914 = n185 & n44887 ;
  assign n27915 = n44874 & n27912 ;
  assign n27916 = n27218 | n27915 ;
  assign n44888 = ~n27914 ;
  assign n27917 = n44888 & n27916 ;
  assign n44889 = ~n27917 ;
  assign n27918 = n186 & n44889 ;
  assign n27919 = n528 | n27918 ;
  assign n44890 = ~n27919 ;
  assign n27920 = n27903 & n44890 ;
  assign n27921 = n27136 | n27920 ;
  assign n44891 = ~n27905 ;
  assign n27922 = n44891 & n27921 ;
  assign n44892 = ~n27922 ;
  assign n27923 = n188 & n44892 ;
  assign n26991 = n26968 | n26981 ;
  assign n44893 = ~n26991 ;
  assign n27221 = n44893 & n134 ;
  assign n27222 = n26430 | n27221 ;
  assign n44894 = ~n26981 ;
  assign n26992 = n26430 & n44894 ;
  assign n26993 = n44443 & n26992 ;
  assign n27223 = n26993 & n134 ;
  assign n44895 = ~n27223 ;
  assign n27224 = n27222 & n44895 ;
  assign n27906 = n413 | n27905 ;
  assign n44896 = ~n27906 ;
  assign n27924 = n44896 & n27921 ;
  assign n27925 = n27224 | n27924 ;
  assign n44897 = ~n27923 ;
  assign n27926 = n44897 & n27925 ;
  assign n44898 = ~n27926 ;
  assign n27927 = n189 & n44898 ;
  assign n44899 = ~n27927 ;
  assign n27929 = n27227 & n44899 ;
  assign n27935 = n44880 & n27916 ;
  assign n27936 = n27220 | n27935 ;
  assign n44900 = ~n27918 ;
  assign n27937 = n44900 & n27936 ;
  assign n44901 = ~n27937 ;
  assign n27938 = n187 & n44901 ;
  assign n27939 = n44890 & n27936 ;
  assign n27940 = n27136 | n27939 ;
  assign n44902 = ~n27938 ;
  assign n27941 = n44902 & n27940 ;
  assign n44903 = ~n27941 ;
  assign n27942 = n413 & n44903 ;
  assign n27943 = n189 | n27942 ;
  assign n44904 = ~n27943 ;
  assign n27944 = n27925 & n44904 ;
  assign n44905 = ~n27944 ;
  assign n27956 = n27929 & n44905 ;
  assign n44906 = ~n26476 ;
  assign n27240 = n44906 & n134 ;
  assign n44907 = ~n27240 ;
  assign n27241 = n27028 & n44907 ;
  assign n27248 = n26476 | n27028 ;
  assign n27250 = n192 & n27248 ;
  assign n44908 = ~n27241 ;
  assign n27251 = n44908 & n27250 ;
  assign n27027 = n27008 | n27021 ;
  assign n44909 = ~n27027 ;
  assign n27231 = n44909 & n134 ;
  assign n27232 = n26440 | n27231 ;
  assign n44910 = ~n27021 ;
  assign n27025 = n26440 & n44910 ;
  assign n27026 = n44459 & n27025 ;
  assign n27236 = n27026 & n134 ;
  assign n44911 = ~n27236 ;
  assign n27237 = n27232 & n44911 ;
  assign n27945 = n27227 | n27944 ;
  assign n27946 = n44899 & n27945 ;
  assign n44912 = ~n27946 ;
  assign n27947 = n190 & n44912 ;
  assign n44913 = ~n27001 ;
  assign n27011 = n26434 & n44913 ;
  assign n27012 = n44451 & n27011 ;
  assign n27116 = n27012 & n134 ;
  assign n27013 = n26988 | n27001 ;
  assign n44914 = ~n27013 ;
  assign n27228 = n44914 & n134 ;
  assign n27229 = n26434 | n27228 ;
  assign n44915 = ~n27116 ;
  assign n27230 = n44915 & n27229 ;
  assign n27928 = n190 | n27927 ;
  assign n44916 = ~n27928 ;
  assign n27948 = n44916 & n27945 ;
  assign n27949 = n27230 | n27948 ;
  assign n44917 = ~n27947 ;
  assign n27950 = n44917 & n27949 ;
  assign n44918 = ~n27950 ;
  assign n27951 = n287 & n44918 ;
  assign n44919 = ~n27951 ;
  assign n27952 = n27237 & n44919 ;
  assign n27010 = n27004 | n27005 ;
  assign n44920 = ~n27010 ;
  assign n27166 = n44920 & n134 ;
  assign n27167 = n26437 | n27166 ;
  assign n44921 = ~n27019 ;
  assign n27265 = n26437 & n44921 ;
  assign n44922 = ~n27005 ;
  assign n27266 = n44922 & n27265 ;
  assign n27267 = n134 & n27266 ;
  assign n44923 = ~n27267 ;
  assign n27268 = n27167 & n44923 ;
  assign n27959 = n44896 & n27940 ;
  assign n27960 = n27224 | n27959 ;
  assign n44924 = ~n27942 ;
  assign n27961 = n44924 & n27960 ;
  assign n44925 = ~n27961 ;
  assign n27962 = n189 & n44925 ;
  assign n27963 = n44904 & n27960 ;
  assign n27964 = n27227 | n27963 ;
  assign n44926 = ~n27962 ;
  assign n27965 = n44926 & n27964 ;
  assign n44927 = ~n27965 ;
  assign n27966 = n190 & n44927 ;
  assign n27967 = n287 | n27966 ;
  assign n44928 = ~n27967 ;
  assign n27968 = n27949 & n44928 ;
  assign n27969 = n27268 | n27968 ;
  assign n27970 = n27952 & n27969 ;
  assign n27971 = n27251 | n27970 ;
  assign n44929 = ~n27248 ;
  assign n27249 = n134 & n44929 ;
  assign n27261 = n27023 | n27249 ;
  assign n27262 = n27237 | n27261 ;
  assign n27974 = n44919 & n27969 ;
  assign n27975 = n27262 | n27974 ;
  assign n27976 = n31336 & n27975 ;
  assign n133 = n27971 | n27976 ;
  assign n28104 = n27956 & n133 ;
  assign n27957 = n27927 | n27944 ;
  assign n44930 = ~n27957 ;
  assign n28150 = n44930 & n133 ;
  assign n28151 = n27227 | n28150 ;
  assign n44931 = ~n28104 ;
  assign n28152 = n44931 & n28151 ;
  assign n260 = x6 | x7 ;
  assign n261 = x8 | n260 ;
  assign n28061 = x8 & n133 ;
  assign n44932 = ~n28061 ;
  assign n28072 = n261 & n44932 ;
  assign n44933 = ~n28072 ;
  assign n28073 = n134 & n44933 ;
  assign n26447 = n261 & n44477 ;
  assign n27263 = n26447 & n44478 ;
  assign n27264 = n44479 & n27263 ;
  assign n28062 = n27264 & n44932 ;
  assign n44934 = ~n257 ;
  assign n28068 = n44934 & n133 ;
  assign n44935 = ~x8 ;
  assign n28200 = n44935 & n133 ;
  assign n44936 = ~n28200 ;
  assign n28201 = x9 & n44936 ;
  assign n28202 = n28068 | n28201 ;
  assign n28212 = n28062 | n28202 ;
  assign n44937 = ~n28073 ;
  assign n28213 = n44937 & n28212 ;
  assign n44938 = ~n28213 ;
  assign n28214 = n26442 & n44938 ;
  assign n262 = n44935 & n260 ;
  assign n44939 = ~n133 ;
  assign n28217 = x8 & n44939 ;
  assign n28218 = n262 | n28217 ;
  assign n44940 = ~n28218 ;
  assign n28219 = n134 & n44940 ;
  assign n28220 = n26442 | n28219 ;
  assign n44941 = ~n28220 ;
  assign n28221 = n28212 & n44941 ;
  assign n44942 = ~n27251 ;
  assign n27253 = n134 & n44942 ;
  assign n44943 = ~n27970 ;
  assign n28230 = n27253 & n44943 ;
  assign n44944 = ~n27976 ;
  assign n28231 = n44944 & n28230 ;
  assign n28232 = n28068 | n28231 ;
  assign n28233 = x10 & n28232 ;
  assign n28234 = x10 | n28231 ;
  assign n28235 = n28068 | n28234 ;
  assign n44945 = ~n28233 ;
  assign n28236 = n44945 & n28235 ;
  assign n28237 = n28221 | n28236 ;
  assign n44946 = ~n28214 ;
  assign n28238 = n44946 & n28237 ;
  assign n44947 = ~n28238 ;
  assign n28239 = n25517 & n44947 ;
  assign n28215 = n25517 | n28214 ;
  assign n44948 = ~n28215 ;
  assign n28241 = n44948 & n28237 ;
  assign n28257 = n27246 | n27306 ;
  assign n44949 = ~n28257 ;
  assign n28258 = n27235 & n44949 ;
  assign n28259 = n133 & n28258 ;
  assign n28260 = n133 & n44949 ;
  assign n28261 = n27235 | n28260 ;
  assign n44950 = ~n28259 ;
  assign n28262 = n44950 & n28261 ;
  assign n28265 = n28241 | n28262 ;
  assign n44951 = ~n28239 ;
  assign n28266 = n44951 & n28265 ;
  assign n44952 = ~n28266 ;
  assign n28267 = n137 & n44952 ;
  assign n27334 = n27311 | n27312 ;
  assign n44953 = ~n27334 ;
  assign n28063 = n44953 & n133 ;
  assign n28064 = n27260 | n28063 ;
  assign n44954 = ~n27312 ;
  assign n27332 = n27260 & n44954 ;
  assign n27333 = n44484 & n27332 ;
  assign n28210 = n27333 & n133 ;
  assign n44955 = ~n28210 ;
  assign n28211 = n28064 & n44955 ;
  assign n28240 = n137 | n28239 ;
  assign n44956 = ~n28240 ;
  assign n28268 = n44956 & n28265 ;
  assign n28269 = n28211 | n28268 ;
  assign n44957 = ~n28267 ;
  assign n28270 = n44957 & n28269 ;
  assign n44958 = ~n28270 ;
  assign n28271 = n138 & n44958 ;
  assign n27331 = n27315 | n27318 ;
  assign n44959 = ~n27331 ;
  assign n28058 = n44959 & n133 ;
  assign n28059 = n27239 | n28058 ;
  assign n27317 = n27239 & n44489 ;
  assign n44960 = ~n27318 ;
  assign n27330 = n27317 & n44960 ;
  assign n28208 = n27330 & n133 ;
  assign n44961 = ~n28208 ;
  assign n28209 = n28059 & n44961 ;
  assign n28216 = n135 & n44938 ;
  assign n28074 = n135 | n28073 ;
  assign n44962 = ~n28074 ;
  assign n28223 = n44962 & n28212 ;
  assign n28245 = n28223 | n28236 ;
  assign n44963 = ~n28216 ;
  assign n28246 = n44963 & n28245 ;
  assign n44964 = ~n28246 ;
  assign n28247 = n136 & n44964 ;
  assign n28248 = n44948 & n28245 ;
  assign n28275 = n28248 | n28262 ;
  assign n44965 = ~n28247 ;
  assign n28276 = n44965 & n28275 ;
  assign n44966 = ~n28276 ;
  assign n28277 = n137 & n44966 ;
  assign n28278 = n138 | n28277 ;
  assign n44967 = ~n28278 ;
  assign n28279 = n28269 & n44967 ;
  assign n28280 = n28209 | n28279 ;
  assign n44968 = ~n28271 ;
  assign n28281 = n44968 & n28280 ;
  assign n44969 = ~n28281 ;
  assign n28282 = n139 & n44969 ;
  assign n44970 = ~n27322 ;
  assign n27328 = n27104 & n44970 ;
  assign n27329 = n44496 & n27328 ;
  assign n28053 = n27329 & n133 ;
  assign n27358 = n27322 | n27342 ;
  assign n44971 = ~n27358 ;
  assign n28081 = n44971 & n133 ;
  assign n28082 = n27104 | n28081 ;
  assign n44972 = ~n28053 ;
  assign n28083 = n44972 & n28082 ;
  assign n28272 = n139 | n28271 ;
  assign n44973 = ~n28272 ;
  assign n28283 = n44973 & n28280 ;
  assign n28284 = n28083 | n28283 ;
  assign n44974 = ~n28282 ;
  assign n28285 = n44974 & n28284 ;
  assign n44975 = ~n28285 ;
  assign n28286 = n22030 & n44975 ;
  assign n27357 = n27325 | n27344 ;
  assign n44976 = ~n27357 ;
  assign n28049 = n44976 & n133 ;
  assign n28050 = n27243 | n28049 ;
  assign n27326 = n27243 & n44507 ;
  assign n44977 = ~n27344 ;
  assign n27356 = n27326 & n44977 ;
  assign n28051 = n27356 & n133 ;
  assign n44978 = ~n28051 ;
  assign n28052 = n28050 & n44978 ;
  assign n28296 = n44956 & n28275 ;
  assign n28297 = n28211 | n28296 ;
  assign n44979 = ~n28277 ;
  assign n28298 = n44979 & n28297 ;
  assign n44980 = ~n28298 ;
  assign n28299 = n138 & n44980 ;
  assign n28300 = n44967 & n28297 ;
  assign n28301 = n28209 | n28300 ;
  assign n44981 = ~n28299 ;
  assign n28302 = n44981 & n28301 ;
  assign n44982 = ~n28302 ;
  assign n28303 = n22661 & n44982 ;
  assign n28304 = n140 | n28303 ;
  assign n44983 = ~n28304 ;
  assign n28305 = n28284 & n44983 ;
  assign n28306 = n28052 | n28305 ;
  assign n44984 = ~n28286 ;
  assign n28307 = n44984 & n28306 ;
  assign n44985 = ~n28307 ;
  assign n28308 = n141 & n44985 ;
  assign n27382 = n27348 | n27366 ;
  assign n44986 = ~n27382 ;
  assign n27985 = n44986 & n133 ;
  assign n27986 = n27301 | n27985 ;
  assign n44987 = ~n27348 ;
  assign n27354 = n27301 & n44987 ;
  assign n27355 = n44513 & n27354 ;
  assign n28030 = n27355 & n133 ;
  assign n44988 = ~n28030 ;
  assign n28031 = n27986 & n44988 ;
  assign n28287 = n141 | n28286 ;
  assign n44989 = ~n28287 ;
  assign n28309 = n44989 & n28306 ;
  assign n28310 = n28031 | n28309 ;
  assign n44990 = ~n28308 ;
  assign n28311 = n44990 & n28310 ;
  assign n44991 = ~n28311 ;
  assign n28312 = n142 & n44991 ;
  assign n27381 = n27351 | n27368 ;
  assign n44992 = ~n27381 ;
  assign n28084 = n44992 & n133 ;
  assign n28085 = n27093 | n28084 ;
  assign n27353 = n27093 & n44523 ;
  assign n44993 = ~n27368 ;
  assign n27380 = n27353 & n44993 ;
  assign n28089 = n27380 & n133 ;
  assign n44994 = ~n28089 ;
  assign n28090 = n28085 & n44994 ;
  assign n28320 = n44973 & n28301 ;
  assign n28321 = n28083 | n28320 ;
  assign n44995 = ~n28303 ;
  assign n28322 = n44995 & n28321 ;
  assign n44996 = ~n28322 ;
  assign n28323 = n140 & n44996 ;
  assign n28324 = n44983 & n28321 ;
  assign n28325 = n28052 | n28324 ;
  assign n44997 = ~n28323 ;
  assign n28326 = n44997 & n28325 ;
  assign n44998 = ~n28326 ;
  assign n28327 = n141 & n44998 ;
  assign n28328 = n142 | n28327 ;
  assign n44999 = ~n28328 ;
  assign n28329 = n28310 & n44999 ;
  assign n28330 = n28090 | n28329 ;
  assign n45000 = ~n28312 ;
  assign n28331 = n45000 & n28330 ;
  assign n45001 = ~n28331 ;
  assign n28332 = n143 & n45001 ;
  assign n27406 = n27372 | n27390 ;
  assign n45002 = ~n27406 ;
  assign n27981 = n45002 & n133 ;
  assign n27982 = n27294 | n27981 ;
  assign n45003 = ~n27372 ;
  assign n27378 = n27294 & n45003 ;
  assign n27379 = n44529 & n27378 ;
  assign n28116 = n27379 & n133 ;
  assign n45004 = ~n28116 ;
  assign n28117 = n27982 & n45004 ;
  assign n28313 = n143 | n28312 ;
  assign n45005 = ~n28313 ;
  assign n28333 = n45005 & n28330 ;
  assign n28334 = n28117 | n28333 ;
  assign n45006 = ~n28332 ;
  assign n28335 = n45006 & n28334 ;
  assign n45007 = ~n28335 ;
  assign n28336 = n18797 & n45007 ;
  assign n27404 = n27375 | n27392 ;
  assign n45008 = ~n27404 ;
  assign n28012 = n45008 & n133 ;
  assign n28013 = n27115 | n28012 ;
  assign n27377 = n27115 & n44539 ;
  assign n45009 = ~n27392 ;
  assign n27405 = n27377 & n45009 ;
  assign n28099 = n27405 & n133 ;
  assign n45010 = ~n28099 ;
  assign n28100 = n28013 & n45010 ;
  assign n28344 = n44989 & n28325 ;
  assign n28345 = n28031 | n28344 ;
  assign n45011 = ~n28327 ;
  assign n28346 = n45011 & n28345 ;
  assign n45012 = ~n28346 ;
  assign n28347 = n142 & n45012 ;
  assign n28348 = n44999 & n28345 ;
  assign n28349 = n28090 | n28348 ;
  assign n45013 = ~n28347 ;
  assign n28350 = n45013 & n28349 ;
  assign n45014 = ~n28350 ;
  assign n28351 = n19362 & n45014 ;
  assign n28352 = n144 | n28351 ;
  assign n45015 = ~n28352 ;
  assign n28353 = n28334 & n45015 ;
  assign n28354 = n28100 | n28353 ;
  assign n45016 = ~n28336 ;
  assign n28355 = n45016 & n28354 ;
  assign n45017 = ~n28355 ;
  assign n28356 = n145 & n45017 ;
  assign n45018 = ~n27396 ;
  assign n27402 = n27287 & n45018 ;
  assign n27403 = n44545 & n27402 ;
  assign n27996 = n27403 & n133 ;
  assign n27430 = n27396 | n27414 ;
  assign n45019 = ~n27430 ;
  assign n28076 = n45019 & n133 ;
  assign n28077 = n27287 | n28076 ;
  assign n45020 = ~n27996 ;
  assign n28078 = n45020 & n28077 ;
  assign n28337 = n145 | n28336 ;
  assign n45021 = ~n28337 ;
  assign n28357 = n45021 & n28354 ;
  assign n28358 = n28078 | n28357 ;
  assign n45022 = ~n28356 ;
  assign n28359 = n45022 & n28358 ;
  assign n45023 = ~n28359 ;
  assign n28360 = n146 & n45023 ;
  assign n27429 = n27399 | n27416 ;
  assign n45024 = ~n27429 ;
  assign n27987 = n45024 & n133 ;
  assign n27988 = n27280 | n27987 ;
  assign n27401 = n27280 & n44555 ;
  assign n45025 = ~n27416 ;
  assign n27428 = n27401 & n45025 ;
  assign n28106 = n27428 & n133 ;
  assign n45026 = ~n28106 ;
  assign n28107 = n27988 & n45026 ;
  assign n28368 = n45005 & n28349 ;
  assign n28369 = n28117 | n28368 ;
  assign n45027 = ~n28351 ;
  assign n28370 = n45027 & n28369 ;
  assign n45028 = ~n28370 ;
  assign n28371 = n144 & n45028 ;
  assign n28372 = n45015 & n28369 ;
  assign n28373 = n28100 | n28372 ;
  assign n45029 = ~n28371 ;
  assign n28374 = n45029 & n28373 ;
  assign n45030 = ~n28374 ;
  assign n28375 = n145 & n45030 ;
  assign n28376 = n146 | n28375 ;
  assign n45031 = ~n28376 ;
  assign n28377 = n28358 & n45031 ;
  assign n28378 = n28107 | n28377 ;
  assign n45032 = ~n28360 ;
  assign n28379 = n45032 & n28378 ;
  assign n45033 = ~n28379 ;
  assign n28380 = n147 & n45033 ;
  assign n27454 = n27420 | n27438 ;
  assign n45034 = ~n27454 ;
  assign n28112 = n45034 & n133 ;
  assign n28113 = n27274 | n28112 ;
  assign n45035 = ~n27420 ;
  assign n27426 = n27274 & n45035 ;
  assign n27427 = n44561 & n27426 ;
  assign n28114 = n27427 & n133 ;
  assign n45036 = ~n28114 ;
  assign n28115 = n28113 & n45036 ;
  assign n28361 = n147 | n28360 ;
  assign n45037 = ~n28361 ;
  assign n28381 = n45037 & n28378 ;
  assign n28382 = n28115 | n28381 ;
  assign n45038 = ~n28380 ;
  assign n28383 = n45038 & n28382 ;
  assign n45039 = ~n28383 ;
  assign n28384 = n15807 & n45039 ;
  assign n27424 = n27145 & n44571 ;
  assign n45040 = ~n27440 ;
  assign n27452 = n27424 & n45040 ;
  assign n28105 = n27452 & n133 ;
  assign n27453 = n27423 | n27440 ;
  assign n45041 = ~n27453 ;
  assign n28118 = n45041 & n133 ;
  assign n28119 = n27145 | n28118 ;
  assign n45042 = ~n28105 ;
  assign n28120 = n45042 & n28119 ;
  assign n28392 = n45021 & n28373 ;
  assign n28393 = n28078 | n28392 ;
  assign n45043 = ~n28375 ;
  assign n28394 = n45043 & n28393 ;
  assign n45044 = ~n28394 ;
  assign n28395 = n146 & n45044 ;
  assign n28396 = n45031 & n28393 ;
  assign n28397 = n28107 | n28396 ;
  assign n45045 = ~n28395 ;
  assign n28398 = n45045 & n28397 ;
  assign n45046 = ~n28398 ;
  assign n28399 = n16322 & n45046 ;
  assign n28400 = n148 | n28399 ;
  assign n45047 = ~n28400 ;
  assign n28401 = n28382 & n45047 ;
  assign n28402 = n28120 | n28401 ;
  assign n45048 = ~n28384 ;
  assign n28403 = n45048 & n28402 ;
  assign n45049 = ~n28403 ;
  assign n28404 = n149 & n45049 ;
  assign n45050 = ~n27444 ;
  assign n27450 = n27155 & n45050 ;
  assign n27451 = n44577 & n27450 ;
  assign n28035 = n27451 & n133 ;
  assign n27478 = n27444 | n27462 ;
  assign n45051 = ~n27478 ;
  assign n28069 = n45051 & n133 ;
  assign n28070 = n27155 | n28069 ;
  assign n45052 = ~n28035 ;
  assign n28071 = n45052 & n28070 ;
  assign n28385 = n149 | n28384 ;
  assign n45053 = ~n28385 ;
  assign n28405 = n45053 & n28402 ;
  assign n28406 = n28071 | n28405 ;
  assign n45054 = ~n28404 ;
  assign n28407 = n45054 & n28406 ;
  assign n45055 = ~n28407 ;
  assign n28408 = n150 & n45055 ;
  assign n27449 = n27157 & n44587 ;
  assign n45056 = ~n27464 ;
  assign n27476 = n27449 & n45056 ;
  assign n28060 = n27476 & n133 ;
  assign n27477 = n27447 | n27464 ;
  assign n45057 = ~n27477 ;
  assign n28121 = n45057 & n133 ;
  assign n28122 = n27157 | n28121 ;
  assign n45058 = ~n28060 ;
  assign n28123 = n45058 & n28122 ;
  assign n28416 = n45037 & n28397 ;
  assign n28417 = n28115 | n28416 ;
  assign n45059 = ~n28399 ;
  assign n28418 = n45059 & n28417 ;
  assign n45060 = ~n28418 ;
  assign n28419 = n148 & n45060 ;
  assign n28420 = n45047 & n28417 ;
  assign n28421 = n28120 | n28420 ;
  assign n45061 = ~n28419 ;
  assign n28422 = n45061 & n28421 ;
  assign n45062 = ~n28422 ;
  assign n28423 = n149 & n45062 ;
  assign n28424 = n150 | n28423 ;
  assign n45063 = ~n28424 ;
  assign n28425 = n28406 & n45063 ;
  assign n28426 = n28123 | n28425 ;
  assign n45064 = ~n28408 ;
  assign n28427 = n45064 & n28426 ;
  assign n45065 = ~n28427 ;
  assign n28428 = n151 & n45065 ;
  assign n27502 = n27468 | n27486 ;
  assign n45066 = ~n27502 ;
  assign n28028 = n45066 & n133 ;
  assign n28029 = n27088 | n28028 ;
  assign n45067 = ~n27468 ;
  assign n27474 = n27088 & n45067 ;
  assign n27475 = n44593 & n27474 ;
  assign n28065 = n27475 & n133 ;
  assign n45068 = ~n28065 ;
  assign n28066 = n28029 & n45068 ;
  assign n28410 = n151 | n28408 ;
  assign n45069 = ~n28410 ;
  assign n28429 = n45069 & n28426 ;
  assign n28430 = n28066 | n28429 ;
  assign n45070 = ~n28428 ;
  assign n28431 = n45070 & n28430 ;
  assign n45071 = ~n28431 ;
  assign n28432 = n13079 & n45071 ;
  assign n27473 = n27082 & n44603 ;
  assign n45072 = ~n27488 ;
  assign n27501 = n27473 & n45072 ;
  assign n28020 = n27501 & n133 ;
  assign n27500 = n27471 | n27488 ;
  assign n45073 = ~n27500 ;
  assign n28021 = n45073 & n133 ;
  assign n28022 = n27082 | n28021 ;
  assign n45074 = ~n28020 ;
  assign n28023 = n45074 & n28022 ;
  assign n28440 = n45053 & n28421 ;
  assign n28441 = n28071 | n28440 ;
  assign n45075 = ~n28423 ;
  assign n28442 = n45075 & n28441 ;
  assign n45076 = ~n28442 ;
  assign n28443 = n150 & n45076 ;
  assign n28444 = n45063 & n28441 ;
  assign n28445 = n28123 | n28444 ;
  assign n45077 = ~n28443 ;
  assign n28446 = n45077 & n28445 ;
  assign n45078 = ~n28446 ;
  assign n28447 = n13662 & n45078 ;
  assign n28448 = n152 | n28447 ;
  assign n45079 = ~n28448 ;
  assign n28449 = n28430 & n45079 ;
  assign n28450 = n28023 | n28449 ;
  assign n45080 = ~n28432 ;
  assign n28451 = n45080 & n28450 ;
  assign n45081 = ~n28451 ;
  assign n28452 = n153 & n45081 ;
  assign n45082 = ~n27492 ;
  assign n27498 = n27080 & n45082 ;
  assign n27499 = n44609 & n27498 ;
  assign n28019 = n27499 & n133 ;
  assign n27526 = n27492 | n27510 ;
  assign n45083 = ~n27526 ;
  assign n28044 = n45083 & n133 ;
  assign n28045 = n27080 | n28044 ;
  assign n45084 = ~n28019 ;
  assign n28046 = n45084 & n28045 ;
  assign n28433 = n153 | n28432 ;
  assign n45085 = ~n28433 ;
  assign n28453 = n45085 & n28450 ;
  assign n28454 = n28046 | n28453 ;
  assign n45086 = ~n28452 ;
  assign n28455 = n45086 & n28454 ;
  assign n45087 = ~n28455 ;
  assign n28456 = n154 & n45087 ;
  assign n27497 = n27075 & n44619 ;
  assign n45088 = ~n27512 ;
  assign n27524 = n27497 & n45088 ;
  assign n28018 = n27524 & n133 ;
  assign n27525 = n27495 | n27512 ;
  assign n45089 = ~n27525 ;
  assign n28024 = n45089 & n133 ;
  assign n28025 = n27075 | n28024 ;
  assign n45090 = ~n28018 ;
  assign n28026 = n45090 & n28025 ;
  assign n28464 = n45069 & n28445 ;
  assign n28465 = n28066 | n28464 ;
  assign n45091 = ~n28447 ;
  assign n28466 = n45091 & n28465 ;
  assign n45092 = ~n28466 ;
  assign n28467 = n152 & n45092 ;
  assign n28468 = n45079 & n28465 ;
  assign n28469 = n28023 | n28468 ;
  assign n45093 = ~n28467 ;
  assign n28470 = n45093 & n28469 ;
  assign n45094 = ~n28470 ;
  assign n28471 = n153 & n45094 ;
  assign n28472 = n154 | n28471 ;
  assign n45095 = ~n28472 ;
  assign n28473 = n28454 & n45095 ;
  assign n28474 = n28026 | n28473 ;
  assign n45096 = ~n28456 ;
  assign n28475 = n45096 & n28474 ;
  assign n45097 = ~n28475 ;
  assign n28476 = n155 & n45097 ;
  assign n27550 = n27516 | n27534 ;
  assign n45098 = ~n27550 ;
  assign n28009 = n45098 & n133 ;
  assign n28010 = n27112 | n28009 ;
  assign n45099 = ~n27516 ;
  assign n27522 = n27112 & n45099 ;
  assign n27523 = n44625 & n27522 ;
  assign n28108 = n27523 & n133 ;
  assign n45100 = ~n28108 ;
  assign n28109 = n28010 & n45100 ;
  assign n28457 = n11067 | n28456 ;
  assign n45101 = ~n28457 ;
  assign n28477 = n45101 & n28474 ;
  assign n28478 = n28109 | n28477 ;
  assign n45102 = ~n28476 ;
  assign n28479 = n45102 & n28478 ;
  assign n45103 = ~n28479 ;
  assign n28480 = n10657 & n45103 ;
  assign n27549 = n27519 | n27536 ;
  assign n45104 = ~n27549 ;
  assign n28016 = n45104 & n133 ;
  assign n28017 = n27129 | n28016 ;
  assign n27520 = n27129 & n44635 ;
  assign n45105 = ~n27536 ;
  assign n27548 = n27520 & n45105 ;
  assign n28056 = n27548 & n133 ;
  assign n45106 = ~n28056 ;
  assign n28057 = n28017 & n45106 ;
  assign n28488 = n45085 & n28469 ;
  assign n28489 = n28046 | n28488 ;
  assign n45107 = ~n28471 ;
  assign n28490 = n45107 & n28489 ;
  assign n45108 = ~n28490 ;
  assign n28491 = n154 & n45108 ;
  assign n28492 = n45095 & n28489 ;
  assign n28493 = n28026 | n28492 ;
  assign n45109 = ~n28491 ;
  assign n28494 = n45109 & n28493 ;
  assign n45110 = ~n28494 ;
  assign n28495 = n11067 & n45110 ;
  assign n28496 = n10657 | n28495 ;
  assign n45111 = ~n28496 ;
  assign n28497 = n28478 & n45111 ;
  assign n28498 = n28057 | n28497 ;
  assign n45112 = ~n28480 ;
  assign n28499 = n45112 & n28498 ;
  assign n45113 = ~n28499 ;
  assign n28500 = n157 & n45113 ;
  assign n45114 = ~n27540 ;
  assign n27546 = n27064 & n45114 ;
  assign n27547 = n44641 & n27546 ;
  assign n28011 = n27547 & n133 ;
  assign n27574 = n27540 | n27558 ;
  assign n45115 = ~n27574 ;
  assign n28096 = n45115 & n133 ;
  assign n28097 = n27064 | n28096 ;
  assign n45116 = ~n28011 ;
  assign n28098 = n45116 & n28097 ;
  assign n28481 = n157 | n28480 ;
  assign n45117 = ~n28481 ;
  assign n28501 = n45117 & n28498 ;
  assign n28505 = n28098 | n28501 ;
  assign n45118 = ~n28500 ;
  assign n28506 = n45118 & n28505 ;
  assign n45119 = ~n28506 ;
  assign n28507 = n158 & n45119 ;
  assign n27545 = n27139 & n44651 ;
  assign n45120 = ~n27560 ;
  assign n27572 = n27545 & n45120 ;
  assign n28005 = n27572 & n133 ;
  assign n27573 = n27543 | n27560 ;
  assign n45121 = ~n27573 ;
  assign n28006 = n45121 & n133 ;
  assign n28007 = n27139 | n28006 ;
  assign n45122 = ~n28005 ;
  assign n28008 = n45122 & n28007 ;
  assign n28512 = n45101 & n28493 ;
  assign n28513 = n28109 | n28512 ;
  assign n45123 = ~n28495 ;
  assign n28514 = n45123 & n28513 ;
  assign n45124 = ~n28514 ;
  assign n28515 = n156 & n45124 ;
  assign n28516 = n45111 & n28513 ;
  assign n28517 = n28057 | n28516 ;
  assign n45125 = ~n28515 ;
  assign n28518 = n45125 & n28517 ;
  assign n45126 = ~n28518 ;
  assign n28519 = n157 & n45126 ;
  assign n28520 = n158 | n28519 ;
  assign n45127 = ~n28520 ;
  assign n28521 = n28505 & n45127 ;
  assign n28522 = n28008 | n28521 ;
  assign n45128 = ~n28507 ;
  assign n28523 = n45128 & n28522 ;
  assign n45129 = ~n28523 ;
  assign n28524 = n159 & n45129 ;
  assign n27598 = n27564 | n27582 ;
  assign n45130 = ~n27598 ;
  assign n28003 = n45130 & n133 ;
  assign n28004 = n27071 | n28003 ;
  assign n45131 = ~n27564 ;
  assign n27570 = n27071 & n45131 ;
  assign n27571 = n44657 & n27570 ;
  assign n28087 = n27571 & n133 ;
  assign n45132 = ~n28087 ;
  assign n28088 = n28004 & n45132 ;
  assign n28509 = n8857 | n28507 ;
  assign n45133 = ~n28509 ;
  assign n28525 = n45133 & n28522 ;
  assign n28526 = n28088 | n28525 ;
  assign n45134 = ~n28524 ;
  assign n28527 = n45134 & n28526 ;
  assign n45135 = ~n28527 ;
  assign n28528 = n8534 & n45135 ;
  assign n27597 = n27567 | n27584 ;
  assign n45136 = ~n27597 ;
  assign n27991 = n45136 & n133 ;
  assign n27992 = n27100 | n27991 ;
  assign n27569 = n27100 & n44667 ;
  assign n45137 = ~n27584 ;
  assign n27596 = n27569 & n45137 ;
  assign n27994 = n27596 & n133 ;
  assign n45138 = ~n27994 ;
  assign n27995 = n27992 & n45138 ;
  assign n28536 = n45117 & n28517 ;
  assign n28537 = n28098 | n28536 ;
  assign n45139 = ~n28519 ;
  assign n28538 = n45139 & n28537 ;
  assign n45140 = ~n28538 ;
  assign n28539 = n158 & n45140 ;
  assign n28540 = n45127 & n28537 ;
  assign n28541 = n28008 | n28540 ;
  assign n45141 = ~n28539 ;
  assign n28542 = n45141 & n28541 ;
  assign n45142 = ~n28542 ;
  assign n28543 = n8857 & n45142 ;
  assign n28544 = n160 | n28543 ;
  assign n45143 = ~n28544 ;
  assign n28545 = n28526 & n45143 ;
  assign n28546 = n27995 | n28545 ;
  assign n45144 = ~n28528 ;
  assign n28547 = n45144 & n28546 ;
  assign n45145 = ~n28547 ;
  assign n28548 = n161 & n45145 ;
  assign n45146 = ~n27588 ;
  assign n27589 = n27142 & n45146 ;
  assign n27590 = n44673 & n27589 ;
  assign n27990 = n27590 & n133 ;
  assign n27622 = n27588 | n27606 ;
  assign n45147 = ~n27622 ;
  assign n27997 = n45147 & n133 ;
  assign n27998 = n27142 | n27997 ;
  assign n45148 = ~n27990 ;
  assign n27999 = n45148 & n27998 ;
  assign n28529 = n161 | n28528 ;
  assign n45149 = ~n28529 ;
  assign n28549 = n45149 & n28546 ;
  assign n28550 = n27999 | n28549 ;
  assign n45150 = ~n28548 ;
  assign n28551 = n45150 & n28550 ;
  assign n45151 = ~n28551 ;
  assign n28552 = n162 & n45151 ;
  assign n27595 = n27151 & n44683 ;
  assign n45152 = ~n27608 ;
  assign n27620 = n27595 & n45152 ;
  assign n27989 = n27620 & n133 ;
  assign n27621 = n27593 | n27608 ;
  assign n45153 = ~n27621 ;
  assign n28032 = n45153 & n133 ;
  assign n28033 = n27151 | n28032 ;
  assign n45154 = ~n27989 ;
  assign n28034 = n45154 & n28033 ;
  assign n28560 = n45133 & n28541 ;
  assign n28561 = n28088 | n28560 ;
  assign n45155 = ~n28543 ;
  assign n28562 = n45155 & n28561 ;
  assign n45156 = ~n28562 ;
  assign n28563 = n160 & n45156 ;
  assign n28564 = n45143 & n28561 ;
  assign n28565 = n27995 | n28564 ;
  assign n45157 = ~n28563 ;
  assign n28566 = n45157 & n28565 ;
  assign n45158 = ~n28566 ;
  assign n28567 = n161 & n45158 ;
  assign n28568 = n162 | n28567 ;
  assign n45159 = ~n28568 ;
  assign n28569 = n28550 & n45159 ;
  assign n28570 = n28034 | n28569 ;
  assign n45160 = ~n28552 ;
  assign n28571 = n45160 & n28570 ;
  assign n45161 = ~n28571 ;
  assign n28572 = n163 & n45161 ;
  assign n45162 = ~n27612 ;
  assign n27618 = n27106 & n45162 ;
  assign n27619 = n44689 & n27618 ;
  assign n27984 = n27619 & n133 ;
  assign n27646 = n27612 | n27630 ;
  assign n45163 = ~n27646 ;
  assign n28039 = n45163 & n133 ;
  assign n28040 = n27106 | n28039 ;
  assign n45164 = ~n27984 ;
  assign n28041 = n45164 & n28040 ;
  assign n28553 = n6889 | n28552 ;
  assign n45165 = ~n28553 ;
  assign n28573 = n45165 & n28570 ;
  assign n28574 = n28041 | n28573 ;
  assign n45166 = ~n28572 ;
  assign n28575 = n45166 & n28574 ;
  assign n45167 = ~n28575 ;
  assign n28576 = n6600 & n45167 ;
  assign n27617 = n27035 & n44699 ;
  assign n45168 = ~n27632 ;
  assign n27644 = n27617 & n45168 ;
  assign n27980 = n27644 & n133 ;
  assign n27645 = n27615 | n27632 ;
  assign n45169 = ~n27645 ;
  assign n28091 = n45169 & n133 ;
  assign n28092 = n27035 | n28091 ;
  assign n45170 = ~n27980 ;
  assign n28093 = n45170 & n28092 ;
  assign n28584 = n45149 & n28565 ;
  assign n28585 = n27999 | n28584 ;
  assign n45171 = ~n28567 ;
  assign n28586 = n45171 & n28585 ;
  assign n45172 = ~n28586 ;
  assign n28587 = n162 & n45172 ;
  assign n28588 = n45159 & n28585 ;
  assign n28589 = n28034 | n28588 ;
  assign n45173 = ~n28587 ;
  assign n28590 = n45173 & n28589 ;
  assign n45174 = ~n28590 ;
  assign n28591 = n6889 & n45174 ;
  assign n28592 = n6600 | n28591 ;
  assign n45175 = ~n28592 ;
  assign n28593 = n28574 & n45175 ;
  assign n28594 = n28093 | n28593 ;
  assign n45176 = ~n28576 ;
  assign n28595 = n45176 & n28594 ;
  assign n45177 = ~n28595 ;
  assign n28596 = n165 & n45177 ;
  assign n27670 = n27636 | n27654 ;
  assign n45178 = ~n27670 ;
  assign n27978 = n45178 & n133 ;
  assign n27979 = n27149 | n27978 ;
  assign n45179 = ~n27636 ;
  assign n27642 = n27149 & n45179 ;
  assign n27643 = n44705 & n27642 ;
  assign n28054 = n27643 & n133 ;
  assign n45180 = ~n28054 ;
  assign n28055 = n27979 & n45180 ;
  assign n28578 = n165 | n28576 ;
  assign n45181 = ~n28578 ;
  assign n28597 = n45181 & n28594 ;
  assign n28598 = n28055 | n28597 ;
  assign n45182 = ~n28596 ;
  assign n28599 = n45182 & n28598 ;
  assign n45183 = ~n28599 ;
  assign n28600 = n166 & n45183 ;
  assign n27641 = n27160 & n44715 ;
  assign n45184 = ~n27656 ;
  assign n27668 = n27641 & n45184 ;
  assign n28027 = n27668 & n133 ;
  assign n27669 = n27639 | n27656 ;
  assign n45185 = ~n27669 ;
  assign n28124 = n45185 & n133 ;
  assign n28125 = n27160 | n28124 ;
  assign n45186 = ~n28027 ;
  assign n28126 = n45186 & n28125 ;
  assign n28608 = n45165 & n28589 ;
  assign n28609 = n28041 | n28608 ;
  assign n45187 = ~n28591 ;
  assign n28610 = n45187 & n28609 ;
  assign n45188 = ~n28610 ;
  assign n28611 = n164 & n45188 ;
  assign n28612 = n45175 & n28609 ;
  assign n28613 = n28093 | n28612 ;
  assign n45189 = ~n28611 ;
  assign n28614 = n45189 & n28613 ;
  assign n45190 = ~n28614 ;
  assign n28615 = n165 & n45190 ;
  assign n28616 = n166 | n28615 ;
  assign n45191 = ~n28616 ;
  assign n28617 = n28598 & n45191 ;
  assign n28618 = n28126 | n28617 ;
  assign n45192 = ~n28600 ;
  assign n28619 = n45192 & n28618 ;
  assign n45193 = ~n28619 ;
  assign n28620 = n167 & n45193 ;
  assign n27694 = n27660 | n27678 ;
  assign n45194 = ~n27694 ;
  assign n28014 = n45194 & n133 ;
  assign n28015 = n27165 | n28014 ;
  assign n45195 = ~n27660 ;
  assign n27661 = n27165 & n45195 ;
  assign n27662 = n44721 & n27661 ;
  assign n28130 = n27662 & n133 ;
  assign n45196 = ~n28130 ;
  assign n28131 = n28015 & n45196 ;
  assign n28602 = n5352 | n28600 ;
  assign n45197 = ~n28602 ;
  assign n28621 = n45197 & n28618 ;
  assign n28622 = n28131 | n28621 ;
  assign n45198 = ~n28620 ;
  assign n28623 = n45198 & n28622 ;
  assign n45199 = ~n28623 ;
  assign n28624 = n4934 & n45199 ;
  assign n27693 = n27665 | n27680 ;
  assign n45200 = ~n27693 ;
  assign n28036 = n45200 & n133 ;
  assign n28037 = n27170 | n28036 ;
  assign n27667 = n27170 & n44731 ;
  assign n45201 = ~n27680 ;
  assign n27692 = n27667 & n45201 ;
  assign n28135 = n27692 & n133 ;
  assign n45202 = ~n28135 ;
  assign n28136 = n28037 & n45202 ;
  assign n28632 = n45181 & n28613 ;
  assign n28633 = n28055 | n28632 ;
  assign n45203 = ~n28615 ;
  assign n28634 = n45203 & n28633 ;
  assign n45204 = ~n28634 ;
  assign n28635 = n166 & n45204 ;
  assign n28636 = n45191 & n28633 ;
  assign n28637 = n28126 | n28636 ;
  assign n45205 = ~n28635 ;
  assign n28638 = n45205 & n28637 ;
  assign n45206 = ~n28638 ;
  assign n28639 = n5352 & n45206 ;
  assign n28640 = n4934 | n28639 ;
  assign n45207 = ~n28640 ;
  assign n28641 = n28622 & n45207 ;
  assign n28642 = n28136 | n28641 ;
  assign n45208 = ~n28624 ;
  assign n28643 = n45208 & n28642 ;
  assign n45209 = ~n28643 ;
  assign n28644 = n169 & n45209 ;
  assign n45210 = ~n27684 ;
  assign n27690 = n27174 & n45210 ;
  assign n27691 = n44737 & n27690 ;
  assign n27983 = n27691 & n133 ;
  assign n27718 = n27684 | n27702 ;
  assign n45211 = ~n27718 ;
  assign n28000 = n45211 & n133 ;
  assign n28001 = n27174 | n28000 ;
  assign n45212 = ~n27983 ;
  assign n28002 = n45212 & n28001 ;
  assign n28625 = n169 | n28624 ;
  assign n45213 = ~n28625 ;
  assign n28645 = n45213 & n28642 ;
  assign n28646 = n28002 | n28645 ;
  assign n45214 = ~n28644 ;
  assign n28647 = n45214 & n28646 ;
  assign n45215 = ~n28647 ;
  assign n28648 = n170 & n45215 ;
  assign n27717 = n27687 | n27704 ;
  assign n45216 = ~n27717 ;
  assign n28079 = n45216 & n133 ;
  assign n28080 = n27177 | n28079 ;
  assign n27688 = n27177 & n44747 ;
  assign n45217 = ~n27704 ;
  assign n27716 = n27688 & n45217 ;
  assign n28094 = n27716 & n133 ;
  assign n45218 = ~n28094 ;
  assign n28095 = n28080 & n45218 ;
  assign n28656 = n45197 & n28637 ;
  assign n28657 = n28131 | n28656 ;
  assign n45219 = ~n28639 ;
  assign n28658 = n45219 & n28657 ;
  assign n45220 = ~n28658 ;
  assign n28659 = n168 & n45220 ;
  assign n28660 = n45207 & n28657 ;
  assign n28661 = n28136 | n28660 ;
  assign n45221 = ~n28659 ;
  assign n28662 = n45221 & n28661 ;
  assign n45222 = ~n28662 ;
  assign n28663 = n169 & n45222 ;
  assign n28664 = n170 | n28663 ;
  assign n45223 = ~n28664 ;
  assign n28665 = n28646 & n45223 ;
  assign n28666 = n28095 | n28665 ;
  assign n45224 = ~n28648 ;
  assign n28667 = n45224 & n28666 ;
  assign n45225 = ~n28667 ;
  assign n28668 = n171 & n45225 ;
  assign n27742 = n27708 | n27726 ;
  assign n45226 = ~n27742 ;
  assign n28137 = n45226 & n133 ;
  assign n28138 = n27180 | n28137 ;
  assign n45227 = ~n27708 ;
  assign n27714 = n27180 & n45227 ;
  assign n27715 = n44753 & n27714 ;
  assign n28139 = n27715 & n133 ;
  assign n45228 = ~n28139 ;
  assign n28140 = n28138 & n45228 ;
  assign n28649 = n3940 | n28648 ;
  assign n45229 = ~n28649 ;
  assign n28669 = n45229 & n28666 ;
  assign n28673 = n28140 | n28669 ;
  assign n45230 = ~n28668 ;
  assign n28674 = n45230 & n28673 ;
  assign n45231 = ~n28674 ;
  assign n28675 = n3631 & n45231 ;
  assign n27741 = n27711 | n27728 ;
  assign n45232 = ~n27741 ;
  assign n28047 = n45232 & n133 ;
  assign n28048 = n27123 | n28047 ;
  assign n27713 = n27123 & n44763 ;
  assign n45233 = ~n27728 ;
  assign n27740 = n27713 & n45233 ;
  assign n28101 = n27740 & n133 ;
  assign n45234 = ~n28101 ;
  assign n28102 = n28048 & n45234 ;
  assign n28680 = n45213 & n28661 ;
  assign n28681 = n28002 | n28680 ;
  assign n45235 = ~n28663 ;
  assign n28682 = n45235 & n28681 ;
  assign n45236 = ~n28682 ;
  assign n28683 = n170 & n45236 ;
  assign n28684 = n45223 & n28681 ;
  assign n28685 = n28095 | n28684 ;
  assign n45237 = ~n28683 ;
  assign n28686 = n45237 & n28685 ;
  assign n45238 = ~n28686 ;
  assign n28687 = n3940 & n45238 ;
  assign n28688 = n3631 | n28687 ;
  assign n45239 = ~n28688 ;
  assign n28689 = n28673 & n45239 ;
  assign n28690 = n28102 | n28689 ;
  assign n45240 = ~n28675 ;
  assign n28691 = n45240 & n28690 ;
  assign n45241 = ~n28691 ;
  assign n28692 = n173 & n45241 ;
  assign n27766 = n27732 | n27750 ;
  assign n45242 = ~n27766 ;
  assign n28132 = n45242 & n133 ;
  assign n28133 = n27186 | n28132 ;
  assign n45243 = ~n27732 ;
  assign n27738 = n27186 & n45243 ;
  assign n27739 = n44769 & n27738 ;
  assign n28141 = n27739 & n133 ;
  assign n45244 = ~n28141 ;
  assign n28142 = n28133 & n45244 ;
  assign n28676 = n173 | n28675 ;
  assign n45245 = ~n28676 ;
  assign n28693 = n45245 & n28690 ;
  assign n28694 = n28142 | n28693 ;
  assign n45246 = ~n28692 ;
  assign n28695 = n45246 & n28694 ;
  assign n45247 = ~n28695 ;
  assign n28696 = n174 & n45247 ;
  assign n27765 = n27735 | n27752 ;
  assign n45248 = ~n27765 ;
  assign n28144 = n45248 & n133 ;
  assign n28145 = n27188 | n28144 ;
  assign n27737 = n27188 & n44779 ;
  assign n45249 = ~n27752 ;
  assign n27764 = n27737 & n45249 ;
  assign n28146 = n27764 & n133 ;
  assign n45250 = ~n28146 ;
  assign n28147 = n28145 & n45250 ;
  assign n28704 = n45229 & n28685 ;
  assign n28705 = n28140 | n28704 ;
  assign n45251 = ~n28687 ;
  assign n28706 = n45251 & n28705 ;
  assign n45252 = ~n28706 ;
  assign n28707 = n172 & n45252 ;
  assign n28708 = n45239 & n28705 ;
  assign n28709 = n28102 | n28708 ;
  assign n45253 = ~n28707 ;
  assign n28710 = n45253 & n28709 ;
  assign n45254 = ~n28710 ;
  assign n28711 = n173 & n45254 ;
  assign n28712 = n174 | n28711 ;
  assign n45255 = ~n28712 ;
  assign n28713 = n28694 & n45255 ;
  assign n28714 = n28147 | n28713 ;
  assign n45256 = ~n28696 ;
  assign n28715 = n45256 & n28714 ;
  assign n45257 = ~n28715 ;
  assign n28716 = n175 & n45257 ;
  assign n27790 = n27756 | n27774 ;
  assign n45258 = ~n27790 ;
  assign n28148 = n45258 & n133 ;
  assign n28149 = n27194 | n28148 ;
  assign n45259 = ~n27756 ;
  assign n27762 = n27194 & n45259 ;
  assign n27763 = n44785 & n27762 ;
  assign n28153 = n27763 & n133 ;
  assign n45260 = ~n28153 ;
  assign n28154 = n28149 & n45260 ;
  assign n28697 = n2753 | n28696 ;
  assign n45261 = ~n28697 ;
  assign n28717 = n45261 & n28714 ;
  assign n28718 = n28154 | n28717 ;
  assign n45262 = ~n28716 ;
  assign n28719 = n45262 & n28718 ;
  assign n45263 = ~n28719 ;
  assign n28720 = n2431 & n45263 ;
  assign n27761 = n27197 & n44795 ;
  assign n45264 = ~n27776 ;
  assign n27788 = n27761 & n45264 ;
  assign n28103 = n27788 & n133 ;
  assign n27789 = n27759 | n27776 ;
  assign n45265 = ~n27789 ;
  assign n28155 = n45265 & n133 ;
  assign n28156 = n27197 | n28155 ;
  assign n45266 = ~n28103 ;
  assign n28157 = n45266 & n28156 ;
  assign n28728 = n45245 & n28709 ;
  assign n28729 = n28142 | n28728 ;
  assign n45267 = ~n28711 ;
  assign n28730 = n45267 & n28729 ;
  assign n45268 = ~n28730 ;
  assign n28731 = n174 & n45268 ;
  assign n28732 = n45255 & n28729 ;
  assign n28733 = n28147 | n28732 ;
  assign n45269 = ~n28731 ;
  assign n28734 = n45269 & n28733 ;
  assign n45270 = ~n28734 ;
  assign n28735 = n2753 & n45270 ;
  assign n28736 = n2431 | n28735 ;
  assign n45271 = ~n28736 ;
  assign n28737 = n28718 & n45271 ;
  assign n28738 = n28157 | n28737 ;
  assign n45272 = ~n28720 ;
  assign n28739 = n45272 & n28738 ;
  assign n45273 = ~n28739 ;
  assign n28740 = n177 & n45273 ;
  assign n45274 = ~n27780 ;
  assign n27786 = n27091 & n45274 ;
  assign n27787 = n44801 & n27786 ;
  assign n28067 = n27787 & n133 ;
  assign n27814 = n27780 | n27798 ;
  assign n45275 = ~n27814 ;
  assign n28158 = n45275 & n133 ;
  assign n28159 = n27091 | n28158 ;
  assign n45276 = ~n28067 ;
  assign n28160 = n45276 & n28159 ;
  assign n28721 = n177 | n28720 ;
  assign n45277 = ~n28721 ;
  assign n28741 = n45277 & n28738 ;
  assign n28742 = n28160 | n28741 ;
  assign n45278 = ~n28740 ;
  assign n28743 = n45278 & n28742 ;
  assign n45279 = ~n28743 ;
  assign n28744 = n178 & n45279 ;
  assign n27785 = n27201 & n44811 ;
  assign n45280 = ~n27800 ;
  assign n27812 = n27785 & n45280 ;
  assign n28042 = n27812 & n133 ;
  assign n27813 = n27783 | n27800 ;
  assign n45281 = ~n27813 ;
  assign n28165 = n45281 & n133 ;
  assign n28166 = n27201 | n28165 ;
  assign n45282 = ~n28042 ;
  assign n28167 = n45282 & n28166 ;
  assign n28752 = n45261 & n28733 ;
  assign n28753 = n28154 | n28752 ;
  assign n45283 = ~n28735 ;
  assign n28754 = n45283 & n28753 ;
  assign n45284 = ~n28754 ;
  assign n28755 = n176 & n45284 ;
  assign n28756 = n45271 & n28753 ;
  assign n28757 = n28157 | n28756 ;
  assign n45285 = ~n28755 ;
  assign n28758 = n45285 & n28757 ;
  assign n45286 = ~n28758 ;
  assign n28759 = n177 & n45286 ;
  assign n28760 = n178 | n28759 ;
  assign n45287 = ~n28760 ;
  assign n28761 = n28742 & n45287 ;
  assign n28762 = n28167 | n28761 ;
  assign n45288 = ~n28744 ;
  assign n28763 = n45288 & n28762 ;
  assign n45289 = ~n28763 ;
  assign n28764 = n179 & n45289 ;
  assign n27838 = n27804 | n27822 ;
  assign n45290 = ~n27838 ;
  assign n28168 = n45290 & n133 ;
  assign n28169 = n27204 | n28168 ;
  assign n45291 = ~n27804 ;
  assign n27810 = n27204 & n45291 ;
  assign n27811 = n44817 & n27810 ;
  assign n28170 = n27811 & n133 ;
  assign n45292 = ~n28170 ;
  assign n28171 = n28169 & n45292 ;
  assign n28745 = n1707 | n28744 ;
  assign n45293 = ~n28745 ;
  assign n28765 = n45293 & n28762 ;
  assign n28766 = n28171 | n28765 ;
  assign n45294 = ~n28764 ;
  assign n28767 = n45294 & n28766 ;
  assign n45295 = ~n28767 ;
  assign n28768 = n1487 & n45295 ;
  assign n27809 = n27208 & n44827 ;
  assign n45296 = ~n27824 ;
  assign n27836 = n27809 & n45296 ;
  assign n28143 = n27836 & n133 ;
  assign n27837 = n27807 | n27824 ;
  assign n45297 = ~n27837 ;
  assign n28172 = n45297 & n133 ;
  assign n28173 = n27208 | n28172 ;
  assign n45298 = ~n28143 ;
  assign n28174 = n45298 & n28173 ;
  assign n28776 = n45277 & n28757 ;
  assign n28777 = n28160 | n28776 ;
  assign n45299 = ~n28759 ;
  assign n28778 = n45299 & n28777 ;
  assign n45300 = ~n28778 ;
  assign n28779 = n178 & n45300 ;
  assign n28780 = n45287 & n28777 ;
  assign n28781 = n28167 | n28780 ;
  assign n45301 = ~n28779 ;
  assign n28782 = n45301 & n28781 ;
  assign n45302 = ~n28782 ;
  assign n28783 = n1707 & n45302 ;
  assign n28784 = n1487 | n28783 ;
  assign n45303 = ~n28784 ;
  assign n28785 = n28766 & n45303 ;
  assign n28786 = n28174 | n28785 ;
  assign n45304 = ~n28768 ;
  assign n28787 = n45304 & n28786 ;
  assign n45305 = ~n28787 ;
  assign n28788 = n181 & n45305 ;
  assign n45306 = ~n27828 ;
  assign n27834 = n27125 & n45306 ;
  assign n27835 = n44833 & n27834 ;
  assign n28038 = n27835 & n133 ;
  assign n27862 = n27828 | n27846 ;
  assign n45307 = ~n27862 ;
  assign n28175 = n45307 & n133 ;
  assign n28176 = n27125 | n28175 ;
  assign n45308 = ~n28038 ;
  assign n28177 = n45308 & n28176 ;
  assign n28769 = n181 | n28768 ;
  assign n45309 = ~n28769 ;
  assign n28789 = n45309 & n28786 ;
  assign n28790 = n28177 | n28789 ;
  assign n45310 = ~n28788 ;
  assign n28791 = n45310 & n28790 ;
  assign n45311 = ~n28791 ;
  assign n28792 = n182 & n45311 ;
  assign n27833 = n27192 & n44843 ;
  assign n45312 = ~n27848 ;
  assign n27860 = n27833 & n45312 ;
  assign n28161 = n27860 & n133 ;
  assign n27861 = n27831 | n27848 ;
  assign n45313 = ~n27861 ;
  assign n28178 = n45313 & n133 ;
  assign n28179 = n27192 | n28178 ;
  assign n45314 = ~n28161 ;
  assign n28180 = n45314 & n28179 ;
  assign n28800 = n45293 & n28781 ;
  assign n28801 = n28171 | n28800 ;
  assign n45315 = ~n28783 ;
  assign n28802 = n45315 & n28801 ;
  assign n45316 = ~n28802 ;
  assign n28803 = n180 & n45316 ;
  assign n28804 = n45303 & n28801 ;
  assign n28805 = n28174 | n28804 ;
  assign n45317 = ~n28803 ;
  assign n28806 = n45317 & n28805 ;
  assign n45318 = ~n28806 ;
  assign n28807 = n181 & n45318 ;
  assign n28808 = n182 | n28807 ;
  assign n45319 = ~n28808 ;
  assign n28809 = n28790 & n45319 ;
  assign n28810 = n28180 | n28809 ;
  assign n45320 = ~n28792 ;
  assign n28811 = n45320 & n28810 ;
  assign n45321 = ~n28811 ;
  assign n28812 = n183 & n45321 ;
  assign n45322 = ~n27852 ;
  assign n27853 = n27153 & n45322 ;
  assign n27854 = n44849 & n27853 ;
  assign n28043 = n27854 & n133 ;
  assign n27886 = n27852 | n27870 ;
  assign n45323 = ~n27886 ;
  assign n28127 = n45323 & n133 ;
  assign n28128 = n27153 | n28127 ;
  assign n45324 = ~n28043 ;
  assign n28129 = n45324 & n28128 ;
  assign n28793 = n183 | n28792 ;
  assign n45325 = ~n28793 ;
  assign n28813 = n45325 & n28810 ;
  assign n28814 = n28129 | n28813 ;
  assign n45326 = ~n28812 ;
  assign n28815 = n45326 & n28814 ;
  assign n45327 = ~n28815 ;
  assign n28816 = n838 & n45327 ;
  assign n27885 = n27857 | n27872 ;
  assign n45328 = ~n27885 ;
  assign n28181 = n45328 & n133 ;
  assign n28182 = n27212 | n28181 ;
  assign n27859 = n27212 & n44859 ;
  assign n45329 = ~n27872 ;
  assign n27884 = n27859 & n45329 ;
  assign n28183 = n27884 & n133 ;
  assign n45330 = ~n28183 ;
  assign n28184 = n28182 & n45330 ;
  assign n28824 = n45309 & n28805 ;
  assign n28825 = n28177 | n28824 ;
  assign n45331 = ~n28807 ;
  assign n28826 = n45331 & n28825 ;
  assign n45332 = ~n28826 ;
  assign n28827 = n182 & n45332 ;
  assign n28828 = n45319 & n28825 ;
  assign n28829 = n28180 | n28828 ;
  assign n45333 = ~n28827 ;
  assign n28830 = n45333 & n28829 ;
  assign n45334 = ~n28830 ;
  assign n28831 = n996 & n45334 ;
  assign n28832 = n838 | n28831 ;
  assign n45335 = ~n28832 ;
  assign n28833 = n28814 & n45335 ;
  assign n28834 = n28184 | n28833 ;
  assign n45336 = ~n28816 ;
  assign n28835 = n45336 & n28834 ;
  assign n45337 = ~n28835 ;
  assign n28836 = n185 & n45337 ;
  assign n27910 = n27876 | n27894 ;
  assign n45338 = ~n27910 ;
  assign n28185 = n45338 & n133 ;
  assign n28186 = n27214 | n28185 ;
  assign n45339 = ~n27876 ;
  assign n27882 = n27214 & n45339 ;
  assign n27883 = n44865 & n27882 ;
  assign n28189 = n27883 & n133 ;
  assign n45340 = ~n28189 ;
  assign n28190 = n28186 & n45340 ;
  assign n28817 = n185 | n28816 ;
  assign n45341 = ~n28817 ;
  assign n28837 = n45341 & n28834 ;
  assign n28838 = n28190 | n28837 ;
  assign n45342 = ~n28836 ;
  assign n28839 = n45342 & n28838 ;
  assign n45343 = ~n28839 ;
  assign n28840 = n186 & n45343 ;
  assign n27909 = n27879 | n27896 ;
  assign n45344 = ~n27909 ;
  assign n28110 = n45344 & n133 ;
  assign n28111 = n27218 | n28110 ;
  assign n27881 = n27218 & n44875 ;
  assign n45345 = ~n27896 ;
  assign n27908 = n27881 & n45345 ;
  assign n28187 = n27908 & n133 ;
  assign n45346 = ~n28187 ;
  assign n28188 = n28111 & n45346 ;
  assign n28848 = n45325 & n28829 ;
  assign n28849 = n28129 | n28848 ;
  assign n45347 = ~n28831 ;
  assign n28850 = n45347 & n28849 ;
  assign n45348 = ~n28850 ;
  assign n28851 = n184 & n45348 ;
  assign n28852 = n45335 & n28849 ;
  assign n28853 = n28184 | n28852 ;
  assign n45349 = ~n28851 ;
  assign n28854 = n45349 & n28853 ;
  assign n45350 = ~n28854 ;
  assign n28855 = n185 & n45350 ;
  assign n28856 = n186 | n28855 ;
  assign n45351 = ~n28856 ;
  assign n28857 = n28838 & n45351 ;
  assign n28858 = n28188 | n28857 ;
  assign n45352 = ~n28840 ;
  assign n28859 = n45352 & n28858 ;
  assign n45353 = ~n28859 ;
  assign n28860 = n187 & n45353 ;
  assign n45354 = ~n27900 ;
  assign n27901 = n27220 & n45354 ;
  assign n27902 = n44881 & n27901 ;
  assign n27993 = n27902 & n133 ;
  assign n27934 = n27900 | n27918 ;
  assign n45355 = ~n27934 ;
  assign n28162 = n45355 & n133 ;
  assign n28163 = n27220 | n28162 ;
  assign n45356 = ~n27993 ;
  assign n28164 = n45356 & n28163 ;
  assign n28842 = n528 | n28840 ;
  assign n45357 = ~n28842 ;
  assign n28861 = n45357 & n28858 ;
  assign n28862 = n28164 | n28861 ;
  assign n45358 = ~n28860 ;
  assign n28863 = n45358 & n28862 ;
  assign n45359 = ~n28863 ;
  assign n28864 = n413 & n45359 ;
  assign n27907 = n27136 & n44891 ;
  assign n45360 = ~n27920 ;
  assign n27932 = n27907 & n45360 ;
  assign n28086 = n27932 & n133 ;
  assign n27933 = n27905 | n27920 ;
  assign n45361 = ~n27933 ;
  assign n28191 = n45361 & n133 ;
  assign n28192 = n27136 | n28191 ;
  assign n45362 = ~n28086 ;
  assign n28193 = n45362 & n28192 ;
  assign n28872 = n45341 & n28853 ;
  assign n28873 = n28190 | n28872 ;
  assign n45363 = ~n28855 ;
  assign n28874 = n45363 & n28873 ;
  assign n45364 = ~n28874 ;
  assign n28875 = n186 & n45364 ;
  assign n28876 = n45351 & n28873 ;
  assign n28877 = n28188 | n28876 ;
  assign n45365 = ~n28875 ;
  assign n28878 = n45365 & n28877 ;
  assign n45366 = ~n28878 ;
  assign n28879 = n528 & n45366 ;
  assign n28880 = n413 | n28879 ;
  assign n45367 = ~n28880 ;
  assign n28881 = n28862 & n45367 ;
  assign n28882 = n28193 | n28881 ;
  assign n45368 = ~n28864 ;
  assign n28883 = n45368 & n28882 ;
  assign n45369 = ~n28883 ;
  assign n28884 = n189 & n45369 ;
  assign n27958 = n27924 | n27942 ;
  assign n45370 = ~n27958 ;
  assign n28194 = n45370 & n133 ;
  assign n28195 = n27224 | n28194 ;
  assign n45371 = ~n27924 ;
  assign n27930 = n27224 & n45371 ;
  assign n27931 = n44897 & n27930 ;
  assign n28196 = n27931 & n133 ;
  assign n45372 = ~n28196 ;
  assign n28197 = n28195 & n45372 ;
  assign n28865 = n189 | n28864 ;
  assign n45373 = ~n28865 ;
  assign n28885 = n45373 & n28882 ;
  assign n28886 = n28197 | n28885 ;
  assign n45374 = ~n28884 ;
  assign n28887 = n45374 & n28886 ;
  assign n45375 = ~n28887 ;
  assign n28888 = n190 & n45375 ;
  assign n28895 = n45357 & n28877 ;
  assign n28896 = n28164 | n28895 ;
  assign n45376 = ~n28879 ;
  assign n28897 = n45376 & n28896 ;
  assign n45377 = ~n28897 ;
  assign n28898 = n188 & n45377 ;
  assign n28899 = n45367 & n28896 ;
  assign n28900 = n28193 | n28899 ;
  assign n45378 = ~n28898 ;
  assign n28901 = n45378 & n28900 ;
  assign n45379 = ~n28901 ;
  assign n28902 = n189 & n45379 ;
  assign n28903 = n190 | n28902 ;
  assign n45380 = ~n28903 ;
  assign n28904 = n28886 & n45380 ;
  assign n28909 = n28888 | n28904 ;
  assign n27973 = n27951 | n27968 ;
  assign n45381 = ~n27973 ;
  assign n28198 = n45381 & n133 ;
  assign n28199 = n27268 | n28198 ;
  assign n27953 = n27268 & n44919 ;
  assign n45382 = ~n27968 ;
  assign n27972 = n27953 & n45382 ;
  assign n28206 = n27972 & n133 ;
  assign n45383 = ~n28206 ;
  assign n28207 = n28199 & n45383 ;
  assign n28224 = n27237 | n27974 ;
  assign n45384 = ~n28224 ;
  assign n28225 = n133 & n45384 ;
  assign n28249 = n27970 | n28225 ;
  assign n28250 = n28207 | n28249 ;
  assign n28905 = n28152 | n28904 ;
  assign n45385 = ~n28888 ;
  assign n28910 = n45385 & n28905 ;
  assign n45386 = ~n28910 ;
  assign n28911 = n191 & n45386 ;
  assign n45387 = ~n27948 ;
  assign n27954 = n27230 & n45387 ;
  assign n27955 = n44917 & n27954 ;
  assign n28134 = n27955 & n133 ;
  assign n28253 = n27948 | n27966 ;
  assign n45388 = ~n28253 ;
  assign n28254 = n133 & n45388 ;
  assign n28255 = n27230 | n28254 ;
  assign n45389 = ~n28134 ;
  assign n28256 = n45389 & n28255 ;
  assign n28891 = n191 | n28888 ;
  assign n45390 = ~n28891 ;
  assign n28934 = n45390 & n28905 ;
  assign n28935 = n28256 | n28934 ;
  assign n45391 = ~n28911 ;
  assign n28936 = n45391 & n28935 ;
  assign n28937 = n28250 | n28936 ;
  assign n28938 = n31336 & n28937 ;
  assign n45392 = ~n27237 ;
  assign n28204 = n45392 & n133 ;
  assign n45393 = ~n28204 ;
  assign n28205 = n27974 & n45393 ;
  assign n28226 = n192 & n28224 ;
  assign n45394 = ~n28205 ;
  assign n28227 = n45394 & n28226 ;
  assign n28915 = n28207 & n45391 ;
  assign n28939 = n28915 & n28935 ;
  assign n28940 = n28227 | n28939 ;
  assign n132 = n28938 | n28940 ;
  assign n45395 = ~n28909 ;
  assign n29519 = n45395 & n132 ;
  assign n29520 = n28152 | n29519 ;
  assign n28889 = n28152 & n45385 ;
  assign n45396 = ~n28904 ;
  assign n28908 = n28889 & n45396 ;
  assign n29740 = n28908 & n132 ;
  assign n45397 = ~n29740 ;
  assign n29741 = n29520 & n45397 ;
  assign n28869 = n28860 | n28861 ;
  assign n45398 = ~n28869 ;
  assign n29010 = n45398 & n132 ;
  assign n29011 = n28164 | n29010 ;
  assign n45399 = ~n28861 ;
  assign n28867 = n28164 & n45399 ;
  assign n28868 = n45358 & n28867 ;
  assign n29682 = n28868 & n132 ;
  assign n45400 = ~n29682 ;
  assign n29683 = n29011 & n45400 ;
  assign n28797 = n28788 | n28789 ;
  assign n45401 = ~n28797 ;
  assign n28958 = n45401 & n132 ;
  assign n28959 = n28177 | n28958 ;
  assign n45402 = ~n28789 ;
  assign n28795 = n28177 & n45402 ;
  assign n28796 = n45310 & n28795 ;
  assign n29076 = n28796 & n132 ;
  assign n45403 = ~n29076 ;
  assign n29077 = n28959 & n45403 ;
  assign n45404 = ~n28741 ;
  assign n28747 = n28160 & n45404 ;
  assign n28748 = n45278 & n28747 ;
  assign n29057 = n28748 & n132 ;
  assign n28749 = n28740 | n28741 ;
  assign n45405 = ~n28749 ;
  assign n29431 = n45405 & n132 ;
  assign n29432 = n28160 | n29431 ;
  assign n45406 = ~n29057 ;
  assign n29433 = n45406 & n29432 ;
  assign n28701 = n28692 | n28693 ;
  assign n45407 = ~n28701 ;
  assign n29049 = n45407 & n132 ;
  assign n29050 = n28142 | n29049 ;
  assign n45408 = ~n28693 ;
  assign n28699 = n28142 & n45408 ;
  assign n28700 = n45246 & n28699 ;
  assign n29064 = n28700 & n132 ;
  assign n45409 = ~n29064 ;
  assign n29065 = n29050 & n45409 ;
  assign n45410 = ~n28645 ;
  assign n28651 = n28002 & n45410 ;
  assign n28652 = n45214 & n28651 ;
  assign n28957 = n28652 & n132 ;
  assign n28653 = n28644 | n28645 ;
  assign n45411 = ~n28653 ;
  assign n29143 = n45411 & n132 ;
  assign n29144 = n28002 | n29143 ;
  assign n45412 = ~n28957 ;
  assign n29145 = n45412 & n29144 ;
  assign n45413 = ~n28621 ;
  assign n28627 = n28131 & n45413 ;
  assign n28628 = n45198 & n28627 ;
  assign n28986 = n28628 & n132 ;
  assign n28629 = n28620 | n28621 ;
  assign n45414 = ~n28629 ;
  assign n29157 = n45414 & n132 ;
  assign n29158 = n28131 | n29157 ;
  assign n45415 = ~n28986 ;
  assign n29159 = n45415 & n29158 ;
  assign n28605 = n28596 | n28597 ;
  assign n45416 = ~n28605 ;
  assign n28946 = n45416 & n132 ;
  assign n28947 = n28055 | n28946 ;
  assign n45417 = ~n28597 ;
  assign n28603 = n28055 & n45417 ;
  assign n28604 = n45182 & n28603 ;
  assign n29019 = n28604 & n132 ;
  assign n45418 = ~n29019 ;
  assign n29020 = n28947 & n45418 ;
  assign n45419 = ~n28573 ;
  assign n28579 = n28041 & n45419 ;
  assign n28580 = n45166 & n28579 ;
  assign n28991 = n28580 & n132 ;
  assign n28581 = n28572 | n28573 ;
  assign n45420 = ~n28581 ;
  assign n29022 = n45420 & n132 ;
  assign n29023 = n28041 | n29022 ;
  assign n45421 = ~n28991 ;
  assign n29024 = n45421 & n29023 ;
  assign n45422 = ~n28549 ;
  assign n28555 = n27999 & n45422 ;
  assign n28556 = n45150 & n28555 ;
  assign n28987 = n28556 & n132 ;
  assign n28557 = n28548 | n28549 ;
  assign n45423 = ~n28557 ;
  assign n29040 = n45423 & n132 ;
  assign n29041 = n27999 | n29040 ;
  assign n45424 = ~n28987 ;
  assign n29042 = n45424 & n29041 ;
  assign n28530 = n27995 & n45144 ;
  assign n45425 = ~n28545 ;
  assign n28558 = n28530 & n45425 ;
  assign n28942 = n28558 & n132 ;
  assign n28559 = n28528 | n28545 ;
  assign n45426 = ~n28559 ;
  assign n29154 = n45426 & n132 ;
  assign n29155 = n27995 | n29154 ;
  assign n45427 = ~n28942 ;
  assign n29156 = n45427 & n29155 ;
  assign n263 = x4 | x5 ;
  assign n45428 = ~x6 ;
  assign n265 = n45428 & n263 ;
  assign n28890 = n287 | n28888 ;
  assign n45429 = ~n28890 ;
  assign n28906 = n45429 & n28905 ;
  assign n28907 = n28256 | n28906 ;
  assign n28912 = n28907 & n45391 ;
  assign n28913 = n28250 | n28912 ;
  assign n28914 = n31336 & n28913 ;
  assign n28916 = n28907 & n28915 ;
  assign n28917 = n28227 | n28916 ;
  assign n28918 = n28914 | n28917 ;
  assign n45430 = ~n28918 ;
  assign n28919 = x6 & n45430 ;
  assign n28920 = n265 | n28919 ;
  assign n45431 = ~n28920 ;
  assign n28921 = n133 & n45431 ;
  assign n45432 = ~n260 ;
  assign n29033 = n45432 & n132 ;
  assign n29084 = n45428 & n132 ;
  assign n45433 = ~n29084 ;
  assign n29085 = x7 & n45433 ;
  assign n29086 = n29033 | n29085 ;
  assign n264 = x6 | n263 ;
  assign n27252 = n264 & n44942 ;
  assign n28251 = n27252 & n44943 ;
  assign n28252 = n44944 & n28251 ;
  assign n29051 = x6 & n132 ;
  assign n45434 = ~n29051 ;
  assign n29087 = n28252 & n45434 ;
  assign n29088 = n29086 | n29087 ;
  assign n45435 = ~n28921 ;
  assign n29089 = n45435 & n29088 ;
  assign n45436 = ~n29089 ;
  assign n29090 = n134 & n45436 ;
  assign n45437 = ~n28227 ;
  assign n28229 = n133 & n45437 ;
  assign n45438 = ~n28916 ;
  assign n28927 = n28229 & n45438 ;
  assign n45439 = ~n28914 ;
  assign n28928 = n45439 & n28927 ;
  assign n28929 = x8 | n28928 ;
  assign n29034 = n28929 | n29033 ;
  assign n29071 = n28928 | n29033 ;
  assign n29072 = x8 & n29071 ;
  assign n45440 = ~n29072 ;
  assign n29073 = n29034 & n45440 ;
  assign n29052 = n264 & n45434 ;
  assign n45441 = ~n29052 ;
  assign n29053 = n133 & n45441 ;
  assign n29054 = n134 | n29053 ;
  assign n45442 = ~n29054 ;
  assign n29092 = n45442 & n29088 ;
  assign n29093 = n29073 | n29092 ;
  assign n45443 = ~n29090 ;
  assign n29094 = n45443 & n29093 ;
  assign n45444 = ~n29094 ;
  assign n29095 = n135 & n45444 ;
  assign n28075 = n28062 | n28073 ;
  assign n45445 = ~n28075 ;
  assign n28203 = n45445 & n28202 ;
  assign n28994 = n28203 & n132 ;
  assign n29068 = n45445 & n132 ;
  assign n29069 = n28202 | n29068 ;
  assign n45446 = ~n28994 ;
  assign n29070 = n45446 & n29069 ;
  assign n29091 = n135 | n29090 ;
  assign n28922 = n134 | n28921 ;
  assign n45447 = ~n28922 ;
  assign n29101 = n45447 & n29088 ;
  assign n29102 = n29073 | n29101 ;
  assign n45448 = ~n29091 ;
  assign n29103 = n45448 & n29102 ;
  assign n29106 = n29070 | n29103 ;
  assign n45449 = ~n29095 ;
  assign n29107 = n45449 & n29106 ;
  assign n45450 = ~n29107 ;
  assign n29108 = n136 & n45450 ;
  assign n45451 = ~n28221 ;
  assign n28243 = n45451 & n28236 ;
  assign n28244 = n44963 & n28243 ;
  assign n29021 = n28244 & n132 ;
  assign n28222 = n28216 | n28221 ;
  assign n45452 = ~n28222 ;
  assign n29078 = n45452 & n132 ;
  assign n29079 = n28236 | n29078 ;
  assign n45453 = ~n29021 ;
  assign n29080 = n45453 & n29079 ;
  assign n29097 = n26442 & n45444 ;
  assign n29098 = n25517 | n29097 ;
  assign n45454 = ~n29098 ;
  assign n29110 = n45454 & n29106 ;
  assign n29111 = n29080 | n29110 ;
  assign n45455 = ~n29108 ;
  assign n29112 = n45455 & n29111 ;
  assign n45456 = ~n29112 ;
  assign n29113 = n137 & n45456 ;
  assign n28242 = n28239 | n28241 ;
  assign n45457 = ~n28242 ;
  assign n28996 = n45457 & n132 ;
  assign n28997 = n28262 | n28996 ;
  assign n28263 = n44951 & n28262 ;
  assign n45458 = ~n28241 ;
  assign n28264 = n45458 & n28263 ;
  assign n29012 = n28264 & n132 ;
  assign n45459 = ~n29012 ;
  assign n29013 = n28997 & n45459 ;
  assign n29109 = n137 | n29108 ;
  assign n45460 = ~n29109 ;
  assign n29116 = n45460 & n29111 ;
  assign n29117 = n29013 | n29116 ;
  assign n45461 = ~n29113 ;
  assign n29118 = n45461 & n29117 ;
  assign n45462 = ~n29118 ;
  assign n29119 = n138 & n45462 ;
  assign n45463 = ~n28268 ;
  assign n28274 = n28211 & n45463 ;
  assign n28294 = n28274 & n44979 ;
  assign n28978 = n28294 & n132 ;
  assign n28295 = n28268 | n28277 ;
  assign n45464 = ~n28295 ;
  assign n28988 = n45464 & n132 ;
  assign n28989 = n28211 | n28988 ;
  assign n45465 = ~n28978 ;
  assign n28990 = n45465 & n28989 ;
  assign n29114 = n138 | n29113 ;
  assign n45466 = ~n29114 ;
  assign n29120 = n45466 & n29117 ;
  assign n29121 = n28990 | n29120 ;
  assign n45467 = ~n29119 ;
  assign n29122 = n45467 & n29121 ;
  assign n45468 = ~n29122 ;
  assign n29127 = n139 & n45468 ;
  assign n29125 = n139 | n29119 ;
  assign n45469 = ~n29125 ;
  assign n29126 = n29121 & n45469 ;
  assign n28293 = n28271 | n28279 ;
  assign n45470 = ~n28293 ;
  assign n29074 = n45470 & n132 ;
  assign n29075 = n28209 | n29074 ;
  assign n28273 = n28209 & n44968 ;
  assign n45471 = ~n28279 ;
  assign n28292 = n28273 & n45471 ;
  assign n29166 = n28292 & n132 ;
  assign n45472 = ~n29166 ;
  assign n29167 = n29075 & n45472 ;
  assign n29168 = n29126 | n29167 ;
  assign n45473 = ~n29127 ;
  assign n29169 = n45473 & n29168 ;
  assign n45474 = ~n29169 ;
  assign n29170 = n22030 & n45474 ;
  assign n28291 = n28282 | n28283 ;
  assign n45475 = ~n28291 ;
  assign n29005 = n45475 & n132 ;
  assign n29006 = n28083 | n29005 ;
  assign n45476 = ~n28283 ;
  assign n28289 = n28083 & n45476 ;
  assign n28290 = n44974 & n28289 ;
  assign n29014 = n28290 & n132 ;
  assign n45477 = ~n29014 ;
  assign n29015 = n29006 & n45477 ;
  assign n29123 = n22661 & n45468 ;
  assign n29124 = n140 | n29123 ;
  assign n45478 = ~n29124 ;
  assign n29172 = n45478 & n29168 ;
  assign n29173 = n29015 | n29172 ;
  assign n45479 = ~n29170 ;
  assign n29174 = n45479 & n29173 ;
  assign n45480 = ~n29174 ;
  assign n29175 = n141 & n45480 ;
  assign n28288 = n28052 & n44984 ;
  assign n45481 = ~n28305 ;
  assign n28318 = n28288 & n45481 ;
  assign n29142 = n28318 & n132 ;
  assign n28319 = n28286 | n28305 ;
  assign n45482 = ~n28319 ;
  assign n29146 = n45482 & n132 ;
  assign n29147 = n28052 | n29146 ;
  assign n45483 = ~n29142 ;
  assign n29148 = n45483 & n29147 ;
  assign n29171 = n141 | n29170 ;
  assign n45484 = ~n29171 ;
  assign n29176 = n45484 & n29173 ;
  assign n29177 = n29148 | n29176 ;
  assign n45485 = ~n29175 ;
  assign n29178 = n45485 & n29177 ;
  assign n45486 = ~n29178 ;
  assign n29179 = n142 & n45486 ;
  assign n45487 = ~n28309 ;
  assign n28315 = n28031 & n45487 ;
  assign n28316 = n44990 & n28315 ;
  assign n29009 = n28316 & n132 ;
  assign n28317 = n28308 | n28309 ;
  assign n45488 = ~n28317 ;
  assign n29149 = n45488 & n132 ;
  assign n29150 = n28031 | n29149 ;
  assign n45489 = ~n29009 ;
  assign n29151 = n45489 & n29150 ;
  assign n45490 = ~n29123 ;
  assign n29186 = n45490 & n29168 ;
  assign n45491 = ~n29186 ;
  assign n29187 = n140 & n45491 ;
  assign n45492 = ~n29187 ;
  assign n29188 = n29173 & n45492 ;
  assign n45493 = ~n29188 ;
  assign n29189 = n141 & n45493 ;
  assign n29190 = n142 | n29189 ;
  assign n45494 = ~n29190 ;
  assign n29191 = n29177 & n45494 ;
  assign n29192 = n29151 | n29191 ;
  assign n45495 = ~n29179 ;
  assign n29193 = n45495 & n29192 ;
  assign n45496 = ~n29193 ;
  assign n29194 = n143 & n45496 ;
  assign n28314 = n28090 & n45000 ;
  assign n45497 = ~n28329 ;
  assign n28342 = n28314 & n45497 ;
  assign n28995 = n28342 & n132 ;
  assign n28343 = n28312 | n28329 ;
  assign n45498 = ~n28343 ;
  assign n29058 = n45498 & n132 ;
  assign n29059 = n28090 | n29058 ;
  assign n45499 = ~n28995 ;
  assign n29060 = n45499 & n29059 ;
  assign n29180 = n143 | n29179 ;
  assign n45500 = ~n29180 ;
  assign n29195 = n45500 & n29192 ;
  assign n29196 = n29060 | n29195 ;
  assign n45501 = ~n29194 ;
  assign n29197 = n45501 & n29196 ;
  assign n45502 = ~n29197 ;
  assign n29198 = n18797 & n45502 ;
  assign n45503 = ~n28333 ;
  assign n28339 = n28117 & n45503 ;
  assign n28340 = n45006 & n28339 ;
  assign n29160 = n28340 & n132 ;
  assign n28341 = n28332 | n28333 ;
  assign n45504 = ~n28341 ;
  assign n29161 = n45504 & n132 ;
  assign n29162 = n28117 | n29161 ;
  assign n45505 = ~n29160 ;
  assign n29163 = n45505 & n29162 ;
  assign n45506 = ~n29189 ;
  assign n29207 = n29177 & n45506 ;
  assign n45507 = ~n29207 ;
  assign n29208 = n142 & n45507 ;
  assign n45508 = ~n29208 ;
  assign n29209 = n29192 & n45508 ;
  assign n45509 = ~n29209 ;
  assign n29210 = n19362 & n45509 ;
  assign n29211 = n144 | n29210 ;
  assign n45510 = ~n29211 ;
  assign n29212 = n29196 & n45510 ;
  assign n29213 = n29163 | n29212 ;
  assign n45511 = ~n29198 ;
  assign n29214 = n45511 & n29213 ;
  assign n45512 = ~n29214 ;
  assign n29215 = n145 & n45512 ;
  assign n28338 = n28100 & n45016 ;
  assign n45513 = ~n28353 ;
  assign n28366 = n28338 & n45513 ;
  assign n28961 = n28366 & n132 ;
  assign n28367 = n28336 | n28353 ;
  assign n45514 = ~n28367 ;
  assign n29037 = n45514 & n132 ;
  assign n29038 = n28100 | n29037 ;
  assign n45515 = ~n28961 ;
  assign n29039 = n45515 & n29038 ;
  assign n29199 = n145 | n29198 ;
  assign n45516 = ~n29199 ;
  assign n29216 = n45516 & n29213 ;
  assign n29217 = n29039 | n29216 ;
  assign n45517 = ~n29215 ;
  assign n29218 = n45517 & n29217 ;
  assign n45518 = ~n29218 ;
  assign n29219 = n146 & n45518 ;
  assign n28365 = n28356 | n28357 ;
  assign n45519 = ~n28365 ;
  assign n28998 = n45519 & n132 ;
  assign n28999 = n28078 | n28998 ;
  assign n45520 = ~n28357 ;
  assign n28363 = n28078 & n45520 ;
  assign n28364 = n45022 & n28363 ;
  assign n29140 = n28364 & n132 ;
  assign n45521 = ~n29140 ;
  assign n29141 = n28999 & n45521 ;
  assign n45522 = ~n29210 ;
  assign n29227 = n29196 & n45522 ;
  assign n45523 = ~n29227 ;
  assign n29228 = n144 & n45523 ;
  assign n45524 = ~n29228 ;
  assign n29229 = n29213 & n45524 ;
  assign n45525 = ~n29229 ;
  assign n29230 = n145 & n45525 ;
  assign n29231 = n146 | n29230 ;
  assign n45526 = ~n29231 ;
  assign n29232 = n29217 & n45526 ;
  assign n29233 = n29141 | n29232 ;
  assign n45527 = ~n29219 ;
  assign n29234 = n45527 & n29233 ;
  assign n45528 = ~n29234 ;
  assign n29235 = n147 & n45528 ;
  assign n28391 = n28360 | n28377 ;
  assign n45529 = ~n28391 ;
  assign n29045 = n45529 & n132 ;
  assign n29046 = n28107 | n29045 ;
  assign n28362 = n28107 & n45032 ;
  assign n45530 = ~n28377 ;
  assign n28390 = n28362 & n45530 ;
  assign n29047 = n28390 & n132 ;
  assign n45531 = ~n29047 ;
  assign n29048 = n29046 & n45531 ;
  assign n29220 = n147 | n29219 ;
  assign n45532 = ~n29220 ;
  assign n29236 = n45532 & n29233 ;
  assign n29237 = n29048 | n29236 ;
  assign n45533 = ~n29235 ;
  assign n29238 = n45533 & n29237 ;
  assign n45534 = ~n29238 ;
  assign n29239 = n15807 & n45534 ;
  assign n45535 = ~n28381 ;
  assign n28387 = n28115 & n45535 ;
  assign n28388 = n45038 & n28387 ;
  assign n28974 = n28388 & n132 ;
  assign n28389 = n28380 | n28381 ;
  assign n45536 = ~n28389 ;
  assign n28983 = n45536 & n132 ;
  assign n28984 = n28115 | n28983 ;
  assign n45537 = ~n28974 ;
  assign n28985 = n45537 & n28984 ;
  assign n45538 = ~n29230 ;
  assign n29246 = n29217 & n45538 ;
  assign n45539 = ~n29246 ;
  assign n29247 = n146 & n45539 ;
  assign n45540 = ~n29247 ;
  assign n29248 = n29233 & n45540 ;
  assign n45541 = ~n29248 ;
  assign n29249 = n16322 & n45541 ;
  assign n29250 = n148 | n29249 ;
  assign n45542 = ~n29250 ;
  assign n29251 = n29237 & n45542 ;
  assign n29252 = n28985 | n29251 ;
  assign n45543 = ~n29239 ;
  assign n29253 = n45543 & n29252 ;
  assign n45544 = ~n29253 ;
  assign n29254 = n149 & n45544 ;
  assign n28415 = n28384 | n28401 ;
  assign n45545 = ~n28415 ;
  assign n28981 = n45545 & n132 ;
  assign n28982 = n28120 | n28981 ;
  assign n28386 = n28120 & n45048 ;
  assign n45546 = ~n28401 ;
  assign n28414 = n28386 & n45546 ;
  assign n29043 = n28414 & n132 ;
  assign n45547 = ~n29043 ;
  assign n29044 = n28982 & n45547 ;
  assign n29240 = n149 | n29239 ;
  assign n45548 = ~n29240 ;
  assign n29255 = n45548 & n29252 ;
  assign n29256 = n29044 | n29255 ;
  assign n45549 = ~n29254 ;
  assign n29257 = n45549 & n29256 ;
  assign n45550 = ~n29257 ;
  assign n29258 = n150 & n45550 ;
  assign n28413 = n28404 | n28405 ;
  assign n45551 = ~n28413 ;
  assign n28976 = n45551 & n132 ;
  assign n28977 = n28071 | n28976 ;
  assign n45552 = ~n28405 ;
  assign n28411 = n28071 & n45552 ;
  assign n28412 = n45054 & n28411 ;
  assign n29055 = n28412 & n132 ;
  assign n45553 = ~n29055 ;
  assign n29056 = n28977 & n45553 ;
  assign n45554 = ~n29249 ;
  assign n29266 = n29237 & n45554 ;
  assign n45555 = ~n29266 ;
  assign n29267 = n148 & n45555 ;
  assign n45556 = ~n29267 ;
  assign n29268 = n29252 & n45556 ;
  assign n45557 = ~n29268 ;
  assign n29269 = n149 & n45557 ;
  assign n29270 = n150 | n29269 ;
  assign n45558 = ~n29270 ;
  assign n29271 = n29256 & n45558 ;
  assign n29272 = n29056 | n29271 ;
  assign n45559 = ~n29258 ;
  assign n29273 = n45559 & n29272 ;
  assign n45560 = ~n29273 ;
  assign n29274 = n151 & n45560 ;
  assign n28439 = n28408 | n28425 ;
  assign n45561 = ~n28439 ;
  assign n28949 = n45561 & n132 ;
  assign n28950 = n28123 | n28949 ;
  assign n28409 = n28123 & n45064 ;
  assign n45562 = ~n28425 ;
  assign n28438 = n28409 & n45562 ;
  assign n28972 = n28438 & n132 ;
  assign n45563 = ~n28972 ;
  assign n28973 = n28950 & n45563 ;
  assign n29259 = n151 | n29258 ;
  assign n45564 = ~n29259 ;
  assign n29275 = n45564 & n29272 ;
  assign n29276 = n28973 | n29275 ;
  assign n45565 = ~n29274 ;
  assign n29277 = n45565 & n29276 ;
  assign n45566 = ~n29277 ;
  assign n29278 = n13079 & n45566 ;
  assign n45567 = ~n28429 ;
  assign n28435 = n28066 & n45567 ;
  assign n28436 = n45070 & n28435 ;
  assign n28923 = n28436 & n28918 ;
  assign n28437 = n28428 | n28429 ;
  assign n45568 = ~n28437 ;
  assign n28962 = n45568 & n132 ;
  assign n28963 = n28066 | n28962 ;
  assign n45569 = ~n28923 ;
  assign n28964 = n45569 & n28963 ;
  assign n45570 = ~n29269 ;
  assign n29286 = n29256 & n45570 ;
  assign n45571 = ~n29286 ;
  assign n29287 = n150 & n45571 ;
  assign n45572 = ~n29287 ;
  assign n29288 = n29272 & n45572 ;
  assign n45573 = ~n29288 ;
  assign n29289 = n13662 & n45573 ;
  assign n29290 = n152 | n29289 ;
  assign n45574 = ~n29290 ;
  assign n29291 = n29276 & n45574 ;
  assign n29292 = n28964 | n29291 ;
  assign n45575 = ~n29278 ;
  assign n29293 = n45575 & n29292 ;
  assign n45576 = ~n29293 ;
  assign n29294 = n153 & n45576 ;
  assign n28434 = n28023 & n45080 ;
  assign n45577 = ~n28449 ;
  assign n28462 = n28434 & n45577 ;
  assign n28960 = n28462 & n132 ;
  assign n28463 = n28432 | n28449 ;
  assign n45578 = ~n28463 ;
  assign n29000 = n45578 & n132 ;
  assign n29001 = n28023 | n29000 ;
  assign n45579 = ~n28960 ;
  assign n29002 = n45579 & n29001 ;
  assign n29279 = n153 | n29278 ;
  assign n45580 = ~n29279 ;
  assign n29295 = n45580 & n29292 ;
  assign n29296 = n29002 | n29295 ;
  assign n45581 = ~n29294 ;
  assign n29297 = n45581 & n29296 ;
  assign n45582 = ~n29297 ;
  assign n29298 = n154 & n45582 ;
  assign n28461 = n28452 | n28453 ;
  assign n45583 = ~n28461 ;
  assign n28955 = n45583 & n132 ;
  assign n28956 = n28046 | n28955 ;
  assign n45584 = ~n28453 ;
  assign n28459 = n28046 & n45584 ;
  assign n28460 = n45086 & n28459 ;
  assign n29007 = n28460 & n132 ;
  assign n45585 = ~n29007 ;
  assign n29008 = n28956 & n45585 ;
  assign n45586 = ~n29289 ;
  assign n29306 = n29276 & n45586 ;
  assign n45587 = ~n29306 ;
  assign n29307 = n152 & n45587 ;
  assign n45588 = ~n29307 ;
  assign n29308 = n29292 & n45588 ;
  assign n45589 = ~n29308 ;
  assign n29309 = n153 & n45589 ;
  assign n29310 = n154 | n29309 ;
  assign n45590 = ~n29310 ;
  assign n29311 = n29296 & n45590 ;
  assign n29312 = n29008 | n29311 ;
  assign n45591 = ~n29298 ;
  assign n29313 = n45591 & n29312 ;
  assign n45592 = ~n29313 ;
  assign n29314 = n155 & n45592 ;
  assign n28458 = n28026 & n45096 ;
  assign n45593 = ~n28473 ;
  assign n28486 = n28458 & n45593 ;
  assign n28952 = n28486 & n132 ;
  assign n28487 = n28456 | n28473 ;
  assign n45594 = ~n28487 ;
  assign n28967 = n45594 & n132 ;
  assign n28968 = n28026 | n28967 ;
  assign n45595 = ~n28952 ;
  assign n28969 = n45595 & n28968 ;
  assign n29299 = n11067 | n29298 ;
  assign n45596 = ~n29299 ;
  assign n29315 = n45596 & n29312 ;
  assign n29316 = n28969 | n29315 ;
  assign n45597 = ~n29314 ;
  assign n29317 = n45597 & n29316 ;
  assign n45598 = ~n29317 ;
  assign n29318 = n10657 & n45598 ;
  assign n28485 = n28476 | n28477 ;
  assign n45599 = ~n28485 ;
  assign n29028 = n45599 & n132 ;
  assign n29029 = n28109 | n29028 ;
  assign n45600 = ~n28477 ;
  assign n28483 = n28109 & n45600 ;
  assign n28484 = n45102 & n28483 ;
  assign n29164 = n28484 & n132 ;
  assign n45601 = ~n29164 ;
  assign n29165 = n29029 & n45601 ;
  assign n45602 = ~n29309 ;
  assign n29326 = n29296 & n45602 ;
  assign n45603 = ~n29326 ;
  assign n29327 = n154 & n45603 ;
  assign n45604 = ~n29327 ;
  assign n29328 = n29312 & n45604 ;
  assign n45605 = ~n29328 ;
  assign n29329 = n11067 & n45605 ;
  assign n29330 = n10657 | n29329 ;
  assign n45606 = ~n29330 ;
  assign n29331 = n29316 & n45606 ;
  assign n29332 = n29165 | n29331 ;
  assign n45607 = ~n29318 ;
  assign n29333 = n45607 & n29332 ;
  assign n45608 = ~n29333 ;
  assign n29334 = n157 & n45608 ;
  assign n28482 = n28057 & n45112 ;
  assign n45609 = ~n28497 ;
  assign n28510 = n28482 & n45609 ;
  assign n28951 = n28510 & n132 ;
  assign n28511 = n28480 | n28497 ;
  assign n45610 = ~n28511 ;
  assign n29061 = n45610 & n132 ;
  assign n29062 = n28057 | n29061 ;
  assign n45611 = ~n28951 ;
  assign n29063 = n45611 & n29062 ;
  assign n29319 = n157 | n29318 ;
  assign n45612 = ~n29319 ;
  assign n29335 = n45612 & n29332 ;
  assign n29336 = n29063 | n29335 ;
  assign n45613 = ~n29334 ;
  assign n29337 = n45613 & n29336 ;
  assign n45614 = ~n29337 ;
  assign n29338 = n158 & n45614 ;
  assign n45615 = ~n28501 ;
  assign n28502 = n28098 & n45615 ;
  assign n28503 = n45118 & n28502 ;
  assign n28948 = n28503 & n132 ;
  assign n28504 = n28500 | n28501 ;
  assign n45616 = ~n28504 ;
  assign n29025 = n45616 & n132 ;
  assign n29026 = n28098 | n29025 ;
  assign n45617 = ~n28948 ;
  assign n29027 = n45617 & n29026 ;
  assign n45618 = ~n29329 ;
  assign n29347 = n29316 & n45618 ;
  assign n45619 = ~n29347 ;
  assign n29348 = n156 & n45619 ;
  assign n45620 = ~n29348 ;
  assign n29349 = n29332 & n45620 ;
  assign n45621 = ~n29349 ;
  assign n29350 = n157 & n45621 ;
  assign n29351 = n158 | n29350 ;
  assign n45622 = ~n29351 ;
  assign n29352 = n29336 & n45622 ;
  assign n29353 = n29027 | n29352 ;
  assign n45623 = ~n29338 ;
  assign n29354 = n45623 & n29353 ;
  assign n45624 = ~n29354 ;
  assign n29355 = n159 & n45624 ;
  assign n28508 = n28008 & n45128 ;
  assign n45625 = ~n28521 ;
  assign n28534 = n28508 & n45625 ;
  assign n28925 = n28534 & n28918 ;
  assign n28535 = n28507 | n28521 ;
  assign n45626 = ~n28535 ;
  assign n28943 = n45626 & n132 ;
  assign n28944 = n28008 | n28943 ;
  assign n45627 = ~n28925 ;
  assign n28945 = n45627 & n28944 ;
  assign n29339 = n8857 | n29338 ;
  assign n45628 = ~n29339 ;
  assign n29356 = n45628 & n29353 ;
  assign n29357 = n28945 | n29356 ;
  assign n45629 = ~n29355 ;
  assign n29358 = n45629 & n29357 ;
  assign n45630 = ~n29358 ;
  assign n29359 = n8534 & n45630 ;
  assign n29360 = n161 | n29359 ;
  assign n45631 = ~n28525 ;
  assign n28531 = n28088 & n45631 ;
  assign n28532 = n45134 & n28531 ;
  assign n28924 = n28532 & n28918 ;
  assign n28533 = n28524 | n28525 ;
  assign n45632 = ~n28533 ;
  assign n29016 = n45632 & n132 ;
  assign n29017 = n28088 | n29016 ;
  assign n45633 = ~n28924 ;
  assign n29018 = n45633 & n29017 ;
  assign n45634 = ~n29350 ;
  assign n29367 = n29336 & n45634 ;
  assign n45635 = ~n29367 ;
  assign n29368 = n158 & n45635 ;
  assign n45636 = ~n29368 ;
  assign n29369 = n29353 & n45636 ;
  assign n45637 = ~n29369 ;
  assign n29370 = n8857 & n45637 ;
  assign n29371 = n160 | n29370 ;
  assign n45638 = ~n29371 ;
  assign n29372 = n29357 & n45638 ;
  assign n29373 = n29018 | n29372 ;
  assign n45639 = ~n29360 ;
  assign n29376 = n45639 & n29373 ;
  assign n29378 = n29156 | n29376 ;
  assign n45640 = ~n29370 ;
  assign n29387 = n29357 & n45640 ;
  assign n45641 = ~n29387 ;
  assign n29388 = n160 & n45641 ;
  assign n45642 = ~n29388 ;
  assign n29389 = n29373 & n45642 ;
  assign n45643 = ~n29389 ;
  assign n29390 = n161 & n45643 ;
  assign n29391 = n162 | n29390 ;
  assign n45644 = ~n29391 ;
  assign n29392 = n29378 & n45644 ;
  assign n29393 = n29042 | n29392 ;
  assign n45645 = ~n29390 ;
  assign n29403 = n29378 & n45645 ;
  assign n45646 = ~n29403 ;
  assign n29404 = n162 & n45646 ;
  assign n45647 = ~n29404 ;
  assign n29405 = n29393 & n45647 ;
  assign n45648 = ~n29405 ;
  assign n29406 = n6889 & n45648 ;
  assign n29407 = n6600 | n29406 ;
  assign n45649 = ~n29359 ;
  assign n29374 = n45649 & n29373 ;
  assign n45650 = ~n29374 ;
  assign n29375 = n161 & n45650 ;
  assign n45651 = ~n29375 ;
  assign n29379 = n45651 & n29378 ;
  assign n45652 = ~n29379 ;
  assign n29380 = n162 & n45652 ;
  assign n29381 = n6889 | n29380 ;
  assign n45653 = ~n29381 ;
  assign n29396 = n45653 & n29393 ;
  assign n28554 = n28034 & n45160 ;
  assign n45654 = ~n28569 ;
  assign n28582 = n28554 & n45654 ;
  assign n29036 = n28582 & n132 ;
  assign n28583 = n28552 | n28569 ;
  assign n45655 = ~n28583 ;
  assign n29408 = n45655 & n132 ;
  assign n29409 = n28034 | n29408 ;
  assign n45656 = ~n29036 ;
  assign n29410 = n45656 & n29409 ;
  assign n29411 = n29396 | n29410 ;
  assign n45657 = ~n29407 ;
  assign n29415 = n45657 & n29411 ;
  assign n29416 = n29024 | n29415 ;
  assign n45658 = ~n29406 ;
  assign n29425 = n45658 & n29411 ;
  assign n45659 = ~n29425 ;
  assign n29426 = n164 & n45659 ;
  assign n45660 = ~n29426 ;
  assign n29427 = n29416 & n45660 ;
  assign n45661 = ~n29427 ;
  assign n29428 = n165 & n45661 ;
  assign n29429 = n166 | n29428 ;
  assign n45662 = ~n29380 ;
  assign n29394 = n45662 & n29393 ;
  assign n45663 = ~n29394 ;
  assign n29395 = n163 & n45663 ;
  assign n45664 = ~n29395 ;
  assign n29412 = n45664 & n29411 ;
  assign n45665 = ~n29412 ;
  assign n29413 = n6600 & n45665 ;
  assign n29414 = n165 | n29413 ;
  assign n45666 = ~n29414 ;
  assign n29419 = n45666 & n29416 ;
  assign n28577 = n28093 & n45176 ;
  assign n45667 = ~n28593 ;
  assign n28606 = n28577 & n45667 ;
  assign n29434 = n28606 & n132 ;
  assign n28607 = n28576 | n28593 ;
  assign n45668 = ~n28607 ;
  assign n29439 = n45668 & n132 ;
  assign n29440 = n28093 | n29439 ;
  assign n45669 = ~n29434 ;
  assign n29441 = n45669 & n29440 ;
  assign n29442 = n29419 | n29441 ;
  assign n45670 = ~n29429 ;
  assign n29446 = n45670 & n29442 ;
  assign n29447 = n29020 | n29446 ;
  assign n45671 = ~n29428 ;
  assign n29456 = n45671 & n29442 ;
  assign n45672 = ~n29456 ;
  assign n29457 = n166 & n45672 ;
  assign n45673 = ~n29457 ;
  assign n29458 = n29447 & n45673 ;
  assign n45674 = ~n29458 ;
  assign n29459 = n5352 & n45674 ;
  assign n29460 = n4934 | n29459 ;
  assign n45675 = ~n29413 ;
  assign n29417 = n45675 & n29416 ;
  assign n45676 = ~n29417 ;
  assign n29418 = n165 & n45676 ;
  assign n45677 = ~n29418 ;
  assign n29443 = n45677 & n29442 ;
  assign n45678 = ~n29443 ;
  assign n29444 = n166 & n45678 ;
  assign n29445 = n5352 | n29444 ;
  assign n45679 = ~n29445 ;
  assign n29450 = n45679 & n29447 ;
  assign n28631 = n28600 | n28617 ;
  assign n45680 = ~n28631 ;
  assign n29003 = n45680 & n132 ;
  assign n29004 = n28126 | n29003 ;
  assign n28601 = n28126 & n45192 ;
  assign n45681 = ~n28617 ;
  assign n28630 = n28601 & n45681 ;
  assign n29462 = n28630 & n132 ;
  assign n45682 = ~n29462 ;
  assign n29463 = n29004 & n45682 ;
  assign n29464 = n29450 | n29463 ;
  assign n45683 = ~n29460 ;
  assign n29468 = n45683 & n29464 ;
  assign n29469 = n29159 | n29468 ;
  assign n45684 = ~n29459 ;
  assign n29478 = n45684 & n29464 ;
  assign n45685 = ~n29478 ;
  assign n29479 = n168 & n45685 ;
  assign n45686 = ~n29479 ;
  assign n29480 = n29469 & n45686 ;
  assign n45687 = ~n29480 ;
  assign n29481 = n169 & n45687 ;
  assign n29482 = n170 | n29481 ;
  assign n45688 = ~n29444 ;
  assign n29448 = n45688 & n29447 ;
  assign n45689 = ~n29448 ;
  assign n29449 = n167 & n45689 ;
  assign n45690 = ~n29449 ;
  assign n29465 = n45690 & n29464 ;
  assign n45691 = ~n29465 ;
  assign n29466 = n4934 & n45691 ;
  assign n29467 = n169 | n29466 ;
  assign n45692 = ~n29467 ;
  assign n29472 = n45692 & n29469 ;
  assign n28654 = n28624 | n28641 ;
  assign n45693 = ~n28654 ;
  assign n28979 = n45693 & n132 ;
  assign n28980 = n28136 | n28979 ;
  assign n28626 = n28136 & n45208 ;
  assign n45694 = ~n28641 ;
  assign n28655 = n28626 & n45694 ;
  assign n29484 = n28655 & n132 ;
  assign n45695 = ~n29484 ;
  assign n29485 = n28980 & n45695 ;
  assign n29486 = n29472 | n29485 ;
  assign n45696 = ~n29482 ;
  assign n29490 = n45696 & n29486 ;
  assign n29491 = n29145 | n29490 ;
  assign n45697 = ~n29481 ;
  assign n29501 = n45697 & n29486 ;
  assign n45698 = ~n29501 ;
  assign n29502 = n170 & n45698 ;
  assign n45699 = ~n29502 ;
  assign n29503 = n29491 & n45699 ;
  assign n45700 = ~n29503 ;
  assign n29504 = n3940 & n45700 ;
  assign n45701 = ~n29466 ;
  assign n29470 = n45701 & n29469 ;
  assign n45702 = ~n29470 ;
  assign n29471 = n169 & n45702 ;
  assign n45703 = ~n29471 ;
  assign n29487 = n45703 & n29486 ;
  assign n45704 = ~n29487 ;
  assign n29488 = n170 & n45704 ;
  assign n29489 = n3940 | n29488 ;
  assign n45705 = ~n29489 ;
  assign n29494 = n45705 & n29491 ;
  assign n28650 = n28095 & n45224 ;
  assign n45706 = ~n28665 ;
  assign n28678 = n28650 & n45706 ;
  assign n29035 = n28678 & n132 ;
  assign n28679 = n28648 | n28665 ;
  assign n45707 = ~n28679 ;
  assign n29506 = n45707 & n132 ;
  assign n29507 = n28095 | n29506 ;
  assign n45708 = ~n29035 ;
  assign n29508 = n45708 & n29507 ;
  assign n29509 = n29494 | n29508 ;
  assign n45709 = ~n29504 ;
  assign n29517 = n45709 & n29509 ;
  assign n45710 = ~n29517 ;
  assign n29518 = n172 & n45710 ;
  assign n29505 = n3631 | n29504 ;
  assign n45711 = ~n29505 ;
  assign n29513 = n45711 & n29509 ;
  assign n28672 = n28668 | n28669 ;
  assign n45712 = ~n28672 ;
  assign n28970 = n45712 & n132 ;
  assign n28971 = n28140 | n28970 ;
  assign n45713 = ~n28669 ;
  assign n28670 = n28140 & n45713 ;
  assign n28671 = n45230 & n28670 ;
  assign n29521 = n28671 & n132 ;
  assign n45714 = ~n29521 ;
  assign n29522 = n28971 & n45714 ;
  assign n29523 = n29513 | n29522 ;
  assign n45715 = ~n29518 ;
  assign n29524 = n45715 & n29523 ;
  assign n45716 = ~n29524 ;
  assign n29525 = n173 & n45716 ;
  assign n29526 = n174 | n29525 ;
  assign n45717 = ~n29488 ;
  assign n29492 = n45717 & n29491 ;
  assign n45718 = ~n29492 ;
  assign n29493 = n171 & n45718 ;
  assign n45719 = ~n29493 ;
  assign n29510 = n45719 & n29509 ;
  assign n45720 = ~n29510 ;
  assign n29511 = n3631 & n45720 ;
  assign n29512 = n173 | n29511 ;
  assign n45721 = ~n29512 ;
  assign n29527 = n45721 & n29523 ;
  assign n28703 = n28675 | n28689 ;
  assign n45722 = ~n28703 ;
  assign n29081 = n45722 & n132 ;
  assign n29082 = n28102 | n29081 ;
  assign n28677 = n28102 & n45240 ;
  assign n45723 = ~n28689 ;
  assign n28702 = n28677 & n45723 ;
  assign n29533 = n28702 & n132 ;
  assign n45724 = ~n29533 ;
  assign n29534 = n29082 & n45724 ;
  assign n29535 = n29527 | n29534 ;
  assign n45725 = ~n29526 ;
  assign n29539 = n45725 & n29535 ;
  assign n29540 = n29065 | n29539 ;
  assign n45726 = ~n29525 ;
  assign n29550 = n45726 & n29535 ;
  assign n45727 = ~n29550 ;
  assign n29551 = n174 & n45727 ;
  assign n45728 = ~n29551 ;
  assign n29552 = n29540 & n45728 ;
  assign n45729 = ~n29552 ;
  assign n29553 = n2753 & n45729 ;
  assign n45730 = ~n29511 ;
  assign n29530 = n45730 & n29523 ;
  assign n45731 = ~n29530 ;
  assign n29531 = n173 & n45731 ;
  assign n45732 = ~n29531 ;
  assign n29536 = n45732 & n29535 ;
  assign n45733 = ~n29536 ;
  assign n29537 = n174 & n45733 ;
  assign n29538 = n2753 | n29537 ;
  assign n45734 = ~n29538 ;
  assign n29543 = n45734 & n29540 ;
  assign n28727 = n28696 | n28713 ;
  assign n45735 = ~n28727 ;
  assign n29066 = n45735 & n132 ;
  assign n29067 = n28147 | n29066 ;
  assign n28698 = n28147 & n45256 ;
  assign n45736 = ~n28713 ;
  assign n28726 = n28698 & n45736 ;
  assign n29555 = n28726 & n132 ;
  assign n45737 = ~n29555 ;
  assign n29556 = n29067 & n45737 ;
  assign n29557 = n29543 | n29556 ;
  assign n45738 = ~n29553 ;
  assign n29565 = n45738 & n29557 ;
  assign n45739 = ~n29565 ;
  assign n29566 = n176 & n45739 ;
  assign n29554 = n2431 | n29553 ;
  assign n45740 = ~n29554 ;
  assign n29561 = n45740 & n29557 ;
  assign n28725 = n28716 | n28717 ;
  assign n45741 = ~n28725 ;
  assign n28992 = n45741 & n132 ;
  assign n28993 = n28154 | n28992 ;
  assign n45742 = ~n28717 ;
  assign n28723 = n28154 & n45742 ;
  assign n28724 = n45262 & n28723 ;
  assign n29567 = n28724 & n132 ;
  assign n45743 = ~n29567 ;
  assign n29568 = n28993 & n45743 ;
  assign n29569 = n29561 | n29568 ;
  assign n45744 = ~n29566 ;
  assign n29570 = n45744 & n29569 ;
  assign n45745 = ~n29570 ;
  assign n29571 = n177 & n45745 ;
  assign n29572 = n178 | n29571 ;
  assign n45746 = ~n29537 ;
  assign n29541 = n45746 & n29540 ;
  assign n45747 = ~n29541 ;
  assign n29542 = n175 & n45747 ;
  assign n45748 = ~n29542 ;
  assign n29558 = n45748 & n29557 ;
  assign n45749 = ~n29558 ;
  assign n29559 = n2431 & n45749 ;
  assign n29560 = n177 | n29559 ;
  assign n45750 = ~n29560 ;
  assign n29573 = n45750 & n29569 ;
  assign n28751 = n28720 | n28737 ;
  assign n45751 = ~n28751 ;
  assign n28965 = n45751 & n132 ;
  assign n28966 = n28157 | n28965 ;
  assign n28722 = n28157 & n45272 ;
  assign n45752 = ~n28737 ;
  assign n28750 = n28722 & n45752 ;
  assign n29579 = n28750 & n132 ;
  assign n45753 = ~n29579 ;
  assign n29580 = n28966 & n45753 ;
  assign n29581 = n29573 | n29580 ;
  assign n45754 = ~n29572 ;
  assign n29585 = n45754 & n29581 ;
  assign n29586 = n29433 | n29585 ;
  assign n45755 = ~n29571 ;
  assign n29596 = n45755 & n29581 ;
  assign n45756 = ~n29596 ;
  assign n29597 = n178 & n45756 ;
  assign n45757 = ~n29597 ;
  assign n29598 = n29586 & n45757 ;
  assign n45758 = ~n29598 ;
  assign n29599 = n1707 & n45758 ;
  assign n45759 = ~n29559 ;
  assign n29576 = n45759 & n29569 ;
  assign n45760 = ~n29576 ;
  assign n29577 = n177 & n45760 ;
  assign n45761 = ~n29577 ;
  assign n29582 = n45761 & n29581 ;
  assign n45762 = ~n29582 ;
  assign n29583 = n178 & n45762 ;
  assign n29584 = n1707 | n29583 ;
  assign n45763 = ~n29584 ;
  assign n29589 = n45763 & n29586 ;
  assign n28746 = n28167 & n45288 ;
  assign n45764 = ~n28761 ;
  assign n28774 = n28746 & n45764 ;
  assign n28975 = n28774 & n132 ;
  assign n28775 = n28744 | n28761 ;
  assign n45765 = ~n28775 ;
  assign n29601 = n45765 & n132 ;
  assign n29602 = n28167 | n29601 ;
  assign n45766 = ~n28975 ;
  assign n29603 = n45766 & n29602 ;
  assign n29604 = n29589 | n29603 ;
  assign n45767 = ~n29599 ;
  assign n29612 = n45767 & n29604 ;
  assign n45768 = ~n29612 ;
  assign n29613 = n180 & n45768 ;
  assign n29600 = n1487 | n29599 ;
  assign n45769 = ~n29600 ;
  assign n29608 = n45769 & n29604 ;
  assign n45770 = ~n28765 ;
  assign n28771 = n28171 & n45770 ;
  assign n28772 = n45294 & n28771 ;
  assign n29614 = n28772 & n132 ;
  assign n28773 = n28764 | n28765 ;
  assign n45771 = ~n28773 ;
  assign n29617 = n45771 & n132 ;
  assign n29618 = n28171 | n29617 ;
  assign n45772 = ~n29614 ;
  assign n29619 = n45772 & n29618 ;
  assign n29620 = n29608 | n29619 ;
  assign n45773 = ~n29613 ;
  assign n29621 = n45773 & n29620 ;
  assign n45774 = ~n29621 ;
  assign n29622 = n181 & n45774 ;
  assign n29623 = n182 | n29622 ;
  assign n45775 = ~n29583 ;
  assign n29587 = n45775 & n29586 ;
  assign n45776 = ~n29587 ;
  assign n29588 = n179 & n45776 ;
  assign n45777 = ~n29588 ;
  assign n29605 = n45777 & n29604 ;
  assign n45778 = ~n29605 ;
  assign n29606 = n1487 & n45778 ;
  assign n29607 = n181 | n29606 ;
  assign n45779 = ~n29607 ;
  assign n29624 = n45779 & n29620 ;
  assign n28770 = n28174 & n45304 ;
  assign n45780 = ~n28785 ;
  assign n28798 = n28770 & n45780 ;
  assign n29630 = n28798 & n132 ;
  assign n28799 = n28768 | n28785 ;
  assign n45781 = ~n28799 ;
  assign n29631 = n45781 & n132 ;
  assign n29632 = n28174 | n29631 ;
  assign n45782 = ~n29630 ;
  assign n29633 = n45782 & n29632 ;
  assign n29634 = n29624 | n29633 ;
  assign n45783 = ~n29623 ;
  assign n29638 = n45783 & n29634 ;
  assign n29639 = n29077 | n29638 ;
  assign n45784 = ~n29622 ;
  assign n29649 = n45784 & n29634 ;
  assign n45785 = ~n29649 ;
  assign n29650 = n182 & n45785 ;
  assign n45786 = ~n29650 ;
  assign n29651 = n29639 & n45786 ;
  assign n45787 = ~n29651 ;
  assign n29652 = n996 & n45787 ;
  assign n45788 = ~n29606 ;
  assign n29627 = n45788 & n29620 ;
  assign n45789 = ~n29627 ;
  assign n29628 = n181 & n45789 ;
  assign n45790 = ~n29628 ;
  assign n29635 = n45790 & n29634 ;
  assign n45791 = ~n29635 ;
  assign n29636 = n182 & n45791 ;
  assign n29637 = n183 | n29636 ;
  assign n45792 = ~n29637 ;
  assign n29642 = n45792 & n29639 ;
  assign n28822 = n28792 | n28809 ;
  assign n45793 = ~n28822 ;
  assign n29615 = n45793 & n132 ;
  assign n29616 = n28180 | n29615 ;
  assign n28794 = n28180 & n45320 ;
  assign n45794 = ~n28809 ;
  assign n28823 = n28794 & n45794 ;
  assign n29654 = n28823 & n132 ;
  assign n45795 = ~n29654 ;
  assign n29655 = n29616 & n45795 ;
  assign n29656 = n29642 | n29655 ;
  assign n45796 = ~n29652 ;
  assign n29664 = n45796 & n29656 ;
  assign n45797 = ~n29664 ;
  assign n29665 = n184 & n45797 ;
  assign n29653 = n838 | n29652 ;
  assign n45798 = ~n29653 ;
  assign n29660 = n45798 & n29656 ;
  assign n45799 = ~n28813 ;
  assign n28819 = n28129 & n45799 ;
  assign n28820 = n45326 & n28819 ;
  assign n29668 = n28820 & n132 ;
  assign n28821 = n28812 | n28813 ;
  assign n45800 = ~n28821 ;
  assign n29669 = n45800 & n132 ;
  assign n29670 = n28129 | n29669 ;
  assign n45801 = ~n29668 ;
  assign n29671 = n45801 & n29670 ;
  assign n29672 = n29660 | n29671 ;
  assign n45802 = ~n29665 ;
  assign n29673 = n45802 & n29672 ;
  assign n45803 = ~n29673 ;
  assign n29674 = n185 & n45803 ;
  assign n45804 = ~n29636 ;
  assign n29640 = n45804 & n29639 ;
  assign n45805 = ~n29640 ;
  assign n29641 = n183 & n45805 ;
  assign n45806 = ~n29641 ;
  assign n29657 = n45806 & n29656 ;
  assign n45807 = ~n29657 ;
  assign n29658 = n838 & n45807 ;
  assign n29659 = n185 | n29658 ;
  assign n45808 = ~n29659 ;
  assign n29676 = n45808 & n29672 ;
  assign n28818 = n28184 & n45336 ;
  assign n45809 = ~n28833 ;
  assign n28846 = n28818 & n45809 ;
  assign n29083 = n28846 & n132 ;
  assign n28847 = n28816 | n28833 ;
  assign n45810 = ~n28847 ;
  assign n29686 = n45810 & n132 ;
  assign n29687 = n28184 | n29686 ;
  assign n45811 = ~n29083 ;
  assign n29688 = n45811 & n29687 ;
  assign n29689 = n29676 | n29688 ;
  assign n45812 = ~n29674 ;
  assign n29697 = n45812 & n29689 ;
  assign n45813 = ~n29697 ;
  assign n29698 = n186 & n45813 ;
  assign n29675 = n186 | n29674 ;
  assign n45814 = ~n29675 ;
  assign n29693 = n45814 & n29689 ;
  assign n28845 = n28836 | n28837 ;
  assign n45815 = ~n28845 ;
  assign n29152 = n45815 & n132 ;
  assign n29153 = n28190 | n29152 ;
  assign n45816 = ~n28837 ;
  assign n28843 = n28190 & n45816 ;
  assign n28844 = n45342 & n28843 ;
  assign n29699 = n28844 & n132 ;
  assign n45817 = ~n29699 ;
  assign n29700 = n29153 & n45817 ;
  assign n29701 = n29693 | n29700 ;
  assign n45818 = ~n29698 ;
  assign n29702 = n45818 & n29701 ;
  assign n45819 = ~n29702 ;
  assign n29703 = n528 & n45819 ;
  assign n29704 = n413 | n29703 ;
  assign n28841 = n28188 & n45352 ;
  assign n45820 = ~n28857 ;
  assign n28870 = n28841 & n45820 ;
  assign n28926 = n28870 & n28918 ;
  assign n28871 = n28840 | n28857 ;
  assign n45821 = ~n28871 ;
  assign n29030 = n45821 & n132 ;
  assign n29031 = n28188 | n29030 ;
  assign n45822 = ~n28926 ;
  assign n29032 = n45822 & n29031 ;
  assign n45823 = ~n29658 ;
  assign n29679 = n45823 & n29672 ;
  assign n45824 = ~n29679 ;
  assign n29680 = n185 & n45824 ;
  assign n45825 = ~n29680 ;
  assign n29690 = n45825 & n29689 ;
  assign n45826 = ~n29690 ;
  assign n29691 = n186 & n45826 ;
  assign n29692 = n528 | n29691 ;
  assign n45827 = ~n29692 ;
  assign n29706 = n45827 & n29701 ;
  assign n29707 = n29032 | n29706 ;
  assign n45828 = ~n29704 ;
  assign n29710 = n45828 & n29707 ;
  assign n29711 = n29683 | n29710 ;
  assign n45829 = ~n29691 ;
  assign n29718 = n45829 & n29701 ;
  assign n45830 = ~n29718 ;
  assign n29719 = n187 & n45830 ;
  assign n45831 = ~n29719 ;
  assign n29722 = n29707 & n45831 ;
  assign n45832 = ~n29722 ;
  assign n29723 = n413 & n45832 ;
  assign n45833 = ~n29723 ;
  assign n29725 = n29711 & n45833 ;
  assign n45834 = ~n29725 ;
  assign n29726 = n189 & n45834 ;
  assign n28894 = n28864 | n28881 ;
  assign n45835 = ~n28894 ;
  assign n28953 = n45835 & n132 ;
  assign n28954 = n28193 | n28953 ;
  assign n28866 = n28193 & n45368 ;
  assign n45836 = ~n28881 ;
  assign n28893 = n28866 & n45836 ;
  assign n29666 = n28893 & n132 ;
  assign n45837 = ~n29666 ;
  assign n29667 = n28954 & n45837 ;
  assign n29724 = n189 | n29723 ;
  assign n45838 = ~n29724 ;
  assign n29727 = n29711 & n45838 ;
  assign n29728 = n29667 | n29727 ;
  assign n45839 = ~n29726 ;
  assign n29730 = n45839 & n29728 ;
  assign n45840 = ~n29730 ;
  assign n29731 = n190 & n45840 ;
  assign n45841 = ~n29703 ;
  assign n29708 = n45841 & n29707 ;
  assign n45842 = ~n29708 ;
  assign n29709 = n188 & n45842 ;
  assign n45843 = ~n29709 ;
  assign n29712 = n45843 & n29711 ;
  assign n45844 = ~n29712 ;
  assign n29713 = n189 & n45844 ;
  assign n29714 = n190 | n29713 ;
  assign n45845 = ~n29714 ;
  assign n29729 = n45845 & n29728 ;
  assign n45846 = ~n28885 ;
  assign n28892 = n28197 & n45846 ;
  assign n45847 = ~n28902 ;
  assign n29750 = n28892 & n45847 ;
  assign n29751 = n132 & n29750 ;
  assign n29752 = n28885 | n28902 ;
  assign n45848 = ~n29752 ;
  assign n29753 = n132 & n45848 ;
  assign n29754 = n28197 | n29753 ;
  assign n45849 = ~n29751 ;
  assign n29755 = n45849 & n29754 ;
  assign n29758 = n29729 | n29755 ;
  assign n45850 = ~n29731 ;
  assign n29759 = n45850 & n29758 ;
  assign n45851 = ~n29759 ;
  assign n29760 = n191 & n45851 ;
  assign n29733 = n191 | n29731 ;
  assign n45852 = ~n29733 ;
  assign n29763 = n45852 & n29758 ;
  assign n30007 = n29760 | n29763 ;
  assign n28932 = n28207 | n28912 ;
  assign n45853 = ~n28932 ;
  assign n29684 = n45853 & n132 ;
  assign n29685 = n28916 | n29684 ;
  assign n45854 = ~n28934 ;
  assign n29742 = n28256 & n45854 ;
  assign n29743 = n45391 & n29742 ;
  assign n29744 = n28918 & n29743 ;
  assign n29745 = n28911 | n28934 ;
  assign n45855 = ~n29745 ;
  assign n29746 = n28918 & n45855 ;
  assign n29747 = n28256 | n29746 ;
  assign n45856 = ~n29744 ;
  assign n29748 = n45856 & n29747 ;
  assign n29749 = n29685 | n29748 ;
  assign n29734 = n287 | n29731 ;
  assign n45857 = ~n29734 ;
  assign n30008 = n45857 & n29758 ;
  assign n30009 = n29741 | n30008 ;
  assign n45858 = ~n29760 ;
  assign n30010 = n45858 & n30009 ;
  assign n30011 = n29749 | n30010 ;
  assign n30012 = n31336 & n30011 ;
  assign n28933 = n192 & n28932 ;
  assign n45859 = ~n28207 ;
  assign n29435 = n45859 & n132 ;
  assign n45860 = ~n29435 ;
  assign n29436 = n28912 & n45860 ;
  assign n45861 = ~n29436 ;
  assign n29437 = n28933 & n45861 ;
  assign n29762 = n29748 & n45858 ;
  assign n30013 = n29762 & n30009 ;
  assign n30014 = n29437 | n30013 ;
  assign n30015 = n30012 | n30014 ;
  assign n45862 = ~n30007 ;
  assign n30035 = n45862 & n30015 ;
  assign n30036 = n29741 | n30035 ;
  assign n29761 = n29741 & n45858 ;
  assign n45863 = ~n29763 ;
  assign n30006 = n29761 & n45863 ;
  assign n30037 = n30006 & n30015 ;
  assign n45864 = ~n30037 ;
  assign n30038 = n30036 & n45864 ;
  assign n29764 = n29741 | n29763 ;
  assign n29765 = n45858 & n29764 ;
  assign n29766 = n29749 | n29765 ;
  assign n29767 = n31336 & n29766 ;
  assign n29768 = n29762 & n29764 ;
  assign n29769 = n29437 | n29768 ;
  assign n131 = n29767 | n29769 ;
  assign n45865 = ~x4 ;
  assign n29792 = n45865 & n131 ;
  assign n45866 = ~n29792 ;
  assign n29793 = x5 & n45866 ;
  assign n45867 = ~n263 ;
  assign n29852 = n45867 & n131 ;
  assign n29876 = n29793 | n29852 ;
  assign n266 = x2 | x3 ;
  assign n268 = x4 | n266 ;
  assign n28228 = n268 & n45437 ;
  assign n28930 = n28228 & n45438 ;
  assign n28931 = n45439 & n28930 ;
  assign n29863 = x4 & n131 ;
  assign n45868 = ~n29863 ;
  assign n29900 = n28931 & n45868 ;
  assign n29901 = n29876 | n29900 ;
  assign n267 = n45865 & n266 ;
  assign n45869 = ~n30015 ;
  assign n30016 = x4 & n45869 ;
  assign n30017 = n267 | n30016 ;
  assign n45870 = ~n30017 ;
  assign n30018 = n28918 & n45870 ;
  assign n45871 = ~n30018 ;
  assign n30019 = n29901 & n45871 ;
  assign n45872 = ~n30019 ;
  assign n30020 = n133 & n45872 ;
  assign n29864 = n268 & n45868 ;
  assign n45873 = ~n29864 ;
  assign n29865 = n132 & n45873 ;
  assign n29866 = n133 | n29865 ;
  assign n45874 = ~n29866 ;
  assign n29902 = n45874 & n29901 ;
  assign n45875 = ~n29437 ;
  assign n29438 = n28918 & n45875 ;
  assign n45876 = ~n30013 ;
  assign n30041 = n29438 & n45876 ;
  assign n45877 = ~n30012 ;
  assign n30042 = n45877 & n30041 ;
  assign n30043 = n29852 | n30042 ;
  assign n30044 = x6 & n30043 ;
  assign n30045 = x6 | n30042 ;
  assign n30046 = n29852 | n30045 ;
  assign n45878 = ~n30044 ;
  assign n30047 = n45878 & n30046 ;
  assign n30048 = n29902 | n30047 ;
  assign n45879 = ~n30020 ;
  assign n30049 = n45879 & n30048 ;
  assign n45880 = ~n30049 ;
  assign n30050 = n134 & n45880 ;
  assign n29099 = n28921 | n29087 ;
  assign n45881 = ~n29099 ;
  assign n29100 = n29086 & n45881 ;
  assign n29838 = n29100 & n131 ;
  assign n29882 = n45881 & n131 ;
  assign n29883 = n29086 | n29882 ;
  assign n45882 = ~n29838 ;
  assign n29884 = n45882 & n29883 ;
  assign n45883 = ~n29865 ;
  assign n29903 = n45883 & n29901 ;
  assign n45884 = ~n29903 ;
  assign n29904 = n133 & n45884 ;
  assign n29905 = n134 | n29904 ;
  assign n30024 = n133 | n30018 ;
  assign n45885 = ~n30024 ;
  assign n30025 = n29901 & n45885 ;
  assign n30055 = n30025 | n30047 ;
  assign n45886 = ~n29905 ;
  assign n30056 = n45886 & n30055 ;
  assign n30057 = n29884 | n30056 ;
  assign n45887 = ~n30050 ;
  assign n30058 = n45887 & n30057 ;
  assign n45888 = ~n30058 ;
  assign n30059 = n26442 & n45888 ;
  assign n45889 = ~n29101 ;
  assign n29137 = n29073 & n45889 ;
  assign n29138 = n45443 & n29137 ;
  assign n29828 = n29138 & n131 ;
  assign n29139 = n29090 | n29101 ;
  assign n45890 = ~n29139 ;
  assign n29853 = n45890 & n131 ;
  assign n29854 = n29073 | n29853 ;
  assign n45891 = ~n29828 ;
  assign n29855 = n45891 & n29854 ;
  assign n30052 = n26442 | n30050 ;
  assign n45892 = ~n30052 ;
  assign n30061 = n45892 & n30057 ;
  assign n30062 = n29855 | n30061 ;
  assign n45893 = ~n30059 ;
  assign n30063 = n45893 & n30062 ;
  assign n45894 = ~n30063 ;
  assign n30064 = n136 & n45894 ;
  assign n29096 = n29070 & n45449 ;
  assign n45895 = ~n29103 ;
  assign n29104 = n29096 & n45895 ;
  assign n29832 = n29104 & n131 ;
  assign n29105 = n29095 | n29103 ;
  assign n45896 = ~n29105 ;
  assign n29844 = n45896 & n131 ;
  assign n29845 = n29070 | n29844 ;
  assign n45897 = ~n29832 ;
  assign n29846 = n45897 & n29845 ;
  assign n30060 = n136 | n30059 ;
  assign n45898 = ~n30060 ;
  assign n30065 = n45898 & n30062 ;
  assign n30066 = n29846 | n30065 ;
  assign n45899 = ~n30064 ;
  assign n30067 = n45899 & n30066 ;
  assign n45900 = ~n30067 ;
  assign n30068 = n137 & n45900 ;
  assign n29136 = n29108 | n29110 ;
  assign n45901 = ~n29136 ;
  assign n29871 = n45901 & n131 ;
  assign n29872 = n29080 | n29871 ;
  assign n45902 = ~n29110 ;
  assign n29134 = n29080 & n45902 ;
  assign n29135 = n45455 & n29134 ;
  assign n29894 = n29135 & n131 ;
  assign n45903 = ~n29894 ;
  assign n29895 = n29872 & n45903 ;
  assign n30021 = n134 | n30020 ;
  assign n45904 = ~n30021 ;
  assign n30074 = n45904 & n30055 ;
  assign n30075 = n29884 | n30074 ;
  assign n30076 = n45887 & n30075 ;
  assign n45905 = ~n30076 ;
  assign n30077 = n135 & n45905 ;
  assign n30078 = n45892 & n30075 ;
  assign n30079 = n29855 | n30078 ;
  assign n45906 = ~n30077 ;
  assign n30080 = n45906 & n30079 ;
  assign n45907 = ~n30080 ;
  assign n30081 = n25517 & n45907 ;
  assign n30082 = n137 | n30081 ;
  assign n45908 = ~n30082 ;
  assign n30083 = n30066 & n45908 ;
  assign n30084 = n29895 | n30083 ;
  assign n45909 = ~n30068 ;
  assign n30085 = n45909 & n30084 ;
  assign n45910 = ~n30085 ;
  assign n30086 = n138 & n45910 ;
  assign n29115 = n29013 & n45461 ;
  assign n45911 = ~n29116 ;
  assign n29132 = n29115 & n45911 ;
  assign n29887 = n29132 & n131 ;
  assign n29133 = n29113 | n29116 ;
  assign n45912 = ~n29133 ;
  assign n29890 = n45912 & n131 ;
  assign n29891 = n29013 | n29890 ;
  assign n45913 = ~n29887 ;
  assign n29892 = n45913 & n29891 ;
  assign n30069 = n138 | n30068 ;
  assign n45914 = ~n30069 ;
  assign n30087 = n45914 & n30084 ;
  assign n30088 = n29892 | n30087 ;
  assign n45915 = ~n30086 ;
  assign n30089 = n45915 & n30088 ;
  assign n45916 = ~n30089 ;
  assign n30090 = n22661 & n45916 ;
  assign n29131 = n29119 | n29120 ;
  assign n45917 = ~n29131 ;
  assign n29888 = n45917 & n131 ;
  assign n29889 = n28990 | n29888 ;
  assign n45918 = ~n29120 ;
  assign n29129 = n28990 & n45918 ;
  assign n29130 = n45467 & n29129 ;
  assign n30027 = n29130 & n30015 ;
  assign n45919 = ~n30027 ;
  assign n30028 = n29889 & n45919 ;
  assign n30098 = n45898 & n30079 ;
  assign n30099 = n29846 | n30098 ;
  assign n45920 = ~n30081 ;
  assign n30100 = n45920 & n30099 ;
  assign n45921 = ~n30100 ;
  assign n30101 = n137 & n45921 ;
  assign n30102 = n45908 & n30099 ;
  assign n30103 = n29895 | n30102 ;
  assign n45922 = ~n30101 ;
  assign n30104 = n45922 & n30103 ;
  assign n45923 = ~n30104 ;
  assign n30105 = n138 & n45923 ;
  assign n30106 = n139 | n30105 ;
  assign n45924 = ~n30106 ;
  assign n30107 = n30088 & n45924 ;
  assign n30108 = n30028 | n30107 ;
  assign n45925 = ~n30090 ;
  assign n30109 = n45925 & n30108 ;
  assign n45926 = ~n30109 ;
  assign n30110 = n140 & n45926 ;
  assign n29128 = n29123 | n29126 ;
  assign n45927 = ~n29128 ;
  assign n29786 = n45927 & n131 ;
  assign n29787 = n29167 | n29786 ;
  assign n29184 = n45490 & n29167 ;
  assign n45928 = ~n29126 ;
  assign n29185 = n45928 & n29184 ;
  assign n29908 = n29185 & n131 ;
  assign n45929 = ~n29908 ;
  assign n29909 = n29787 & n45929 ;
  assign n30091 = n140 | n30090 ;
  assign n45930 = ~n30091 ;
  assign n30111 = n45930 & n30108 ;
  assign n30112 = n29909 | n30111 ;
  assign n45931 = ~n30110 ;
  assign n30113 = n45931 & n30112 ;
  assign n45932 = ~n30113 ;
  assign n30114 = n141 & n45932 ;
  assign n29183 = n29170 | n29172 ;
  assign n45933 = ~n29183 ;
  assign n29910 = n45933 & n131 ;
  assign n29911 = n29015 | n29910 ;
  assign n45934 = ~n29172 ;
  assign n29181 = n29015 & n45934 ;
  assign n29182 = n45479 & n29181 ;
  assign n29912 = n29182 & n131 ;
  assign n45935 = ~n29912 ;
  assign n29913 = n29911 & n45935 ;
  assign n30122 = n45914 & n30103 ;
  assign n30123 = n29892 | n30122 ;
  assign n45936 = ~n30105 ;
  assign n30124 = n45936 & n30123 ;
  assign n45937 = ~n30124 ;
  assign n30125 = n139 & n45937 ;
  assign n30126 = n45924 & n30123 ;
  assign n30127 = n30028 | n30126 ;
  assign n45938 = ~n30125 ;
  assign n30128 = n45938 & n30127 ;
  assign n45939 = ~n30128 ;
  assign n30129 = n22030 & n45939 ;
  assign n30130 = n141 | n30129 ;
  assign n45940 = ~n30130 ;
  assign n30131 = n30112 & n45940 ;
  assign n30132 = n29913 | n30131 ;
  assign n45941 = ~n30114 ;
  assign n30133 = n45941 & n30132 ;
  assign n45942 = ~n30133 ;
  assign n30134 = n142 & n45942 ;
  assign n29206 = n29176 | n29189 ;
  assign n45943 = ~n29206 ;
  assign n29898 = n45943 & n131 ;
  assign n29899 = n29148 | n29898 ;
  assign n29204 = n29148 & n45506 ;
  assign n45944 = ~n29176 ;
  assign n29205 = n45944 & n29204 ;
  assign n29915 = n29205 & n131 ;
  assign n45945 = ~n29915 ;
  assign n29916 = n29899 & n45945 ;
  assign n30115 = n142 | n30114 ;
  assign n45946 = ~n30115 ;
  assign n30135 = n45946 & n30132 ;
  assign n30136 = n29916 | n30135 ;
  assign n45947 = ~n30134 ;
  assign n30137 = n45947 & n30136 ;
  assign n45948 = ~n30137 ;
  assign n30138 = n19362 & n45948 ;
  assign n45949 = ~n29191 ;
  assign n29201 = n29151 & n45949 ;
  assign n29202 = n45495 & n29201 ;
  assign n29842 = n29202 & n131 ;
  assign n29203 = n29179 | n29191 ;
  assign n45950 = ~n29203 ;
  assign n29917 = n45950 & n131 ;
  assign n29918 = n29151 | n29917 ;
  assign n45951 = ~n29842 ;
  assign n29919 = n45951 & n29918 ;
  assign n30146 = n45930 & n30127 ;
  assign n30147 = n29909 | n30146 ;
  assign n45952 = ~n30129 ;
  assign n30148 = n45952 & n30147 ;
  assign n45953 = ~n30148 ;
  assign n30149 = n141 & n45953 ;
  assign n30150 = n45940 & n30147 ;
  assign n30151 = n29913 | n30150 ;
  assign n45954 = ~n30149 ;
  assign n30152 = n45954 & n30151 ;
  assign n45955 = ~n30152 ;
  assign n30153 = n142 & n45955 ;
  assign n30154 = n143 | n30153 ;
  assign n45956 = ~n30154 ;
  assign n30155 = n30136 & n45956 ;
  assign n30156 = n29919 | n30155 ;
  assign n45957 = ~n30138 ;
  assign n30157 = n45957 & n30156 ;
  assign n45958 = ~n30157 ;
  assign n30158 = n144 & n45958 ;
  assign n29200 = n29194 | n29195 ;
  assign n45959 = ~n29200 ;
  assign n29794 = n45959 & n131 ;
  assign n29795 = n29060 | n29794 ;
  assign n29225 = n29060 & n45522 ;
  assign n45960 = ~n29195 ;
  assign n29226 = n45960 & n29225 ;
  assign n30031 = n29226 & n30015 ;
  assign n45961 = ~n30031 ;
  assign n30032 = n29795 & n45961 ;
  assign n30139 = n144 | n30138 ;
  assign n45962 = ~n30139 ;
  assign n30159 = n45962 & n30156 ;
  assign n30160 = n30032 | n30159 ;
  assign n45963 = ~n30158 ;
  assign n30161 = n45963 & n30160 ;
  assign n45964 = ~n30161 ;
  assign n30162 = n145 & n45964 ;
  assign n29224 = n29198 | n29212 ;
  assign n45965 = ~n29224 ;
  assign n29834 = n45965 & n131 ;
  assign n29835 = n29163 | n29834 ;
  assign n45966 = ~n29212 ;
  assign n29222 = n29163 & n45966 ;
  assign n29223 = n45511 & n29222 ;
  assign n29906 = n29223 & n131 ;
  assign n45967 = ~n29906 ;
  assign n29907 = n29835 & n45967 ;
  assign n30170 = n45946 & n30151 ;
  assign n30171 = n29916 | n30170 ;
  assign n45968 = ~n30153 ;
  assign n30172 = n45968 & n30171 ;
  assign n45969 = ~n30172 ;
  assign n30173 = n143 & n45969 ;
  assign n30174 = n45956 & n30171 ;
  assign n30175 = n29919 | n30174 ;
  assign n45970 = ~n30173 ;
  assign n30176 = n45970 & n30175 ;
  assign n45971 = ~n30176 ;
  assign n30177 = n18797 & n45971 ;
  assign n30178 = n145 | n30177 ;
  assign n45972 = ~n30178 ;
  assign n30179 = n30160 & n45972 ;
  assign n30180 = n29907 | n30179 ;
  assign n45973 = ~n30162 ;
  assign n30181 = n45973 & n30180 ;
  assign n45974 = ~n30181 ;
  assign n30182 = n146 & n45974 ;
  assign n29244 = n29039 & n45538 ;
  assign n45975 = ~n29216 ;
  assign n29245 = n45975 & n29244 ;
  assign n29851 = n29245 & n131 ;
  assign n29221 = n29215 | n29216 ;
  assign n45976 = ~n29221 ;
  assign n29877 = n45976 & n131 ;
  assign n29878 = n29039 | n29877 ;
  assign n45977 = ~n29851 ;
  assign n29879 = n45977 & n29878 ;
  assign n30163 = n146 | n30162 ;
  assign n45978 = ~n30163 ;
  assign n30183 = n45978 & n30180 ;
  assign n30184 = n29879 | n30183 ;
  assign n45979 = ~n30182 ;
  assign n30185 = n45979 & n30184 ;
  assign n45980 = ~n30185 ;
  assign n30186 = n16322 & n45980 ;
  assign n45981 = ~n29232 ;
  assign n29241 = n29141 & n45981 ;
  assign n29242 = n45527 & n29241 ;
  assign n29782 = n29242 & n131 ;
  assign n29243 = n29219 | n29232 ;
  assign n45982 = ~n29243 ;
  assign n29822 = n45982 & n131 ;
  assign n29823 = n29141 | n29822 ;
  assign n45983 = ~n29782 ;
  assign n29824 = n45983 & n29823 ;
  assign n30194 = n45962 & n30175 ;
  assign n30195 = n30032 | n30194 ;
  assign n45984 = ~n30177 ;
  assign n30196 = n45984 & n30195 ;
  assign n45985 = ~n30196 ;
  assign n30197 = n145 & n45985 ;
  assign n30198 = n45972 & n30195 ;
  assign n30199 = n29907 | n30198 ;
  assign n45986 = ~n30197 ;
  assign n30200 = n45986 & n30199 ;
  assign n45987 = ~n30200 ;
  assign n30201 = n146 & n45987 ;
  assign n30202 = n147 | n30201 ;
  assign n45988 = ~n30202 ;
  assign n30203 = n30184 & n45988 ;
  assign n30204 = n29824 | n30203 ;
  assign n45989 = ~n30186 ;
  assign n30205 = n45989 & n30204 ;
  assign n45990 = ~n30205 ;
  assign n30206 = n148 & n45990 ;
  assign n29263 = n29048 & n45554 ;
  assign n45991 = ~n29236 ;
  assign n29264 = n45991 & n29263 ;
  assign n29817 = n29264 & n131 ;
  assign n29265 = n29236 | n29249 ;
  assign n45992 = ~n29265 ;
  assign n29839 = n45992 & n131 ;
  assign n29840 = n29048 | n29839 ;
  assign n45993 = ~n29817 ;
  assign n29841 = n45993 & n29840 ;
  assign n30187 = n148 | n30186 ;
  assign n45994 = ~n30187 ;
  assign n30207 = n45994 & n30204 ;
  assign n30208 = n29841 | n30207 ;
  assign n45995 = ~n30206 ;
  assign n30209 = n45995 & n30208 ;
  assign n45996 = ~n30209 ;
  assign n30210 = n149 & n45996 ;
  assign n29262 = n29239 | n29251 ;
  assign n45997 = ~n29262 ;
  assign n29811 = n45997 & n131 ;
  assign n29812 = n28985 | n29811 ;
  assign n45998 = ~n29251 ;
  assign n29260 = n28985 & n45998 ;
  assign n29261 = n45543 & n29260 ;
  assign n29813 = n29261 & n131 ;
  assign n45999 = ~n29813 ;
  assign n29814 = n29812 & n45999 ;
  assign n30218 = n45978 & n30199 ;
  assign n30219 = n29879 | n30218 ;
  assign n46000 = ~n30201 ;
  assign n30220 = n46000 & n30219 ;
  assign n46001 = ~n30220 ;
  assign n30221 = n147 & n46001 ;
  assign n30222 = n45988 & n30219 ;
  assign n30223 = n29824 | n30222 ;
  assign n46002 = ~n30221 ;
  assign n30224 = n46002 & n30223 ;
  assign n46003 = ~n30224 ;
  assign n30225 = n15807 & n46003 ;
  assign n30226 = n149 | n30225 ;
  assign n46004 = ~n30226 ;
  assign n30227 = n30208 & n46004 ;
  assign n30228 = n29814 | n30227 ;
  assign n46005 = ~n30210 ;
  assign n30229 = n46005 & n30228 ;
  assign n46006 = ~n30229 ;
  assign n30230 = n150 & n46006 ;
  assign n29285 = n29255 | n29269 ;
  assign n46007 = ~n29285 ;
  assign n29805 = n46007 & n131 ;
  assign n29806 = n29044 | n29805 ;
  assign n29283 = n29044 & n45570 ;
  assign n46008 = ~n29255 ;
  assign n29284 = n46008 & n29283 ;
  assign n29859 = n29284 & n131 ;
  assign n46009 = ~n29859 ;
  assign n29860 = n29806 & n46009 ;
  assign n30211 = n150 | n30210 ;
  assign n46010 = ~n30211 ;
  assign n30231 = n46010 & n30228 ;
  assign n30232 = n29860 | n30231 ;
  assign n46011 = ~n30230 ;
  assign n30233 = n46011 & n30232 ;
  assign n46012 = ~n30233 ;
  assign n30234 = n13662 & n46012 ;
  assign n46013 = ~n29271 ;
  assign n29280 = n29056 & n46013 ;
  assign n29281 = n45559 & n29280 ;
  assign n29773 = n29281 & n131 ;
  assign n29282 = n29258 | n29271 ;
  assign n46014 = ~n29282 ;
  assign n29825 = n46014 & n131 ;
  assign n29826 = n29056 | n29825 ;
  assign n46015 = ~n29773 ;
  assign n29827 = n46015 & n29826 ;
  assign n30242 = n45994 & n30223 ;
  assign n30243 = n29841 | n30242 ;
  assign n46016 = ~n30225 ;
  assign n30244 = n46016 & n30243 ;
  assign n46017 = ~n30244 ;
  assign n30245 = n149 & n46017 ;
  assign n30246 = n46004 & n30243 ;
  assign n30247 = n29814 | n30246 ;
  assign n46018 = ~n30245 ;
  assign n30248 = n46018 & n30247 ;
  assign n46019 = ~n30248 ;
  assign n30249 = n150 & n46019 ;
  assign n30250 = n151 | n30249 ;
  assign n46020 = ~n30250 ;
  assign n30251 = n30232 & n46020 ;
  assign n30252 = n29827 | n30251 ;
  assign n46021 = ~n30234 ;
  assign n30253 = n46021 & n30252 ;
  assign n46022 = ~n30253 ;
  assign n30254 = n152 & n46022 ;
  assign n29305 = n29275 | n29289 ;
  assign n46023 = ~n29305 ;
  assign n29796 = n46023 & n131 ;
  assign n29797 = n28973 | n29796 ;
  assign n29303 = n28973 & n45586 ;
  assign n46024 = ~n29275 ;
  assign n29304 = n46024 & n29303 ;
  assign n29801 = n29304 & n131 ;
  assign n46025 = ~n29801 ;
  assign n29802 = n29797 & n46025 ;
  assign n30235 = n152 | n30234 ;
  assign n46026 = ~n30235 ;
  assign n30255 = n46026 & n30252 ;
  assign n30256 = n29802 | n30255 ;
  assign n46027 = ~n30254 ;
  assign n30257 = n46027 & n30256 ;
  assign n46028 = ~n30257 ;
  assign n30258 = n153 & n46028 ;
  assign n29302 = n29278 | n29291 ;
  assign n46029 = ~n29302 ;
  assign n29819 = n46029 & n131 ;
  assign n29820 = n28964 | n29819 ;
  assign n46030 = ~n29291 ;
  assign n29300 = n28964 & n46030 ;
  assign n29301 = n45575 & n29300 ;
  assign n29869 = n29301 & n131 ;
  assign n46031 = ~n29869 ;
  assign n29870 = n29820 & n46031 ;
  assign n30266 = n46010 & n30247 ;
  assign n30267 = n29860 | n30266 ;
  assign n46032 = ~n30249 ;
  assign n30268 = n46032 & n30267 ;
  assign n46033 = ~n30268 ;
  assign n30269 = n151 & n46033 ;
  assign n30270 = n46020 & n30267 ;
  assign n30271 = n29827 | n30270 ;
  assign n46034 = ~n30269 ;
  assign n30272 = n46034 & n30271 ;
  assign n46035 = ~n30272 ;
  assign n30273 = n13079 & n46035 ;
  assign n30274 = n153 | n30273 ;
  assign n46036 = ~n30274 ;
  assign n30275 = n30256 & n46036 ;
  assign n30276 = n29870 | n30275 ;
  assign n46037 = ~n30258 ;
  assign n30277 = n46037 & n30276 ;
  assign n46038 = ~n30277 ;
  assign n30278 = n154 & n46038 ;
  assign n29323 = n29002 & n45602 ;
  assign n46039 = ~n29295 ;
  assign n29324 = n46039 & n29323 ;
  assign n29785 = n29324 & n131 ;
  assign n29325 = n29295 | n29309 ;
  assign n46040 = ~n29325 ;
  assign n29798 = n46040 & n131 ;
  assign n29799 = n29002 | n29798 ;
  assign n46041 = ~n29785 ;
  assign n29800 = n46041 & n29799 ;
  assign n30259 = n154 | n30258 ;
  assign n46042 = ~n30259 ;
  assign n30279 = n46042 & n30276 ;
  assign n30280 = n29800 | n30279 ;
  assign n46043 = ~n30278 ;
  assign n30281 = n46043 & n30280 ;
  assign n46044 = ~n30281 ;
  assign n30282 = n11067 & n46044 ;
  assign n29322 = n29298 | n29311 ;
  assign n46045 = ~n29322 ;
  assign n29790 = n46045 & n131 ;
  assign n29791 = n29008 | n29790 ;
  assign n46046 = ~n29311 ;
  assign n29320 = n29008 & n46046 ;
  assign n29321 = n45591 & n29320 ;
  assign n29809 = n29321 & n131 ;
  assign n46047 = ~n29809 ;
  assign n29810 = n29791 & n46047 ;
  assign n30290 = n46026 & n30271 ;
  assign n30291 = n29802 | n30290 ;
  assign n46048 = ~n30273 ;
  assign n30292 = n46048 & n30291 ;
  assign n46049 = ~n30292 ;
  assign n30293 = n153 & n46049 ;
  assign n30294 = n46036 & n30291 ;
  assign n30295 = n29870 | n30294 ;
  assign n46050 = ~n30293 ;
  assign n30296 = n46050 & n30295 ;
  assign n46051 = ~n30296 ;
  assign n30297 = n154 & n46051 ;
  assign n30298 = n11067 | n30297 ;
  assign n46052 = ~n30298 ;
  assign n30299 = n30280 & n46052 ;
  assign n30300 = n29810 | n30299 ;
  assign n46053 = ~n30282 ;
  assign n30301 = n46053 & n30300 ;
  assign n46054 = ~n30301 ;
  assign n30302 = n156 & n46054 ;
  assign n29346 = n29315 | n29329 ;
  assign n46055 = ~n29346 ;
  assign n29783 = n46055 & n131 ;
  assign n29784 = n28969 | n29783 ;
  assign n29344 = n28969 & n45618 ;
  assign n46056 = ~n29315 ;
  assign n29345 = n46056 & n29344 ;
  assign n29788 = n29345 & n131 ;
  assign n46057 = ~n29788 ;
  assign n29789 = n29784 & n46057 ;
  assign n30283 = n10657 | n30282 ;
  assign n46058 = ~n30283 ;
  assign n30303 = n46058 & n30300 ;
  assign n30304 = n29789 | n30303 ;
  assign n46059 = ~n30302 ;
  assign n30305 = n46059 & n30304 ;
  assign n46060 = ~n30305 ;
  assign n30306 = n157 & n46060 ;
  assign n29343 = n29318 | n29331 ;
  assign n46061 = ~n29343 ;
  assign n29778 = n46061 & n131 ;
  assign n29779 = n29165 | n29778 ;
  assign n46062 = ~n29331 ;
  assign n29341 = n29165 & n46062 ;
  assign n29342 = n45607 & n29341 ;
  assign n29880 = n29342 & n131 ;
  assign n46063 = ~n29880 ;
  assign n29881 = n29779 & n46063 ;
  assign n30314 = n46042 & n30295 ;
  assign n30315 = n29800 | n30314 ;
  assign n46064 = ~n30297 ;
  assign n30316 = n46064 & n30315 ;
  assign n46065 = ~n30316 ;
  assign n30317 = n155 & n46065 ;
  assign n30318 = n46052 & n30315 ;
  assign n30319 = n29810 | n30318 ;
  assign n46066 = ~n30317 ;
  assign n30320 = n46066 & n30319 ;
  assign n46067 = ~n30320 ;
  assign n30321 = n10657 & n46067 ;
  assign n30322 = n157 | n30321 ;
  assign n46068 = ~n30322 ;
  assign n30323 = n30304 & n46068 ;
  assign n30324 = n29881 | n30323 ;
  assign n46069 = ~n30306 ;
  assign n30325 = n46069 & n30324 ;
  assign n46070 = ~n30325 ;
  assign n30326 = n158 & n46070 ;
  assign n29340 = n29334 | n29335 ;
  assign n46071 = ~n29340 ;
  assign n29774 = n46071 & n131 ;
  assign n29775 = n29063 | n29774 ;
  assign n29365 = n29063 & n45634 ;
  assign n46072 = ~n29335 ;
  assign n29366 = n46072 & n29365 ;
  assign n29836 = n29366 & n131 ;
  assign n46073 = ~n29836 ;
  assign n29837 = n29775 & n46073 ;
  assign n30307 = n158 | n30306 ;
  assign n46074 = ~n30307 ;
  assign n30327 = n46074 & n30324 ;
  assign n30328 = n29837 | n30327 ;
  assign n46075 = ~n30326 ;
  assign n30329 = n46075 & n30328 ;
  assign n46076 = ~n30329 ;
  assign n30330 = n8857 & n46076 ;
  assign n29364 = n29338 | n29352 ;
  assign n46077 = ~n29364 ;
  assign n29815 = n46077 & n131 ;
  assign n29816 = n29027 | n29815 ;
  assign n46078 = ~n29352 ;
  assign n29362 = n29027 & n46078 ;
  assign n29363 = n45623 & n29362 ;
  assign n29867 = n29363 & n131 ;
  assign n46079 = ~n29867 ;
  assign n29868 = n29816 & n46079 ;
  assign n30338 = n46058 & n30319 ;
  assign n30339 = n29789 | n30338 ;
  assign n46080 = ~n30321 ;
  assign n30340 = n46080 & n30339 ;
  assign n46081 = ~n30340 ;
  assign n30341 = n157 & n46081 ;
  assign n30342 = n46068 & n30339 ;
  assign n30343 = n29881 | n30342 ;
  assign n46082 = ~n30341 ;
  assign n30344 = n46082 & n30343 ;
  assign n46083 = ~n30344 ;
  assign n30345 = n158 & n46083 ;
  assign n30346 = n8857 | n30345 ;
  assign n46084 = ~n30346 ;
  assign n30347 = n30328 & n46084 ;
  assign n30348 = n29868 | n30347 ;
  assign n46085 = ~n30330 ;
  assign n30349 = n46085 & n30348 ;
  assign n46086 = ~n30349 ;
  assign n30350 = n160 & n46086 ;
  assign n29361 = n29355 | n29356 ;
  assign n46087 = ~n29361 ;
  assign n29771 = n46087 & n131 ;
  assign n29772 = n28945 | n29771 ;
  assign n29385 = n28945 & n45640 ;
  assign n46088 = ~n29356 ;
  assign n29386 = n46088 & n29385 ;
  assign n29776 = n29386 & n131 ;
  assign n46089 = ~n29776 ;
  assign n29777 = n29772 & n46089 ;
  assign n30331 = n160 | n30330 ;
  assign n46090 = ~n30331 ;
  assign n30351 = n46090 & n30348 ;
  assign n30352 = n29777 | n30351 ;
  assign n46091 = ~n30350 ;
  assign n30353 = n46091 & n30352 ;
  assign n46092 = ~n30353 ;
  assign n30354 = n161 & n46092 ;
  assign n29384 = n29359 | n29372 ;
  assign n46093 = ~n29384 ;
  assign n29780 = n46093 & n131 ;
  assign n29781 = n29018 | n29780 ;
  assign n46094 = ~n29372 ;
  assign n29382 = n29018 & n46094 ;
  assign n29383 = n45649 & n29382 ;
  assign n29896 = n29383 & n131 ;
  assign n46095 = ~n29896 ;
  assign n29897 = n29781 & n46095 ;
  assign n30362 = n46074 & n30343 ;
  assign n30363 = n29837 | n30362 ;
  assign n46096 = ~n30345 ;
  assign n30364 = n46096 & n30363 ;
  assign n46097 = ~n30364 ;
  assign n30365 = n159 & n46097 ;
  assign n30366 = n46084 & n30363 ;
  assign n30367 = n29868 | n30366 ;
  assign n46098 = ~n30365 ;
  assign n30368 = n46098 & n30367 ;
  assign n46099 = ~n30368 ;
  assign n30369 = n8534 & n46099 ;
  assign n30370 = n161 | n30369 ;
  assign n46100 = ~n30370 ;
  assign n30371 = n30352 & n46100 ;
  assign n30372 = n29897 | n30371 ;
  assign n46101 = ~n30354 ;
  assign n30373 = n46101 & n30372 ;
  assign n46102 = ~n30373 ;
  assign n30374 = n162 & n46102 ;
  assign n29401 = n29156 & n45645 ;
  assign n46103 = ~n29376 ;
  assign n29402 = n46103 & n29401 ;
  assign n29920 = n29402 & n131 ;
  assign n29377 = n29375 | n29376 ;
  assign n46104 = ~n29377 ;
  assign n29921 = n46104 & n131 ;
  assign n29922 = n29156 | n29921 ;
  assign n46105 = ~n29920 ;
  assign n29923 = n46105 & n29922 ;
  assign n30355 = n162 | n30354 ;
  assign n46106 = ~n30355 ;
  assign n30375 = n46106 & n30372 ;
  assign n30376 = n29923 | n30375 ;
  assign n46107 = ~n30374 ;
  assign n30377 = n46107 & n30376 ;
  assign n46108 = ~n30377 ;
  assign n30378 = n6889 & n46108 ;
  assign n46109 = ~n29392 ;
  assign n29398 = n29042 & n46109 ;
  assign n29399 = n45662 & n29398 ;
  assign n29924 = n29399 & n131 ;
  assign n29400 = n29380 | n29392 ;
  assign n46110 = ~n29400 ;
  assign n29925 = n46110 & n131 ;
  assign n29926 = n29042 | n29925 ;
  assign n46111 = ~n29924 ;
  assign n29927 = n46111 & n29926 ;
  assign n30386 = n46090 & n30367 ;
  assign n30387 = n29777 | n30386 ;
  assign n46112 = ~n30369 ;
  assign n30388 = n46112 & n30387 ;
  assign n46113 = ~n30388 ;
  assign n30389 = n161 & n46113 ;
  assign n30390 = n46100 & n30387 ;
  assign n30391 = n29897 | n30390 ;
  assign n46114 = ~n30389 ;
  assign n30392 = n46114 & n30391 ;
  assign n46115 = ~n30392 ;
  assign n30393 = n162 & n46115 ;
  assign n30394 = n6889 | n30393 ;
  assign n46116 = ~n30394 ;
  assign n30395 = n30376 & n46116 ;
  assign n30396 = n29927 | n30395 ;
  assign n46117 = ~n30378 ;
  assign n30397 = n46117 & n30396 ;
  assign n46118 = ~n30397 ;
  assign n30398 = n164 & n46118 ;
  assign n29423 = n45658 & n29410 ;
  assign n46119 = ~n29396 ;
  assign n29424 = n46119 & n29423 ;
  assign n29893 = n29424 & n131 ;
  assign n29397 = n29395 | n29396 ;
  assign n46120 = ~n29397 ;
  assign n29930 = n46120 & n131 ;
  assign n29931 = n29410 | n29930 ;
  assign n46121 = ~n29893 ;
  assign n29932 = n46121 & n29931 ;
  assign n30379 = n6600 | n30378 ;
  assign n46122 = ~n30379 ;
  assign n30399 = n46122 & n30396 ;
  assign n30400 = n29932 | n30399 ;
  assign n46123 = ~n30398 ;
  assign n30401 = n46123 & n30400 ;
  assign n46124 = ~n30401 ;
  assign n30402 = n165 & n46124 ;
  assign n46125 = ~n29415 ;
  assign n29420 = n29024 & n46125 ;
  assign n29421 = n45675 & n29420 ;
  assign n29933 = n29421 & n131 ;
  assign n29422 = n29413 | n29415 ;
  assign n46126 = ~n29422 ;
  assign n29937 = n46126 & n131 ;
  assign n29938 = n29024 | n29937 ;
  assign n46127 = ~n29933 ;
  assign n29939 = n46127 & n29938 ;
  assign n30410 = n46106 & n30391 ;
  assign n30411 = n29923 | n30410 ;
  assign n46128 = ~n30393 ;
  assign n30412 = n46128 & n30411 ;
  assign n46129 = ~n30412 ;
  assign n30413 = n163 & n46129 ;
  assign n30414 = n46116 & n30411 ;
  assign n30415 = n29927 | n30414 ;
  assign n46130 = ~n30413 ;
  assign n30416 = n46130 & n30415 ;
  assign n46131 = ~n30416 ;
  assign n30417 = n6600 & n46131 ;
  assign n30418 = n165 | n30417 ;
  assign n46132 = ~n30418 ;
  assign n30419 = n30400 & n46132 ;
  assign n30420 = n29939 | n30419 ;
  assign n46133 = ~n30402 ;
  assign n30421 = n46133 & n30420 ;
  assign n46134 = ~n30421 ;
  assign n30422 = n166 & n46134 ;
  assign n29454 = n45671 & n29441 ;
  assign n46135 = ~n29419 ;
  assign n29455 = n46135 & n29454 ;
  assign n29807 = n29455 & n131 ;
  assign n29430 = n29419 | n29428 ;
  assign n46136 = ~n29430 ;
  assign n29847 = n46136 & n131 ;
  assign n29848 = n29441 | n29847 ;
  assign n46137 = ~n29807 ;
  assign n29849 = n46137 & n29848 ;
  assign n30403 = n166 | n30402 ;
  assign n46138 = ~n30403 ;
  assign n30423 = n46138 & n30420 ;
  assign n30425 = n29849 | n30423 ;
  assign n46139 = ~n30422 ;
  assign n30426 = n46139 & n30425 ;
  assign n46140 = ~n30426 ;
  assign n30427 = n5352 & n46140 ;
  assign n46141 = ~n29446 ;
  assign n29451 = n29020 & n46141 ;
  assign n29452 = n45688 & n29451 ;
  assign n29942 = n29452 & n131 ;
  assign n29453 = n29444 | n29446 ;
  assign n46142 = ~n29453 ;
  assign n29943 = n46142 & n131 ;
  assign n29944 = n29020 | n29943 ;
  assign n46143 = ~n29942 ;
  assign n29945 = n46143 & n29944 ;
  assign n30434 = n46122 & n30415 ;
  assign n30435 = n29932 | n30434 ;
  assign n46144 = ~n30417 ;
  assign n30436 = n46144 & n30435 ;
  assign n46145 = ~n30436 ;
  assign n30437 = n165 & n46145 ;
  assign n30438 = n46132 & n30435 ;
  assign n30439 = n29939 | n30438 ;
  assign n46146 = ~n30437 ;
  assign n30440 = n46146 & n30439 ;
  assign n46147 = ~n30440 ;
  assign n30441 = n166 & n46147 ;
  assign n30442 = n5352 | n30441 ;
  assign n46148 = ~n30442 ;
  assign n30443 = n30425 & n46148 ;
  assign n30444 = n29945 | n30443 ;
  assign n46149 = ~n30427 ;
  assign n30445 = n46149 & n30444 ;
  assign n46150 = ~n30445 ;
  assign n30446 = n168 & n46150 ;
  assign n29461 = n29450 | n29459 ;
  assign n46151 = ~n29461 ;
  assign n29861 = n46151 & n131 ;
  assign n29862 = n29463 | n29861 ;
  assign n29476 = n45684 & n29463 ;
  assign n46152 = ~n29450 ;
  assign n29477 = n46152 & n29476 ;
  assign n29946 = n29477 & n131 ;
  assign n46153 = ~n29946 ;
  assign n29947 = n29862 & n46153 ;
  assign n30428 = n4934 | n30427 ;
  assign n46154 = ~n30428 ;
  assign n30447 = n46154 & n30444 ;
  assign n30448 = n29947 | n30447 ;
  assign n46155 = ~n30446 ;
  assign n30449 = n46155 & n30448 ;
  assign n46156 = ~n30449 ;
  assign n30450 = n169 & n46156 ;
  assign n46157 = ~n29468 ;
  assign n29473 = n29159 & n46157 ;
  assign n29474 = n45701 & n29473 ;
  assign n29856 = n29474 & n131 ;
  assign n29475 = n29466 | n29468 ;
  assign n46158 = ~n29475 ;
  assign n29948 = n46158 & n131 ;
  assign n29949 = n29159 | n29948 ;
  assign n46159 = ~n29856 ;
  assign n29950 = n46159 & n29949 ;
  assign n30458 = n46138 & n30439 ;
  assign n30459 = n29849 | n30458 ;
  assign n46160 = ~n30441 ;
  assign n30460 = n46160 & n30459 ;
  assign n46161 = ~n30460 ;
  assign n30461 = n167 & n46161 ;
  assign n30462 = n46148 & n30459 ;
  assign n30463 = n29945 | n30462 ;
  assign n46162 = ~n30461 ;
  assign n30464 = n46162 & n30463 ;
  assign n46163 = ~n30464 ;
  assign n30465 = n4934 & n46163 ;
  assign n30466 = n169 | n30465 ;
  assign n46164 = ~n30466 ;
  assign n30467 = n30448 & n46164 ;
  assign n30468 = n29950 | n30467 ;
  assign n46165 = ~n30450 ;
  assign n30469 = n46165 & n30468 ;
  assign n46166 = ~n30469 ;
  assign n30470 = n170 & n46166 ;
  assign n29499 = n45697 & n29485 ;
  assign n46167 = ~n29472 ;
  assign n29500 = n46167 & n29499 ;
  assign n29951 = n29500 & n131 ;
  assign n29483 = n29472 | n29481 ;
  assign n46168 = ~n29483 ;
  assign n29955 = n46168 & n131 ;
  assign n29956 = n29485 | n29955 ;
  assign n46169 = ~n29951 ;
  assign n29957 = n46169 & n29956 ;
  assign n30451 = n170 | n30450 ;
  assign n46170 = ~n30451 ;
  assign n30471 = n46170 & n30468 ;
  assign n30472 = n29957 | n30471 ;
  assign n46171 = ~n30470 ;
  assign n30473 = n46171 & n30472 ;
  assign n46172 = ~n30473 ;
  assign n30474 = n3940 & n46172 ;
  assign n29498 = n29488 | n29490 ;
  assign n46173 = ~n29498 ;
  assign n29940 = n46173 & n131 ;
  assign n29941 = n29145 | n29940 ;
  assign n46174 = ~n29490 ;
  assign n29496 = n29145 & n46174 ;
  assign n29497 = n45717 & n29496 ;
  assign n29960 = n29497 & n131 ;
  assign n46175 = ~n29960 ;
  assign n29961 = n29941 & n46175 ;
  assign n30482 = n46154 & n30463 ;
  assign n30483 = n29947 | n30482 ;
  assign n46176 = ~n30465 ;
  assign n30484 = n46176 & n30483 ;
  assign n46177 = ~n30484 ;
  assign n30485 = n169 & n46177 ;
  assign n30486 = n46164 & n30483 ;
  assign n30487 = n29950 | n30486 ;
  assign n46178 = ~n30485 ;
  assign n30488 = n46178 & n30487 ;
  assign n46179 = ~n30488 ;
  assign n30489 = n170 & n46179 ;
  assign n30490 = n3940 | n30489 ;
  assign n46180 = ~n30490 ;
  assign n30491 = n30472 & n46180 ;
  assign n30492 = n29961 | n30491 ;
  assign n46181 = ~n30474 ;
  assign n30493 = n46181 & n30492 ;
  assign n46182 = ~n30493 ;
  assign n30494 = n172 & n46182 ;
  assign n29515 = n45709 & n29508 ;
  assign n46183 = ~n29494 ;
  assign n29516 = n46183 & n29515 ;
  assign n29962 = n29516 & n131 ;
  assign n29495 = n29493 | n29494 ;
  assign n46184 = ~n29495 ;
  assign n29963 = n46184 & n131 ;
  assign n29964 = n29508 | n29963 ;
  assign n46185 = ~n29962 ;
  assign n29965 = n46185 & n29964 ;
  assign n30475 = n3631 | n30474 ;
  assign n46186 = ~n30475 ;
  assign n30495 = n46186 & n30492 ;
  assign n30496 = n29965 | n30495 ;
  assign n46187 = ~n30494 ;
  assign n30497 = n46187 & n30496 ;
  assign n46188 = ~n30497 ;
  assign n30498 = n173 & n46188 ;
  assign n46189 = ~n29513 ;
  assign n29528 = n46189 & n29522 ;
  assign n29529 = n45730 & n29528 ;
  assign n29818 = n29529 & n131 ;
  assign n29514 = n29511 | n29513 ;
  assign n46190 = ~n29514 ;
  assign n29966 = n46190 & n131 ;
  assign n29967 = n29522 | n29966 ;
  assign n46191 = ~n29818 ;
  assign n29968 = n46191 & n29967 ;
  assign n30506 = n46170 & n30487 ;
  assign n30507 = n29957 | n30506 ;
  assign n46192 = ~n30489 ;
  assign n30508 = n46192 & n30507 ;
  assign n46193 = ~n30508 ;
  assign n30509 = n171 & n46193 ;
  assign n30510 = n46180 & n30507 ;
  assign n30511 = n29961 | n30510 ;
  assign n46194 = ~n30509 ;
  assign n30512 = n46194 & n30511 ;
  assign n46195 = ~n30512 ;
  assign n30513 = n3631 & n46195 ;
  assign n30514 = n173 | n30513 ;
  assign n46196 = ~n30514 ;
  assign n30515 = n30496 & n46196 ;
  assign n30516 = n29968 | n30515 ;
  assign n46197 = ~n30498 ;
  assign n30517 = n46197 & n30516 ;
  assign n46198 = ~n30517 ;
  assign n30518 = n174 & n46198 ;
  assign n29548 = n45726 & n29534 ;
  assign n46199 = ~n29527 ;
  assign n29549 = n46199 & n29548 ;
  assign n29808 = n29549 & n131 ;
  assign n29532 = n29527 | n29531 ;
  assign n46200 = ~n29532 ;
  assign n29969 = n46200 & n131 ;
  assign n29970 = n29534 | n29969 ;
  assign n46201 = ~n29808 ;
  assign n29971 = n46201 & n29970 ;
  assign n30499 = n174 | n30498 ;
  assign n46202 = ~n30499 ;
  assign n30519 = n46202 & n30516 ;
  assign n30521 = n29971 | n30519 ;
  assign n46203 = ~n30518 ;
  assign n30522 = n46203 & n30521 ;
  assign n46204 = ~n30522 ;
  assign n30523 = n2753 & n46204 ;
  assign n46205 = ~n29539 ;
  assign n29545 = n29065 & n46205 ;
  assign n29546 = n45746 & n29545 ;
  assign n29972 = n29546 & n131 ;
  assign n29547 = n29537 | n29539 ;
  assign n46206 = ~n29547 ;
  assign n29973 = n46206 & n131 ;
  assign n29974 = n29065 | n29973 ;
  assign n46207 = ~n29972 ;
  assign n29975 = n46207 & n29974 ;
  assign n30530 = n46186 & n30511 ;
  assign n30531 = n29965 | n30530 ;
  assign n46208 = ~n30513 ;
  assign n30532 = n46208 & n30531 ;
  assign n46209 = ~n30532 ;
  assign n30533 = n173 & n46209 ;
  assign n30534 = n46196 & n30531 ;
  assign n30535 = n29968 | n30534 ;
  assign n46210 = ~n30533 ;
  assign n30536 = n46210 & n30535 ;
  assign n46211 = ~n30536 ;
  assign n30537 = n174 & n46211 ;
  assign n30538 = n2753 | n30537 ;
  assign n46212 = ~n30538 ;
  assign n30539 = n30521 & n46212 ;
  assign n30540 = n29975 | n30539 ;
  assign n46213 = ~n30523 ;
  assign n30541 = n46213 & n30540 ;
  assign n46214 = ~n30541 ;
  assign n30542 = n176 & n46214 ;
  assign n29544 = n29542 | n29543 ;
  assign n46215 = ~n29544 ;
  assign n29885 = n46215 & n131 ;
  assign n29886 = n29556 | n29885 ;
  assign n29563 = n45738 & n29556 ;
  assign n46216 = ~n29543 ;
  assign n29564 = n46216 & n29563 ;
  assign n29976 = n29564 & n131 ;
  assign n46217 = ~n29976 ;
  assign n29977 = n29886 & n46217 ;
  assign n30524 = n2431 | n30523 ;
  assign n46218 = ~n30524 ;
  assign n30543 = n46218 & n30540 ;
  assign n30544 = n29977 | n30543 ;
  assign n46219 = ~n30542 ;
  assign n30545 = n46219 & n30544 ;
  assign n46220 = ~n30545 ;
  assign n30546 = n177 & n46220 ;
  assign n29562 = n29559 | n29561 ;
  assign n46221 = ~n29562 ;
  assign n29857 = n46221 & n131 ;
  assign n29858 = n29568 | n29857 ;
  assign n46222 = ~n29561 ;
  assign n29574 = n46222 & n29568 ;
  assign n29575 = n45759 & n29574 ;
  assign n29978 = n29575 & n131 ;
  assign n46223 = ~n29978 ;
  assign n29979 = n29858 & n46223 ;
  assign n30554 = n46202 & n30535 ;
  assign n30555 = n29971 | n30554 ;
  assign n46224 = ~n30537 ;
  assign n30556 = n46224 & n30555 ;
  assign n46225 = ~n30556 ;
  assign n30557 = n175 & n46225 ;
  assign n30558 = n46212 & n30555 ;
  assign n30559 = n29975 | n30558 ;
  assign n46226 = ~n30557 ;
  assign n30560 = n46226 & n30559 ;
  assign n46227 = ~n30560 ;
  assign n30561 = n2431 & n46227 ;
  assign n30562 = n177 | n30561 ;
  assign n46228 = ~n30562 ;
  assign n30563 = n30544 & n46228 ;
  assign n30564 = n29979 | n30563 ;
  assign n46229 = ~n30546 ;
  assign n30565 = n46229 & n30564 ;
  assign n46230 = ~n30565 ;
  assign n30566 = n178 & n46230 ;
  assign n29594 = n45755 & n29580 ;
  assign n46231 = ~n29573 ;
  assign n29595 = n46231 & n29594 ;
  assign n29821 = n29595 & n131 ;
  assign n29578 = n29573 | n29577 ;
  assign n46232 = ~n29578 ;
  assign n29980 = n46232 & n131 ;
  assign n29981 = n29580 | n29980 ;
  assign n46233 = ~n29821 ;
  assign n29982 = n46233 & n29981 ;
  assign n30547 = n178 | n30546 ;
  assign n46234 = ~n30547 ;
  assign n30567 = n46234 & n30564 ;
  assign n30568 = n29982 | n30567 ;
  assign n46235 = ~n30566 ;
  assign n30569 = n46235 & n30568 ;
  assign n46236 = ~n30569 ;
  assign n30570 = n1707 & n46236 ;
  assign n46237 = ~n29585 ;
  assign n29591 = n29433 & n46237 ;
  assign n29592 = n45775 & n29591 ;
  assign n29983 = n29592 & n131 ;
  assign n29593 = n29583 | n29585 ;
  assign n46238 = ~n29593 ;
  assign n29984 = n46238 & n131 ;
  assign n29985 = n29433 | n29984 ;
  assign n46239 = ~n29983 ;
  assign n29986 = n46239 & n29985 ;
  assign n30578 = n46218 & n30559 ;
  assign n30579 = n29977 | n30578 ;
  assign n46240 = ~n30561 ;
  assign n30580 = n46240 & n30579 ;
  assign n46241 = ~n30580 ;
  assign n30581 = n177 & n46241 ;
  assign n30582 = n46228 & n30579 ;
  assign n30583 = n29979 | n30582 ;
  assign n46242 = ~n30581 ;
  assign n30584 = n46242 & n30583 ;
  assign n46243 = ~n30584 ;
  assign n30585 = n178 & n46243 ;
  assign n30586 = n1707 | n30585 ;
  assign n46244 = ~n30586 ;
  assign n30587 = n30568 & n46244 ;
  assign n30588 = n29986 | n30587 ;
  assign n46245 = ~n30570 ;
  assign n30589 = n46245 & n30588 ;
  assign n46246 = ~n30589 ;
  assign n30590 = n180 & n46246 ;
  assign n29590 = n29588 | n29589 ;
  assign n46247 = ~n29590 ;
  assign n29803 = n46247 & n131 ;
  assign n29804 = n29603 | n29803 ;
  assign n29610 = n45767 & n29603 ;
  assign n46248 = ~n29589 ;
  assign n29611 = n46248 & n29610 ;
  assign n30033 = n29611 & n30015 ;
  assign n46249 = ~n30033 ;
  assign n30034 = n29804 & n46249 ;
  assign n30571 = n1487 | n30570 ;
  assign n46250 = ~n30571 ;
  assign n30591 = n46250 & n30588 ;
  assign n30592 = n30034 | n30591 ;
  assign n46251 = ~n30590 ;
  assign n30593 = n46251 & n30592 ;
  assign n46252 = ~n30593 ;
  assign n30594 = n181 & n46252 ;
  assign n46253 = ~n29608 ;
  assign n29625 = n46253 & n29619 ;
  assign n29626 = n45788 & n29625 ;
  assign n29829 = n29626 & n131 ;
  assign n29609 = n29606 | n29608 ;
  assign n46254 = ~n29609 ;
  assign n29934 = n46254 & n131 ;
  assign n29935 = n29619 | n29934 ;
  assign n46255 = ~n29829 ;
  assign n29936 = n46255 & n29935 ;
  assign n30602 = n46234 & n30583 ;
  assign n30603 = n29982 | n30602 ;
  assign n46256 = ~n30585 ;
  assign n30604 = n46256 & n30603 ;
  assign n46257 = ~n30604 ;
  assign n30605 = n179 & n46257 ;
  assign n30606 = n46244 & n30603 ;
  assign n30607 = n29986 | n30606 ;
  assign n46258 = ~n30605 ;
  assign n30608 = n46258 & n30607 ;
  assign n46259 = ~n30608 ;
  assign n30609 = n1487 & n46259 ;
  assign n30610 = n181 | n30609 ;
  assign n46260 = ~n30610 ;
  assign n30611 = n30592 & n46260 ;
  assign n30612 = n29936 | n30611 ;
  assign n46261 = ~n30594 ;
  assign n30613 = n46261 & n30612 ;
  assign n46262 = ~n30613 ;
  assign n30614 = n182 & n46262 ;
  assign n29629 = n29624 | n29628 ;
  assign n46263 = ~n29629 ;
  assign n29928 = n46263 & n131 ;
  assign n29929 = n29633 | n29928 ;
  assign n29647 = n45784 & n29633 ;
  assign n46264 = ~n29624 ;
  assign n29648 = n46264 & n29647 ;
  assign n29987 = n29648 & n131 ;
  assign n46265 = ~n29987 ;
  assign n29988 = n29929 & n46265 ;
  assign n30595 = n182 | n30594 ;
  assign n46266 = ~n30595 ;
  assign n30615 = n46266 & n30612 ;
  assign n30616 = n29988 | n30615 ;
  assign n46267 = ~n30614 ;
  assign n30617 = n46267 & n30616 ;
  assign n46268 = ~n30617 ;
  assign n30618 = n996 & n46268 ;
  assign n46269 = ~n29638 ;
  assign n29645 = n29077 & n46269 ;
  assign n29646 = n45804 & n29645 ;
  assign n29914 = n29646 & n131 ;
  assign n29644 = n29636 | n29638 ;
  assign n46270 = ~n29644 ;
  assign n29952 = n46270 & n131 ;
  assign n29953 = n29077 | n29952 ;
  assign n46271 = ~n29914 ;
  assign n29954 = n46271 & n29953 ;
  assign n30626 = n46250 & n30607 ;
  assign n30627 = n30034 | n30626 ;
  assign n46272 = ~n30609 ;
  assign n30628 = n46272 & n30627 ;
  assign n46273 = ~n30628 ;
  assign n30629 = n181 & n46273 ;
  assign n30630 = n46260 & n30627 ;
  assign n30631 = n29936 | n30630 ;
  assign n46274 = ~n30629 ;
  assign n30632 = n46274 & n30631 ;
  assign n46275 = ~n30632 ;
  assign n30633 = n182 & n46275 ;
  assign n30634 = n183 | n30633 ;
  assign n46276 = ~n30634 ;
  assign n30635 = n30616 & n46276 ;
  assign n30636 = n29954 | n30635 ;
  assign n46277 = ~n30618 ;
  assign n30637 = n46277 & n30636 ;
  assign n46278 = ~n30637 ;
  assign n30638 = n184 & n46278 ;
  assign n29662 = n45796 & n29655 ;
  assign n46279 = ~n29642 ;
  assign n29663 = n46279 & n29662 ;
  assign n29989 = n29663 & n131 ;
  assign n29643 = n29641 | n29642 ;
  assign n46280 = ~n29643 ;
  assign n29990 = n46280 & n131 ;
  assign n29991 = n29655 | n29990 ;
  assign n46281 = ~n29989 ;
  assign n29992 = n46281 & n29991 ;
  assign n30619 = n838 | n30618 ;
  assign n46282 = ~n30619 ;
  assign n30639 = n46282 & n30636 ;
  assign n30640 = n29992 | n30639 ;
  assign n46283 = ~n30638 ;
  assign n30641 = n46283 & n30640 ;
  assign n46284 = ~n30641 ;
  assign n30642 = n185 & n46284 ;
  assign n29661 = n29658 | n29660 ;
  assign n46285 = ~n29661 ;
  assign n29993 = n46285 & n131 ;
  assign n29994 = n29671 | n29993 ;
  assign n46286 = ~n29660 ;
  assign n29677 = n46286 & n29671 ;
  assign n29678 = n45823 & n29677 ;
  assign n30039 = n29678 & n30015 ;
  assign n46287 = ~n30039 ;
  assign n30040 = n29994 & n46287 ;
  assign n30650 = n46266 & n30631 ;
  assign n30651 = n29988 | n30650 ;
  assign n46288 = ~n30633 ;
  assign n30652 = n46288 & n30651 ;
  assign n46289 = ~n30652 ;
  assign n30653 = n183 & n46289 ;
  assign n30654 = n46276 & n30651 ;
  assign n30655 = n29954 | n30654 ;
  assign n46290 = ~n30653 ;
  assign n30656 = n46290 & n30655 ;
  assign n46291 = ~n30656 ;
  assign n30657 = n838 & n46291 ;
  assign n30658 = n185 | n30657 ;
  assign n46292 = ~n30658 ;
  assign n30659 = n30640 & n46292 ;
  assign n30660 = n30040 | n30659 ;
  assign n46293 = ~n30642 ;
  assign n30661 = n46293 & n30660 ;
  assign n46294 = ~n30661 ;
  assign n30662 = n186 & n46294 ;
  assign n29695 = n45812 & n29688 ;
  assign n46295 = ~n29676 ;
  assign n29696 = n46295 & n29695 ;
  assign n29843 = n29696 & n131 ;
  assign n29681 = n29676 | n29680 ;
  assign n46296 = ~n29681 ;
  assign n29995 = n46296 & n131 ;
  assign n29996 = n29688 | n29995 ;
  assign n46297 = ~n29843 ;
  assign n29997 = n46297 & n29996 ;
  assign n30643 = n186 | n30642 ;
  assign n46298 = ~n30643 ;
  assign n30663 = n46298 & n30660 ;
  assign n30664 = n29997 | n30663 ;
  assign n46299 = ~n30662 ;
  assign n30665 = n46299 & n30664 ;
  assign n46300 = ~n30665 ;
  assign n30666 = n528 & n46300 ;
  assign n46301 = ~n29693 ;
  assign n29716 = n46301 & n29700 ;
  assign n29717 = n45829 & n29716 ;
  assign n29998 = n29717 & n131 ;
  assign n29694 = n29691 | n29693 ;
  assign n46302 = ~n29694 ;
  assign n29999 = n46302 & n131 ;
  assign n30000 = n29700 | n29999 ;
  assign n46303 = ~n29998 ;
  assign n30001 = n46303 & n30000 ;
  assign n30674 = n46282 & n30655 ;
  assign n30675 = n29992 | n30674 ;
  assign n46304 = ~n30657 ;
  assign n30676 = n46304 & n30675 ;
  assign n46305 = ~n30676 ;
  assign n30677 = n185 & n46305 ;
  assign n30678 = n46292 & n30675 ;
  assign n30679 = n30040 | n30678 ;
  assign n46306 = ~n30677 ;
  assign n30680 = n46306 & n30679 ;
  assign n46307 = ~n30680 ;
  assign n30681 = n186 & n46307 ;
  assign n30682 = n528 | n30681 ;
  assign n46308 = ~n30682 ;
  assign n30683 = n30664 & n46308 ;
  assign n30684 = n30001 | n30683 ;
  assign n46309 = ~n30666 ;
  assign n30685 = n46309 & n30684 ;
  assign n46310 = ~n30685 ;
  assign n30686 = n188 & n46310 ;
  assign n29721 = n29706 | n29719 ;
  assign n46311 = ~n29721 ;
  assign n29830 = n46311 & n131 ;
  assign n29831 = n29032 | n29830 ;
  assign n29705 = n29032 & n45841 ;
  assign n46312 = ~n29706 ;
  assign n29720 = n29705 & n46312 ;
  assign n30029 = n29720 & n30015 ;
  assign n46313 = ~n30029 ;
  assign n30030 = n29831 & n46313 ;
  assign n30667 = n413 | n30666 ;
  assign n46314 = ~n30667 ;
  assign n30687 = n46314 & n30684 ;
  assign n30688 = n30030 | n30687 ;
  assign n46315 = ~n30686 ;
  assign n30689 = n46315 & n30688 ;
  assign n46316 = ~n30689 ;
  assign n30690 = n189 & n46316 ;
  assign n29739 = n29710 | n29723 ;
  assign n46317 = ~n29739 ;
  assign n29958 = n46317 & n131 ;
  assign n29959 = n29683 | n29958 ;
  assign n46318 = ~n29710 ;
  assign n29737 = n29683 & n46318 ;
  assign n29738 = n45833 & n29737 ;
  assign n30002 = n29738 & n131 ;
  assign n46319 = ~n30002 ;
  assign n30003 = n29959 & n46319 ;
  assign n30698 = n46298 & n30679 ;
  assign n30699 = n29997 | n30698 ;
  assign n46320 = ~n30681 ;
  assign n30700 = n46320 & n30699 ;
  assign n46321 = ~n30700 ;
  assign n30701 = n187 & n46321 ;
  assign n30702 = n46308 & n30699 ;
  assign n30703 = n30001 | n30702 ;
  assign n46322 = ~n30701 ;
  assign n30704 = n46322 & n30703 ;
  assign n46323 = ~n30704 ;
  assign n30705 = n413 & n46323 ;
  assign n30706 = n189 | n30705 ;
  assign n46324 = ~n30706 ;
  assign n30707 = n30688 & n46324 ;
  assign n30708 = n30003 | n30707 ;
  assign n46325 = ~n30690 ;
  assign n30709 = n46325 & n30708 ;
  assign n46326 = ~n30709 ;
  assign n30710 = n190 & n46326 ;
  assign n46327 = ~n29713 ;
  assign n29715 = n29667 & n46327 ;
  assign n46328 = ~n29727 ;
  assign n29735 = n29715 & n46328 ;
  assign n29850 = n29735 & n131 ;
  assign n29736 = n29726 | n29727 ;
  assign n46329 = ~n29736 ;
  assign n29873 = n46329 & n131 ;
  assign n29874 = n29667 | n29873 ;
  assign n46330 = ~n29850 ;
  assign n29875 = n46330 & n29874 ;
  assign n30691 = n190 | n30690 ;
  assign n46331 = ~n30691 ;
  assign n30711 = n46331 & n30708 ;
  assign n30712 = n29875 | n30711 ;
  assign n46332 = ~n30710 ;
  assign n30713 = n46332 & n30712 ;
  assign n46333 = ~n30713 ;
  assign n30714 = n287 & n46333 ;
  assign n30722 = n46314 & n30703 ;
  assign n30723 = n30030 | n30722 ;
  assign n46334 = ~n30705 ;
  assign n30724 = n46334 & n30723 ;
  assign n46335 = ~n30724 ;
  assign n30725 = n189 & n46335 ;
  assign n30726 = n46324 & n30723 ;
  assign n30727 = n30003 | n30726 ;
  assign n46336 = ~n30725 ;
  assign n30728 = n46336 & n30727 ;
  assign n46337 = ~n30728 ;
  assign n30729 = n190 & n46337 ;
  assign n30730 = n287 | n30729 ;
  assign n46338 = ~n30730 ;
  assign n30731 = n30712 & n46338 ;
  assign n46339 = ~n29729 ;
  assign n29756 = n46339 & n29755 ;
  assign n29757 = n45850 & n29756 ;
  assign n30004 = n29757 & n131 ;
  assign n29732 = n29729 | n29731 ;
  assign n46340 = ~n29732 ;
  assign n30005 = n46340 & n131 ;
  assign n30746 = n29755 | n30005 ;
  assign n46341 = ~n30004 ;
  assign n30747 = n46341 & n30746 ;
  assign n30750 = n30731 | n30747 ;
  assign n46342 = ~n30714 ;
  assign n30751 = n46342 & n30750 ;
  assign n30752 = n30038 | n30751 ;
  assign n30753 = n192 & n30752 ;
  assign n30738 = n29748 | n30010 ;
  assign n46343 = ~n30738 ;
  assign n30739 = n131 & n46343 ;
  assign n30740 = n30013 | n30739 ;
  assign n30741 = n30038 | n30740 ;
  assign n30754 = n30741 | n30751 ;
  assign n30755 = n31336 & n30754 ;
  assign n46344 = ~n29748 ;
  assign n29833 = n46344 & n131 ;
  assign n46345 = ~n29833 ;
  assign n30737 = n46345 & n30010 ;
  assign n30742 = n192 & n30738 ;
  assign n46346 = ~n30737 ;
  assign n30743 = n46346 & n30742 ;
  assign n30715 = n30038 & n46342 ;
  assign n30756 = n30715 & n30750 ;
  assign n30757 = n30743 | n30756 ;
  assign n130 = n30755 | n30757 ;
  assign n46347 = ~n30038 ;
  assign n30996 = n46347 & n130 ;
  assign n46348 = ~n30996 ;
  assign n30997 = n30751 & n46348 ;
  assign n46349 = ~n30997 ;
  assign n30998 = n30753 & n46349 ;
  assign n46350 = ~n30729 ;
  assign n30733 = n29875 & n46350 ;
  assign n46351 = ~n30711 ;
  assign n30734 = n46351 & n30733 ;
  assign n30872 = n30734 & n130 ;
  assign n30716 = n30710 | n30711 ;
  assign n46352 = ~n30716 ;
  assign n30876 = n46352 & n130 ;
  assign n30877 = n29875 | n30876 ;
  assign n46353 = ~n30872 ;
  assign n30878 = n46353 & n30877 ;
  assign n30720 = n30030 & n46334 ;
  assign n46354 = ~n30687 ;
  assign n30721 = n46354 & n30720 ;
  assign n30861 = n30721 & n130 ;
  assign n30692 = n30686 | n30687 ;
  assign n46355 = ~n30692 ;
  assign n30881 = n46355 & n130 ;
  assign n30882 = n30030 | n30881 ;
  assign n46356 = ~n30861 ;
  assign n30883 = n46356 & n30882 ;
  assign n30696 = n29997 & n46320 ;
  assign n46357 = ~n30663 ;
  assign n30697 = n46357 & n30696 ;
  assign n30826 = n30697 & n130 ;
  assign n30668 = n30662 | n30663 ;
  assign n46358 = ~n30668 ;
  assign n30831 = n46358 & n130 ;
  assign n30832 = n29997 | n30831 ;
  assign n46359 = ~n30826 ;
  assign n30833 = n46359 & n30832 ;
  assign n30644 = n30638 | n30639 ;
  assign n46360 = ~n30644 ;
  assign n30851 = n46360 & n130 ;
  assign n30852 = n29992 | n30851 ;
  assign n30672 = n29992 & n46304 ;
  assign n46361 = ~n30639 ;
  assign n30673 = n46361 & n30672 ;
  assign n30866 = n30673 & n130 ;
  assign n46362 = ~n30866 ;
  assign n30867 = n30852 & n46362 ;
  assign n30648 = n29988 & n46288 ;
  assign n46363 = ~n30615 ;
  assign n30649 = n46363 & n30648 ;
  assign n30825 = n30649 & n130 ;
  assign n30620 = n30614 | n30615 ;
  assign n46364 = ~n30620 ;
  assign n30841 = n46364 & n130 ;
  assign n30842 = n29988 | n30841 ;
  assign n46365 = ~n30825 ;
  assign n30843 = n46365 & n30842 ;
  assign n30624 = n30034 & n46272 ;
  assign n46366 = ~n30591 ;
  assign n30625 = n46366 & n30624 ;
  assign n30808 = n30625 & n130 ;
  assign n30596 = n30590 | n30591 ;
  assign n46367 = ~n30596 ;
  assign n30812 = n46367 & n130 ;
  assign n30813 = n30034 | n30812 ;
  assign n46368 = ~n30808 ;
  assign n30814 = n46368 & n30813 ;
  assign n30600 = n29982 & n46256 ;
  assign n46369 = ~n30567 ;
  assign n30601 = n46369 & n30600 ;
  assign n30880 = n30601 & n130 ;
  assign n30572 = n30566 | n30567 ;
  assign n46370 = ~n30572 ;
  assign n30900 = n46370 & n130 ;
  assign n30901 = n29982 | n30900 ;
  assign n46371 = ~n30880 ;
  assign n30902 = n46371 & n30901 ;
  assign n30548 = n30542 | n30543 ;
  assign n46372 = ~n30548 ;
  assign n30764 = n46372 & n130 ;
  assign n30765 = n29977 | n30764 ;
  assign n30576 = n29977 & n46240 ;
  assign n46373 = ~n30543 ;
  assign n30577 = n46373 & n30576 ;
  assign n30781 = n30577 & n130 ;
  assign n46374 = ~n30781 ;
  assign n30782 = n30765 & n46374 ;
  assign n30520 = n30518 | n30519 ;
  assign n46375 = ~n30520 ;
  assign n30760 = n46375 & n130 ;
  assign n30761 = n29971 | n30760 ;
  assign n30552 = n29971 & n46224 ;
  assign n46376 = ~n30519 ;
  assign n30553 = n46376 & n30552 ;
  assign n30846 = n30553 & n130 ;
  assign n46377 = ~n30846 ;
  assign n30847 = n30761 & n46377 ;
  assign n30528 = n29965 & n46208 ;
  assign n46378 = ~n30495 ;
  assign n30529 = n46378 & n30528 ;
  assign n30821 = n30529 & n130 ;
  assign n30500 = n30494 | n30495 ;
  assign n46379 = ~n30500 ;
  assign n30897 = n46379 & n130 ;
  assign n30898 = n29965 | n30897 ;
  assign n46380 = ~n30821 ;
  assign n30899 = n46380 & n30898 ;
  assign n30476 = n30470 | n30471 ;
  assign n46381 = ~n30476 ;
  assign n30788 = n46381 & n130 ;
  assign n30789 = n29957 | n30788 ;
  assign n30504 = n29957 & n46192 ;
  assign n46382 = ~n30471 ;
  assign n30505 = n46382 & n30504 ;
  assign n30905 = n30505 & n130 ;
  assign n46383 = ~n30905 ;
  assign n30906 = n30789 & n46383 ;
  assign n30480 = n29947 & n46176 ;
  assign n46384 = ~n30447 ;
  assign n30481 = n46384 & n30480 ;
  assign n30845 = n30481 & n130 ;
  assign n30452 = n30446 | n30447 ;
  assign n46385 = ~n30452 ;
  assign n30853 = n46385 & n130 ;
  assign n30854 = n29947 | n30853 ;
  assign n46386 = ~n30845 ;
  assign n30855 = n46386 & n30854 ;
  assign n30424 = n30422 | n30423 ;
  assign n46387 = ~n30424 ;
  assign n30913 = n46387 & n130 ;
  assign n30914 = n29849 | n30913 ;
  assign n30456 = n29849 & n46160 ;
  assign n46388 = ~n30423 ;
  assign n30457 = n46388 & n30456 ;
  assign n30917 = n30457 & n130 ;
  assign n46389 = ~n30917 ;
  assign n30918 = n30914 & n46389 ;
  assign n30404 = n30398 | n30399 ;
  assign n46390 = ~n30404 ;
  assign n30829 = n46390 & n130 ;
  assign n30830 = n29932 | n30829 ;
  assign n30432 = n29932 & n46144 ;
  assign n46391 = ~n30399 ;
  assign n30433 = n46391 & n30432 ;
  assign n30837 = n30433 & n130 ;
  assign n46392 = ~n30837 ;
  assign n30838 = n30830 & n46392 ;
  assign n30380 = n30374 | n30375 ;
  assign n46393 = ~n30380 ;
  assign n30804 = n46393 & n130 ;
  assign n30805 = n29923 | n30804 ;
  assign n30408 = n29923 & n46128 ;
  assign n46394 = ~n30375 ;
  assign n30409 = n46394 & n30408 ;
  assign n30839 = n30409 & n130 ;
  assign n46395 = ~n30839 ;
  assign n30840 = n30805 & n46395 ;
  assign n30384 = n29777 & n46112 ;
  assign n46396 = ~n30351 ;
  assign n30385 = n46396 & n30384 ;
  assign n30772 = n30385 & n130 ;
  assign n30356 = n30350 | n30351 ;
  assign n46397 = ~n30356 ;
  assign n30801 = n46397 & n130 ;
  assign n30802 = n29777 | n30801 ;
  assign n46398 = ~n30772 ;
  assign n30803 = n46398 & n30802 ;
  assign n30332 = n30326 | n30327 ;
  assign n46399 = ~n30332 ;
  assign n30799 = n46399 & n130 ;
  assign n30800 = n29837 | n30799 ;
  assign n30360 = n29837 & n46096 ;
  assign n46400 = ~n30327 ;
  assign n30361 = n46400 & n30360 ;
  assign n30910 = n30361 & n130 ;
  assign n46401 = ~n30910 ;
  assign n30911 = n30800 & n46401 ;
  assign n30336 = n29789 & n46080 ;
  assign n46402 = ~n30303 ;
  assign n30337 = n46402 & n30336 ;
  assign n30795 = n30337 & n130 ;
  assign n30308 = n30302 | n30303 ;
  assign n46403 = ~n30308 ;
  assign n30796 = n46403 & n130 ;
  assign n30797 = n29789 | n30796 ;
  assign n46404 = ~n30795 ;
  assign n30798 = n46404 & n30797 ;
  assign n30312 = n29800 & n46064 ;
  assign n46405 = ~n30279 ;
  assign n30313 = n46405 & n30312 ;
  assign n30790 = n30313 & n130 ;
  assign n30284 = n30278 | n30279 ;
  assign n46406 = ~n30284 ;
  assign n30792 = n46406 & n130 ;
  assign n30793 = n29800 | n30792 ;
  assign n46407 = ~n30790 ;
  assign n30794 = n46407 & n30793 ;
  assign n30260 = n30254 | n30255 ;
  assign n46408 = ~n30260 ;
  assign n30859 = n46408 & n130 ;
  assign n30860 = n29802 | n30859 ;
  assign n30288 = n29802 & n46048 ;
  assign n46409 = ~n30255 ;
  assign n30289 = n46409 & n30288 ;
  assign n30870 = n30289 & n130 ;
  assign n46410 = ~n30870 ;
  assign n30871 = n30860 & n46410 ;
  assign n30264 = n29860 & n46032 ;
  assign n46411 = ~n30231 ;
  assign n30265 = n46411 & n30264 ;
  assign n30780 = n30265 & n130 ;
  assign n30236 = n30230 | n30231 ;
  assign n46412 = ~n30236 ;
  assign n30785 = n46412 & n130 ;
  assign n30786 = n29860 | n30785 ;
  assign n46413 = ~n30780 ;
  assign n30787 = n46413 & n30786 ;
  assign n30212 = n30206 | n30207 ;
  assign n46414 = ~n30212 ;
  assign n30766 = n46414 & n130 ;
  assign n30767 = n29841 | n30766 ;
  assign n30240 = n29841 & n46016 ;
  assign n46415 = ~n30207 ;
  assign n30241 = n46415 & n30240 ;
  assign n30862 = n30241 & n130 ;
  assign n46416 = ~n30862 ;
  assign n30863 = n30767 & n46416 ;
  assign n30188 = n30182 | n30183 ;
  assign n46417 = ~n30188 ;
  assign n30777 = n46417 & n130 ;
  assign n30778 = n29879 | n30777 ;
  assign n30216 = n29879 & n46000 ;
  assign n46418 = ~n30183 ;
  assign n30217 = n46418 & n30216 ;
  assign n30868 = n30217 & n130 ;
  assign n46419 = ~n30868 ;
  assign n30869 = n30778 & n46419 ;
  assign n30192 = n30032 & n45984 ;
  assign n46420 = ~n30159 ;
  assign n30193 = n46420 & n30192 ;
  assign n30864 = n30193 & n130 ;
  assign n30164 = n30158 | n30159 ;
  assign n46421 = ~n30164 ;
  assign n30891 = n46421 & n130 ;
  assign n30892 = n30032 | n30891 ;
  assign n46422 = ~n30864 ;
  assign n30893 = n46422 & n30892 ;
  assign n30140 = n30134 | n30135 ;
  assign n46423 = ~n30140 ;
  assign n30773 = n46423 & n130 ;
  assign n30774 = n29916 | n30773 ;
  assign n30168 = n29916 & n45968 ;
  assign n46424 = ~n30135 ;
  assign n30169 = n46424 & n30168 ;
  assign n30823 = n30169 & n130 ;
  assign n46425 = ~n30823 ;
  assign n30824 = n30774 & n46425 ;
  assign n30116 = n30110 | n30111 ;
  assign n46426 = ~n30116 ;
  assign n30770 = n46426 & n130 ;
  assign n30771 = n29909 | n30770 ;
  assign n30144 = n29909 & n45952 ;
  assign n46427 = ~n30111 ;
  assign n30145 = n46427 & n30144 ;
  assign n30835 = n30145 & n130 ;
  assign n46428 = ~n30835 ;
  assign n30836 = n30771 & n46428 ;
  assign n30092 = n30086 | n30087 ;
  assign n46429 = ~n30092 ;
  assign n30768 = n46429 & n130 ;
  assign n30769 = n29892 | n30768 ;
  assign n30120 = n29892 & n45936 ;
  assign n46430 = ~n30087 ;
  assign n30121 = n46430 & n30120 ;
  assign n30889 = n30121 & n130 ;
  assign n46431 = ~n30889 ;
  assign n30890 = n30769 & n46431 ;
  assign n30070 = n30064 | n30065 ;
  assign n46432 = ~n30070 ;
  assign n30819 = n46432 & n130 ;
  assign n30820 = n29846 | n30819 ;
  assign n30096 = n29846 & n45920 ;
  assign n46433 = ~n30065 ;
  assign n30097 = n46433 & n30096 ;
  assign n30857 = n30097 & n130 ;
  assign n46434 = ~n30857 ;
  assign n30858 = n30820 & n46434 ;
  assign n30051 = n29884 & n45887 ;
  assign n46435 = ~n30056 ;
  assign n30735 = n30051 & n46435 ;
  assign n30763 = n30735 & n130 ;
  assign n30736 = n30050 | n30056 ;
  assign n46436 = ~n30736 ;
  assign n30999 = n46436 & n130 ;
  assign n31000 = n29884 | n30999 ;
  assign n46437 = ~n30763 ;
  assign n31001 = n46437 & n31000 ;
  assign n30022 = n29900 | n30018 ;
  assign n46438 = ~n30022 ;
  assign n30023 = n29876 & n46438 ;
  assign n30759 = n30023 & n130 ;
  assign n30894 = n46438 & n130 ;
  assign n30895 = n29876 | n30894 ;
  assign n46439 = ~n30759 ;
  assign n30896 = n46439 & n30895 ;
  assign n46440 = ~n266 ;
  assign n30762 = n46440 & n130 ;
  assign n46441 = ~n30743 ;
  assign n30744 = n131 & n46441 ;
  assign n46442 = ~n30756 ;
  assign n31012 = n30744 & n46442 ;
  assign n46443 = ~n30755 ;
  assign n31013 = n46443 & n31012 ;
  assign n31014 = n30762 | n31013 ;
  assign n31015 = x4 & n31014 ;
  assign n31016 = x4 | n31013 ;
  assign n31017 = n30762 | n31016 ;
  assign n46444 = ~n31015 ;
  assign n31018 = n46444 & n31017 ;
  assign n46445 = ~x2 ;
  assign n30903 = n46445 & n130 ;
  assign n46446 = ~n30903 ;
  assign n30904 = x3 & n46446 ;
  assign n30907 = n30762 | n30904 ;
  assign n269 = x0 | x1 ;
  assign n270 = n46445 & n269 ;
  assign n30745 = x2 & n46441 ;
  assign n31005 = n30745 & n46442 ;
  assign n31006 = n46443 & n31005 ;
  assign n31007 = n270 | n31006 ;
  assign n31008 = n30907 & n31007 ;
  assign n31009 = n30762 | n31007 ;
  assign n31010 = n30904 | n31009 ;
  assign n31019 = n45869 & n31010 ;
  assign n31020 = n31008 | n31019 ;
  assign n31021 = n31018 & n31020 ;
  assign n46447 = ~n131 ;
  assign n31011 = n46447 & n31010 ;
  assign n31023 = n31008 | n31011 ;
  assign n31024 = n31018 | n31023 ;
  assign n46448 = ~n132 ;
  assign n31025 = n46448 & n31024 ;
  assign n31026 = n31021 | n31025 ;
  assign n31027 = n30896 & n31026 ;
  assign n46449 = ~n30025 ;
  assign n30053 = n46449 & n30047 ;
  assign n46450 = ~n29904 ;
  assign n30054 = n46450 & n30053 ;
  assign n30844 = n30054 & n130 ;
  assign n30026 = n29904 | n30025 ;
  assign n46451 = ~n30026 ;
  assign n31002 = n46451 & n130 ;
  assign n31003 = n30047 | n31002 ;
  assign n46452 = ~n30844 ;
  assign n31004 = n46452 & n31003 ;
  assign n31022 = n30896 | n31021 ;
  assign n31028 = n31022 | n31025 ;
  assign n31029 = n44939 & n31028 ;
  assign n31030 = n31004 | n31029 ;
  assign n31031 = n31027 | n31030 ;
  assign n31032 = n44481 & n31031 ;
  assign n31033 = n31027 | n31029 ;
  assign n31034 = n31004 & n31033 ;
  assign n31035 = n31032 | n31034 ;
  assign n31036 = n31001 & n31035 ;
  assign n46453 = ~n30061 ;
  assign n30072 = n29855 & n46453 ;
  assign n30073 = n45893 & n30072 ;
  assign n30873 = n30073 & n130 ;
  assign n30071 = n30059 | n30061 ;
  assign n46454 = ~n30071 ;
  assign n30921 = n46454 & n130 ;
  assign n30922 = n29855 | n30921 ;
  assign n46455 = ~n30873 ;
  assign n30923 = n46455 & n30922 ;
  assign n31037 = n31001 | n31034 ;
  assign n31038 = n31032 | n31037 ;
  assign n31039 = n44023 & n31038 ;
  assign n31040 = n30923 | n31039 ;
  assign n31041 = n31036 | n31040 ;
  assign n46456 = ~n136 ;
  assign n31042 = n46456 & n31041 ;
  assign n31043 = n31036 | n31039 ;
  assign n31044 = n30923 & n31043 ;
  assign n31045 = n31042 | n31044 ;
  assign n31046 = n30858 & n31045 ;
  assign n46457 = ~n30083 ;
  assign n30094 = n29895 & n46457 ;
  assign n30095 = n45909 & n30094 ;
  assign n30791 = n30095 & n130 ;
  assign n30093 = n30068 | n30083 ;
  assign n46458 = ~n30093 ;
  assign n30928 = n46458 & n130 ;
  assign n30929 = n29895 | n30928 ;
  assign n46459 = ~n30791 ;
  assign n30930 = n46459 & n30929 ;
  assign n31047 = n30858 | n31044 ;
  assign n31048 = n31042 | n31047 ;
  assign n31049 = n43132 & n31048 ;
  assign n31050 = n30930 | n31049 ;
  assign n31051 = n31046 | n31050 ;
  assign n31052 = n42704 & n31051 ;
  assign n31053 = n31046 | n31049 ;
  assign n31054 = n30930 & n31053 ;
  assign n31055 = n31052 | n31054 ;
  assign n31056 = n30890 & n31055 ;
  assign n30117 = n30090 | n30107 ;
  assign n46460 = ~n30117 ;
  assign n30933 = n46460 & n130 ;
  assign n30934 = n30028 | n30933 ;
  assign n46461 = ~n30107 ;
  assign n30118 = n30028 & n46461 ;
  assign n30119 = n45925 & n30118 ;
  assign n30937 = n30119 & n130 ;
  assign n46462 = ~n30937 ;
  assign n30938 = n30934 & n46462 ;
  assign n31057 = n30890 | n31054 ;
  assign n31058 = n31052 | n31057 ;
  assign n31059 = n42281 & n31058 ;
  assign n31060 = n30938 | n31059 ;
  assign n31061 = n31056 | n31060 ;
  assign n46463 = ~n140 ;
  assign n31062 = n46463 & n31061 ;
  assign n31063 = n31056 | n31059 ;
  assign n31064 = n30938 & n31063 ;
  assign n31065 = n31062 | n31064 ;
  assign n31066 = n30836 & n31065 ;
  assign n46464 = ~n30131 ;
  assign n30142 = n29913 & n46464 ;
  assign n30143 = n45941 & n30142 ;
  assign n30879 = n30143 & n130 ;
  assign n30141 = n30114 | n30131 ;
  assign n46465 = ~n30141 ;
  assign n30939 = n46465 & n130 ;
  assign n30940 = n29913 | n30939 ;
  assign n46466 = ~n30879 ;
  assign n30941 = n46466 & n30940 ;
  assign n31067 = n30836 | n31064 ;
  assign n31068 = n31062 | n31067 ;
  assign n31069 = n41464 & n31068 ;
  assign n31070 = n30941 | n31069 ;
  assign n31071 = n31066 | n31070 ;
  assign n31072 = n41064 & n31071 ;
  assign n31073 = n31066 | n31069 ;
  assign n31074 = n30941 & n31073 ;
  assign n31075 = n31072 | n31074 ;
  assign n31076 = n30824 & n31075 ;
  assign n30165 = n30138 | n30155 ;
  assign n46467 = ~n30165 ;
  assign n30915 = n46467 & n130 ;
  assign n30916 = n29919 | n30915 ;
  assign n46468 = ~n30155 ;
  assign n30166 = n29919 & n46468 ;
  assign n30167 = n45957 & n30166 ;
  assign n30942 = n30167 & n130 ;
  assign n46469 = ~n30942 ;
  assign n30943 = n30916 & n46469 ;
  assign n31077 = n30824 | n31074 ;
  assign n31078 = n31072 | n31077 ;
  assign n31079 = n40664 & n31078 ;
  assign n31080 = n30943 | n31079 ;
  assign n31081 = n31076 | n31080 ;
  assign n46470 = ~n144 ;
  assign n31082 = n46470 & n31081 ;
  assign n31083 = n31076 | n31079 ;
  assign n31084 = n30943 & n31083 ;
  assign n31085 = n31082 | n31084 ;
  assign n31086 = n30893 & n31085 ;
  assign n30189 = n30162 | n30179 ;
  assign n46471 = ~n30189 ;
  assign n30815 = n46471 & n130 ;
  assign n30816 = n29907 | n30815 ;
  assign n46472 = ~n30179 ;
  assign n30190 = n29907 & n46472 ;
  assign n30191 = n45973 & n30190 ;
  assign n30817 = n30191 & n130 ;
  assign n46473 = ~n30817 ;
  assign n30818 = n30816 & n46473 ;
  assign n31087 = n30893 | n31084 ;
  assign n31088 = n31082 | n31087 ;
  assign n31089 = n39906 & n31088 ;
  assign n31090 = n30818 | n31089 ;
  assign n31091 = n31086 | n31090 ;
  assign n31092 = n39535 & n31091 ;
  assign n31093 = n31086 | n31089 ;
  assign n31094 = n30818 & n31093 ;
  assign n31095 = n31092 | n31094 ;
  assign n31096 = n30869 & n31095 ;
  assign n30213 = n30186 | n30203 ;
  assign n46474 = ~n30213 ;
  assign n30935 = n46474 & n130 ;
  assign n30936 = n29824 | n30935 ;
  assign n46475 = ~n30203 ;
  assign n30214 = n29824 & n46475 ;
  assign n30215 = n45989 & n30214 ;
  assign n30947 = n30215 & n130 ;
  assign n46476 = ~n30947 ;
  assign n30948 = n30936 & n46476 ;
  assign n31097 = n30869 | n31094 ;
  assign n31098 = n31092 | n31097 ;
  assign n31099 = n39174 & n31098 ;
  assign n31100 = n30948 | n31099 ;
  assign n31101 = n31096 | n31100 ;
  assign n46477 = ~n148 ;
  assign n31102 = n46477 & n31101 ;
  assign n31103 = n31096 | n31099 ;
  assign n31104 = n30948 & n31103 ;
  assign n31105 = n31102 | n31104 ;
  assign n31106 = n30863 & n31105 ;
  assign n30237 = n30210 | n30227 ;
  assign n46478 = ~n30237 ;
  assign n30874 = n46478 & n130 ;
  assign n30875 = n29814 | n30874 ;
  assign n46479 = ~n30227 ;
  assign n30238 = n29814 & n46479 ;
  assign n30239 = n46005 & n30238 ;
  assign n30949 = n30239 & n130 ;
  assign n46480 = ~n30949 ;
  assign n30950 = n30875 & n46480 ;
  assign n31107 = n30863 | n31104 ;
  assign n31108 = n31102 | n31107 ;
  assign n31109 = n38485 & n31108 ;
  assign n31110 = n30950 | n31109 ;
  assign n31111 = n31106 | n31110 ;
  assign n31112 = n38149 & n31111 ;
  assign n31113 = n31106 | n31109 ;
  assign n31114 = n30950 & n31113 ;
  assign n31115 = n31112 | n31114 ;
  assign n31116 = n30787 & n31115 ;
  assign n30261 = n30234 | n30251 ;
  assign n46481 = ~n30261 ;
  assign n30775 = n46481 & n130 ;
  assign n30776 = n29827 | n30775 ;
  assign n46482 = ~n30251 ;
  assign n30262 = n29827 & n46482 ;
  assign n30263 = n46021 & n30262 ;
  assign n30827 = n30263 & n130 ;
  assign n46483 = ~n30827 ;
  assign n30828 = n30776 & n46483 ;
  assign n31117 = n30787 | n31114 ;
  assign n31118 = n31112 | n31117 ;
  assign n31119 = n37821 & n31118 ;
  assign n31120 = n30828 | n31119 ;
  assign n31121 = n31116 | n31120 ;
  assign n46484 = ~n152 ;
  assign n31122 = n46484 & n31121 ;
  assign n31123 = n31116 | n31119 ;
  assign n31124 = n30828 & n31123 ;
  assign n31125 = n31122 | n31124 ;
  assign n31126 = n30871 & n31125 ;
  assign n30287 = n30258 | n30275 ;
  assign n46485 = ~n30287 ;
  assign n30931 = n46485 & n130 ;
  assign n30932 = n29870 | n30931 ;
  assign n46486 = ~n30275 ;
  assign n30285 = n29870 & n46486 ;
  assign n30286 = n46037 & n30285 ;
  assign n30951 = n30286 & n130 ;
  assign n46487 = ~n30951 ;
  assign n30952 = n30932 & n46487 ;
  assign n31127 = n30871 | n31124 ;
  assign n31128 = n31122 | n31127 ;
  assign n31129 = n37194 & n31128 ;
  assign n31130 = n30952 | n31129 ;
  assign n31131 = n31126 | n31130 ;
  assign n31132 = n36891 & n31131 ;
  assign n31133 = n31126 | n31129 ;
  assign n31134 = n30952 & n31133 ;
  assign n31135 = n31132 | n31134 ;
  assign n31136 = n30794 & n31135 ;
  assign n46488 = ~n30299 ;
  assign n30310 = n29810 & n46488 ;
  assign n30311 = n46053 & n30310 ;
  assign n30809 = n30311 & n130 ;
  assign n30309 = n30282 | n30299 ;
  assign n46489 = ~n30309 ;
  assign n30924 = n46489 & n130 ;
  assign n30925 = n29810 | n30924 ;
  assign n46490 = ~n30809 ;
  assign n30926 = n46490 & n30925 ;
  assign n31137 = n30794 | n31134 ;
  assign n31138 = n31132 | n31137 ;
  assign n31139 = n36600 & n31138 ;
  assign n31140 = n30926 | n31139 ;
  assign n31141 = n31136 | n31140 ;
  assign n46491 = ~n156 ;
  assign n31142 = n46491 & n31141 ;
  assign n31143 = n31136 | n31139 ;
  assign n31144 = n30926 & n31143 ;
  assign n31145 = n31142 | n31144 ;
  assign n31146 = n30798 & n31145 ;
  assign n30333 = n30306 | n30323 ;
  assign n46492 = ~n30333 ;
  assign n30848 = n46492 & n130 ;
  assign n30849 = n29881 | n30848 ;
  assign n46493 = ~n30323 ;
  assign n30334 = n29881 & n46493 ;
  assign n30335 = n46069 & n30334 ;
  assign n30884 = n30335 & n130 ;
  assign n46494 = ~n30884 ;
  assign n30885 = n30849 & n46494 ;
  assign n31147 = n30798 | n31144 ;
  assign n31148 = n31142 | n31147 ;
  assign n31149 = n36042 & n31148 ;
  assign n31150 = n30885 | n31149 ;
  assign n31151 = n31146 | n31150 ;
  assign n31152 = n35770 & n31151 ;
  assign n31153 = n31146 | n31149 ;
  assign n31154 = n30885 & n31153 ;
  assign n31155 = n31152 | n31154 ;
  assign n31156 = n30911 & n31155 ;
  assign n30357 = n30330 | n30347 ;
  assign n46495 = ~n30357 ;
  assign n30806 = n46495 & n130 ;
  assign n30807 = n29868 | n30806 ;
  assign n46496 = ~n30347 ;
  assign n30358 = n29868 & n46496 ;
  assign n30359 = n46085 & n30358 ;
  assign n30953 = n30359 & n130 ;
  assign n46497 = ~n30953 ;
  assign n30954 = n30807 & n46497 ;
  assign n31157 = n30911 | n31154 ;
  assign n31158 = n31152 | n31157 ;
  assign n31159 = n35503 & n31158 ;
  assign n31160 = n30954 | n31159 ;
  assign n31161 = n31156 | n31160 ;
  assign n46498 = ~n160 ;
  assign n31162 = n46498 & n31161 ;
  assign n31163 = n31156 | n31159 ;
  assign n31164 = n30954 & n31163 ;
  assign n31165 = n31162 | n31164 ;
  assign n31166 = n30803 & n31165 ;
  assign n46499 = ~n30371 ;
  assign n30382 = n29897 & n46499 ;
  assign n30383 = n46101 & n30382 ;
  assign n30912 = n30383 & n130 ;
  assign n30381 = n30354 | n30371 ;
  assign n46500 = ~n30381 ;
  assign n30944 = n46500 & n130 ;
  assign n30945 = n29897 | n30944 ;
  assign n46501 = ~n30912 ;
  assign n30946 = n46501 & n30945 ;
  assign n31167 = n30803 | n31164 ;
  assign n31168 = n31162 | n31167 ;
  assign n31169 = n35001 & n31168 ;
  assign n31170 = n30946 | n31169 ;
  assign n31171 = n31166 | n31170 ;
  assign n31172 = n34762 & n31171 ;
  assign n31173 = n31166 | n31169 ;
  assign n31174 = n30946 & n31173 ;
  assign n31175 = n31172 | n31174 ;
  assign n31176 = n30840 & n31175 ;
  assign n46502 = ~n30395 ;
  assign n30406 = n29927 & n46502 ;
  assign n30407 = n46117 & n30406 ;
  assign n30927 = n30407 & n130 ;
  assign n30405 = n30378 | n30395 ;
  assign n46503 = ~n30405 ;
  assign n30955 = n46503 & n130 ;
  assign n30956 = n29927 | n30955 ;
  assign n46504 = ~n30927 ;
  assign n30957 = n46504 & n30956 ;
  assign n31177 = n30840 | n31174 ;
  assign n31178 = n31172 | n31177 ;
  assign n31179 = n34532 & n31178 ;
  assign n31180 = n30957 | n31179 ;
  assign n31181 = n31176 | n31180 ;
  assign n46505 = ~n164 ;
  assign n31182 = n46505 & n31181 ;
  assign n31183 = n31176 | n31179 ;
  assign n31184 = n30957 & n31183 ;
  assign n31185 = n31182 | n31184 ;
  assign n31186 = n30838 & n31185 ;
  assign n46506 = ~n30419 ;
  assign n30430 = n29939 & n46506 ;
  assign n30431 = n46133 & n30430 ;
  assign n30822 = n30431 & n130 ;
  assign n30429 = n30402 | n30419 ;
  assign n46507 = ~n30429 ;
  assign n30886 = n46507 & n130 ;
  assign n30887 = n29939 | n30886 ;
  assign n46508 = ~n30822 ;
  assign n30888 = n46508 & n30887 ;
  assign n31187 = n30838 | n31184 ;
  assign n31188 = n31182 | n31187 ;
  assign n31189 = n34101 & n31188 ;
  assign n31190 = n30888 | n31189 ;
  assign n31191 = n31186 | n31190 ;
  assign n31192 = n33894 & n31191 ;
  assign n31193 = n31186 | n31189 ;
  assign n31194 = n30888 & n31193 ;
  assign n31195 = n31192 | n31194 ;
  assign n31196 = n30918 & n31195 ;
  assign n30453 = n30427 | n30443 ;
  assign n46509 = ~n30453 ;
  assign n30958 = n46509 & n130 ;
  assign n30959 = n29945 | n30958 ;
  assign n46510 = ~n30443 ;
  assign n30454 = n29945 & n46510 ;
  assign n30455 = n46149 & n30454 ;
  assign n30960 = n30455 & n130 ;
  assign n46511 = ~n30960 ;
  assign n30961 = n30959 & n46511 ;
  assign n31197 = n30918 | n31194 ;
  assign n31198 = n31192 | n31197 ;
  assign n31199 = n33697 & n31198 ;
  assign n31200 = n30961 | n31199 ;
  assign n31201 = n31196 | n31200 ;
  assign n46512 = ~n168 ;
  assign n31202 = n46512 & n31201 ;
  assign n31203 = n31196 | n31199 ;
  assign n31204 = n30961 & n31203 ;
  assign n31205 = n31202 | n31204 ;
  assign n31206 = n30855 & n31205 ;
  assign n30479 = n30450 | n30467 ;
  assign n46513 = ~n30479 ;
  assign n30962 = n46513 & n130 ;
  assign n30963 = n29950 | n30962 ;
  assign n46514 = ~n30467 ;
  assign n30477 = n29950 & n46514 ;
  assign n30478 = n46165 & n30477 ;
  assign n30964 = n30478 & n130 ;
  assign n46515 = ~n30964 ;
  assign n30965 = n30963 & n46515 ;
  assign n31207 = n30855 | n31204 ;
  assign n31208 = n31202 | n31207 ;
  assign n31209 = n33337 & n31208 ;
  assign n31210 = n30965 | n31209 ;
  assign n31211 = n31206 | n31210 ;
  assign n31212 = n33162 & n31211 ;
  assign n31213 = n31206 | n31209 ;
  assign n31214 = n30965 & n31213 ;
  assign n31215 = n31212 | n31214 ;
  assign n31216 = n30906 & n31215 ;
  assign n46516 = ~n30491 ;
  assign n30502 = n29961 & n46516 ;
  assign n30503 = n46181 & n30502 ;
  assign n30919 = n30503 & n130 ;
  assign n30501 = n30474 | n30491 ;
  assign n46517 = ~n30501 ;
  assign n30966 = n46517 & n130 ;
  assign n30967 = n29961 | n30966 ;
  assign n46518 = ~n30919 ;
  assign n30968 = n46518 & n30967 ;
  assign n31217 = n30906 | n31214 ;
  assign n31218 = n31212 | n31217 ;
  assign n31219 = n32993 & n31218 ;
  assign n31220 = n30968 | n31219 ;
  assign n31221 = n31216 | n31220 ;
  assign n46519 = ~n172 ;
  assign n31222 = n46519 & n31221 ;
  assign n31223 = n31216 | n31219 ;
  assign n31224 = n30968 & n31223 ;
  assign n31225 = n31222 | n31224 ;
  assign n31226 = n30899 & n31225 ;
  assign n30525 = n30498 | n30515 ;
  assign n46520 = ~n30525 ;
  assign n30969 = n46520 & n130 ;
  assign n30970 = n29968 | n30969 ;
  assign n46521 = ~n30515 ;
  assign n30526 = n29968 & n46521 ;
  assign n30527 = n46197 & n30526 ;
  assign n30971 = n30527 & n130 ;
  assign n46522 = ~n30971 ;
  assign n30972 = n30970 & n46522 ;
  assign n31227 = n30899 | n31224 ;
  assign n31228 = n31222 | n31227 ;
  assign n31229 = n32693 & n31228 ;
  assign n31230 = n30972 | n31229 ;
  assign n31231 = n31226 | n31230 ;
  assign n31232 = n32554 & n31231 ;
  assign n31233 = n31226 | n31229 ;
  assign n31234 = n30972 & n31233 ;
  assign n31235 = n31232 | n31234 ;
  assign n31236 = n30847 & n31235 ;
  assign n46523 = ~n30539 ;
  assign n30550 = n29975 & n46523 ;
  assign n30551 = n46213 & n30550 ;
  assign n30920 = n30551 & n130 ;
  assign n30549 = n30523 | n30539 ;
  assign n46524 = ~n30549 ;
  assign n30975 = n46524 & n130 ;
  assign n30976 = n29975 | n30975 ;
  assign n46525 = ~n30920 ;
  assign n30977 = n46525 & n30976 ;
  assign n31237 = n30847 | n31234 ;
  assign n31238 = n31232 | n31237 ;
  assign n31239 = n32418 & n31238 ;
  assign n31240 = n30977 | n31239 ;
  assign n31241 = n31236 | n31240 ;
  assign n46526 = ~n176 ;
  assign n31242 = n46526 & n31241 ;
  assign n31243 = n31236 | n31239 ;
  assign n31244 = n30977 & n31243 ;
  assign n31245 = n31242 | n31244 ;
  assign n31246 = n30782 & n31245 ;
  assign n46527 = ~n30563 ;
  assign n30574 = n29979 & n46527 ;
  assign n30575 = n46229 & n30574 ;
  assign n30856 = n30575 & n130 ;
  assign n30573 = n30546 | n30563 ;
  assign n46528 = ~n30573 ;
  assign n30978 = n46528 & n130 ;
  assign n30979 = n29979 | n30978 ;
  assign n46529 = ~n30856 ;
  assign n30980 = n46529 & n30979 ;
  assign n31247 = n30782 | n31244 ;
  assign n31248 = n31242 | n31247 ;
  assign n31249 = n32175 & n31248 ;
  assign n31250 = n30980 | n31249 ;
  assign n31251 = n31246 | n31250 ;
  assign n31252 = n32065 & n31251 ;
  assign n31253 = n31246 | n31249 ;
  assign n31254 = n30980 & n31253 ;
  assign n31255 = n31252 | n31254 ;
  assign n31256 = n30902 & n31255 ;
  assign n46530 = ~n30587 ;
  assign n30597 = n29986 & n46530 ;
  assign n30598 = n46245 & n30597 ;
  assign n30865 = n30598 & n130 ;
  assign n30599 = n30570 | n30587 ;
  assign n46531 = ~n30599 ;
  assign n30981 = n46531 & n130 ;
  assign n30982 = n29986 | n30981 ;
  assign n46532 = ~n30865 ;
  assign n30983 = n46532 & n30982 ;
  assign n31257 = n30902 | n31254 ;
  assign n31258 = n31252 | n31257 ;
  assign n31259 = n31951 & n31258 ;
  assign n31260 = n30983 | n31259 ;
  assign n31261 = n31256 | n31260 ;
  assign n46533 = ~n180 ;
  assign n31262 = n46533 & n31261 ;
  assign n31263 = n31256 | n31259 ;
  assign n31264 = n30983 & n31263 ;
  assign n31265 = n31262 | n31264 ;
  assign n31266 = n30814 & n31265 ;
  assign n46534 = ~n30611 ;
  assign n30622 = n29936 & n46534 ;
  assign n30623 = n46261 & n30622 ;
  assign n30850 = n30623 & n130 ;
  assign n30621 = n30594 | n30611 ;
  assign n46535 = ~n30621 ;
  assign n30984 = n46535 & n130 ;
  assign n30985 = n29936 | n30984 ;
  assign n46536 = ~n30850 ;
  assign n30986 = n46536 & n30985 ;
  assign n31267 = n30814 | n31264 ;
  assign n31268 = n31262 | n31267 ;
  assign n31269 = n31788 & n31268 ;
  assign n31270 = n30986 | n31269 ;
  assign n31271 = n31266 | n31270 ;
  assign n31272 = n31705 & n31271 ;
  assign n31273 = n31266 | n31269 ;
  assign n31274 = n30986 & n31273 ;
  assign n31275 = n31272 | n31274 ;
  assign n31276 = n30843 & n31275 ;
  assign n46537 = ~n30635 ;
  assign n30645 = n29954 & n46537 ;
  assign n30646 = n46277 & n30645 ;
  assign n30779 = n30646 & n130 ;
  assign n30647 = n30618 | n30635 ;
  assign n46538 = ~n30647 ;
  assign n30990 = n46538 & n130 ;
  assign n30991 = n29954 | n30990 ;
  assign n46539 = ~n30779 ;
  assign n30992 = n46539 & n30991 ;
  assign n31277 = n30843 | n31274 ;
  assign n31278 = n31272 | n31277 ;
  assign n31279 = n31624 & n31278 ;
  assign n31280 = n30992 | n31279 ;
  assign n31281 = n31276 | n31280 ;
  assign n46540 = ~n184 ;
  assign n31282 = n46540 & n31281 ;
  assign n31283 = n31276 | n31279 ;
  assign n31284 = n30992 & n31283 ;
  assign n31285 = n31282 | n31284 ;
  assign n31286 = n30867 & n31285 ;
  assign n46541 = ~n30659 ;
  assign n30670 = n30040 & n46541 ;
  assign n30671 = n46293 & n30670 ;
  assign n30973 = n30671 & n130 ;
  assign n30669 = n30642 | n30659 ;
  assign n46542 = ~n30669 ;
  assign n30987 = n46542 & n130 ;
  assign n30988 = n30040 | n30987 ;
  assign n46543 = ~n30973 ;
  assign n30989 = n46543 & n30988 ;
  assign n31287 = n30867 | n31284 ;
  assign n31288 = n31282 | n31287 ;
  assign n31289 = n31523 & n31288 ;
  assign n31290 = n30989 | n31289 ;
  assign n31291 = n31286 | n31290 ;
  assign n31292 = n31468 & n31291 ;
  assign n31293 = n31286 | n31289 ;
  assign n31294 = n30989 & n31293 ;
  assign n31295 = n31292 | n31294 ;
  assign n31296 = n30833 & n31295 ;
  assign n30693 = n30666 | n30683 ;
  assign n46544 = ~n30693 ;
  assign n30908 = n46544 & n130 ;
  assign n30909 = n30001 | n30908 ;
  assign n46545 = ~n30683 ;
  assign n30694 = n30001 & n46545 ;
  assign n30695 = n46309 & n30694 ;
  assign n30993 = n30695 & n130 ;
  assign n46546 = ~n30993 ;
  assign n30994 = n30909 & n46546 ;
  assign n31297 = n30833 | n31294 ;
  assign n31298 = n31292 | n31297 ;
  assign n31299 = n31420 & n31298 ;
  assign n31300 = n30994 | n31299 ;
  assign n31301 = n31296 | n31300 ;
  assign n46547 = ~n188 ;
  assign n31302 = n46547 & n31301 ;
  assign n31303 = n31296 | n31299 ;
  assign n31304 = n30994 & n31303 ;
  assign n31305 = n31302 | n31304 ;
  assign n31306 = n30883 & n31305 ;
  assign n30717 = n30690 | n30707 ;
  assign n46548 = ~n30717 ;
  assign n30783 = n46548 & n130 ;
  assign n30784 = n30003 | n30783 ;
  assign n46549 = ~n30707 ;
  assign n30718 = n30003 & n46549 ;
  assign n30719 = n46325 & n30718 ;
  assign n30810 = n30719 & n130 ;
  assign n46550 = ~n30810 ;
  assign n30811 = n30784 & n46550 ;
  assign n31307 = n30883 | n31304 ;
  assign n31308 = n31302 | n31307 ;
  assign n31309 = n31383 & n31308 ;
  assign n31310 = n30811 | n31309 ;
  assign n31311 = n31306 | n31310 ;
  assign n31312 = n31357 & n31311 ;
  assign n31313 = n31306 | n31309 ;
  assign n31314 = n30811 & n31313 ;
  assign n31315 = n31312 | n31314 ;
  assign n31316 = n30878 & n31315 ;
  assign n31317 = n30878 | n31314 ;
  assign n31318 = n31312 | n31317 ;
  assign n46551 = ~n191 ;
  assign n31319 = n46551 & n31318 ;
  assign n31320 = n31316 | n31319 ;
  assign n46552 = ~n30731 ;
  assign n30748 = n46552 & n30747 ;
  assign n30749 = n46342 & n30748 ;
  assign n30834 = n30749 & n130 ;
  assign n30732 = n30714 | n30731 ;
  assign n46553 = ~n30732 ;
  assign n30995 = n46553 & n130 ;
  assign n31322 = n30747 | n30995 ;
  assign n46554 = ~n30834 ;
  assign n31323 = n46554 & n31322 ;
  assign n31324 = n31320 & n31323 ;
  assign n31325 = n30998 | n31324 ;
  assign n46555 = ~n30752 ;
  assign n30974 = n46555 & n130 ;
  assign n31321 = n30756 | n30974 ;
  assign n31326 = n31321 | n31323 ;
  assign n31327 = n31319 | n31326 ;
  assign n31328 = n31316 | n31327 ;
  assign n31329 = n31336 & n31328 ;
  assign n129 = n31325 | n31329 ;
  assign y0 = n129 ;
  assign y1 = n130 ;
  assign y2 = n131 ;
  assign y3 = n132 ;
  assign y4 = n133 ;
  assign y5 = n134 ;
  assign y6 = n135 ;
  assign y7 = n136 ;
  assign y8 = n137 ;
  assign y9 = n138 ;
  assign y10 = n139 ;
  assign y11 = n140 ;
  assign y12 = n141 ;
  assign y13 = n142 ;
  assign y14 = n143 ;
  assign y15 = n144 ;
  assign y16 = n145 ;
  assign y17 = n146 ;
  assign y18 = n147 ;
  assign y19 = n148 ;
  assign y20 = n149 ;
  assign y21 = n150 ;
  assign y22 = n151 ;
  assign y23 = n152 ;
  assign y24 = n153 ;
  assign y25 = n154 ;
  assign y26 = n155 ;
  assign y27 = n156 ;
  assign y28 = n157 ;
  assign y29 = n158 ;
  assign y30 = n159 ;
  assign y31 = n160 ;
  assign y32 = n161 ;
  assign y33 = n162 ;
  assign y34 = n163 ;
  assign y35 = n164 ;
  assign y36 = n165 ;
  assign y37 = n166 ;
  assign y38 = n167 ;
  assign y39 = n168 ;
  assign y40 = n169 ;
  assign y41 = n170 ;
  assign y42 = n171 ;
  assign y43 = n172 ;
  assign y44 = n173 ;
  assign y45 = n174 ;
  assign y46 = n175 ;
  assign y47 = n176 ;
  assign y48 = n177 ;
  assign y49 = n178 ;
  assign y50 = n179 ;
  assign y51 = n180 ;
  assign y52 = n181 ;
  assign y53 = n182 ;
  assign y54 = n183 ;
  assign y55 = n184 ;
  assign y56 = n185 ;
  assign y57 = n186 ;
  assign y58 = n187 ;
  assign y59 = n188 ;
  assign y60 = n189 ;
  assign y61 = n190 ;
  assign y62 = n191 ;
  assign y63 = n192 ;
endmodule
