module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 ;
  assign n12 = ~x6 & x10 ;
  assign n13 = x7 & n12 ;
  assign n14 = x9 & x10 ;
  assign n15 = x8 & n14 ;
  assign n16 = x3 ^ x2 ^ 1'b0 ;
  assign n17 = ~x9 & n16 ;
  assign n18 = ~x8 & n17 ;
  assign n19 = x10 | n18 ;
  assign n20 = ~x7 & n19 ;
  assign n21 = n15 | n20 ;
  assign n22 = x6 & n21 ;
  assign n23 = n13 | n22 ;
  assign n24 = x7 | x8 ;
  assign n25 = ~x1 & x2 ;
  assign n26 = ~n24 & n25 ;
  assign n27 = x9 | n26 ;
  assign n28 = x4 & ~x8 ;
  assign n29 = ~x3 & n28 ;
  assign n30 = x4 | x7 ;
  assign n31 = ~n29 & n30 ;
  assign n32 = x2 | n31 ;
  assign n33 = x1 & ~n32 ;
  assign n34 = n27 | n33 ;
  assign n35 = ~x6 & n34 ;
  assign n36 = x5 & n35 ;
  assign n37 = x6 & x9 ;
  assign n38 = ~x5 & n37 ;
  assign n39 = n36 | n38 ;
  assign n40 = x1 & ~x2 ;
  assign n41 = x5 & ~x7 ;
  assign n42 = n40 & n41 ;
  assign n43 = ~x4 & x7 ;
  assign n44 = n42 | n43 ;
  assign n45 = x3 & n44 ;
  assign n46 = x3 & x4 ;
  assign n47 = x7 & ~n46 ;
  assign n48 = n47 ^ n30 ^ x4 ;
  assign n49 = n45 | n48 ;
  assign n50 = ~x8 & n49 ;
  assign n51 = ~x4 & x8 ;
  assign n52 = ~x4 & x5 ;
  assign n53 = ( x4 & n51 ) | ( x4 & n52 ) | ( n51 & n52 ) ;
  assign n54 = n50 | n53 ;
  assign n55 = x1 & x4 ;
  assign n56 = x0 | n55 ;
  assign n57 = ( x0 & n51 ) | ( x0 & n55 ) | ( n51 & n55 ) ;
  assign n58 = n56 & ~n57 ;
  assign n59 = ~x6 & n58 ;
  assign n60 = ~x7 & n59 ;
  assign n61 = x4 & x8 ;
  assign n62 = n60 | n61 ;
  assign n63 = ~x5 & n62 ;
  assign n64 = n54 | n63 ;
  assign n65 = ~x9 & n64 ;
  assign n66 = n39 | n65 ;
  assign n67 = ~x10 & n66 ;
  assign n68 = n23 | n67 ;
  assign n69 = x8 & ~x9 ;
  assign n70 = x6 & x10 ;
  assign n71 = x7 & n70 ;
  assign n72 = n69 & n71 ;
  assign n73 = x6 & ~x9 ;
  assign n74 = x4 & ~x6 ;
  assign n75 = x3 & ~x6 ;
  assign n76 = ~x2 & n75 ;
  assign n77 = x3 & x6 ;
  assign n78 = x2 & n46 ;
  assign n79 = ( n76 & n77 ) | ( n76 & n78 ) | ( n77 & n78 ) ;
  assign n80 = ( n73 & n74 ) | ( n73 & n79 ) | ( n74 & n79 ) ;
  assign n81 = x10 | n80 ;
  assign n82 = ~x4 & n73 ;
  assign n83 = x5 & ~x6 ;
  assign n84 = ~x1 & n83 ;
  assign n85 = ( ~x3 & n82 ) | ( ~x3 & n84 ) | ( n82 & n84 ) ;
  assign n86 = n81 | n85 ;
  assign n87 = ~x3 & n83 ;
  assign n88 = n82 | n87 ;
  assign n89 = ~x2 & n88 ;
  assign n90 = n86 | n89 ;
  assign n91 = ~x7 & n90 ;
  assign n92 = n12 | n91 ;
  assign n93 = ~x8 & n92 ;
  assign n94 = n72 | n93 ;
  assign n96 = ~x7 & x9 ;
  assign n95 = x4 & n69 ;
  assign n97 = n96 ^ n95 ^ n69 ;
  assign n98 = ~x6 & n97 ;
  assign n99 = x7 & ~x9 ;
  assign n100 = n99 ^ n95 ^ x7 ;
  assign n101 = x6 & n100 ;
  assign n102 = n28 & n99 ;
  assign n103 = x6 | x7 ;
  assign n104 = x4 | n103 ;
  assign n105 = x4 | x9 ;
  assign n106 = n105 ^ n95 ^ x9 ;
  assign n107 = n104 & ~n106 ;
  assign n108 = x2 & ~n107 ;
  assign n109 = x1 & n108 ;
  assign n110 = n102 | n109 ;
  assign n111 = x3 & n110 ;
  assign n112 = n101 | n111 ;
  assign n113 = x5 & n112 ;
  assign n114 = n98 | n113 ;
  assign n115 = ~x9 & n47 ;
  assign n116 = ~x8 & n115 ;
  assign n117 = n96 | n116 ;
  assign n118 = x1 & x2 ;
  assign n119 = x0 & ~n118 ;
  assign n120 = ~x0 & x2 ;
  assign n121 = n119 | n120 ;
  assign n122 = x7 | n121 ;
  assign n123 = x4 & ~n122 ;
  assign n124 = n69 | n123 ;
  assign n125 = x2 | x7 ;
  assign n126 = n105 & n125 ;
  assign n127 = x1 | n126 ;
  assign n128 = ~n124 & n127 ;
  assign n129 = x6 | n128 ;
  assign n130 = ~n117 & n129 ;
  assign n131 = x5 | n130 ;
  assign n132 = ~n114 & n131 ;
  assign n133 = x10 | n132 ;
  assign n134 = ~n94 & n133 ;
  assign n135 = x5 & x7 ;
  assign n136 = x8 & ~n135 ;
  assign n137 = x10 | n136 ;
  assign n138 = x9 & n137 ;
  assign n139 = ~x8 & x9 ;
  assign n140 = x5 & n139 ;
  assign n141 = x8 & x10 ;
  assign n142 = n140 | n141 ;
  assign n143 = x7 & n142 ;
  assign n144 = x6 & n143 ;
  assign n145 = n138 | n144 ;
  assign n146 = x6 & ~x7 ;
  assign n147 = ~x2 & n146 ;
  assign n148 = ~x6 & x7 ;
  assign n149 = x3 & n148 ;
  assign n150 = n147 | n149 ;
  assign n151 = x5 & n150 ;
  assign n152 = x4 & n151 ;
  assign n153 = ~x5 & x6 ;
  assign n154 = x6 & x7 ;
  assign n155 = ( n43 & n153 ) | ( n43 & n154 ) | ( n153 & n154 ) ;
  assign n156 = n152 | n155 ;
  assign n157 = x2 & n153 ;
  assign n158 = n84 | n157 ;
  assign n159 = x4 & n158 ;
  assign n160 = x3 & n159 ;
  assign n161 = ~x3 & x5 ;
  assign n162 = x3 & n52 ;
  assign n163 = x5 & x6 ;
  assign n164 = ( n161 & n162 ) | ( n161 & n163 ) | ( n162 & n163 ) ;
  assign n165 = n160 | n164 ;
  assign n166 = n76 | n161 ;
  assign n167 = x4 & n166 ;
  assign n168 = x0 & x1 ;
  assign n169 = x4 & ~n168 ;
  assign n170 = x3 & n169 ;
  assign n171 = x4 | x6 ;
  assign n172 = ~n170 & n171 ;
  assign n173 = x5 | n172 ;
  assign n174 = x0 & ~x3 ;
  assign n175 = n74 & n174 ;
  assign n176 = n162 | n175 ;
  assign n177 = x1 & n176 ;
  assign n178 = n173 & ~n177 ;
  assign n179 = x2 & ~n178 ;
  assign n180 = n167 | n179 ;
  assign n181 = ~x7 & n180 ;
  assign n182 = n165 | n181 ;
  assign n183 = ~x8 & n182 ;
  assign n184 = n156 | n183 ;
  assign n185 = ~x9 & n184 ;
  assign n186 = x4 & x6 ;
  assign n187 = ( n41 & n148 ) | ( n41 & n186 ) | ( n148 & n186 ) ;
  assign n188 = ( x8 & n148 ) | ( x8 & n187 ) | ( n148 & n187 ) ;
  assign n189 = n185 | n188 ;
  assign n190 = ~x10 & n189 ;
  assign n191 = n145 | n190 ;
  assign n192 = x4 | x8 ;
  assign n193 = x5 | n192 ;
  assign n194 = n103 | n193 ;
  assign n195 = ~x2 & n154 ;
  assign n196 = x5 & n61 ;
  assign n197 = n195 & n196 ;
  assign n198 = n194 & ~n197 ;
  assign n199 = x9 | n198 ;
  assign n200 = x10 | n199 ;
  assign n201 = x3 | n200 ;
  assign n202 = x5 | x6 ;
  assign n203 = n168 & ~n202 ;
  assign n204 = n187 | n203 ;
  assign n205 = x3 & n204 ;
  assign n206 = x2 & n205 ;
  assign n207 = x4 | n146 ;
  assign n208 = ( n40 & n83 ) | ( n40 & n84 ) | ( n83 & n84 ) ;
  assign n209 = x9 | n208 ;
  assign n210 = x7 & ~n163 ;
  assign n211 = n209 | n210 ;
  assign n212 = ( ~x3 & x7 ) | ( ~x3 & n87 ) | ( x7 & n87 ) ;
  assign n213 = n211 | n212 ;
  assign n214 = n207 & ~n213 ;
  assign n215 = ~n206 & n214 ;
  assign n216 = x8 | n215 ;
  assign n217 = ( x2 & x8 ) | ( x2 & n16 ) | ( x8 & n16 ) ;
  assign n218 = x6 & n217 ;
  assign n219 = x5 & n218 ;
  assign n220 = x7 & n219 ;
  assign n221 = ~x9 & n220 ;
  assign n222 = x4 & n221 ;
  assign n223 = ( x9 & n96 ) | ( x9 & n210 ) | ( n96 & n210 ) ;
  assign n224 = n222 | n223 ;
  assign n225 = n216 & ~n224 ;
  assign n226 = x10 | n225 ;
  assign n227 = x9 | x10 ;
  assign n228 = n78 & n163 ;
  assign n229 = n228 ^ n83 ^ x6 ;
  assign n230 = ~x7 & n229 ;
  assign n231 = ~x8 & n230 ;
  assign n232 = n227 | n231 ;
  assign n233 = x6 & x8 ;
  assign n234 = n135 & n233 ;
  assign n235 = x1 & x3 ;
  assign n236 = x0 & n235 ;
  assign n237 = x5 | x7 ;
  assign n238 = x8 | n237 ;
  assign n239 = n236 & ~n238 ;
  assign n240 = n234 | n239 ;
  assign n241 = x2 & n240 ;
  assign n242 = ( n75 & n77 ) | ( n75 & n234 ) | ( n77 & n234 ) ;
  assign n243 = n241 | n242 ;
  assign n244 = x4 & n243 ;
  assign n245 = n232 | n244 ;
  assign n246 = x9 | n228 ;
  assign n247 = x10 | n246 ;
  assign n248 = n24 | n247 ;
  assign y0 = n68 ;
  assign y1 = n134 ;
  assign y2 = n191 ;
  assign y3 = n201 ;
  assign y4 = n226 ;
  assign y5 = n245 ;
  assign y6 = n248 ;
endmodule
