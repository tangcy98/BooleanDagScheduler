module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 ;
  assign n25 = x0 | x1 ;
  assign n26 = x2 & n25 ;
  assign n27 = n26 ^ n25 ^ x2 ;
  assign n28 = x3 | n27 ;
  assign n29 = x4 | n28 ;
  assign n30 = x5 | n29 ;
  assign n31 = x6 | n30 ;
  assign n32 = x7 | n31 ;
  assign n33 = x8 | n32 ;
  assign n34 = x9 | n33 ;
  assign n35 = x10 | n34 ;
  assign n36 = x11 | n35 ;
  assign n37 = x12 | n36 ;
  assign n38 = x13 | n37 ;
  assign n39 = x14 | n38 ;
  assign n40 = ~x22 & n37 ;
  assign n41 = ( ~x22 & n39 ) | ( ~x22 & n40 ) | ( n39 & n40 ) ;
  assign n42 = n41 ^ x15 ^ 1'b0 ;
  assign n43 = x15 | n39 ;
  assign n44 = x16 | n43 ;
  assign n45 = x17 | n44 ;
  assign n46 = x18 | n45 ;
  assign n47 = x19 | n46 ;
  assign n48 = x20 | n47 ;
  assign n49 = n48 ^ x21 ^ 1'b0 ;
  assign n50 = n49 ^ x22 ^ 1'b0 ;
  assign n51 = ( x21 & n49 ) | ( x21 & n50 ) | ( n49 & n50 ) ;
  assign n52 = n47 ^ x20 ^ 1'b0 ;
  assign n53 = n52 ^ x22 ^ 1'b0 ;
  assign n54 = ( x20 & n52 ) | ( x20 & n53 ) | ( n52 & n53 ) ;
  assign n55 = n51 & ~n54 ;
  assign n56 = ~n42 & n55 ;
  assign n57 = ~x22 & n46 ;
  assign n58 = n57 ^ x19 ^ 1'b0 ;
  assign n59 = ~x22 & n44 ;
  assign n60 = n59 ^ x17 ^ 1'b0 ;
  assign n61 = ( ~x22 & n59 ) | ( ~x22 & n60 ) | ( n59 & n60 ) ;
  assign n62 = n61 ^ x18 ^ 1'b0 ;
  assign n63 = n58 & ~n62 ;
  assign n64 = ~x22 & n43 ;
  assign n65 = n64 ^ x16 ^ 1'b0 ;
  assign n66 = ~n60 & n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = n56 & n67 ;
  assign n69 = n42 & n55 ;
  assign n70 = n58 & n62 ;
  assign n71 = n66 & n70 ;
  assign n72 = n69 & n71 ;
  assign n73 = n68 | n72 ;
  assign n74 = n58 | n62 ;
  assign n75 = n66 & ~n74 ;
  assign n76 = n51 | n54 ;
  assign n77 = n42 & ~n76 ;
  assign n78 = n75 & n77 ;
  assign n79 = n60 & ~n65 ;
  assign n80 = ~n58 & n62 ;
  assign n81 = n79 & n80 ;
  assign n82 = ~n51 & n54 ;
  assign n83 = ~n42 & n82 ;
  assign n84 = n81 & n83 ;
  assign n85 = n60 | n65 ;
  assign n86 = n63 & ~n85 ;
  assign n87 = n83 & n86 ;
  assign n88 = n84 | n87 ;
  assign n89 = n78 | n88 ;
  assign n90 = n60 & n65 ;
  assign n91 = n80 & n90 ;
  assign n92 = n77 & n91 ;
  assign n93 = n63 & n90 ;
  assign n94 = n77 & n93 ;
  assign n95 = ( ~n89 & n92 ) | ( ~n89 & n94 ) | ( n92 & n94 ) ;
  assign n96 = n89 | n95 ;
  assign n97 = n73 | n96 ;
  assign n98 = n51 & n54 ;
  assign n99 = ~n42 & n98 ;
  assign n100 = n67 & n99 ;
  assign n101 = n63 & n79 ;
  assign n102 = n99 & n101 ;
  assign n103 = ( ~n97 & n100 ) | ( ~n97 & n102 ) | ( n100 & n102 ) ;
  assign n104 = n97 | n103 ;
  assign n105 = n69 & n91 ;
  assign n106 = n70 & ~n85 ;
  assign n107 = n69 & n106 ;
  assign n108 = ( ~n104 & n105 ) | ( ~n104 & n107 ) | ( n105 & n107 ) ;
  assign n109 = n104 | n108 ;
  assign n110 = n70 & n79 ;
  assign n111 = n69 & n110 ;
  assign n112 = n80 & ~n85 ;
  assign n113 = n83 & n112 ;
  assign n114 = ( ~n109 & n111 ) | ( ~n109 & n113 ) | ( n111 & n113 ) ;
  assign n115 = n109 | n114 ;
  assign n116 = n83 & n110 ;
  assign n117 = n42 | n76 ;
  assign n118 = n110 & ~n117 ;
  assign n119 = ( ~n115 & n116 ) | ( ~n115 & n118 ) | ( n116 & n118 ) ;
  assign n120 = n115 | n119 ;
  assign n121 = n42 & n98 ;
  assign n122 = n93 & n121 ;
  assign n123 = n93 & n99 ;
  assign n124 = n81 & n99 ;
  assign n125 = n69 & n86 ;
  assign n126 = n124 | n125 ;
  assign n127 = n123 | n126 ;
  assign n128 = n122 | n127 ;
  assign n129 = n70 & n90 ;
  assign n130 = n83 & n129 ;
  assign n131 = n81 & ~n117 ;
  assign n132 = ( ~n128 & n130 ) | ( ~n128 & n131 ) | ( n130 & n131 ) ;
  assign n133 = n128 | n132 ;
  assign n134 = n71 & n77 ;
  assign n135 = ~n74 & n90 ;
  assign n136 = n77 & n135 ;
  assign n137 = n56 & n110 ;
  assign n138 = n71 & n83 ;
  assign n139 = n137 | n138 ;
  assign n140 = n136 | n139 ;
  assign n141 = n134 | n140 ;
  assign n142 = n83 & n101 ;
  assign n143 = n42 & n82 ;
  assign n144 = n91 & n143 ;
  assign n145 = n142 | n144 ;
  assign n146 = ~n117 & n129 ;
  assign n147 = ~n74 & n79 ;
  assign n148 = n56 & n147 ;
  assign n149 = n101 & n121 ;
  assign n150 = n101 & ~n117 ;
  assign n151 = n149 | n150 ;
  assign n152 = n148 | n151 ;
  assign n153 = n146 | n152 ;
  assign n154 = n145 | n153 ;
  assign n155 = n66 & n80 ;
  assign n156 = n69 & n155 ;
  assign n157 = n67 & n69 ;
  assign n158 = n106 & n121 ;
  assign n159 = n157 | n158 ;
  assign n160 = n69 & n147 ;
  assign n161 = n69 & n75 ;
  assign n162 = n160 | n161 ;
  assign n163 = n67 & n77 ;
  assign n164 = n112 & ~n117 ;
  assign n165 = n163 | n164 ;
  assign n166 = n162 | n165 ;
  assign n167 = n159 | n166 ;
  assign n168 = n81 & n121 ;
  assign n169 = n121 & n129 ;
  assign n170 = ( ~n167 & n168 ) | ( ~n167 & n169 ) | ( n168 & n169 ) ;
  assign n171 = n167 | n170 ;
  assign n172 = ( ~n154 & n156 ) | ( ~n154 & n171 ) | ( n156 & n171 ) ;
  assign n173 = n154 | n172 ;
  assign n174 = n69 & n129 ;
  assign n175 = n75 & n143 ;
  assign n176 = ( ~n173 & n174 ) | ( ~n173 & n175 ) | ( n174 & n175 ) ;
  assign n177 = n173 | n176 ;
  assign n178 = n67 & ~n117 ;
  assign n179 = ~n117 & n147 ;
  assign n180 = ( ~n177 & n178 ) | ( ~n177 & n179 ) | ( n178 & n179 ) ;
  assign n181 = n177 | n180 ;
  assign n182 = n77 & n112 ;
  assign n183 = n77 & n129 ;
  assign n184 = ( ~n181 & n182 ) | ( ~n181 & n183 ) | ( n182 & n183 ) ;
  assign n185 = n181 | n184 ;
  assign n186 = n141 | n185 ;
  assign n187 = n56 & n71 ;
  assign n188 = n86 & n143 ;
  assign n189 = ( ~n186 & n187 ) | ( ~n186 & n188 ) | ( n187 & n188 ) ;
  assign n190 = n186 | n189 ;
  assign n191 = n133 | n190 ;
  assign n192 = n120 | n191 ;
  assign n193 = n91 & n121 ;
  assign n194 = n99 & n112 ;
  assign n195 = n75 & n99 ;
  assign n196 = n194 | n195 ;
  assign n197 = ( ~n192 & n193 ) | ( ~n192 & n196 ) | ( n193 & n196 ) ;
  assign n198 = n192 | n197 ;
  assign n199 = n56 & n91 ;
  assign n200 = n56 & n75 ;
  assign n201 = ( ~n198 & n199 ) | ( ~n198 & n200 ) | ( n199 & n200 ) ;
  assign n202 = n198 | n201 ;
  assign n203 = n110 & n143 ;
  assign n204 = n74 | n85 ;
  assign n205 = n69 & ~n204 ;
  assign n206 = ( ~n202 & n203 ) | ( ~n202 & n205 ) | ( n203 & n205 ) ;
  assign n207 = n202 | n206 ;
  assign n208 = n106 & n143 ;
  assign n209 = n75 & n83 ;
  assign n210 = ( ~n207 & n208 ) | ( ~n207 & n209 ) | ( n208 & n209 ) ;
  assign n211 = n207 | n210 ;
  assign n212 = n106 & ~n117 ;
  assign n213 = n77 & n106 ;
  assign n214 = ( ~n211 & n212 ) | ( ~n211 & n213 ) | ( n212 & n213 ) ;
  assign n215 = n211 | n214 ;
  assign n2419 = x0 & ~x22 ;
  assign n2420 = n2419 ^ x1 ^ 1'b0 ;
  assign n537 = x2 & x22 ;
  assign n538 = ~x22 & n27 ;
  assign n539 = ~n26 & n538 ;
  assign n540 = n537 | n539 ;
  assign n2421 = n2420 ^ n540 ^ 1'b0 ;
  assign n2422 = x0 & ~n2421 ;
  assign n405 = n99 & n155 ;
  assign n890 = n194 | n405 ;
  assign n263 = n83 & n106 ;
  assign n891 = ( n116 & n263 ) | ( n116 & ~n890 ) | ( n263 & ~n890 ) ;
  assign n892 = n890 | n891 ;
  assign n384 = n56 & n81 ;
  assign n510 = n130 | n384 ;
  assign n445 = n56 & n106 ;
  assign n242 = n102 | n123 ;
  assign n394 = n99 & n135 ;
  assign n814 = n107 | n394 ;
  assign n815 = n242 | n814 ;
  assign n816 = n149 | n815 ;
  assign n349 = n121 & n135 ;
  assign n817 = ( n72 & n349 ) | ( n72 & ~n816 ) | ( n349 & ~n816 ) ;
  assign n818 = n816 | n817 ;
  assign n819 = n187 | n818 ;
  assign n820 = n445 | n819 ;
  assign n2685 = n510 | n820 ;
  assign n2686 = n892 | n2685 ;
  assign n305 = n69 & n81 ;
  assign n799 = n199 | n305 ;
  assign n347 = n99 & n106 ;
  assign n829 = n122 | n347 ;
  assign n309 = n56 & n129 ;
  assign n830 = ( n158 & n309 ) | ( n158 & ~n829 ) | ( n309 & ~n829 ) ;
  assign n831 = n829 | n830 ;
  assign n832 = ( n111 & n137 ) | ( n111 & ~n831 ) | ( n137 & ~n831 ) ;
  assign n833 = n831 | n832 ;
  assign n2687 = ( n799 & n833 ) | ( n799 & ~n2686 ) | ( n833 & ~n2686 ) ;
  assign n2688 = n2686 | n2687 ;
  assign n299 = n121 & n155 ;
  assign n300 = n105 | n299 ;
  assign n321 = n56 & n112 ;
  assign n322 = n56 & n155 ;
  assign n323 = n321 | n322 ;
  assign n378 = n77 & n110 ;
  assign n379 = n83 & ~n204 ;
  assign n380 = n378 | n379 ;
  assign n414 = n143 & ~n204 ;
  assign n423 = n69 & n112 ;
  assign n491 = n156 | n423 ;
  assign n492 = n414 | n491 ;
  assign n493 = n134 | n213 ;
  assign n494 = n492 | n493 ;
  assign n495 = n380 | n494 ;
  assign n496 = n323 | n495 ;
  assign n497 = ( n118 & n146 ) | ( n118 & ~n496 ) | ( n146 & ~n496 ) ;
  assign n498 = n496 | n497 ;
  assign n296 = n71 & ~n117 ;
  assign n499 = ( n183 & n296 ) | ( n183 & ~n498 ) | ( n296 & ~n498 ) ;
  assign n500 = n498 | n499 ;
  assign n2689 = ( n300 & n500 ) | ( n300 & ~n2688 ) | ( n500 & ~n2688 ) ;
  assign n2690 = n2688 | n2689 ;
  assign n273 = n93 & n143 ;
  assign n515 = n83 & n93 ;
  assign n516 = n273 | n515 ;
  assign n268 = n71 & n143 ;
  assign n517 = n208 | n268 ;
  assign n518 = n138 | n517 ;
  assign n519 = n516 | n518 ;
  assign n520 = n203 | n519 ;
  assign n462 = n135 & n143 ;
  assign n325 = n112 & n143 ;
  assign n753 = n209 | n325 ;
  assign n781 = n175 | n753 ;
  assign n293 = n83 & n147 ;
  assign n301 = n83 & n135 ;
  assign n782 = ( n293 & n301 ) | ( n293 & ~n781 ) | ( n301 & ~n781 ) ;
  assign n783 = n781 | n782 ;
  assign n784 = n462 | n783 ;
  assign n559 = n143 & n147 ;
  assign n785 = ( n113 & n559 ) | ( n113 & ~n784 ) | ( n559 & ~n784 ) ;
  assign n786 = n784 | n785 ;
  assign n2691 = ( n520 & n786 ) | ( n520 & ~n2690 ) | ( n786 & ~n2690 ) ;
  assign n2692 = n2690 | n2691 ;
  assign n250 = n67 & n121 ;
  assign n381 = n112 & n121 ;
  assign n2693 = n250 | n381 ;
  assign n2694 = ( n124 & ~n2692 ) | ( n124 & n2693 ) | ( ~n2692 & n2693 ) ;
  assign n2695 = n2692 | n2694 ;
  assign n233 = n69 & n135 ;
  assign n451 = n69 & n93 ;
  assign n376 = n56 & n135 ;
  assign n363 = n71 & n121 ;
  assign n404 = n67 & n143 ;
  assign n572 = n107 | n404 ;
  assign n573 = ( n130 & n163 ) | ( n130 & ~n572 ) | ( n163 & ~n572 ) ;
  assign n574 = n572 | n573 ;
  assign n1944 = n124 | n574 ;
  assign n1945 = n68 | n1944 ;
  assign n283 = n83 & n91 ;
  assign n1946 = ( n161 & n283 ) | ( n161 & ~n1945 ) | ( n283 & ~n1945 ) ;
  assign n1947 = n1945 | n1946 ;
  assign n240 = n83 & n155 ;
  assign n1948 = ( n179 & n240 ) | ( n179 & ~n1947 ) | ( n240 & ~n1947 ) ;
  assign n1949 = n1947 | n1948 ;
  assign n315 = n86 & n99 ;
  assign n316 = n56 & n93 ;
  assign n317 = n315 | n316 ;
  assign n1950 = n84 | n347 ;
  assign n1951 = n183 | n1950 ;
  assign n1952 = n317 | n1951 ;
  assign n1953 = ( n100 & n518 ) | ( n100 & ~n1952 ) | ( n518 & ~n1952 ) ;
  assign n1954 = n1952 | n1953 ;
  assign n304 = n99 & n110 ;
  assign n1955 = ( n304 & n394 ) | ( n304 & ~n1954 ) | ( n394 & ~n1954 ) ;
  assign n1956 = n1954 | n1955 ;
  assign n1957 = ( n113 & n209 ) | ( n113 & ~n1956 ) | ( n209 & ~n1956 ) ;
  assign n1958 = n1956 | n1957 ;
  assign n1959 = ( n146 & n164 ) | ( n146 & ~n1958 ) | ( n164 & ~n1958 ) ;
  assign n1960 = n1958 | n1959 ;
  assign n274 = n91 & ~n117 ;
  assign n275 = n274 ^ n273 ^ n136 ;
  assign n313 = n117 | n204 ;
  assign n314 = ~n157 & n313 ;
  assign n580 = n56 & n101 ;
  assign n974 = n168 | n580 ;
  assign n975 = n301 | n974 ;
  assign n1961 = n378 | n462 ;
  assign n284 = n143 & n155 ;
  assign n235 = n56 & n86 ;
  assign n698 = n111 | n235 ;
  assign n1538 = n284 | n698 ;
  assign n1539 = n116 | n1538 ;
  assign n256 = n99 & n147 ;
  assign n1962 = n322 ^ n256 ^ n174 ;
  assign n1963 = n1539 | n1962 ;
  assign n1964 = n1961 | n1963 ;
  assign n319 = n99 & ~n204 ;
  assign n362 = n309 | n319 ;
  assign n426 = n77 & n155 ;
  assign n560 = n160 | n426 ;
  assign n1965 = ( n362 & n560 ) | ( n362 & ~n1964 ) | ( n560 & ~n1964 ) ;
  assign n1966 = n1964 | n1965 ;
  assign n484 = n69 & n101 ;
  assign n331 = n86 & ~n117 ;
  assign n485 = n484 ^ n331 ^ n137 ;
  assign n486 = n156 | n485 ;
  assign n487 = n142 | n486 ;
  assign n278 = n77 & n86 ;
  assign n1967 = n250 | n278 ;
  assign n1968 = n349 | n1967 ;
  assign n1969 = ( n487 & ~n1966 ) | ( n487 & n1968 ) | ( ~n1966 & n1968 ) ;
  assign n1970 = n1966 | n1969 ;
  assign n1971 = ( n169 & n299 ) | ( n169 & ~n1970 ) | ( n299 & ~n1970 ) ;
  assign n1972 = n1970 | n1971 ;
  assign n1973 = ( n72 & n559 ) | ( n72 & ~n1972 ) | ( n559 & ~n1972 ) ;
  assign n1974 = n1972 | n1973 ;
  assign n1975 = n123 | n1974 ;
  assign n1976 = ( n94 & n182 ) | ( n94 & ~n1975 ) | ( n182 & ~n1975 ) ;
  assign n1977 = n1975 | n1976 ;
  assign n1978 = n975 | n1977 ;
  assign n1979 = ( n275 & n314 ) | ( n275 & ~n1978 ) | ( n314 & ~n1978 ) ;
  assign n1980 = ~n275 & n1979 ;
  assign n1981 = ( n1949 & ~n1960 ) | ( n1949 & n1980 ) | ( ~n1960 & n1980 ) ;
  assign n1982 = ~n1949 & n1981 ;
  assign n1983 = ( ~n196 & n363 ) | ( ~n196 & n1982 ) | ( n363 & n1982 ) ;
  assign n1984 = ~n363 & n1983 ;
  assign n1985 = ( ~n376 & n451 ) | ( ~n376 & n1984 ) | ( n451 & n1984 ) ;
  assign n1986 = ~n451 & n1985 ;
  assign n1987 = ( n105 & ~n233 ) | ( n105 & n1986 ) | ( ~n233 & n1986 ) ;
  assign n1988 = ~n105 & n1987 ;
  assign n535 = ~x22 & n31 ;
  assign n545 = n535 ^ x7 ^ 1'b0 ;
  assign n800 = n317 | n799 ;
  assign n237 = n100 | n124 ;
  assign n801 = ( n237 & n300 ) | ( n237 & ~n800 ) | ( n300 & ~n800 ) ;
  assign n802 = n800 | n801 ;
  assign n258 = n86 & n121 ;
  assign n803 = ( n258 & n405 ) | ( n258 & ~n802 ) | ( n405 & ~n802 ) ;
  assign n804 = n802 | n803 ;
  assign n805 = n484 | n580 ;
  assign n806 = ( n451 & ~n804 ) | ( n451 & n805 ) | ( ~n804 & n805 ) ;
  assign n807 = n804 | n806 ;
  assign n730 = n235 ^ n193 ^ n125 ;
  assign n236 = n91 & n99 ;
  assign n808 = n194 | n236 ;
  assign n809 = ( n68 & n168 ) | ( n68 & ~n808 ) | ( n168 & ~n808 ) ;
  assign n810 = n808 | n809 ;
  assign n811 = n730 | n810 ;
  assign n812 = ( n157 & n381 ) | ( n157 & ~n811 ) | ( n381 & ~n811 ) ;
  assign n813 = n811 | n812 ;
  assign n320 = n174 | n319 ;
  assign n821 = n320 | n820 ;
  assign n822 = n813 | n821 ;
  assign n238 = n71 & n99 ;
  assign n823 = ( n195 & n238 ) | ( n195 & ~n822 ) | ( n238 & ~n822 ) ;
  assign n824 = n822 | n823 ;
  assign n825 = ( n304 & n363 ) | ( n304 & ~n824 ) | ( n363 & ~n824 ) ;
  assign n826 = n824 | n825 ;
  assign n234 = n121 & ~n204 ;
  assign n827 = ( n234 & n250 ) | ( n234 & ~n826 ) | ( n250 & ~n826 ) ;
  assign n828 = n826 | n827 ;
  assign n243 = n110 & n121 ;
  assign n389 = n75 & n121 ;
  assign n390 = n243 | n389 ;
  assign n834 = n390 | n833 ;
  assign n835 = n828 | n834 ;
  assign n836 = n807 | n835 ;
  assign n367 = n99 & n129 ;
  assign n837 = ( n256 & n367 ) | ( n256 & ~n836 ) | ( n367 & ~n836 ) ;
  assign n838 = n836 | n837 ;
  assign n303 = n121 & n147 ;
  assign n839 = ( n169 & n303 ) | ( n169 & ~n838 ) | ( n303 & ~n838 ) ;
  assign n840 = n838 | n839 ;
  assign n1695 = n545 & n840 ;
  assign n345 = n236 | n258 ;
  assign n595 = n345 | n384 ;
  assign n596 = n580 | n595 ;
  assign n597 = ( n240 & n445 ) | ( n240 & ~n596 ) | ( n445 & ~n596 ) ;
  assign n598 = n596 | n597 ;
  assign n599 = n321 | n426 ;
  assign n600 = n182 | n599 ;
  assign n310 = n129 & n143 ;
  assign n601 = n296 | n310 ;
  assign n602 = n600 | n601 ;
  assign n603 = n598 | n602 ;
  assign n253 = n77 & n81 ;
  assign n604 = n188 | n253 ;
  assign n605 = ( n394 & ~n603 ) | ( n394 & n604 ) | ( ~n603 & n604 ) ;
  assign n606 = n603 | n605 ;
  assign n607 = ( n116 & n235 ) | ( n116 & ~n606 ) | ( n235 & ~n606 ) ;
  assign n608 = n606 | n607 ;
  assign n609 = ( n178 & n274 ) | ( n178 & ~n608 ) | ( n274 & ~n608 ) ;
  assign n610 = n608 | n609 ;
  assign n611 = n105 | n193 ;
  assign n612 = ( n273 & n301 ) | ( n273 & ~n611 ) | ( n301 & ~n611 ) ;
  assign n613 = n611 | n612 ;
  assign n475 = n93 & ~n117 ;
  assign n614 = ( n183 & n475 ) | ( n183 & ~n613 ) | ( n475 & ~n613 ) ;
  assign n615 = n613 | n614 ;
  assign n370 = n81 & n143 ;
  assign n616 = n234 | n381 ;
  assign n617 = n370 | n616 ;
  assign n618 = n160 | n200 ;
  assign n619 = n72 | n618 ;
  assign n620 = n617 | n619 ;
  assign n621 = n615 | n620 ;
  assign n622 = n610 | n621 ;
  assign n623 = n195 | n319 ;
  assign n624 = ( n113 & n349 ) | ( n113 & ~n623 ) | ( n349 & ~n623 ) ;
  assign n625 = n623 | n624 ;
  assign n626 = ( n138 & n212 ) | ( n138 & ~n625 ) | ( n212 & ~n625 ) ;
  assign n627 = n625 | n626 ;
  assign n288 = n77 & ~n204 ;
  assign n628 = ( n150 & n288 ) | ( n150 & ~n627 ) | ( n288 & ~n627 ) ;
  assign n629 = n627 | n628 ;
  assign n630 = n157 | n451 ;
  assign n631 = n142 | n630 ;
  assign n632 = n78 | n631 ;
  assign n633 = n175 | n315 ;
  assign n364 = n67 & n83 ;
  assign n634 = ( n84 & n364 ) | ( n84 & ~n633 ) | ( n364 & ~n633 ) ;
  assign n635 = n633 | n634 ;
  assign n636 = ( n331 & n378 ) | ( n331 & ~n635 ) | ( n378 & ~n635 ) ;
  assign n637 = n635 | n636 ;
  assign n638 = n492 | n637 ;
  assign n639 = n632 | n638 ;
  assign n640 = ( n100 & n144 ) | ( n100 & ~n639 ) | ( n144 & ~n639 ) ;
  assign n641 = n639 | n640 ;
  assign n642 = ( n208 & n559 ) | ( n208 & ~n641 ) | ( n559 & ~n641 ) ;
  assign n643 = n641 | n642 ;
  assign n232 = n77 & n147 ;
  assign n644 = ( n118 & n232 ) | ( n118 & ~n643 ) | ( n232 & ~n643 ) ;
  assign n645 = n643 | n644 ;
  assign n646 = ( ~n622 & n629 ) | ( ~n622 & n645 ) | ( n629 & n645 ) ;
  assign n647 = n622 | n646 ;
  assign n648 = ( n137 & n194 ) | ( n137 & ~n647 ) | ( n194 & ~n647 ) ;
  assign n649 = n647 | n648 ;
  assign n650 = ( n111 & n136 ) | ( n111 & ~n649 ) | ( n136 & ~n649 ) ;
  assign n651 = n649 | n650 ;
  assign n564 = n75 & ~n117 ;
  assign n239 = n116 | n238 ;
  assign n711 = n138 | n205 ;
  assign n712 = n239 | n711 ;
  assign n713 = n274 | n712 ;
  assign n714 = ( n94 & n232 ) | ( n94 & ~n713 ) | ( n232 & ~n713 ) ;
  assign n715 = n713 | n714 ;
  assign n302 = n87 | n301 ;
  assign n306 = n305 ^ n304 ^ n303 ;
  assign n307 = n302 | n306 ;
  assign n308 = n300 | n307 ;
  assign n311 = ( ~n308 & n309 ) | ( ~n308 & n310 ) | ( n309 & n310 ) ;
  assign n312 = n308 | n311 ;
  assign n716 = n263 | n370 ;
  assign n717 = n212 | n316 ;
  assign n718 = n195 | n717 ;
  assign n719 = ( n288 & n580 ) | ( n288 & ~n718 ) | ( n580 & ~n718 ) ;
  assign n720 = n718 | n719 ;
  assign n721 = n716 | n720 ;
  assign n722 = n312 | n721 ;
  assign n723 = n715 | n722 ;
  assign n724 = ( n123 & n367 ) | ( n123 & ~n723 ) | ( n367 & ~n723 ) ;
  assign n725 = n723 | n724 ;
  assign n726 = ( n107 & n144 ) | ( n107 & ~n725 ) | ( n144 & ~n725 ) ;
  assign n727 = n725 | n726 ;
  assign n728 = ( n92 & n175 ) | ( n92 & ~n727 ) | ( n175 & ~n727 ) ;
  assign n729 = n727 | n728 ;
  assign n731 = n149 | n730 ;
  assign n732 = n142 | n731 ;
  assign n437 = ~n117 & n135 ;
  assign n733 = ( n146 & n437 ) | ( n146 & ~n732 ) | ( n437 & ~n732 ) ;
  assign n734 = n732 | n733 ;
  assign n735 = n100 | n199 ;
  assign n365 = n363 | n364 ;
  assign n463 = n183 | n462 ;
  assign n464 = n136 | n463 ;
  assign n736 = n365 | n464 ;
  assign n737 = n735 | n736 ;
  assign n738 = n734 | n737 ;
  assign n279 = n148 | n278 ;
  assign n280 = ( n130 & n178 ) | ( n130 & ~n279 ) | ( n178 & ~n279 ) ;
  assign n281 = n279 | n280 ;
  assign n739 = ( n281 & n349 ) | ( n281 & ~n738 ) | ( n349 & ~n738 ) ;
  assign n740 = n738 | n739 ;
  assign n741 = ( n68 & n240 ) | ( n68 & ~n740 ) | ( n240 & ~n740 ) ;
  assign n742 = n740 | n741 ;
  assign n743 = n234 | n321 ;
  assign n744 = n445 | n743 ;
  assign n745 = ( n111 & n484 ) | ( n111 & ~n744 ) | ( n484 & ~n744 ) ;
  assign n746 = n744 | n745 ;
  assign n747 = ( n78 & n213 ) | ( n78 & ~n746 ) | ( n213 & ~n746 ) ;
  assign n748 = n746 | n747 ;
  assign n749 = n169 | n515 ;
  assign n750 = n378 | n749 ;
  assign n751 = n243 | n381 ;
  assign n752 = n331 | n751 ;
  assign n452 = n168 | n451 ;
  assign n453 = n423 | n452 ;
  assign n754 = n453 | n753 ;
  assign n755 = n752 | n754 ;
  assign n756 = n750 | n755 ;
  assign n757 = ( n314 & n748 ) | ( n314 & ~n756 ) | ( n748 & ~n756 ) ;
  assign n758 = ~n748 & n757 ;
  assign n759 = ( n729 & ~n742 ) | ( n729 & n758 ) | ( ~n742 & n758 ) ;
  assign n760 = ~n729 & n759 ;
  assign n761 = ( ~n160 & n174 ) | ( ~n160 & n760 ) | ( n174 & n760 ) ;
  assign n762 = ~n174 & n761 ;
  assign n763 = ( ~n179 & n564 ) | ( ~n179 & n762 ) | ( n564 & n762 ) ;
  assign n764 = ~n564 & n763 ;
  assign n668 = n370 | n515 ;
  assign n669 = n316 | n668 ;
  assign n670 = n423 | n669 ;
  assign n671 = n475 | n670 ;
  assign n350 = n174 | n200 ;
  assign n672 = n304 | n347 ;
  assign n673 = ( n268 & n367 ) | ( n268 & ~n672 ) | ( n367 & ~n672 ) ;
  assign n674 = n672 | n673 ;
  assign n675 = n350 | n674 ;
  assign n257 = n169 | n196 ;
  assign n259 = ( n187 & ~n257 ) | ( n187 & n258 ) | ( ~n257 & n258 ) ;
  assign n260 = n257 | n259 ;
  assign n676 = ( n260 & n281 ) | ( n260 & ~n675 ) | ( n281 & ~n675 ) ;
  assign n677 = n675 | n676 ;
  assign n678 = ( n256 & n363 ) | ( n256 & ~n677 ) | ( n363 & ~n677 ) ;
  assign n679 = n677 | n678 ;
  assign n680 = ( n168 & n414 ) | ( n168 & ~n679 ) | ( n414 & ~n679 ) ;
  assign n681 = n679 | n680 ;
  assign n682 = ( n139 & n163 ) | ( n139 & ~n681 ) | ( n163 & ~n681 ) ;
  assign n683 = n681 | n682 ;
  assign n684 = n315 | n683 ;
  assign n685 = n158 | n684 ;
  assign n686 = ( n274 & n331 ) | ( n274 & ~n685 ) | ( n331 & ~n685 ) ;
  assign n687 = n685 | n686 ;
  assign n688 = n671 | n687 ;
  assign n689 = n237 | n688 ;
  assign n690 = n233 | n404 ;
  assign n691 = n273 | n690 ;
  assign n692 = n243 | n691 ;
  assign n693 = n580 | n692 ;
  assign n694 = ( n445 & n462 ) | ( n445 & ~n693 ) | ( n462 & ~n693 ) ;
  assign n695 = n693 | n694 ;
  assign n696 = ( n113 & n283 ) | ( n113 & ~n695 ) | ( n283 & ~n695 ) ;
  assign n697 = n695 | n696 ;
  assign n266 = n77 & n101 ;
  assign n267 = n183 | n266 ;
  assign n699 = n150 | n698 ;
  assign n700 = n267 | n699 ;
  assign n701 = ( n199 & n238 ) | ( n199 & ~n700 ) | ( n238 & ~n700 ) ;
  assign n702 = n700 | n701 ;
  assign n703 = ( n205 & n301 ) | ( n205 & ~n702 ) | ( n301 & ~n702 ) ;
  assign n704 = n702 | n703 ;
  assign n705 = ( ~n689 & n697 ) | ( ~n689 & n704 ) | ( n697 & n704 ) ;
  assign n706 = n689 | n705 ;
  assign n382 = n303 | n381 ;
  assign n383 = n380 | n382 ;
  assign n385 = ( n122 & ~n383 ) | ( n122 & n384 ) | ( ~n383 & n384 ) ;
  assign n386 = n383 | n385 ;
  assign n387 = ( n92 & n322 ) | ( n92 & ~n386 ) | ( n322 & ~n386 ) ;
  assign n388 = n386 | n387 ;
  assign n707 = ( n68 & n388 ) | ( n68 & ~n706 ) | ( n388 & ~n706 ) ;
  assign n708 = n706 | n707 ;
  assign n709 = ( n146 & n364 ) | ( n146 & ~n708 ) | ( n364 & ~n708 ) ;
  assign n710 = n708 | n709 ;
  assign n765 = n764 ^ n710 ^ 1'b0 ;
  assign n766 = ~n710 & n764 ;
  assign n767 = n651 | n766 ;
  assign n769 = ~n765 & n767 ;
  assign n770 = ( n651 & n764 ) | ( n651 & n769 ) | ( n764 & n769 ) ;
  assign n1796 = n1695 ^ n770 ^ 1'b0 ;
  assign n536 = ~x22 & n29 ;
  assign n541 = n536 ^ x5 ^ 1'b0 ;
  assign n542 = n541 ^ n540 ^ 1'b0 ;
  assign n543 = ( ~x22 & n536 ) | ( ~x22 & n542 ) | ( n536 & n542 ) ;
  assign n544 = n543 ^ x6 ^ 1'b0 ;
  assign n546 = n545 ^ n544 ^ 1'b0 ;
  assign n547 = ( ~x22 & n535 ) | ( ~x22 & n546 ) | ( n535 & n546 ) ;
  assign n548 = n547 ^ x8 ^ 1'b0 ;
  assign n1795 = n548 & ~n840 ;
  assign n1797 = n1796 ^ n1795 ^ n548 ;
  assign n216 = n38 ^ x14 ^ 1'b0 ;
  assign n217 = n216 ^ x22 ^ 1'b0 ;
  assign n218 = ( x14 & n216 ) | ( x14 & n217 ) | ( n216 & n217 ) ;
  assign n768 = n765 & n767 ;
  assign n1692 = n218 & n768 ;
  assign n774 = n765 | n770 ;
  assign n1693 = ( n218 & n770 ) | ( n218 & n774 ) | ( n770 & n774 ) ;
  assign n1694 = ~n1692 & n1693 ;
  assign n558 = n125 | n238 ;
  assign n391 = n242 | n390 ;
  assign n392 = n145 | n391 ;
  assign n393 = n388 | n392 ;
  assign n395 = ( n194 & ~n393 ) | ( n194 & n394 ) | ( ~n393 & n394 ) ;
  assign n396 = n393 | n395 ;
  assign n397 = ( n156 & n304 ) | ( n156 & ~n396 ) | ( n304 & ~n396 ) ;
  assign n398 = n396 | n397 ;
  assign n399 = ~n117 & n155 ;
  assign n400 = ( n283 & ~n398 ) | ( n283 & n399 ) | ( ~n398 & n399 ) ;
  assign n401 = n398 | n400 ;
  assign n402 = n169 | n401 ;
  assign n403 = n331 | n402 ;
  assign n241 = n203 | n240 ;
  assign n561 = n161 | n437 ;
  assign n562 = n560 | n561 ;
  assign n563 = n241 | n562 ;
  assign n565 = ( n150 & ~n563 ) | ( n150 & n564 ) | ( ~n563 & n564 ) ;
  assign n566 = n563 | n565 ;
  assign n567 = n208 | n566 ;
  assign n568 = n559 | n567 ;
  assign n569 = n403 | n568 ;
  assign n570 = n558 | n569 ;
  assign n571 = n159 | n570 ;
  assign n351 = ( n51 & n152 ) | ( n51 & n256 ) | ( n152 & n256 ) ;
  assign n575 = n363 ^ n263 ^ n212 ;
  assign n576 = n347 ^ n310 ^ n250 ;
  assign n577 = n575 | n576 ;
  assign n578 = n351 | n577 ;
  assign n579 = n574 | n578 ;
  assign n581 = ( n349 & ~n579 ) | ( n349 & n580 ) | ( ~n579 & n580 ) ;
  assign n582 = n579 | n581 ;
  assign n583 = ( n111 & n187 ) | ( n111 & ~n582 ) | ( n187 & ~n582 ) ;
  assign n584 = n582 | n583 ;
  assign n585 = ( n118 & n301 ) | ( n118 & ~n584 ) | ( n301 & ~n584 ) ;
  assign n586 = n584 | n585 ;
  assign n587 = ( n73 & ~n571 ) | ( n73 & n586 ) | ( ~n571 & n586 ) ;
  assign n588 = n571 | n587 ;
  assign n589 = ( n141 & n414 ) | ( n141 & ~n588 ) | ( n414 & ~n588 ) ;
  assign n590 = n588 | n589 ;
  assign n441 = n325 | n367 ;
  assign n591 = ( n293 & n441 ) | ( n293 & ~n590 ) | ( n441 & ~n590 ) ;
  assign n592 = n590 | n591 ;
  assign n593 = ( n78 & n94 ) | ( n78 & ~n592 ) | ( n94 & ~n592 ) ;
  assign n594 = n592 | n593 ;
  assign n652 = n651 ^ n594 ^ 1'b0 ;
  assign n433 = n130 | n188 ;
  assign n434 = n379 | n433 ;
  assign n244 = n92 | n243 ;
  assign n245 = n242 | n244 ;
  assign n246 = n241 | n245 ;
  assign n247 = n239 | n246 ;
  assign n248 = n237 | n247 ;
  assign n249 = n236 | n248 ;
  assign n251 = ( n193 & ~n249 ) | ( n193 & n250 ) | ( ~n249 & n250 ) ;
  assign n252 = n249 | n251 ;
  assign n254 = ( n111 & ~n252 ) | ( n111 & n253 ) | ( ~n252 & n253 ) ;
  assign n255 = n252 | n254 ;
  assign n435 = n255 | n258 ;
  assign n436 = n113 | n435 ;
  assign n438 = n107 | n437 ;
  assign n439 = n436 | n438 ;
  assign n440 = n434 | n439 ;
  assign n442 = n87 | n441 ;
  assign n443 = ( n266 & n364 ) | ( n266 & ~n442 ) | ( n364 & ~n442 ) ;
  assign n444 = n442 | n443 ;
  assign n446 = ( n56 & n376 ) | ( n56 & n445 ) | ( n376 & n445 ) ;
  assign n447 = ( n268 & n322 ) | ( n268 & ~n446 ) | ( n322 & ~n446 ) ;
  assign n448 = n446 | n447 ;
  assign n449 = ( ~n440 & n444 ) | ( ~n440 & n448 ) | ( n444 & n448 ) ;
  assign n450 = n440 | n449 ;
  assign n454 = n315 | n453 ;
  assign n455 = n233 | n454 ;
  assign n456 = ( n212 & n310 ) | ( n212 & ~n455 ) | ( n310 & ~n455 ) ;
  assign n457 = n455 | n456 ;
  assign n458 = n131 | n232 ;
  assign n459 = n405 | n458 ;
  assign n460 = ( n146 & n299 ) | ( n146 & ~n459 ) | ( n299 & ~n459 ) ;
  assign n461 = n459 | n460 ;
  assign n465 = n122 | n169 ;
  assign n466 = n149 | n465 ;
  assign n467 = n464 | n466 ;
  assign n468 = n187 ^ n94 ^ n72 ;
  assign n469 = n467 | n468 ;
  assign n470 = n461 | n469 ;
  assign n348 = n321 | n347 ;
  assign n471 = n348 | n363 ;
  assign n472 = n158 | n471 ;
  assign n473 = ( n316 & n414 ) | ( n316 & ~n472 ) | ( n414 & ~n472 ) ;
  assign n474 = n472 | n473 ;
  assign n476 = ( n404 & ~n474 ) | ( n404 & n475 ) | ( ~n474 & n475 ) ;
  assign n477 = n474 | n476 ;
  assign n478 = ( n304 & ~n470 ) | ( n304 & n477 ) | ( ~n470 & n477 ) ;
  assign n479 = n470 | n478 ;
  assign n480 = ( n179 & n384 ) | ( n179 & ~n479 ) | ( n384 & ~n479 ) ;
  assign n481 = n479 | n480 ;
  assign n482 = ( ~n450 & n457 ) | ( ~n450 & n481 ) | ( n457 & n481 ) ;
  assign n483 = n450 | n482 ;
  assign n488 = ( n274 & ~n483 ) | ( n274 & n487 ) | ( ~n483 & n487 ) ;
  assign n489 = n483 | n488 ;
  assign n653 = n594 & n651 ;
  assign n654 = n489 & ~n653 ;
  assign n655 = n652 & ~n654 ;
  assign n656 = ( ~n489 & n651 ) | ( ~n489 & n655 ) | ( n651 & n655 ) ;
  assign n657 = n652 | n656 ;
  assign n658 = n652 | n654 ;
  assign n219 = ~x22 & n35 ;
  assign n221 = ~x22 & n33 ;
  assign n222 = n221 ^ x9 ^ 1'b0 ;
  assign n223 = ( ~x22 & n221 ) | ( ~x22 & n222 ) | ( n221 & n222 ) ;
  assign n224 = n223 ^ x10 ^ 1'b0 ;
  assign n220 = n219 ^ x11 ^ 1'b0 ;
  assign n225 = n224 ^ n220 ^ 1'b0 ;
  assign n226 = ( ~x22 & n219 ) | ( ~x22 & n225 ) | ( n219 & n225 ) ;
  assign n227 = n226 ^ x12 ^ 1'b0 ;
  assign n1697 = n657 ^ n227 ^ 1'b0 ;
  assign n1698 = ( n657 & n658 ) | ( n657 & ~n1697 ) | ( n658 & ~n1697 ) ;
  assign n229 = n40 ^ x13 ^ 1'b0 ;
  assign n1699 = n1698 ^ n229 ^ 1'b0 ;
  assign n1700 = ( n229 & ~n655 ) | ( n229 & n1699 ) | ( ~n655 & n1699 ) ;
  assign n1701 = ( n1698 & ~n1699 ) | ( n1698 & n1700 ) | ( ~n1699 & n1700 ) ;
  assign n664 = n652 & ~n656 ;
  assign n1702 = ( n229 & n664 ) | ( n229 & ~n1701 ) | ( n664 & ~n1701 ) ;
  assign n1703 = n1702 ^ n1701 ^ 1'b0 ;
  assign n1704 = ( n1701 & ~n1702 ) | ( n1701 & n1703 ) | ( ~n1702 & n1703 ) ;
  assign n1798 = ( n1694 & ~n1695 ) | ( n1694 & n1704 ) | ( ~n1695 & n1704 ) ;
  assign n907 = n175 | n384 ;
  assign n908 = n209 | n907 ;
  assign n909 = n158 | n376 ;
  assign n910 = ( n296 & n364 ) | ( n296 & ~n909 ) | ( n364 & ~n909 ) ;
  assign n911 = n909 | n910 ;
  assign n912 = n205 ^ n179 ^ n137 ;
  assign n913 = n911 | n912 ;
  assign n914 = n908 | n913 ;
  assign n915 = ( n241 & n260 ) | ( n241 & ~n914 ) | ( n260 & ~n914 ) ;
  assign n916 = n914 | n915 ;
  assign n917 = ( n199 & n367 ) | ( n199 & ~n916 ) | ( n367 & ~n916 ) ;
  assign n918 = n916 | n917 ;
  assign n919 = ( n266 & n310 ) | ( n266 & ~n918 ) | ( n310 & ~n918 ) ;
  assign n920 = n918 | n919 ;
  assign n921 = n348 | n716 ;
  assign n922 = ( n193 & n560 ) | ( n193 & ~n921 ) | ( n560 & ~n921 ) ;
  assign n923 = n921 | n922 ;
  assign n924 = n68 | n923 ;
  assign n925 = ( n188 & n423 ) | ( n188 & ~n924 ) | ( n423 & ~n924 ) ;
  assign n926 = n924 | n925 ;
  assign n927 = ( n94 & n208 ) | ( n94 & ~n926 ) | ( n208 & ~n926 ) ;
  assign n928 = n926 | n927 ;
  assign n328 = n101 & n143 ;
  assign n859 = n325 | n805 ;
  assign n860 = n378 | n859 ;
  assign n861 = n516 | n860 ;
  assign n862 = n328 | n861 ;
  assign n511 = n148 | n233 ;
  assign n929 = n278 | n511 ;
  assign n930 = ( n234 & n363 ) | ( n234 & ~n929 ) | ( n363 & ~n929 ) ;
  assign n931 = n929 | n930 ;
  assign n932 = ( n144 & n445 ) | ( n144 & ~n931 ) | ( n445 & ~n931 ) ;
  assign n933 = n931 | n932 ;
  assign n934 = ( n288 & n293 ) | ( n288 & ~n933 ) | ( n293 & ~n933 ) ;
  assign n935 = n933 | n934 ;
  assign n936 = n126 | n165 ;
  assign n937 = ( n382 & n461 ) | ( n382 & ~n936 ) | ( n461 & ~n936 ) ;
  assign n938 = n936 | n937 ;
  assign n939 = ( n314 & n935 ) | ( n314 & ~n938 ) | ( n935 & ~n938 ) ;
  assign n940 = ~n935 & n939 ;
  assign n941 = ( ~n862 & n928 ) | ( ~n862 & n940 ) | ( n928 & n940 ) ;
  assign n942 = ~n928 & n941 ;
  assign n943 = ( n394 & ~n920 ) | ( n394 & n942 ) | ( ~n920 & n942 ) ;
  assign n944 = ~n394 & n943 ;
  assign n945 = ( n111 & ~n559 ) | ( n111 & n944 ) | ( ~n559 & n944 ) ;
  assign n946 = ~n111 & n945 ;
  assign n947 = ( n138 & ~n274 ) | ( n138 & n946 ) | ( ~n274 & n946 ) ;
  assign n948 = ~n138 & n947 ;
  assign n346 = n134 | n345 ;
  assign n858 = n346 | n752 ;
  assign n863 = ( n300 & ~n858 ) | ( n300 & n862 ) | ( ~n858 & n862 ) ;
  assign n864 = n858 | n863 ;
  assign n865 = ( n171 & n304 ) | ( n171 & ~n864 ) | ( n304 & ~n864 ) ;
  assign n866 = n864 | n865 ;
  assign n867 = ( n102 & n367 ) | ( n102 & ~n866 ) | ( n367 & ~n866 ) ;
  assign n868 = n866 | n867 ;
  assign n282 = n56 & ~n204 ;
  assign n869 = ( n282 & n404 ) | ( n282 & ~n868 ) | ( n404 & ~n868 ) ;
  assign n870 = n868 | n869 ;
  assign n871 = ( n301 & n399 ) | ( n301 & ~n870 ) | ( n399 & ~n870 ) ;
  assign n872 = n870 | n871 ;
  assign n873 = n362 | n717 ;
  assign n874 = ( n234 & n389 ) | ( n234 & ~n873 ) | ( n389 & ~n873 ) ;
  assign n875 = n873 | n874 ;
  assign n876 = ( n68 & n384 ) | ( n68 & ~n875 ) | ( n384 & ~n875 ) ;
  assign n877 = n875 | n876 ;
  assign n878 = ( n78 & n274 ) | ( n78 & ~n877 ) | ( n274 & ~n877 ) ;
  assign n879 = n877 | n878 ;
  assign n880 = n468 | n699 ;
  assign n881 = n313 & ~n880 ;
  assign n882 = ( n491 & ~n879 ) | ( n491 & n881 ) | ( ~n879 & n881 ) ;
  assign n883 = ~n491 & n882 ;
  assign n884 = ( ~n125 & n451 ) | ( ~n125 & n883 ) | ( n451 & n883 ) ;
  assign n885 = ~n451 & n884 ;
  assign n886 = ( ~n288 & n564 ) | ( ~n288 & n885 ) | ( n564 & n885 ) ;
  assign n887 = ~n564 & n886 ;
  assign n888 = ( n92 & ~n182 ) | ( n92 & n887 ) | ( ~n182 & n887 ) ;
  assign n889 = ~n92 & n888 ;
  assign n893 = n601 | n892 ;
  assign n894 = n518 | n893 ;
  assign n375 = n233 | n284 ;
  assign n895 = n113 | n375 ;
  assign n896 = n293 | n895 ;
  assign n897 = ( n283 & n379 ) | ( n283 & ~n896 ) | ( n379 & ~n896 ) ;
  assign n898 = n896 | n897 ;
  assign n899 = ( n145 & ~n894 ) | ( n145 & n898 ) | ( ~n894 & n898 ) ;
  assign n900 = n894 | n899 ;
  assign n901 = ( n237 & n889 ) | ( n237 & ~n900 ) | ( n889 & ~n900 ) ;
  assign n902 = ~n237 & n901 ;
  assign n903 = ( n123 & ~n872 ) | ( n123 & n902 ) | ( ~n872 & n902 ) ;
  assign n904 = ~n123 & n903 ;
  assign n905 = ( ~n209 & n349 ) | ( ~n209 & n904 ) | ( n349 & n904 ) ;
  assign n906 = ~n349 & n905 ;
  assign n949 = n948 ^ n906 ^ 1'b0 ;
  assign n950 = n906 & n948 ;
  assign n951 = n764 & ~n950 ;
  assign n952 = n949 | n951 ;
  assign n953 = n952 ^ n950 ^ n764 ;
  assign n1587 = ~n948 & n953 ;
  assign n1588 = ( n764 & n948 ) | ( n764 & n1587 ) | ( n948 & n1587 ) ;
  assign n1589 = n544 & n840 ;
  assign n1590 = n1589 ^ n1588 ^ n1587 ;
  assign n1674 = ( n1588 & n1589 ) | ( n1588 & n1590 ) | ( n1589 & n1590 ) ;
  assign n506 = n200 | n376 ;
  assign n507 = n328 | n506 ;
  assign n508 = ( n116 & n310 ) | ( n116 & ~n507 ) | ( n310 & ~n507 ) ;
  assign n509 = n507 | n508 ;
  assign n512 = n510 | n511 ;
  assign n513 = n162 | n512 ;
  assign n514 = n509 | n513 ;
  assign n521 = ( n282 & ~n514 ) | ( n282 & n520 ) | ( ~n514 & n520 ) ;
  assign n522 = n514 | n521 ;
  assign n523 = ( n205 & n263 ) | ( n205 & ~n522 ) | ( n263 & ~n522 ) ;
  assign n524 = n522 | n523 ;
  assign n285 = n283 | n284 ;
  assign n286 = n84 | n285 ;
  assign n787 = n145 | n286 ;
  assign n788 = n370 | n787 ;
  assign n789 = ( n188 & n404 ) | ( n188 & ~n788 ) | ( n404 & ~n788 ) ;
  assign n790 = n788 | n789 ;
  assign n791 = ( n87 & n364 ) | ( n87 & ~n790 ) | ( n364 & ~n790 ) ;
  assign n792 = n790 | n791 ;
  assign n793 = n524 | n792 ;
  assign n794 = ( n323 & n491 ) | ( n323 & ~n793 ) | ( n491 & ~n793 ) ;
  assign n795 = n793 | n794 ;
  assign n796 = n786 | n795 ;
  assign n797 = n240 | n796 ;
  assign n501 = n212 | n500 ;
  assign n502 = ( n94 & n475 ) | ( n94 & ~n501 ) | ( n475 & ~n501 ) ;
  assign n503 = n501 | n502 ;
  assign n504 = n266 | n503 ;
  assign n505 = n278 | n504 ;
  assign n525 = ( n150 & ~n505 ) | ( n150 & n524 ) | ( ~n505 & n524 ) ;
  assign n526 = n505 | n525 ;
  assign n527 = ( n163 & n178 ) | ( n163 & ~n526 ) | ( n178 & ~n526 ) ;
  assign n528 = n526 | n527 ;
  assign n798 = n797 ^ n528 ^ 1'b0 ;
  assign n841 = n528 & n797 ;
  assign n842 = n840 & ~n841 ;
  assign n843 = n798 & ~n842 ;
  assign n844 = ( n797 & ~n840 ) | ( n797 & n843 ) | ( ~n840 & n843 ) ;
  assign n845 = n798 | n844 ;
  assign n846 = n798 | n842 ;
  assign n1675 = n845 ^ n548 ^ 1'b0 ;
  assign n1676 = ( n845 & n846 ) | ( n845 & ~n1675 ) | ( n846 & ~n1675 ) ;
  assign n1677 = n1676 ^ n222 ^ 1'b0 ;
  assign n1678 = ( n222 & ~n843 ) | ( n222 & n1677 ) | ( ~n843 & n1677 ) ;
  assign n1679 = ( n1676 & ~n1677 ) | ( n1676 & n1678 ) | ( ~n1677 & n1678 ) ;
  assign n852 = n798 & ~n844 ;
  assign n1680 = ( n222 & n852 ) | ( n222 & ~n1679 ) | ( n852 & ~n1679 ) ;
  assign n1681 = n1680 ^ n1679 ^ 1'b0 ;
  assign n1682 = ( n1679 & ~n1680 ) | ( n1679 & n1681 ) | ( ~n1680 & n1681 ) ;
  assign n352 = n350 | n351 ;
  assign n353 = ( n238 & n299 ) | ( n238 & ~n352 ) | ( n299 & ~n352 ) ;
  assign n354 = n352 | n353 ;
  assign n355 = ( n183 & n253 ) | ( n183 & ~n354 ) | ( n253 & ~n354 ) ;
  assign n356 = n354 | n355 ;
  assign n357 = n349 | n356 ;
  assign n358 = n161 | n357 ;
  assign n359 = n348 | n358 ;
  assign n360 = n346 | n359 ;
  assign n361 = n282 | n296 ;
  assign n366 = n362 | n365 ;
  assign n368 = ( n158 & ~n366 ) | ( n158 & n367 ) | ( ~n366 & n367 ) ;
  assign n369 = n366 | n368 ;
  assign n371 = ( n160 & ~n369 ) | ( n160 & n370 ) | ( ~n369 & n370 ) ;
  assign n372 = n369 | n371 ;
  assign n373 = ( ~n360 & n361 ) | ( ~n360 & n372 ) | ( n361 & n372 ) ;
  assign n374 = n360 | n373 ;
  assign n377 = n213 | n376 ;
  assign n406 = n234 | n405 ;
  assign n407 = n193 | n406 ;
  assign n408 = n404 | n407 ;
  assign n409 = n403 | n408 ;
  assign n410 = n377 | n409 ;
  assign n272 = n118 | n182 ;
  assign n411 = n237 | n272 ;
  assign n412 = ( n168 & n250 ) | ( n168 & ~n411 ) | ( n250 & ~n411 ) ;
  assign n413 = n411 | n412 ;
  assign n415 = ( n188 & ~n413 ) | ( n188 & n414 ) | ( ~n413 & n414 ) ;
  assign n416 = n413 | n415 ;
  assign n417 = ( n84 & n131 ) | ( n84 & ~n416 ) | ( n131 & ~n416 ) ;
  assign n418 = n416 | n417 ;
  assign n419 = n195 | n315 ;
  assign n420 = n87 | n419 ;
  assign n421 = ( ~n410 & n418 ) | ( ~n410 & n420 ) | ( n418 & n420 ) ;
  assign n422 = n410 | n421 ;
  assign n424 = ( n205 & ~n422 ) | ( n205 & n423 ) | ( ~n422 & n423 ) ;
  assign n425 = n422 | n424 ;
  assign n427 = ( n164 & ~n425 ) | ( n164 & n426 ) | ( ~n425 & n426 ) ;
  assign n428 = n425 | n427 ;
  assign n429 = ( ~n374 & n375 ) | ( ~n374 & n428 ) | ( n375 & n428 ) ;
  assign n430 = n374 | n429 ;
  assign n431 = ( n146 & n274 ) | ( n146 & ~n430 ) | ( n274 & ~n430 ) ;
  assign n432 = n430 | n431 ;
  assign n490 = n489 ^ n432 ^ 1'b0 ;
  assign n529 = n432 & n489 ;
  assign n530 = n528 & ~n529 ;
  assign n531 = n490 & ~n530 ;
  assign n532 = ( n489 & ~n528 ) | ( n489 & n531 ) | ( ~n528 & n531 ) ;
  assign n533 = n490 | n532 ;
  assign n534 = n490 | n530 ;
  assign n1683 = n534 ^ n224 ^ 1'b0 ;
  assign n1684 = ( n533 & n534 ) | ( n533 & n1683 ) | ( n534 & n1683 ) ;
  assign n1685 = n1684 ^ n220 ^ 1'b0 ;
  assign n1686 = ( n220 & ~n531 ) | ( n220 & n1685 ) | ( ~n531 & n1685 ) ;
  assign n1687 = ( n1684 & ~n1685 ) | ( n1684 & n1686 ) | ( ~n1685 & n1686 ) ;
  assign n554 = n490 & ~n532 ;
  assign n1688 = ( n220 & n554 ) | ( n220 & ~n1687 ) | ( n554 & ~n1687 ) ;
  assign n1689 = n1688 ^ n1687 ^ 1'b0 ;
  assign n1690 = ( n1687 & ~n1688 ) | ( n1687 & n1689 ) | ( ~n1688 & n1689 ) ;
  assign n1799 = ( n1674 & n1682 ) | ( n1674 & n1690 ) | ( n1682 & n1690 ) ;
  assign n1891 = ( ~n1797 & n1798 ) | ( ~n1797 & n1799 ) | ( n1798 & n1799 ) ;
  assign n1882 = n533 ^ n227 ^ 1'b0 ;
  assign n1883 = ( n533 & n534 ) | ( n533 & ~n1882 ) | ( n534 & ~n1882 ) ;
  assign n1884 = n1883 ^ n229 ^ 1'b0 ;
  assign n1885 = ( n229 & ~n531 ) | ( n229 & n1884 ) | ( ~n531 & n1884 ) ;
  assign n1886 = ( n1883 & ~n1884 ) | ( n1883 & n1885 ) | ( ~n1884 & n1885 ) ;
  assign n1887 = ( n229 & n554 ) | ( n229 & ~n1886 ) | ( n554 & ~n1886 ) ;
  assign n1888 = n1887 ^ n1886 ^ 1'b0 ;
  assign n1889 = ( n1886 & ~n1887 ) | ( n1886 & n1888 ) | ( ~n1887 & n1888 ) ;
  assign n1880 = n222 & n840 ;
  assign n1876 = n218 & ~n657 ;
  assign n1877 = n218 | n654 ;
  assign n1878 = ( ~n655 & n1876 ) | ( ~n655 & n1877 ) | ( n1876 & n1877 ) ;
  assign n1879 = ~n1876 & n1878 ;
  assign n1881 = n1880 ^ n1879 ^ 1'b0 ;
  assign n1890 = n1889 ^ n1881 ^ 1'b0 ;
  assign n1801 = n845 ^ n222 ^ 1'b0 ;
  assign n1802 = ( n845 & n846 ) | ( n845 & ~n1801 ) | ( n846 & ~n1801 ) ;
  assign n1803 = n1802 ^ n224 ^ 1'b0 ;
  assign n1804 = ( n224 & ~n843 ) | ( n224 & n1803 ) | ( ~n843 & n1803 ) ;
  assign n1805 = ( n1802 & ~n1803 ) | ( n1802 & n1804 ) | ( ~n1803 & n1804 ) ;
  assign n1806 = ( n224 & n852 ) | ( n224 & ~n1805 ) | ( n852 & ~n1805 ) ;
  assign n1807 = n1806 ^ n1805 ^ 1'b0 ;
  assign n1808 = ( n1805 & ~n1806 ) | ( n1805 & n1807 ) | ( ~n1806 & n1807 ) ;
  assign n1809 = n533 ^ n220 ^ 1'b0 ;
  assign n1810 = ( n533 & n534 ) | ( n533 & ~n1809 ) | ( n534 & ~n1809 ) ;
  assign n1811 = n1810 ^ n227 ^ 1'b0 ;
  assign n1812 = ( n227 & ~n531 ) | ( n227 & n1811 ) | ( ~n531 & n1811 ) ;
  assign n1813 = ( n1810 & ~n1811 ) | ( n1810 & n1812 ) | ( ~n1811 & n1812 ) ;
  assign n1814 = ( n227 & n554 ) | ( n227 & ~n1813 ) | ( n554 & ~n1813 ) ;
  assign n1815 = n1814 ^ n1813 ^ 1'b0 ;
  assign n1816 = ( n1813 & ~n1814 ) | ( n1813 & n1815 ) | ( ~n1814 & n1815 ) ;
  assign n1817 = n657 ^ n229 ^ 1'b0 ;
  assign n1818 = ( n657 & n658 ) | ( n657 & ~n1817 ) | ( n658 & ~n1817 ) ;
  assign n1819 = n1818 ^ n218 ^ 1'b0 ;
  assign n1820 = ( n218 & ~n655 ) | ( n218 & n1819 ) | ( ~n655 & n1819 ) ;
  assign n1821 = ( n1818 & ~n1819 ) | ( n1818 & n1820 ) | ( ~n1819 & n1820 ) ;
  assign n1822 = ( n218 & n664 ) | ( n218 & ~n1821 ) | ( n664 & ~n1821 ) ;
  assign n1823 = n1822 ^ n1821 ^ 1'b0 ;
  assign n1824 = ( n1821 & ~n1822 ) | ( n1821 & n1823 ) | ( ~n1822 & n1823 ) ;
  assign n1874 = ( n1808 & n1816 ) | ( n1808 & n1824 ) | ( n1816 & n1824 ) ;
  assign n1865 = n845 ^ n224 ^ 1'b0 ;
  assign n1866 = ( n845 & n846 ) | ( n845 & ~n1865 ) | ( n846 & ~n1865 ) ;
  assign n1867 = n1866 ^ n220 ^ 1'b0 ;
  assign n1868 = ( n220 & ~n843 ) | ( n220 & n1867 ) | ( ~n843 & n1867 ) ;
  assign n1869 = ( n1866 & ~n1867 ) | ( n1866 & n1868 ) | ( ~n1867 & n1868 ) ;
  assign n1870 = ( n220 & n852 ) | ( n220 & ~n1869 ) | ( n852 & ~n1869 ) ;
  assign n1871 = n1870 ^ n1869 ^ 1'b0 ;
  assign n1872 = ( n1869 & ~n1870 ) | ( n1869 & n1871 ) | ( ~n1870 & n1871 ) ;
  assign n1861 = n548 & ~n1796 ;
  assign n1862 = n840 & n1861 ;
  assign n1863 = ~n770 & n1695 ;
  assign n1864 = n1862 | n1863 ;
  assign n1873 = n1872 ^ n1864 ^ 1'b0 ;
  assign n1875 = n1874 ^ n1873 ^ 1'b0 ;
  assign n1892 = n1891 ^ n1890 ^ n1875 ;
  assign n1800 = n1799 ^ n1798 ^ n1797 ;
  assign n1825 = n1824 ^ n1816 ^ n1808 ;
  assign n1691 = n1690 ^ n1682 ^ n1674 ;
  assign n1696 = n1695 ^ n1694 ^ 1'b0 ;
  assign n1705 = n1704 ^ n1696 ^ 1'b0 ;
  assign n771 = n765 & ~n770 ;
  assign n1559 = n768 ^ n229 ^ 1'b0 ;
  assign n1560 = ( n768 & n771 ) | ( n768 & ~n1559 ) | ( n771 & ~n1559 ) ;
  assign n1561 = ( n218 & n774 ) | ( n218 & ~n1560 ) | ( n774 & ~n1560 ) ;
  assign n1562 = ~n1560 & n1561 ;
  assign n1563 = ( n218 & n769 ) | ( n218 & ~n1562 ) | ( n769 & ~n1562 ) ;
  assign n1564 = n1563 ^ n1562 ^ 1'b0 ;
  assign n1565 = ( n1562 & ~n1563 ) | ( n1562 & n1564 ) | ( ~n1563 & n1564 ) ;
  assign n1566 = n845 ^ n545 ^ 1'b0 ;
  assign n1567 = ( n845 & n846 ) | ( n845 & ~n1566 ) | ( n846 & ~n1566 ) ;
  assign n1568 = n1567 ^ n548 ^ 1'b0 ;
  assign n1569 = ( n548 & ~n843 ) | ( n548 & n1568 ) | ( ~n843 & n1568 ) ;
  assign n1570 = ( n1567 & ~n1568 ) | ( n1567 & n1569 ) | ( ~n1568 & n1569 ) ;
  assign n1571 = ( n548 & n852 ) | ( n548 & ~n1570 ) | ( n852 & ~n1570 ) ;
  assign n1572 = n1571 ^ n1570 ^ 1'b0 ;
  assign n1573 = ( n1570 & ~n1571 ) | ( n1570 & n1572 ) | ( ~n1571 & n1572 ) ;
  assign n1574 = n534 ^ n222 ^ 1'b0 ;
  assign n1575 = ( n533 & n534 ) | ( n533 & n1574 ) | ( n534 & n1574 ) ;
  assign n1576 = n1575 ^ n224 ^ 1'b0 ;
  assign n1577 = ( n224 & ~n531 ) | ( n224 & n1576 ) | ( ~n531 & n1576 ) ;
  assign n1578 = ( n1575 & ~n1576 ) | ( n1575 & n1577 ) | ( ~n1576 & n1577 ) ;
  assign n1579 = ( n224 & n554 ) | ( n224 & ~n1578 ) | ( n554 & ~n1578 ) ;
  assign n1580 = n1579 ^ n1578 ^ 1'b0 ;
  assign n1581 = ( n1578 & ~n1579 ) | ( n1578 & n1580 ) | ( ~n1579 & n1580 ) ;
  assign n1706 = ( n1565 & n1573 ) | ( n1565 & n1581 ) | ( n1573 & n1581 ) ;
  assign n1826 = ( n1691 & ~n1705 ) | ( n1691 & n1706 ) | ( ~n1705 & n1706 ) ;
  assign n1893 = ( ~n1800 & n1825 ) | ( ~n1800 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1827 = n1826 ^ n1825 ^ n1800 ;
  assign n1707 = n1706 ^ n1705 ^ n1691 ;
  assign n1582 = n1581 ^ n1573 ^ n1565 ;
  assign n856 = n538 ^ x3 ^ 1'b0 ;
  assign n1038 = n856 ^ n540 ^ 1'b0 ;
  assign n1039 = ( ~x22 & n538 ) | ( ~x22 & n1038 ) | ( n538 & n1038 ) ;
  assign n1040 = n1039 ^ x4 ^ 1'b0 ;
  assign n1041 = n840 & n1040 ;
  assign n961 = n949 & ~n951 ;
  assign n1042 = n218 & n961 ;
  assign n954 = n949 | n953 ;
  assign n1043 = n952 ^ n229 ^ 1'b0 ;
  assign n1044 = ( n952 & n954 ) | ( n952 & ~n1043 ) | ( n954 & ~n1043 ) ;
  assign n958 = n949 & ~n953 ;
  assign n1045 = ~n218 & n958 ;
  assign n1046 = ( n1042 & n1044 ) | ( n1042 & ~n1045 ) | ( n1044 & ~n1045 ) ;
  assign n1047 = ~n1042 & n1046 ;
  assign n1048 = ( ~n948 & n1041 ) | ( ~n948 & n1047 ) | ( n1041 & n1047 ) ;
  assign n1049 = n845 ^ n544 ^ 1'b0 ;
  assign n1050 = ( n845 & n846 ) | ( n845 & ~n1049 ) | ( n846 & ~n1049 ) ;
  assign n1051 = n1050 ^ n545 ^ 1'b0 ;
  assign n1052 = ( n545 & ~n843 ) | ( n545 & n1051 ) | ( ~n843 & n1051 ) ;
  assign n1053 = ( n1050 & ~n1051 ) | ( n1050 & n1052 ) | ( ~n1051 & n1052 ) ;
  assign n1054 = ( n545 & n852 ) | ( n545 & ~n1053 ) | ( n852 & ~n1053 ) ;
  assign n1055 = n1054 ^ n1053 ^ 1'b0 ;
  assign n1056 = ( n1053 & ~n1054 ) | ( n1053 & n1055 ) | ( ~n1054 & n1055 ) ;
  assign n1058 = n657 ^ n222 ^ 1'b0 ;
  assign n1059 = ( n657 & n658 ) | ( n657 & ~n1058 ) | ( n658 & ~n1058 ) ;
  assign n1060 = n1059 ^ n224 ^ 1'b0 ;
  assign n1061 = ( n224 & ~n655 ) | ( n224 & n1060 ) | ( ~n655 & n1060 ) ;
  assign n1062 = ( n1059 & ~n1060 ) | ( n1059 & n1061 ) | ( ~n1060 & n1061 ) ;
  assign n1063 = ( n224 & n664 ) | ( n224 & ~n1062 ) | ( n664 & ~n1062 ) ;
  assign n1064 = n1063 ^ n1062 ^ 1'b0 ;
  assign n1065 = ( n1062 & ~n1063 ) | ( n1062 & n1064 ) | ( ~n1063 & n1064 ) ;
  assign n1066 = n768 ^ n220 ^ 1'b0 ;
  assign n1067 = ( n768 & n771 ) | ( n768 & ~n1066 ) | ( n771 & ~n1066 ) ;
  assign n1068 = ( n227 & n774 ) | ( n227 & ~n1067 ) | ( n774 & ~n1067 ) ;
  assign n1069 = ~n1067 & n1068 ;
  assign n1070 = ( n227 & n769 ) | ( n227 & ~n1069 ) | ( n769 & ~n1069 ) ;
  assign n1071 = n1070 ^ n1069 ^ 1'b0 ;
  assign n1072 = ( n1069 & ~n1070 ) | ( n1069 & n1071 ) | ( ~n1070 & n1071 ) ;
  assign n1073 = n545 ^ n533 ^ 1'b0 ;
  assign n1074 = ( n533 & n534 ) | ( n533 & ~n1073 ) | ( n534 & ~n1073 ) ;
  assign n1075 = n1074 ^ n548 ^ 1'b0 ;
  assign n1076 = ( ~n531 & n548 ) | ( ~n531 & n1075 ) | ( n548 & n1075 ) ;
  assign n1077 = ( n1074 & ~n1075 ) | ( n1074 & n1076 ) | ( ~n1075 & n1076 ) ;
  assign n1078 = ( n548 & n554 ) | ( n548 & ~n1077 ) | ( n554 & ~n1077 ) ;
  assign n1079 = n1078 ^ n1077 ^ 1'b0 ;
  assign n1080 = ( n1077 & ~n1078 ) | ( n1077 & n1079 ) | ( ~n1078 & n1079 ) ;
  assign n1081 = ( n1065 & n1072 ) | ( n1065 & n1080 ) | ( n1072 & n1080 ) ;
  assign n1583 = ( n1048 & n1056 ) | ( n1048 & n1081 ) | ( n1056 & n1081 ) ;
  assign n549 = n548 ^ n533 ^ 1'b0 ;
  assign n550 = ( n533 & n534 ) | ( n533 & ~n549 ) | ( n534 & ~n549 ) ;
  assign n551 = n550 ^ n222 ^ 1'b0 ;
  assign n552 = ( n222 & ~n531 ) | ( n222 & n551 ) | ( ~n531 & n551 ) ;
  assign n553 = ( n550 & ~n551 ) | ( n550 & n552 ) | ( ~n551 & n552 ) ;
  assign n555 = ( n222 & ~n553 ) | ( n222 & n554 ) | ( ~n553 & n554 ) ;
  assign n556 = n555 ^ n553 ^ 1'b0 ;
  assign n557 = ( n553 & ~n555 ) | ( n553 & n556 ) | ( ~n555 & n556 ) ;
  assign n659 = n657 ^ n224 ^ 1'b0 ;
  assign n660 = ( n657 & n658 ) | ( n657 & ~n659 ) | ( n658 & ~n659 ) ;
  assign n661 = n660 ^ n220 ^ 1'b0 ;
  assign n662 = ( n220 & ~n655 ) | ( n220 & n661 ) | ( ~n655 & n661 ) ;
  assign n663 = ( n660 & ~n661 ) | ( n660 & n662 ) | ( ~n661 & n662 ) ;
  assign n665 = ( n220 & ~n663 ) | ( n220 & n664 ) | ( ~n663 & n664 ) ;
  assign n666 = n665 ^ n663 ^ 1'b0 ;
  assign n667 = ( n663 & ~n665 ) | ( n663 & n666 ) | ( ~n665 & n666 ) ;
  assign n772 = n768 ^ n227 ^ 1'b0 ;
  assign n773 = ( n768 & n771 ) | ( n768 & ~n772 ) | ( n771 & ~n772 ) ;
  assign n775 = ( n229 & ~n773 ) | ( n229 & n774 ) | ( ~n773 & n774 ) ;
  assign n776 = ~n773 & n775 ;
  assign n777 = ( n229 & n769 ) | ( n229 & ~n776 ) | ( n769 & ~n776 ) ;
  assign n778 = n777 ^ n776 ^ 1'b0 ;
  assign n779 = ( n776 & ~n777 ) | ( n776 & n778 ) | ( ~n777 & n778 ) ;
  assign n1584 = ( n557 & n667 ) | ( n557 & n779 ) | ( n667 & n779 ) ;
  assign n1708 = ( n1582 & n1583 ) | ( n1582 & n1584 ) | ( n1583 & n1584 ) ;
  assign n1031 = n218 & ~n952 ;
  assign n1032 = n218 & ~n949 ;
  assign n1033 = ( n953 & ~n1031 ) | ( n953 & n1032 ) | ( ~n1031 & n1032 ) ;
  assign n1034 = ~n1031 & n1033 ;
  assign n1035 = n541 & n840 ;
  assign n1586 = ( ~n948 & n1034 ) | ( ~n948 & n1035 ) | ( n1034 & n1035 ) ;
  assign n1591 = n657 ^ n220 ^ 1'b0 ;
  assign n1592 = ( n657 & n658 ) | ( n657 & ~n1591 ) | ( n658 & ~n1591 ) ;
  assign n1593 = n1592 ^ n227 ^ 1'b0 ;
  assign n1594 = ( n227 & ~n655 ) | ( n227 & n1593 ) | ( ~n655 & n1593 ) ;
  assign n1595 = ( n1592 & ~n1593 ) | ( n1592 & n1594 ) | ( ~n1593 & n1594 ) ;
  assign n1596 = ( n227 & n664 ) | ( n227 & ~n1595 ) | ( n664 & ~n1595 ) ;
  assign n1597 = n1596 ^ n1595 ^ 1'b0 ;
  assign n1598 = ( n1595 & ~n1596 ) | ( n1595 & n1597 ) | ( ~n1596 & n1597 ) ;
  assign n1709 = ( n1586 & ~n1590 ) | ( n1586 & n1598 ) | ( ~n1590 & n1598 ) ;
  assign n1828 = ( ~n1707 & n1708 ) | ( ~n1707 & n1709 ) | ( n1708 & n1709 ) ;
  assign n1710 = n1709 ^ n1708 ^ n1707 ;
  assign n1585 = n1584 ^ n1583 ^ n1582 ;
  assign n1599 = n1598 ^ n1590 ^ n1586 ;
  assign n780 = n779 ^ n667 ^ n557 ;
  assign n847 = n845 ^ n541 ^ 1'b0 ;
  assign n848 = ( n845 & n846 ) | ( n845 & ~n847 ) | ( n846 & ~n847 ) ;
  assign n849 = n848 ^ n544 ^ 1'b0 ;
  assign n850 = ( n544 & ~n843 ) | ( n544 & n849 ) | ( ~n843 & n849 ) ;
  assign n851 = ( n848 & ~n849 ) | ( n848 & n850 ) | ( ~n849 & n850 ) ;
  assign n853 = ( n544 & ~n851 ) | ( n544 & n852 ) | ( ~n851 & n852 ) ;
  assign n854 = n853 ^ n851 ^ 1'b0 ;
  assign n855 = ( n851 & ~n853 ) | ( n851 & n854 ) | ( ~n853 & n854 ) ;
  assign n857 = n840 & n856 ;
  assign n955 = n952 ^ n227 ^ 1'b0 ;
  assign n956 = ( n952 & n954 ) | ( n952 & ~n955 ) | ( n954 & ~n955 ) ;
  assign n957 = n956 ^ n229 ^ 1'b0 ;
  assign n959 = ( n229 & n957 ) | ( n229 & ~n958 ) | ( n957 & ~n958 ) ;
  assign n960 = ( n956 & ~n957 ) | ( n956 & n959 ) | ( ~n957 & n959 ) ;
  assign n962 = ( n229 & ~n960 ) | ( n229 & n961 ) | ( ~n960 & n961 ) ;
  assign n963 = n962 ^ n960 ^ 1'b0 ;
  assign n964 = ( n960 & ~n962 ) | ( n960 & n963 ) | ( ~n962 & n963 ) ;
  assign n965 = n299 | n561 ;
  assign n966 = n316 | n965 ;
  assign n967 = ( n157 & n160 ) | ( n157 & ~n966 ) | ( n160 & ~n966 ) ;
  assign n968 = n966 | n967 ;
  assign n969 = ( n130 & n310 ) | ( n130 & ~n968 ) | ( n310 & ~n968 ) ;
  assign n970 = n968 | n969 ;
  assign n971 = ( n179 & n274 ) | ( n179 & ~n970 ) | ( n274 & ~n970 ) ;
  assign n972 = n970 | n971 ;
  assign n973 = n390 | n448 ;
  assign n976 = ( n698 & ~n973 ) | ( n698 & n975 ) | ( ~n973 & n975 ) ;
  assign n977 = n973 | n976 ;
  assign n978 = ( n315 & n361 ) | ( n315 & ~n977 ) | ( n361 & ~n977 ) ;
  assign n979 = n977 | n978 ;
  assign n980 = ( n187 & n234 ) | ( n187 & ~n979 ) | ( n234 & ~n979 ) ;
  assign n981 = n979 | n980 ;
  assign n982 = ( n146 & n462 ) | ( n146 & ~n981 ) | ( n462 & ~n981 ) ;
  assign n983 = n981 | n982 ;
  assign n984 = ~n233 & n313 ;
  assign n985 = ~n205 & n984 ;
  assign n986 = ( ~n364 & n414 ) | ( ~n364 & n985 ) | ( n414 & n985 ) ;
  assign n987 = ~n414 & n986 ;
  assign n988 = ( n142 & ~n379 ) | ( n142 & n987 ) | ( ~n379 & n987 ) ;
  assign n989 = ~n142 & n988 ;
  assign n990 = ( n92 & ~n213 ) | ( n92 & n989 ) | ( ~n213 & n989 ) ;
  assign n991 = ~n92 & n990 ;
  assign n992 = ~n272 & n991 ;
  assign n993 = ( n818 & ~n983 ) | ( n818 & n992 ) | ( ~n983 & n992 ) ;
  assign n994 = ~n818 & n993 ;
  assign n995 = ( n347 & ~n972 ) | ( n347 & n994 ) | ( ~n972 & n994 ) ;
  assign n996 = ~n347 & n995 ;
  assign n997 = ( n325 & ~n405 ) | ( n325 & n996 ) | ( ~n405 & n996 ) ;
  assign n998 = ~n325 & n997 ;
  assign n999 = ( ~n284 & n564 ) | ( ~n284 & n998 ) | ( n564 & n998 ) ;
  assign n1000 = ~n564 & n999 ;
  assign n1001 = ( ~n164 & n426 ) | ( ~n164 & n1000 ) | ( n426 & n1000 ) ;
  assign n1002 = ~n426 & n1001 ;
  assign n1003 = n948 | n1002 ;
  assign n1004 = ( n218 & n948 ) | ( n218 & n1003 ) | ( n948 & n1003 ) ;
  assign n1005 = ( n857 & n964 ) | ( n857 & ~n1004 ) | ( n964 & ~n1004 ) ;
  assign n1006 = n658 ^ n548 ^ 1'b0 ;
  assign n1007 = ( n657 & n658 ) | ( n657 & n1006 ) | ( n658 & n1006 ) ;
  assign n1008 = n1007 ^ n222 ^ 1'b0 ;
  assign n1009 = ( n222 & ~n655 ) | ( n222 & n1008 ) | ( ~n655 & n1008 ) ;
  assign n1010 = ( n1007 & ~n1008 ) | ( n1007 & n1009 ) | ( ~n1008 & n1009 ) ;
  assign n1011 = ( n222 & n664 ) | ( n222 & ~n1010 ) | ( n664 & ~n1010 ) ;
  assign n1012 = n1011 ^ n1010 ^ 1'b0 ;
  assign n1013 = ( n1010 & ~n1011 ) | ( n1010 & n1012 ) | ( ~n1011 & n1012 ) ;
  assign n1014 = n768 ^ n224 ^ 1'b0 ;
  assign n1015 = ( n768 & n771 ) | ( n768 & ~n1014 ) | ( n771 & ~n1014 ) ;
  assign n1016 = ( n220 & n774 ) | ( n220 & ~n1015 ) | ( n774 & ~n1015 ) ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1018 = ( n220 & n769 ) | ( n220 & ~n1017 ) | ( n769 & ~n1017 ) ;
  assign n1019 = n1018 ^ n1017 ^ 1'b0 ;
  assign n1020 = ( n1017 & ~n1018 ) | ( n1017 & n1019 ) | ( ~n1018 & n1019 ) ;
  assign n1021 = n544 ^ n533 ^ 1'b0 ;
  assign n1022 = ( n533 & n534 ) | ( n533 & ~n1021 ) | ( n534 & ~n1021 ) ;
  assign n1023 = n1022 ^ n545 ^ 1'b0 ;
  assign n1024 = ( ~n531 & n545 ) | ( ~n531 & n1023 ) | ( n545 & n1023 ) ;
  assign n1025 = ( n1022 & ~n1023 ) | ( n1022 & n1024 ) | ( ~n1023 & n1024 ) ;
  assign n1026 = ( n545 & n554 ) | ( n545 & ~n1025 ) | ( n554 & ~n1025 ) ;
  assign n1027 = n1026 ^ n1025 ^ 1'b0 ;
  assign n1028 = ( n1025 & ~n1026 ) | ( n1025 & n1027 ) | ( ~n1026 & n1027 ) ;
  assign n1029 = ( n1013 & n1020 ) | ( n1013 & n1028 ) | ( n1020 & n1028 ) ;
  assign n1030 = ( n855 & n1005 ) | ( n855 & n1029 ) | ( n1005 & n1029 ) ;
  assign n1036 = n1035 ^ n1034 ^ n948 ;
  assign n1600 = ( n780 & n1030 ) | ( n780 & ~n1036 ) | ( n1030 & ~n1036 ) ;
  assign n1711 = ( n1585 & ~n1599 ) | ( n1585 & n1600 ) | ( ~n1599 & n1600 ) ;
  assign n1601 = n1600 ^ n1599 ^ n1585 ;
  assign n1037 = n1036 ^ n1030 ^ n780 ;
  assign n1057 = n1056 ^ n1048 ^ 1'b0 ;
  assign n1082 = n1081 ^ n1057 ^ 1'b0 ;
  assign n1083 = n229 | n948 ;
  assign n1084 = n1002 & n1083 ;
  assign n1085 = n948 & ~n1002 ;
  assign n1086 = ~n218 & n1085 ;
  assign n1087 = n1084 | n1086 ;
  assign n1088 = n1003 & ~n1087 ;
  assign n1089 = ( n218 & n1087 ) | ( n218 & ~n1088 ) | ( n1087 & ~n1088 ) ;
  assign n1090 = n852 & n856 ;
  assign n1091 = ( n842 & n846 ) | ( n842 & n856 ) | ( n846 & n856 ) ;
  assign n1092 = ~n1090 & n1091 ;
  assign n1093 = n842 & n1092 ;
  assign n1094 = ~n1089 & n1093 ;
  assign n1095 = n1040 ^ n845 ^ 1'b0 ;
  assign n1096 = ( n845 & n846 ) | ( n845 & ~n1095 ) | ( n846 & ~n1095 ) ;
  assign n1097 = n1096 ^ n541 ^ 1'b0 ;
  assign n1098 = ( n541 & ~n843 ) | ( n541 & n1097 ) | ( ~n843 & n1097 ) ;
  assign n1099 = ( n1096 & ~n1097 ) | ( n1096 & n1098 ) | ( ~n1097 & n1098 ) ;
  assign n1100 = ( n541 & n852 ) | ( n541 & ~n1099 ) | ( n852 & ~n1099 ) ;
  assign n1101 = n1100 ^ n1099 ^ 1'b0 ;
  assign n1102 = ( n1099 & ~n1100 ) | ( n1099 & n1101 ) | ( ~n1100 & n1101 ) ;
  assign n1103 = n658 ^ n545 ^ 1'b0 ;
  assign n1104 = ( n657 & n658 ) | ( n657 & n1103 ) | ( n658 & n1103 ) ;
  assign n1105 = n1104 ^ n548 ^ 1'b0 ;
  assign n1106 = ( n548 & ~n655 ) | ( n548 & n1105 ) | ( ~n655 & n1105 ) ;
  assign n1107 = ( n1104 & ~n1105 ) | ( n1104 & n1106 ) | ( ~n1105 & n1106 ) ;
  assign n1108 = ( n548 & n664 ) | ( n548 & ~n1107 ) | ( n664 & ~n1107 ) ;
  assign n1109 = n1108 ^ n1107 ^ 1'b0 ;
  assign n1110 = ( n1107 & ~n1108 ) | ( n1107 & n1109 ) | ( ~n1108 & n1109 ) ;
  assign n1111 = n541 ^ n533 ^ 1'b0 ;
  assign n1112 = ( n533 & n534 ) | ( n533 & ~n1111 ) | ( n534 & ~n1111 ) ;
  assign n1113 = n1112 ^ n544 ^ 1'b0 ;
  assign n1114 = ( ~n531 & n544 ) | ( ~n531 & n1113 ) | ( n544 & n1113 ) ;
  assign n1115 = ( n1112 & ~n1113 ) | ( n1112 & n1114 ) | ( ~n1113 & n1114 ) ;
  assign n1116 = ( n544 & n554 ) | ( n544 & ~n1115 ) | ( n554 & ~n1115 ) ;
  assign n1117 = n1116 ^ n1115 ^ 1'b0 ;
  assign n1118 = ( n1115 & ~n1116 ) | ( n1115 & n1117 ) | ( ~n1116 & n1117 ) ;
  assign n1119 = n768 ^ n222 ^ 1'b0 ;
  assign n1120 = ( n768 & n771 ) | ( n768 & ~n1119 ) | ( n771 & ~n1119 ) ;
  assign n1121 = ( n224 & n774 ) | ( n224 & ~n1120 ) | ( n774 & ~n1120 ) ;
  assign n1122 = ~n1120 & n1121 ;
  assign n1123 = ( n224 & n769 ) | ( n224 & ~n1122 ) | ( n769 & ~n1122 ) ;
  assign n1124 = n1123 ^ n1122 ^ 1'b0 ;
  assign n1125 = ( n1122 & ~n1123 ) | ( n1122 & n1124 ) | ( ~n1123 & n1124 ) ;
  assign n1126 = ( n1110 & n1118 ) | ( n1110 & n1125 ) | ( n1118 & n1125 ) ;
  assign n1127 = ( n1094 & n1102 ) | ( n1094 & n1126 ) | ( n1102 & n1126 ) ;
  assign n1128 = n1047 ^ n1041 ^ n948 ;
  assign n1129 = n1080 ^ n1072 ^ n1065 ;
  assign n1130 = ( n1127 & ~n1128 ) | ( n1127 & n1129 ) | ( ~n1128 & n1129 ) ;
  assign n1602 = ( ~n1037 & n1082 ) | ( ~n1037 & n1130 ) | ( n1082 & n1130 ) ;
  assign n1131 = n1130 ^ n1082 ^ n1037 ;
  assign n1132 = n952 ^ n220 ^ 1'b0 ;
  assign n1133 = ( n952 & n954 ) | ( n952 & ~n1132 ) | ( n954 & ~n1132 ) ;
  assign n1134 = n1133 ^ n227 ^ 1'b0 ;
  assign n1135 = ( n227 & ~n958 ) | ( n227 & n1134 ) | ( ~n958 & n1134 ) ;
  assign n1136 = ( n1133 & ~n1134 ) | ( n1133 & n1135 ) | ( ~n1134 & n1135 ) ;
  assign n1137 = ( n227 & n961 ) | ( n227 & ~n1136 ) | ( n961 & ~n1136 ) ;
  assign n1138 = n1137 ^ n1136 ^ 1'b0 ;
  assign n1139 = ( n1136 & ~n1137 ) | ( n1136 & n1138 ) | ( ~n1137 & n1138 ) ;
  assign n1140 = n856 ^ n845 ^ 1'b0 ;
  assign n1141 = ( n845 & n846 ) | ( n845 & ~n1140 ) | ( n846 & ~n1140 ) ;
  assign n1142 = n1141 ^ n1040 ^ 1'b0 ;
  assign n1143 = ( ~n843 & n1040 ) | ( ~n843 & n1142 ) | ( n1040 & n1142 ) ;
  assign n1144 = ( n1141 & ~n1142 ) | ( n1141 & n1143 ) | ( ~n1142 & n1143 ) ;
  assign n1145 = ( n852 & n1040 ) | ( n852 & ~n1144 ) | ( n1040 & ~n1144 ) ;
  assign n1146 = n1145 ^ n1144 ^ 1'b0 ;
  assign n1147 = ( n1144 & ~n1145 ) | ( n1144 & n1146 ) | ( ~n1145 & n1146 ) ;
  assign n1148 = n1093 ^ n1089 ^ 1'b0 ;
  assign n1149 = ( n1139 & n1147 ) | ( n1139 & ~n1148 ) | ( n1147 & ~n1148 ) ;
  assign n1150 = n1004 ^ n857 ^ 1'b0 ;
  assign n1151 = n1150 ^ n964 ^ 1'b0 ;
  assign n1152 = n1028 ^ n1020 ^ n1013 ;
  assign n1153 = ( n1149 & ~n1151 ) | ( n1149 & n1152 ) | ( ~n1151 & n1152 ) ;
  assign n1154 = n1005 ^ n855 ^ 1'b0 ;
  assign n1155 = n1154 ^ n1029 ^ 1'b0 ;
  assign n1156 = n1129 ^ n1128 ^ n1127 ;
  assign n1157 = ( n1153 & n1155 ) | ( n1153 & ~n1156 ) | ( n1155 & ~n1156 ) ;
  assign n1159 = n1151 ^ n1149 ^ 1'b0 ;
  assign n1160 = n1159 ^ n1152 ^ 1'b0 ;
  assign n1161 = n220 | n948 ;
  assign n1162 = n1002 & n1161 ;
  assign n1163 = ~n227 & n1085 ;
  assign n1164 = n1162 | n1163 ;
  assign n1165 = n1003 & ~n1164 ;
  assign n1166 = ( n227 & n1164 ) | ( n227 & ~n1165 ) | ( n1164 & ~n1165 ) ;
  assign n1167 = n490 & n856 ;
  assign n1168 = n1167 ^ n534 ^ n531 ;
  assign n1169 = n530 & n1168 ;
  assign n1170 = ~n1166 & n1169 ;
  assign n1171 = n768 ^ n548 ^ 1'b0 ;
  assign n1172 = ( n768 & n771 ) | ( n768 & ~n1171 ) | ( n771 & ~n1171 ) ;
  assign n1173 = ( n222 & n774 ) | ( n222 & ~n1172 ) | ( n774 & ~n1172 ) ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = ( n222 & n769 ) | ( n222 & ~n1174 ) | ( n769 & ~n1174 ) ;
  assign n1176 = n1175 ^ n1174 ^ 1'b0 ;
  assign n1177 = ( n1174 & ~n1175 ) | ( n1174 & n1176 ) | ( ~n1175 & n1176 ) ;
  assign n1178 = n657 ^ n544 ^ 1'b0 ;
  assign n1179 = ( n657 & n658 ) | ( n657 & ~n1178 ) | ( n658 & ~n1178 ) ;
  assign n1180 = n1179 ^ n545 ^ 1'b0 ;
  assign n1181 = ( n545 & ~n655 ) | ( n545 & n1180 ) | ( ~n655 & n1180 ) ;
  assign n1182 = ( n1179 & ~n1180 ) | ( n1179 & n1181 ) | ( ~n1180 & n1181 ) ;
  assign n1183 = ( n545 & n664 ) | ( n545 & ~n1182 ) | ( n664 & ~n1182 ) ;
  assign n1184 = n1183 ^ n1182 ^ 1'b0 ;
  assign n1185 = ( n1182 & ~n1183 ) | ( n1182 & n1184 ) | ( ~n1183 & n1184 ) ;
  assign n1186 = ( n1170 & n1177 ) | ( n1170 & n1185 ) | ( n1177 & n1185 ) ;
  assign n1187 = n227 | n948 ;
  assign n1188 = n1002 & n1187 ;
  assign n1189 = ~n229 & n1085 ;
  assign n1190 = n1188 | n1189 ;
  assign n1191 = n1003 & ~n1190 ;
  assign n1192 = ( n229 & n1190 ) | ( n229 & ~n1191 ) | ( n1190 & ~n1191 ) ;
  assign n1193 = n952 ^ n224 ^ 1'b0 ;
  assign n1194 = ( n952 & n954 ) | ( n952 & ~n1193 ) | ( n954 & ~n1193 ) ;
  assign n1195 = n1194 ^ n220 ^ 1'b0 ;
  assign n1196 = ( n220 & ~n958 ) | ( n220 & n1195 ) | ( ~n958 & n1195 ) ;
  assign n1197 = ( n1194 & ~n1195 ) | ( n1194 & n1196 ) | ( ~n1195 & n1196 ) ;
  assign n1198 = ( n220 & n961 ) | ( n220 & ~n1197 ) | ( n961 & ~n1197 ) ;
  assign n1199 = n1198 ^ n1197 ^ 1'b0 ;
  assign n1200 = ( n1197 & ~n1198 ) | ( n1197 & n1199 ) | ( ~n1198 & n1199 ) ;
  assign n1201 = n1040 ^ n533 ^ 1'b0 ;
  assign n1202 = ( n533 & n534 ) | ( n533 & ~n1201 ) | ( n534 & ~n1201 ) ;
  assign n1203 = n1202 ^ n541 ^ 1'b0 ;
  assign n1204 = ( ~n531 & n541 ) | ( ~n531 & n1203 ) | ( n541 & n1203 ) ;
  assign n1205 = ( n1202 & ~n1203 ) | ( n1202 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = ( n541 & n554 ) | ( n541 & ~n1205 ) | ( n554 & ~n1205 ) ;
  assign n1207 = n1206 ^ n1205 ^ 1'b0 ;
  assign n1208 = ( n1205 & ~n1206 ) | ( n1205 & n1207 ) | ( ~n1206 & n1207 ) ;
  assign n1209 = ( ~n1192 & n1200 ) | ( ~n1192 & n1208 ) | ( n1200 & n1208 ) ;
  assign n1210 = n1125 ^ n1118 ^ n1110 ;
  assign n1211 = ( n1186 & n1209 ) | ( n1186 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = n1102 ^ n1094 ^ 1'b0 ;
  assign n1213 = n1212 ^ n1126 ^ 1'b0 ;
  assign n1214 = ( ~n1160 & n1211 ) | ( ~n1160 & n1213 ) | ( n1211 & n1213 ) ;
  assign n1215 = n952 ^ n222 ^ 1'b0 ;
  assign n1216 = ( n952 & n954 ) | ( n952 & ~n1215 ) | ( n954 & ~n1215 ) ;
  assign n1217 = n1216 ^ n224 ^ 1'b0 ;
  assign n1218 = ( n224 & ~n958 ) | ( n224 & n1217 ) | ( ~n958 & n1217 ) ;
  assign n1219 = ( n1216 & ~n1217 ) | ( n1216 & n1218 ) | ( ~n1217 & n1218 ) ;
  assign n1220 = ( n224 & n961 ) | ( n224 & ~n1219 ) | ( n961 & ~n1219 ) ;
  assign n1221 = n1220 ^ n1219 ^ 1'b0 ;
  assign n1222 = ( n1219 & ~n1220 ) | ( n1219 & n1221 ) | ( ~n1220 & n1221 ) ;
  assign n1223 = n657 ^ n541 ^ 1'b0 ;
  assign n1224 = ( n657 & n658 ) | ( n657 & ~n1223 ) | ( n658 & ~n1223 ) ;
  assign n1225 = n1224 ^ n544 ^ 1'b0 ;
  assign n1226 = ( n544 & ~n655 ) | ( n544 & n1225 ) | ( ~n655 & n1225 ) ;
  assign n1227 = ( n1224 & ~n1225 ) | ( n1224 & n1226 ) | ( ~n1225 & n1226 ) ;
  assign n1228 = ( n544 & n664 ) | ( n544 & ~n1227 ) | ( n664 & ~n1227 ) ;
  assign n1229 = n1228 ^ n1227 ^ 1'b0 ;
  assign n1230 = ( n1227 & ~n1228 ) | ( n1227 & n1229 ) | ( ~n1228 & n1229 ) ;
  assign n1231 = n768 ^ n545 ^ 1'b0 ;
  assign n1232 = ( n768 & n771 ) | ( n768 & ~n1231 ) | ( n771 & ~n1231 ) ;
  assign n1233 = ( n548 & n774 ) | ( n548 & ~n1232 ) | ( n774 & ~n1232 ) ;
  assign n1234 = ~n1232 & n1233 ;
  assign n1235 = ( n548 & n769 ) | ( n548 & ~n1234 ) | ( n769 & ~n1234 ) ;
  assign n1236 = n1235 ^ n1234 ^ 1'b0 ;
  assign n1237 = ( n1234 & ~n1235 ) | ( n1234 & n1236 ) | ( ~n1235 & n1236 ) ;
  assign n1238 = ( n1222 & n1230 ) | ( n1222 & n1237 ) | ( n1230 & n1237 ) ;
  assign n1239 = ~n1093 & n1238 ;
  assign n1240 = n1091 & n1239 ;
  assign n1241 = n1238 ^ n1092 ^ n842 ;
  assign n1242 = n1185 ^ n1177 ^ n1170 ;
  assign n1243 = n1241 & n1242 ;
  assign n1244 = n1240 | n1243 ;
  assign n1245 = n1148 ^ n1147 ^ n1139 ;
  assign n1246 = n1210 ^ n1209 ^ n1186 ;
  assign n1247 = ( n1244 & ~n1245 ) | ( n1244 & n1246 ) | ( ~n1245 & n1246 ) ;
  assign n1248 = n1245 ^ n1244 ^ 1'b0 ;
  assign n1249 = ~n1246 & n1248 ;
  assign n1250 = n1246 & ~n1248 ;
  assign n1251 = n224 | n948 ;
  assign n1252 = n1002 & n1251 ;
  assign n1253 = ~n220 & n1085 ;
  assign n1254 = n1252 | n1253 ;
  assign n1255 = n1003 & ~n1254 ;
  assign n1256 = ( n220 & n1254 ) | ( n220 & ~n1255 ) | ( n1254 & ~n1255 ) ;
  assign n1257 = n952 ^ n548 ^ 1'b0 ;
  assign n1258 = ( n952 & n954 ) | ( n952 & ~n1257 ) | ( n954 & ~n1257 ) ;
  assign n1259 = n1258 ^ n222 ^ 1'b0 ;
  assign n1260 = ( n222 & ~n958 ) | ( n222 & n1259 ) | ( ~n958 & n1259 ) ;
  assign n1261 = ( n1258 & ~n1259 ) | ( n1258 & n1260 ) | ( ~n1259 & n1260 ) ;
  assign n1262 = ( n222 & n961 ) | ( n222 & ~n1261 ) | ( n961 & ~n1261 ) ;
  assign n1263 = n1262 ^ n1261 ^ 1'b0 ;
  assign n1264 = ( n1261 & ~n1262 ) | ( n1261 & n1263 ) | ( ~n1262 & n1263 ) ;
  assign n1265 = n768 ^ n544 ^ 1'b0 ;
  assign n1266 = ( n768 & n771 ) | ( n768 & ~n1265 ) | ( n771 & ~n1265 ) ;
  assign n1267 = ( n545 & n774 ) | ( n545 & ~n1266 ) | ( n774 & ~n1266 ) ;
  assign n1268 = ~n1266 & n1267 ;
  assign n1269 = ( n545 & n769 ) | ( n545 & ~n1268 ) | ( n769 & ~n1268 ) ;
  assign n1270 = n1269 ^ n1268 ^ 1'b0 ;
  assign n1271 = ( n1268 & ~n1269 ) | ( n1268 & n1270 ) | ( ~n1269 & n1270 ) ;
  assign n1272 = ( ~n1256 & n1264 ) | ( ~n1256 & n1271 ) | ( n1264 & n1271 ) ;
  assign n1273 = n856 ^ n533 ^ 1'b0 ;
  assign n1274 = ( n533 & n534 ) | ( n533 & ~n1273 ) | ( n534 & ~n1273 ) ;
  assign n1275 = n1274 ^ n1040 ^ 1'b0 ;
  assign n1276 = ( ~n531 & n1040 ) | ( ~n531 & n1275 ) | ( n1040 & n1275 ) ;
  assign n1277 = ( n1274 & ~n1275 ) | ( n1274 & n1276 ) | ( ~n1275 & n1276 ) ;
  assign n1278 = ( n554 & n1040 ) | ( n554 & ~n1277 ) | ( n1040 & ~n1277 ) ;
  assign n1279 = n1278 ^ n1277 ^ 1'b0 ;
  assign n1280 = ( n1277 & ~n1278 ) | ( n1277 & n1279 ) | ( ~n1278 & n1279 ) ;
  assign n1281 = n1169 ^ n1166 ^ 1'b0 ;
  assign n1282 = ( n1272 & n1280 ) | ( n1272 & ~n1281 ) | ( n1280 & ~n1281 ) ;
  assign n1283 = n1242 ^ n1241 ^ 1'b0 ;
  assign n1284 = n1208 ^ n1200 ^ n1192 ;
  assign n1285 = ( n1282 & n1283 ) | ( n1282 & ~n1284 ) | ( n1283 & ~n1284 ) ;
  assign n1286 = n952 ^ n545 ^ 1'b0 ;
  assign n1287 = ( n952 & n954 ) | ( n952 & ~n1286 ) | ( n954 & ~n1286 ) ;
  assign n1288 = n1287 ^ n548 ^ 1'b0 ;
  assign n1289 = ( n548 & ~n958 ) | ( n548 & n1288 ) | ( ~n958 & n1288 ) ;
  assign n1290 = ( n1287 & ~n1288 ) | ( n1287 & n1289 ) | ( ~n1288 & n1289 ) ;
  assign n1291 = ( n548 & n961 ) | ( n548 & ~n1290 ) | ( n961 & ~n1290 ) ;
  assign n1292 = n1291 ^ n1290 ^ 1'b0 ;
  assign n1293 = ( n1290 & ~n1291 ) | ( n1290 & n1292 ) | ( ~n1291 & n1292 ) ;
  assign n1294 = n768 ^ n541 ^ 1'b0 ;
  assign n1295 = ( n768 & n771 ) | ( n768 & ~n1294 ) | ( n771 & ~n1294 ) ;
  assign n1296 = ( n544 & n774 ) | ( n544 & ~n1295 ) | ( n774 & ~n1295 ) ;
  assign n1297 = ~n1295 & n1296 ;
  assign n1298 = ( n544 & n769 ) | ( n544 & ~n1297 ) | ( n769 & ~n1297 ) ;
  assign n1299 = n1298 ^ n1297 ^ 1'b0 ;
  assign n1300 = ( n1297 & ~n1298 ) | ( n1297 & n1299 ) | ( ~n1298 & n1299 ) ;
  assign n1301 = n856 ^ n657 ^ 1'b0 ;
  assign n1302 = ( n657 & n658 ) | ( n657 & ~n1301 ) | ( n658 & ~n1301 ) ;
  assign n1303 = n1302 ^ n1040 ^ 1'b0 ;
  assign n1304 = ( ~n655 & n1040 ) | ( ~n655 & n1303 ) | ( n1040 & n1303 ) ;
  assign n1305 = ( n1302 & ~n1303 ) | ( n1302 & n1304 ) | ( ~n1303 & n1304 ) ;
  assign n1306 = ( n664 & n1040 ) | ( n664 & ~n1305 ) | ( n1040 & ~n1305 ) ;
  assign n1307 = n1306 ^ n1305 ^ 1'b0 ;
  assign n1308 = ( n1305 & ~n1306 ) | ( n1305 & n1307 ) | ( ~n1306 & n1307 ) ;
  assign n1309 = ( n1293 & n1300 ) | ( n1293 & n1308 ) | ( n1300 & n1308 ) ;
  assign n1310 = n1271 ^ n1264 ^ n1256 ;
  assign n1322 = n1040 ^ n657 ^ 1'b0 ;
  assign n1323 = ( n657 & n658 ) | ( n657 & ~n1322 ) | ( n658 & ~n1322 ) ;
  assign n1324 = n1323 ^ n541 ^ 1'b0 ;
  assign n1325 = ( n541 & ~n655 ) | ( n541 & n1324 ) | ( ~n655 & n1324 ) ;
  assign n1326 = ( n1323 & ~n1324 ) | ( n1323 & n1325 ) | ( ~n1324 & n1325 ) ;
  assign n1327 = ( n541 & n664 ) | ( n541 & ~n1326 ) | ( n664 & ~n1326 ) ;
  assign n1328 = n1327 ^ n1326 ^ 1'b0 ;
  assign n1329 = ( n1326 & ~n1327 ) | ( n1326 & n1328 ) | ( ~n1327 & n1328 ) ;
  assign n1311 = n222 | n948 ;
  assign n1312 = n1002 & n1311 ;
  assign n1313 = ~n224 & n1085 ;
  assign n1314 = n1312 | n1313 ;
  assign n1315 = n1003 & ~n1314 ;
  assign n1316 = ( n224 & n1314 ) | ( n224 & ~n1315 ) | ( n1314 & ~n1315 ) ;
  assign n1317 = n664 & n856 ;
  assign n1318 = ( n654 & n658 ) | ( n654 & n856 ) | ( n658 & n856 ) ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1320 = n654 & n1319 ;
  assign n1321 = ~n1316 & n1320 ;
  assign n1330 = n1329 ^ n1321 ^ n1167 ;
  assign n1331 = ( n1309 & ~n1310 ) | ( n1309 & n1330 ) | ( ~n1310 & n1330 ) ;
  assign n1332 = ~n548 & n1085 ;
  assign n1333 = n548 & ~n1003 ;
  assign n1334 = n545 | n948 ;
  assign n1335 = n1002 & n1334 ;
  assign n1336 = ( ~n1332 & n1333 ) | ( ~n1332 & n1335 ) | ( n1333 & n1335 ) ;
  assign n1337 = n1332 | n1336 ;
  assign n1338 = ~n765 & n856 ;
  assign n1339 = n1338 ^ n774 ^ n771 ;
  assign n1340 = n770 & n1339 ;
  assign n1341 = ~n1337 & n1340 ;
  assign n1342 = ~n1320 & n1341 ;
  assign n1343 = n1318 & n1342 ;
  assign n1344 = n952 ^ n541 ^ 1'b0 ;
  assign n1345 = ( n952 & n954 ) | ( n952 & ~n1344 ) | ( n954 & ~n1344 ) ;
  assign n1346 = n1345 ^ n544 ^ 1'b0 ;
  assign n1347 = ( n544 & ~n958 ) | ( n544 & n1346 ) | ( ~n958 & n1346 ) ;
  assign n1348 = ( n1345 & ~n1346 ) | ( n1345 & n1347 ) | ( ~n1346 & n1347 ) ;
  assign n1349 = ( n544 & n961 ) | ( n544 & ~n1348 ) | ( n961 & ~n1348 ) ;
  assign n1350 = n1349 ^ n1348 ^ 1'b0 ;
  assign n1351 = ( n1348 & ~n1349 ) | ( n1348 & n1350 ) | ( ~n1349 & n1350 ) ;
  assign n1352 = n856 ^ n768 ^ 1'b0 ;
  assign n1353 = ( n768 & n771 ) | ( n768 & ~n1352 ) | ( n771 & ~n1352 ) ;
  assign n1354 = ( n774 & n1040 ) | ( n774 & ~n1353 ) | ( n1040 & ~n1353 ) ;
  assign n1355 = ~n1353 & n1354 ;
  assign n1356 = ( n769 & n1040 ) | ( n769 & ~n1355 ) | ( n1040 & ~n1355 ) ;
  assign n1357 = n1356 ^ n1355 ^ 1'b0 ;
  assign n1358 = ( n1355 & ~n1356 ) | ( n1355 & n1357 ) | ( ~n1356 & n1357 ) ;
  assign n1359 = n1340 ^ n1337 ^ 1'b0 ;
  assign n1360 = ( n1351 & n1358 ) | ( n1351 & ~n1359 ) | ( n1358 & ~n1359 ) ;
  assign n1361 = n1341 ^ n1319 ^ n654 ;
  assign n1362 = n1360 & n1361 ;
  assign n1363 = n1343 | n1362 ;
  assign n1364 = n961 & n1040 ;
  assign n1365 = n856 & ~n952 ;
  assign n1366 = n856 & n961 ;
  assign n1367 = ( n856 & n953 ) | ( n856 & n954 ) | ( n953 & n954 ) ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = n953 & n1368 ;
  assign n1370 = ~n541 & n1085 ;
  assign n1371 = n541 & ~n1003 ;
  assign n1372 = n948 | n1040 ;
  assign n1373 = n1002 & n1372 ;
  assign n1374 = ( ~n1370 & n1371 ) | ( ~n1370 & n1373 ) | ( n1371 & n1373 ) ;
  assign n1375 = n1370 | n1374 ;
  assign n1376 = ~n1002 & n1040 ;
  assign n1377 = n856 | n948 ;
  assign n1378 = n1376 | n1377 ;
  assign n1379 = n1375 & n1378 ;
  assign n1380 = ( n1367 & n1369 ) | ( n1367 & ~n1379 ) | ( n1369 & ~n1379 ) ;
  assign n1381 = ~n1369 & n1380 ;
  assign n1382 = ( n1375 & n1378 ) | ( n1375 & ~n1381 ) | ( n1378 & ~n1381 ) ;
  assign n1383 = ~n1381 & n1382 ;
  assign n1384 = n541 | n948 ;
  assign n1385 = n1002 & n1384 ;
  assign n1386 = ~n544 & n1085 ;
  assign n1387 = n1385 | n1386 ;
  assign n1388 = n1003 & ~n1387 ;
  assign n1389 = ( n544 & n1387 ) | ( n544 & ~n1388 ) | ( n1387 & ~n1388 ) ;
  assign n1390 = n1389 ^ n1369 ^ 1'b0 ;
  assign n1391 = n1383 & n1390 ;
  assign n1392 = n856 | n954 ;
  assign n1393 = ( n1365 & ~n1391 ) | ( n1365 & n1392 ) | ( ~n1391 & n1392 ) ;
  assign n1394 = ~n1365 & n1393 ;
  assign n1395 = n958 & ~n1040 ;
  assign n1396 = ( n1364 & n1394 ) | ( n1364 & ~n1395 ) | ( n1394 & ~n1395 ) ;
  assign n1397 = ~n1364 & n1396 ;
  assign n1398 = ( n1383 & n1390 ) | ( n1383 & ~n1397 ) | ( n1390 & ~n1397 ) ;
  assign n1399 = ~n1397 & n1398 ;
  assign n1400 = n1338 & ~n1399 ;
  assign n1409 = n544 | n948 ;
  assign n1410 = n1002 & n1409 ;
  assign n1411 = ~n545 & n1085 ;
  assign n1412 = n1410 | n1411 ;
  assign n1413 = n1003 & ~n1412 ;
  assign n1414 = ( n545 & n1412 ) | ( n545 & ~n1413 ) | ( n1412 & ~n1413 ) ;
  assign n1401 = n1040 ^ n952 ^ 1'b0 ;
  assign n1402 = ( n952 & n954 ) | ( n952 & ~n1401 ) | ( n954 & ~n1401 ) ;
  assign n1403 = n1402 ^ n541 ^ 1'b0 ;
  assign n1404 = ( n541 & ~n958 ) | ( n541 & n1403 ) | ( ~n958 & n1403 ) ;
  assign n1405 = ( n1402 & ~n1403 ) | ( n1402 & n1404 ) | ( ~n1403 & n1404 ) ;
  assign n1406 = ( n541 & n961 ) | ( n541 & ~n1405 ) | ( n961 & ~n1405 ) ;
  assign n1407 = n1406 ^ n1405 ^ 1'b0 ;
  assign n1408 = ( n1405 & ~n1406 ) | ( n1405 & n1407 ) | ( ~n1406 & n1407 ) ;
  assign n1415 = n1414 ^ n1408 ^ 1'b0 ;
  assign n1416 = n1369 & ~n1389 ;
  assign n1417 = n1415 & ~n1416 ;
  assign n1418 = ~n1415 & n1416 ;
  assign n1419 = ~n1338 & n1399 ;
  assign n1420 = n1418 | n1419 ;
  assign n1421 = ( ~n1400 & n1417 ) | ( ~n1400 & n1420 ) | ( n1417 & n1420 ) ;
  assign n1422 = ~n1400 & n1421 ;
  assign n1423 = n1359 ^ n1358 ^ n1351 ;
  assign n1424 = ( n1408 & ~n1414 ) | ( n1408 & n1416 ) | ( ~n1414 & n1416 ) ;
  assign n1425 = ( n1422 & n1423 ) | ( n1422 & ~n1424 ) | ( n1423 & ~n1424 ) ;
  assign n1426 = n1361 ^ n1360 ^ 1'b0 ;
  assign n1427 = ~n1425 & n1426 ;
  assign n1428 = n1040 ^ n768 ^ 1'b0 ;
  assign n1429 = ( n768 & n771 ) | ( n768 & ~n1428 ) | ( n771 & ~n1428 ) ;
  assign n1430 = ( n541 & n774 ) | ( n541 & ~n1429 ) | ( n774 & ~n1429 ) ;
  assign n1431 = ~n1429 & n1430 ;
  assign n1432 = ( n541 & n769 ) | ( n541 & ~n1431 ) | ( n769 & ~n1431 ) ;
  assign n1433 = n1432 ^ n1431 ^ 1'b0 ;
  assign n1434 = ( n1431 & ~n1432 ) | ( n1431 & n1433 ) | ( ~n1432 & n1433 ) ;
  assign n1441 = n952 ^ n544 ^ 1'b0 ;
  assign n1442 = ( n952 & n954 ) | ( n952 & ~n1441 ) | ( n954 & ~n1441 ) ;
  assign n1443 = n1442 ^ n545 ^ 1'b0 ;
  assign n1444 = ( n545 & ~n958 ) | ( n545 & n1443 ) | ( ~n958 & n1443 ) ;
  assign n1445 = ( n1442 & ~n1443 ) | ( n1442 & n1444 ) | ( ~n1443 & n1444 ) ;
  assign n1446 = ( n545 & n961 ) | ( n545 & ~n1445 ) | ( n961 & ~n1445 ) ;
  assign n1447 = n1446 ^ n1445 ^ 1'b0 ;
  assign n1448 = ( n1445 & ~n1446 ) | ( n1445 & n1447 ) | ( ~n1446 & n1447 ) ;
  assign n1435 = n548 | n948 ;
  assign n1436 = n1002 & n1435 ;
  assign n1437 = ~n222 & n1085 ;
  assign n1438 = n1436 | n1437 ;
  assign n1439 = n1003 & ~n1438 ;
  assign n1440 = ( n222 & n1438 ) | ( n222 & ~n1439 ) | ( n1438 & ~n1439 ) ;
  assign n1449 = n1448 ^ n1440 ^ 1'b0 ;
  assign n1450 = ~n1434 & n1449 ;
  assign n1451 = n1434 & ~n1449 ;
  assign n1452 = n1425 & ~n1426 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = ( ~n1427 & n1450 ) | ( ~n1427 & n1453 ) | ( n1450 & n1453 ) ;
  assign n1455 = ~n1427 & n1454 ;
  assign n1458 = n1320 ^ n1316 ^ 1'b0 ;
  assign n1457 = ( n1434 & ~n1440 ) | ( n1434 & n1448 ) | ( ~n1440 & n1448 ) ;
  assign n1456 = n1308 ^ n1300 ^ n1293 ;
  assign n1459 = n1458 ^ n1457 ^ n1456 ;
  assign n1460 = ( ~n1363 & n1455 ) | ( ~n1363 & n1459 ) | ( n1455 & n1459 ) ;
  assign n1461 = ( n1456 & n1457 ) | ( n1456 & ~n1458 ) | ( n1457 & ~n1458 ) ;
  assign n1462 = n1330 ^ n1310 ^ n1309 ;
  assign n1463 = ( n1460 & ~n1461 ) | ( n1460 & n1462 ) | ( ~n1461 & n1462 ) ;
  assign n1464 = ~n1331 & n1463 ;
  assign n1466 = ( n1167 & n1321 ) | ( n1167 & n1329 ) | ( n1321 & n1329 ) ;
  assign n1465 = n1237 ^ n1230 ^ n1222 ;
  assign n1467 = n1466 ^ n1465 ^ 1'b0 ;
  assign n1468 = n1281 ^ n1280 ^ n1272 ;
  assign n1469 = ~n1467 & n1468 ;
  assign n1470 = n1467 & ~n1468 ;
  assign n1471 = ( ~n1464 & n1469 ) | ( ~n1464 & n1470 ) | ( n1469 & n1470 ) ;
  assign n1472 = n1464 | n1471 ;
  assign n1473 = n1472 ^ n1463 ^ 1'b0 ;
  assign n1474 = ( ~n1331 & n1463 ) | ( ~n1331 & n1473 ) | ( n1463 & n1473 ) ;
  assign n1475 = ( n1472 & ~n1473 ) | ( n1472 & n1474 ) | ( ~n1473 & n1474 ) ;
  assign n1476 = ( n1465 & n1466 ) | ( n1465 & ~n1468 ) | ( n1466 & ~n1468 ) ;
  assign n1477 = n1284 ^ n1283 ^ n1282 ;
  assign n1478 = ( n1475 & ~n1476 ) | ( n1475 & n1477 ) | ( ~n1476 & n1477 ) ;
  assign n1479 = ~n1285 & n1478 ;
  assign n1480 = ( ~n1249 & n1250 ) | ( ~n1249 & n1479 ) | ( n1250 & n1479 ) ;
  assign n1481 = n1249 | n1480 ;
  assign n1482 = n1481 ^ n1478 ^ 1'b0 ;
  assign n1483 = ( ~n1285 & n1478 ) | ( ~n1285 & n1482 ) | ( n1478 & n1482 ) ;
  assign n1484 = ( n1481 & ~n1482 ) | ( n1481 & n1483 ) | ( ~n1482 & n1483 ) ;
  assign n1485 = n1213 ^ n1211 ^ n1160 ;
  assign n1486 = ( ~n1247 & n1484 ) | ( ~n1247 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = n1156 ^ n1155 ^ n1153 ;
  assign n1488 = ( ~n1214 & n1486 ) | ( ~n1214 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1604 = ( n1131 & ~n1157 ) | ( n1131 & n1488 ) | ( ~n1157 & n1488 ) ;
  assign n1713 = ( n1601 & ~n1602 ) | ( n1601 & n1604 ) | ( ~n1602 & n1604 ) ;
  assign n1830 = ( n1710 & ~n1711 ) | ( n1710 & n1713 ) | ( ~n1711 & n1713 ) ;
  assign n1895 = ( n1827 & ~n1828 ) | ( n1827 & n1830 ) | ( ~n1828 & n1830 ) ;
  assign n2013 = ( n1892 & ~n1893 ) | ( n1892 & n1895 ) | ( ~n1893 & n1895 ) ;
  assign n2011 = ( n1875 & ~n1890 ) | ( n1875 & n1891 ) | ( ~n1890 & n1891 ) ;
  assign n2009 = ( n1864 & n1872 ) | ( n1864 & n1874 ) | ( n1872 & n1874 ) ;
  assign n2007 = ( n1879 & ~n1880 ) | ( n1879 & n1889 ) | ( ~n1880 & n1889 ) ;
  assign n1999 = n533 ^ n229 ^ 1'b0 ;
  assign n2000 = ( n533 & n534 ) | ( n533 & ~n1999 ) | ( n534 & ~n1999 ) ;
  assign n2001 = n2000 ^ n218 ^ 1'b0 ;
  assign n2002 = ( n218 & ~n531 ) | ( n218 & n2001 ) | ( ~n531 & n2001 ) ;
  assign n2003 = ( n2000 & ~n2001 ) | ( n2000 & n2002 ) | ( ~n2001 & n2002 ) ;
  assign n2004 = ( n218 & n554 ) | ( n218 & ~n2003 ) | ( n554 & ~n2003 ) ;
  assign n2005 = n2004 ^ n2003 ^ 1'b0 ;
  assign n2006 = ( n2003 & ~n2004 ) | ( n2003 & n2005 ) | ( ~n2004 & n2005 ) ;
  assign n1991 = n846 ^ n220 ^ 1'b0 ;
  assign n1992 = ( n845 & n846 ) | ( n845 & n1991 ) | ( n846 & n1991 ) ;
  assign n1993 = n1992 ^ n227 ^ 1'b0 ;
  assign n1994 = ( n227 & ~n843 ) | ( n227 & n1993 ) | ( ~n843 & n1993 ) ;
  assign n1995 = ( n1992 & ~n1993 ) | ( n1992 & n1994 ) | ( ~n1993 & n1994 ) ;
  assign n1996 = ( n227 & n852 ) | ( n227 & ~n1995 ) | ( n852 & ~n1995 ) ;
  assign n1997 = n1996 ^ n1995 ^ 1'b0 ;
  assign n1998 = ( n1995 & ~n1996 ) | ( n1995 & n1997 ) | ( ~n1996 & n1997 ) ;
  assign n2008 = n2007 ^ n2006 ^ n1998 ;
  assign n1989 = n224 & n840 ;
  assign n1990 = n1989 ^ n1880 ^ n654 ;
  assign n2010 = n2009 ^ n2008 ^ n1990 ;
  assign n2012 = n2011 ^ n2010 ^ 1'b0 ;
  assign n2014 = n2013 ^ n2012 ^ 1'b0 ;
  assign n261 = n164 | n179 ;
  assign n262 = n209 | n261 ;
  assign n264 = ( n134 & ~n262 ) | ( n134 & n263 ) | ( ~n262 & n263 ) ;
  assign n265 = n262 | n264 ;
  assign n269 = n94 | n268 ;
  assign n270 = n267 | n269 ;
  assign n271 = n265 | n270 ;
  assign n276 = ( ~n271 & n272 ) | ( ~n271 & n275 ) | ( n272 & n275 ) ;
  assign n277 = n271 | n276 ;
  assign n287 = n282 | n286 ;
  assign n289 = ( n78 & ~n287 ) | ( n78 & n288 ) | ( ~n287 & n288 ) ;
  assign n290 = n287 | n289 ;
  assign n291 = ( ~n277 & n281 ) | ( ~n277 & n290 ) | ( n281 & n290 ) ;
  assign n292 = n277 | n291 ;
  assign n294 = ( n113 & ~n292 ) | ( n113 & n293 ) | ( ~n292 & n293 ) ;
  assign n295 = n292 | n294 ;
  assign n297 = ( n163 & ~n295 ) | ( n163 & n296 ) | ( ~n295 & n296 ) ;
  assign n298 = n295 | n297 ;
  assign n318 = n73 | n317 ;
  assign n324 = n320 | n323 ;
  assign n326 = ( n188 & ~n324 ) | ( n188 & n325 ) | ( ~n324 & n325 ) ;
  assign n327 = n324 | n326 ;
  assign n329 = ( n146 & ~n327 ) | ( n146 & n328 ) | ( ~n327 & n328 ) ;
  assign n330 = n327 | n329 ;
  assign n332 = n144 | n331 ;
  assign n333 = ( ~n318 & n330 ) | ( ~n318 & n332 ) | ( n330 & n332 ) ;
  assign n334 = n318 | n333 ;
  assign n335 = ( n312 & n314 ) | ( n312 & ~n334 ) | ( n314 & ~n334 ) ;
  assign n336 = ~n312 & n335 ;
  assign n337 = ( n260 & ~n298 ) | ( n260 & n336 ) | ( ~n298 & n336 ) ;
  assign n338 = ~n260 & n337 ;
  assign n339 = ( n255 & ~n256 ) | ( n255 & n338 ) | ( ~n256 & n338 ) ;
  assign n340 = ~n255 & n339 ;
  assign n341 = ( n234 & ~n235 ) | ( n234 & n340 ) | ( ~n235 & n340 ) ;
  assign n342 = ~n234 & n341 ;
  assign n343 = ( n232 & ~n233 ) | ( n232 & n342 ) | ( ~n233 & n342 ) ;
  assign n344 = ~n232 & n343 ;
  assign n1158 = n1157 ^ n1131 ^ 1'b0 ;
  assign n1489 = n1488 ^ n1158 ^ 1'b0 ;
  assign n1490 = n269 | n350 ;
  assign n1491 = n600 | n716 ;
  assign n1492 = n735 | n1491 ;
  assign n1493 = ( n87 & n404 ) | ( n87 & ~n1492 ) | ( n404 & ~n1492 ) ;
  assign n1494 = n1492 | n1493 ;
  assign n1495 = ( n266 & n399 ) | ( n266 & ~n1494 ) | ( n399 & ~n1494 ) ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = ( n380 & ~n1490 ) | ( n380 & n1496 ) | ( ~n1490 & n1496 ) ;
  assign n1498 = n1490 | n1497 ;
  assign n1499 = n309 | n363 ;
  assign n1500 = n148 | n1499 ;
  assign n1501 = ( n253 & n284 ) | ( n253 & ~n1500 ) | ( n284 & ~n1500 ) ;
  assign n1502 = n1500 | n1501 ;
  assign n1503 = n133 | n1502 ;
  assign n1504 = n376 | n1503 ;
  assign n1505 = ( n113 & n161 ) | ( n113 & ~n1504 ) | ( n161 & ~n1504 ) ;
  assign n1506 = n1504 | n1505 ;
  assign n1507 = ( n92 & n274 ) | ( n92 & ~n1506 ) | ( n274 & ~n1506 ) ;
  assign n1508 = n1506 | n1507 ;
  assign n1509 = ( n141 & ~n1498 ) | ( n141 & n1508 ) | ( ~n1498 & n1508 ) ;
  assign n1510 = n1498 | n1509 ;
  assign n1511 = ( n315 & n405 ) | ( n315 & ~n1510 ) | ( n405 & ~n1510 ) ;
  assign n1512 = n1510 | n1511 ;
  assign n1513 = ( n250 & n484 ) | ( n250 & ~n1512 ) | ( n484 & ~n1512 ) ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = ( n157 & n328 ) | ( n157 & ~n1514 ) | ( n328 & ~n1514 ) ;
  assign n1516 = n1514 | n1515 ;
  assign n1517 = ( n178 & n283 ) | ( n178 & ~n1516 ) | ( n283 & ~n1516 ) ;
  assign n1518 = n1516 | n1517 ;
  assign n1519 = n1487 ^ n1486 ^ n1214 ;
  assign n1520 = n1247 & ~n1485 ;
  assign n1521 = ~n1247 & n1485 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = n1522 ^ n1484 ^ 1'b0 ;
  assign n1524 = n619 | n911 ;
  assign n1525 = ( n272 & n720 ) | ( n272 & ~n1524 ) | ( n720 & ~n1524 ) ;
  assign n1526 = n1524 | n1525 ;
  assign n1527 = n105 | n370 ;
  assign n1528 = n178 | n1527 ;
  assign n1529 = n466 | n1528 ;
  assign n1530 = ( n711 & n810 ) | ( n711 & ~n1529 ) | ( n810 & ~n1529 ) ;
  assign n1531 = n1529 | n1530 ;
  assign n1532 = ( n87 & n233 ) | ( n87 & ~n1531 ) | ( n233 & ~n1531 ) ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = ( n163 & n399 ) | ( n163 & ~n1533 ) | ( n399 & ~n1533 ) ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = ( n632 & ~n1526 ) | ( n632 & n1535 ) | ( ~n1526 & n1535 ) ;
  assign n1537 = n1526 | n1536 ;
  assign n1540 = n458 | n1539 ;
  assign n1541 = ( n492 & n908 ) | ( n492 & ~n1540 ) | ( n908 & ~n1540 ) ;
  assign n1542 = n1540 | n1541 ;
  assign n1543 = n319 | n406 ;
  assign n1544 = ( n208 & n379 ) | ( n208 & ~n1543 ) | ( n379 & ~n1543 ) ;
  assign n1545 = n1543 | n1544 ;
  assign n1546 = ( n674 & ~n1542 ) | ( n674 & n1545 ) | ( ~n1542 & n1545 ) ;
  assign n1547 = n1542 | n1546 ;
  assign n1548 = ( n92 & n604 ) | ( n92 & ~n1547 ) | ( n604 & ~n1547 ) ;
  assign n1549 = n1547 | n1548 ;
  assign n1550 = ( n187 & ~n1537 ) | ( n187 & n1549 ) | ( ~n1537 & n1549 ) ;
  assign n1551 = n1537 | n1550 ;
  assign n1552 = ( n293 & n484 ) | ( n293 & ~n1551 ) | ( n484 & ~n1551 ) ;
  assign n1553 = n1551 | n1552 ;
  assign n1554 = ( n164 & n515 ) | ( n164 & ~n1553 ) | ( n515 & ~n1553 ) ;
  assign n1555 = n1553 | n1554 ;
  assign n1556 = n1523 & ~n1555 ;
  assign n1557 = ( ~n1518 & n1519 ) | ( ~n1518 & n1556 ) | ( n1519 & n1556 ) ;
  assign n1558 = ( n344 & n1489 ) | ( n344 & n1557 ) | ( n1489 & n1557 ) ;
  assign n1603 = n1602 ^ n1601 ^ 1'b0 ;
  assign n1605 = n1604 ^ n1603 ^ 1'b0 ;
  assign n1606 = n330 | n438 ;
  assign n1607 = n1535 | n1606 ;
  assign n1608 = ( n645 & n674 ) | ( n645 & ~n1607 ) | ( n674 & ~n1607 ) ;
  assign n1609 = n1607 | n1608 ;
  assign n1610 = ( n241 & n258 ) | ( n241 & ~n1609 ) | ( n258 & ~n1609 ) ;
  assign n1611 = n1609 | n1610 ;
  assign n1612 = ( n137 & n349 ) | ( n137 & ~n1611 ) | ( n349 & ~n1611 ) ;
  assign n1613 = n1611 | n1612 ;
  assign n1614 = ( n125 & n462 ) | ( n125 & ~n1613 ) | ( n462 & ~n1613 ) ;
  assign n1615 = n1613 | n1614 ;
  assign n1616 = ( n131 & n564 ) | ( n131 & ~n1615 ) | ( n564 & ~n1615 ) ;
  assign n1617 = n1615 | n1616 ;
  assign n1618 = ( n94 & n213 ) | ( n94 & ~n1617 ) | ( n213 & ~n1617 ) ;
  assign n1619 = n1617 | n1618 ;
  assign n1673 = ( n1558 & n1605 ) | ( n1558 & ~n1619 ) | ( n1605 & ~n1619 ) ;
  assign n1712 = n1711 ^ n1710 ^ 1'b0 ;
  assign n1714 = n1713 ^ n1712 ^ 1'b0 ;
  assign n1715 = n237 | n309 ;
  assign n1716 = n187 | n1715 ;
  assign n1717 = ( n105 & n328 ) | ( n105 & ~n1716 ) | ( n328 & ~n1716 ) ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = ( n179 & n378 ) | ( n179 & ~n1718 ) | ( n378 & ~n1718 ) ;
  assign n1720 = n1718 | n1719 ;
  assign n1721 = n153 | n272 ;
  assign n1722 = n898 | n1721 ;
  assign n1723 = n487 | n1722 ;
  assign n1724 = ( n111 & n316 ) | ( n111 & ~n1723 ) | ( n316 & ~n1723 ) ;
  assign n1725 = n1723 | n1724 ;
  assign n1726 = ( n163 & n203 ) | ( n163 & ~n1725 ) | ( n203 & ~n1725 ) ;
  assign n1727 = n1725 | n1726 ;
  assign n1728 = n244 | n1727 ;
  assign n1729 = n580 | n1728 ;
  assign n1730 = n516 | n1729 ;
  assign n1731 = n174 | n268 ;
  assign n1732 = n131 | n1731 ;
  assign n1733 = n136 | n389 ;
  assign n1734 = n1732 | n1733 ;
  assign n1735 = n715 | n1734 ;
  assign n1736 = ( n199 & n394 ) | ( n199 & ~n1735 ) | ( n394 & ~n1735 ) ;
  assign n1737 = n1735 | n1736 ;
  assign n1738 = ( n322 & n384 ) | ( n322 & ~n1737 ) | ( n384 & ~n1737 ) ;
  assign n1739 = n1737 | n1738 ;
  assign n1740 = ( n364 & n423 ) | ( n364 & ~n1739 ) | ( n423 & ~n1739 ) ;
  assign n1741 = n1739 | n1740 ;
  assign n1742 = ( n604 & ~n1730 ) | ( n604 & n1741 ) | ( ~n1730 & n1741 ) ;
  assign n1743 = n1730 | n1742 ;
  assign n1744 = n1720 | n1743 ;
  assign n1745 = ( n299 & n367 ) | ( n299 & ~n1744 ) | ( n367 & ~n1744 ) ;
  assign n1746 = n1744 | n1745 ;
  assign n1747 = ( n169 & n451 ) | ( n169 & ~n1746 ) | ( n451 & ~n1746 ) ;
  assign n1748 = n1746 | n1747 ;
  assign n1749 = ( n130 & n296 ) | ( n130 & ~n1748 ) | ( n296 & ~n1748 ) ;
  assign n1750 = n1748 | n1749 ;
  assign n1794 = ( n1673 & n1714 ) | ( n1673 & ~n1750 ) | ( n1714 & ~n1750 ) ;
  assign n1829 = n1828 ^ n1827 ^ 1'b0 ;
  assign n1831 = n1830 ^ n1829 ^ 1'b0 ;
  assign n1832 = n203 | n236 ;
  assign n1833 = n384 ^ n232 ^ n118 ;
  assign n1834 = n390 | n1833 ;
  assign n1835 = n1832 | n1834 ;
  assign n1836 = ( n377 & n860 ) | ( n377 & ~n1835 ) | ( n860 & ~n1835 ) ;
  assign n1837 = n1835 | n1836 ;
  assign n1838 = ( n300 & n1496 ) | ( n300 & ~n1837 ) | ( n1496 & ~n1837 ) ;
  assign n1839 = n1837 | n1838 ;
  assign n1840 = ( n683 & n734 ) | ( n683 & ~n1839 ) | ( n734 & ~n1839 ) ;
  assign n1841 = n1839 | n1840 ;
  assign n1842 = ( n123 & n290 ) | ( n123 & ~n1841 ) | ( n290 & ~n1841 ) ;
  assign n1843 = n1841 | n1842 ;
  assign n1844 = ( n156 & n175 ) | ( n156 & ~n1843 ) | ( n175 & ~n1843 ) ;
  assign n1845 = n1843 | n1844 ;
  assign n1860 = ( n1794 & n1831 ) | ( n1794 & ~n1845 ) | ( n1831 & ~n1845 ) ;
  assign n1894 = n1893 ^ n1892 ^ 1'b0 ;
  assign n1896 = n1895 ^ n1894 ^ 1'b0 ;
  assign n1897 = n165 | n237 ;
  assign n1898 = n748 | n1897 ;
  assign n1899 = ( n151 & n361 ) | ( n151 & ~n1898 ) | ( n361 & ~n1898 ) ;
  assign n1900 = n1898 | n1899 ;
  assign n1901 = ( n161 & n315 ) | ( n161 & ~n1900 ) | ( n315 & ~n1900 ) ;
  assign n1902 = n1900 | n1901 ;
  assign n1903 = ( n130 & n273 ) | ( n130 & ~n1902 ) | ( n273 & ~n1902 ) ;
  assign n1904 = n1902 | n1903 ;
  assign n1905 = n118 | n729 ;
  assign n1906 = n399 | n1905 ;
  assign n1907 = n156 | n258 ;
  assign n1908 = n203 | n1907 ;
  assign n1909 = ( n266 & n426 ) | ( n266 & ~n1908 ) | ( n426 & ~n1908 ) ;
  assign n1910 = n1908 | n1909 ;
  assign n1911 = n1906 | n1910 ;
  assign n1912 = n1904 | n1911 ;
  assign n1913 = n122 | n236 ;
  assign n1914 = ( n157 & n414 ) | ( n157 & ~n1913 ) | ( n414 & ~n1913 ) ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = ( n283 & n462 ) | ( n283 & ~n1915 ) | ( n462 & ~n1915 ) ;
  assign n1917 = n1915 | n1916 ;
  assign n1918 = ( n142 & n475 ) | ( n142 & ~n1917 ) | ( n475 & ~n1917 ) ;
  assign n1919 = n1917 | n1918 ;
  assign n1920 = ( n256 & ~n1912 ) | ( n256 & n1919 ) | ( ~n1912 & n1919 ) ;
  assign n1921 = n1912 | n1920 ;
  assign n1922 = ( n194 & n389 ) | ( n194 & ~n1921 ) | ( n389 & ~n1921 ) ;
  assign n1923 = n1921 | n1922 ;
  assign n1924 = ( n188 & n349 ) | ( n188 & ~n1923 ) | ( n349 & ~n1923 ) ;
  assign n1925 = n1923 | n1924 ;
  assign n1926 = ( n178 & n517 ) | ( n178 & ~n1925 ) | ( n517 & ~n1925 ) ;
  assign n1927 = n1925 | n1926 ;
  assign n2015 = ( n1860 & n1896 ) | ( n1860 & ~n1927 ) | ( n1896 & ~n1927 ) ;
  assign n2016 = ( n1988 & n2014 ) | ( n1988 & n2015 ) | ( n2014 & n2015 ) ;
  assign n2017 = n493 | n1528 ;
  assign n2018 = n1951 | n2017 ;
  assign n2019 = ( n244 & n457 ) | ( n244 & ~n2018 ) | ( n457 & ~n2018 ) ;
  assign n2020 = n2018 | n2019 ;
  assign n2021 = n200 | n711 ;
  assign n2022 = ( n240 & n273 ) | ( n240 & ~n2021 ) | ( n273 & ~n2021 ) ;
  assign n2023 = n2021 | n2022 ;
  assign n2024 = ( n232 & n263 ) | ( n232 & ~n2023 ) | ( n263 & ~n2023 ) ;
  assign n2025 = n2023 | n2024 ;
  assign n2026 = n408 | n444 ;
  assign n2027 = n2025 | n2026 ;
  assign n2028 = ( n122 & n187 ) | ( n122 & ~n2027 ) | ( n187 & ~n2027 ) ;
  assign n2029 = n2027 | n2028 ;
  assign n2030 = ( n78 & n157 ) | ( n78 & ~n2029 ) | ( n157 & ~n2029 ) ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = ( n361 & ~n2020 ) | ( n361 & n2031 ) | ( ~n2020 & n2031 ) ;
  assign n2033 = n2020 | n2032 ;
  assign n2034 = ( n303 & n1974 ) | ( n303 & ~n2033 ) | ( n1974 & ~n2033 ) ;
  assign n2035 = n2033 | n2034 ;
  assign n2036 = ( n125 & n131 ) | ( n125 & ~n2035 ) | ( n131 & ~n2035 ) ;
  assign n2037 = n2035 | n2036 ;
  assign n2056 = ( ~n1990 & n2008 ) | ( ~n1990 & n2009 ) | ( n2008 & n2009 ) ;
  assign n2054 = ( ~n654 & n1880 ) | ( ~n654 & n1989 ) | ( n1880 & n1989 ) ;
  assign n2053 = ( n1998 & n2006 ) | ( n1998 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2044 = n846 ^ n227 ^ 1'b0 ;
  assign n2045 = ( n845 & n846 ) | ( n845 & n2044 ) | ( n846 & n2044 ) ;
  assign n2046 = n2045 ^ n229 ^ 1'b0 ;
  assign n2047 = ( n229 & ~n843 ) | ( n229 & n2046 ) | ( ~n843 & n2046 ) ;
  assign n2048 = ( n2045 & ~n2046 ) | ( n2045 & n2047 ) | ( ~n2046 & n2047 ) ;
  assign n2049 = ( n229 & n852 ) | ( n229 & ~n2048 ) | ( n852 & ~n2048 ) ;
  assign n2050 = n2049 ^ n2048 ^ 1'b0 ;
  assign n2051 = ( n2048 & ~n2049 ) | ( n2048 & n2050 ) | ( ~n2049 & n2050 ) ;
  assign n2043 = n220 & n840 ;
  assign n2039 = n218 | n530 ;
  assign n2040 = n218 & ~n533 ;
  assign n2041 = ( n531 & n2039 ) | ( n531 & ~n2040 ) | ( n2039 & ~n2040 ) ;
  assign n2042 = ~n531 & n2041 ;
  assign n2052 = n2051 ^ n2043 ^ n2042 ;
  assign n2055 = n2054 ^ n2053 ^ n2052 ;
  assign n2057 = n2056 ^ n2055 ^ 1'b0 ;
  assign n2038 = ( n2010 & ~n2011 ) | ( n2010 & n2013 ) | ( ~n2011 & n2013 ) ;
  assign n2058 = n2057 ^ n2038 ^ 1'b0 ;
  assign n2155 = ( n2016 & ~n2037 ) | ( n2016 & n2058 ) | ( ~n2037 & n2058 ) ;
  assign n2170 = ( n2038 & n2055 ) | ( n2038 & ~n2056 ) | ( n2055 & ~n2056 ) ;
  assign n2168 = ( ~n2052 & n2053 ) | ( ~n2052 & n2054 ) | ( n2053 & n2054 ) ;
  assign n2159 = n845 ^ n229 ^ 1'b0 ;
  assign n2160 = ( n845 & n846 ) | ( n845 & ~n2159 ) | ( n846 & ~n2159 ) ;
  assign n2161 = n2160 ^ n218 ^ 1'b0 ;
  assign n2162 = ( n218 & ~n843 ) | ( n218 & n2161 ) | ( ~n843 & n2161 ) ;
  assign n2163 = ( n2160 & ~n2161 ) | ( n2160 & n2162 ) | ( ~n2161 & n2162 ) ;
  assign n2164 = ( n218 & n852 ) | ( n218 & ~n2163 ) | ( n852 & ~n2163 ) ;
  assign n2165 = n2164 ^ n2163 ^ 1'b0 ;
  assign n2166 = ( n2163 & ~n2164 ) | ( n2163 & n2165 ) | ( ~n2164 & n2165 ) ;
  assign n2158 = ( n2042 & ~n2043 ) | ( n2042 & n2051 ) | ( ~n2043 & n2051 ) ;
  assign n2156 = n227 & n840 ;
  assign n2157 = n2156 ^ n2043 ^ n530 ;
  assign n2167 = n2166 ^ n2158 ^ n2157 ;
  assign n2169 = n2168 ^ n2167 ^ 1'b0 ;
  assign n2171 = n2170 ^ n2169 ^ 1'b0 ;
  assign n2172 = n239 | n575 ;
  assign n2173 = ( n306 & n380 ) | ( n306 & ~n2172 ) | ( n380 & ~n2172 ) ;
  assign n2174 = n2172 | n2173 ;
  assign n2175 = ( n362 & n632 ) | ( n362 & ~n2174 ) | ( n632 & ~n2174 ) ;
  assign n2176 = n2174 | n2175 ;
  assign n2177 = ( n418 & n697 ) | ( n418 & ~n2176 ) | ( n697 & ~n2176 ) ;
  assign n2178 = n2176 | n2177 ;
  assign n2179 = ( n161 & n920 ) | ( n161 & ~n2178 ) | ( n920 & ~n2178 ) ;
  assign n2180 = n2178 | n2179 ;
  assign n2181 = ( n208 & n293 ) | ( n208 & ~n2180 ) | ( n293 & ~n2180 ) ;
  assign n2182 = n2180 | n2181 ;
  assign n2183 = ( n136 & n475 ) | ( n136 & ~n2182 ) | ( n475 & ~n2182 ) ;
  assign n2184 = n2182 | n2183 ;
  assign n2204 = ( n2155 & n2171 ) | ( n2155 & ~n2184 ) | ( n2171 & ~n2184 ) ;
  assign n2205 = n242 | n558 ;
  assign n2206 = ( n615 & n799 ) | ( n615 & ~n2205 ) | ( n799 & ~n2205 ) ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = n1949 | n2207 ;
  assign n2209 = n200 | n322 ;
  assign n2210 = n293 | n2209 ;
  assign n2211 = ( n213 & n399 ) | ( n213 & ~n2210 ) | ( n399 & ~n2210 ) ;
  assign n2212 = n2210 | n2211 ;
  assign n2213 = n601 | n2212 ;
  assign n2214 = n137 | n2213 ;
  assign n2215 = ( n445 & n451 ) | ( n445 & ~n2214 ) | ( n451 & ~n2214 ) ;
  assign n2216 = n2214 | n2215 ;
  assign n2217 = ( n515 & n559 ) | ( n515 & ~n2216 ) | ( n559 & ~n2216 ) ;
  assign n2218 = n2216 | n2217 ;
  assign n2219 = ( n78 & n437 ) | ( n78 & ~n2218 ) | ( n437 & ~n2218 ) ;
  assign n2220 = n2218 | n2219 ;
  assign n2221 = ( n1549 & ~n2208 ) | ( n1549 & n2220 ) | ( ~n2208 & n2220 ) ;
  assign n2222 = n2208 | n2221 ;
  assign n2223 = ( n349 & n1967 ) | ( n349 & ~n2222 ) | ( n1967 & ~n2222 ) ;
  assign n2224 = n2222 | n2223 ;
  assign n2225 = ( n256 & n258 ) | ( n256 & ~n2224 ) | ( n258 & ~n2224 ) ;
  assign n2226 = n2224 | n2225 ;
  assign n2227 = ( n144 & n321 ) | ( n144 & ~n2226 ) | ( n321 & ~n2226 ) ;
  assign n2228 = n2226 | n2227 ;
  assign n2229 = ( n146 & n182 ) | ( n146 & ~n2228 ) | ( n182 & ~n2228 ) ;
  assign n2230 = n2228 | n2229 ;
  assign n2240 = ( n2167 & ~n2168 ) | ( n2167 & n2170 ) | ( ~n2168 & n2170 ) ;
  assign n2237 = ( ~n530 & n2043 ) | ( ~n530 & n2156 ) | ( n2043 & n2156 ) ;
  assign n2236 = n229 & n840 ;
  assign n2232 = n218 & ~n845 ;
  assign n2233 = n218 & ~n798 ;
  assign n2234 = ( n842 & ~n2232 ) | ( n842 & n2233 ) | ( ~n2232 & n2233 ) ;
  assign n2235 = ~n2232 & n2234 ;
  assign n2238 = n2237 ^ n2236 ^ n2235 ;
  assign n2231 = ( ~n2157 & n2158 ) | ( ~n2157 & n2166 ) | ( n2158 & n2166 ) ;
  assign n2239 = n2238 ^ n2231 ^ 1'b0 ;
  assign n2241 = n2240 ^ n2239 ^ 1'b0 ;
  assign n2245 = ( n2204 & ~n2230 ) | ( n2204 & n2241 ) | ( ~n2230 & n2241 ) ;
  assign n230 = n229 ^ n218 ^ 1'b0 ;
  assign n2248 = n841 ^ n230 ^ 1'b0 ;
  assign n2249 = n840 & ~n2248 ;
  assign n2247 = ( n2235 & ~n2236 ) | ( n2235 & n2237 ) | ( ~n2236 & n2237 ) ;
  assign n2246 = ( ~n2231 & n2238 ) | ( ~n2231 & n2240 ) | ( n2238 & n2240 ) ;
  assign n2250 = n2249 ^ n2247 ^ n2246 ;
  assign n2251 = n510 | n1729 ;
  assign n2252 = n235 | n564 ;
  assign n2253 = n102 | n288 ;
  assign n2254 = ( ~n2251 & n2252 ) | ( ~n2251 & n2253 ) | ( n2252 & n2253 ) ;
  assign n2255 = n2251 | n2254 ;
  assign n2256 = n315 | n394 ;
  assign n2257 = n158 | n2256 ;
  assign n2258 = ( n125 & n209 ) | ( n125 & ~n2257 ) | ( n209 & ~n2257 ) ;
  assign n2259 = n2257 | n2258 ;
  assign n2260 = ( n377 & ~n2255 ) | ( n377 & n2259 ) | ( ~n2255 & n2259 ) ;
  assign n2261 = n2255 | n2260 ;
  assign n2262 = n199 | n1962 ;
  assign n2263 = n475 | n2262 ;
  assign n2264 = ( n399 & ~n2261 ) | ( n399 & n2263 ) | ( ~n2261 & n2263 ) ;
  assign n2265 = n2261 | n2264 ;
  assign n2266 = ( n157 & n313 ) | ( n157 & ~n2265 ) | ( n313 & ~n2265 ) ;
  assign n2267 = ~n157 & n2266 ;
  assign n2268 = ( ~n312 & n928 ) | ( ~n312 & n2267 ) | ( n928 & n2267 ) ;
  assign n2269 = ~n928 & n2268 ;
  assign n2270 = ( n250 & ~n405 ) | ( n250 & n2269 ) | ( ~n405 & n2269 ) ;
  assign n2271 = ~n250 & n2270 ;
  assign n2389 = ( n2245 & n2250 ) | ( n2245 & n2271 ) | ( n2250 & n2271 ) ;
  assign n2390 = n493 | n908 ;
  assign n2391 = ( n983 & n1496 ) | ( n983 & ~n2390 ) | ( n1496 & ~n2390 ) ;
  assign n2392 = n2390 | n2391 ;
  assign n2393 = n194 | n576 ;
  assign n2394 = ( n122 & n394 ) | ( n122 & ~n2393 ) | ( n394 & ~n2393 ) ;
  assign n2395 = n2393 | n2394 ;
  assign n2396 = ( n150 & n316 ) | ( n150 & ~n2395 ) | ( n316 & ~n2395 ) ;
  assign n2397 = n2395 | n2396 ;
  assign n2398 = ( n356 & ~n2392 ) | ( n356 & n2397 ) | ( ~n2392 & n2397 ) ;
  assign n2399 = n2392 | n2398 ;
  assign n2400 = ( n68 & n241 ) | ( n68 & ~n2399 ) | ( n241 & ~n2399 ) ;
  assign n2401 = n2399 | n2400 ;
  assign n2402 = ( n274 & n749 ) | ( n274 & ~n2401 ) | ( n749 & ~n2401 ) ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = ( n131 & n163 ) | ( n131 & ~n2403 ) | ( n163 & ~n2403 ) ;
  assign n2405 = n2403 | n2404 ;
  assign n2424 = n2389 & ~n2405 ;
  assign n2425 = n637 | n1732 ;
  assign n2426 = ( n244 & n610 ) | ( n244 & ~n2425 ) | ( n610 & ~n2425 ) ;
  assign n2427 = n2425 | n2426 ;
  assign n2428 = n305 | n405 ;
  assign n2429 = n559 | n2428 ;
  assign n2430 = n484 ^ n389 ^ n367 ;
  assign n2431 = ( n423 & n515 ) | ( n423 & ~n2430 ) | ( n515 & ~n2430 ) ;
  assign n2432 = n2430 | n2431 ;
  assign n2433 = n160 | n558 ;
  assign n2434 = n399 | n2433 ;
  assign n2435 = n2432 | n2434 ;
  assign n2436 = n1968 | n2435 ;
  assign n2437 = ( n137 & n319 ) | ( n137 & ~n2436 ) | ( n319 & ~n2436 ) ;
  assign n2438 = n2436 | n2437 ;
  assign n2439 = ( n148 & n282 ) | ( n148 & ~n2438 ) | ( n282 & ~n2438 ) ;
  assign n2440 = n2438 | n2439 ;
  assign n2441 = ( n209 & n273 ) | ( n209 & ~n2440 ) | ( n273 & ~n2440 ) ;
  assign n2442 = n2440 | n2441 ;
  assign n2443 = ( n87 & n293 ) | ( n87 & ~n2442 ) | ( n293 & ~n2442 ) ;
  assign n2444 = n2442 | n2443 ;
  assign n2445 = ( n118 & n213 ) | ( n118 & ~n2444 ) | ( n213 & ~n2444 ) ;
  assign n2446 = n2444 | n2445 ;
  assign n2447 = ( ~n2427 & n2429 ) | ( ~n2427 & n2446 ) | ( n2429 & n2446 ) ;
  assign n2448 = n2427 | n2447 ;
  assign n2449 = ( n102 & n363 ) | ( n102 & ~n2448 ) | ( n363 & ~n2448 ) ;
  assign n2450 = n2448 | n2449 ;
  assign n2451 = ( n122 & n168 ) | ( n122 & ~n2450 ) | ( n168 & ~n2450 ) ;
  assign n2452 = n2450 | n2451 ;
  assign n2453 = ( n107 & n205 ) | ( n107 & ~n2452 ) | ( n205 & ~n2452 ) ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = ( n134 & n284 ) | ( n134 & ~n2454 ) | ( n284 & ~n2454 ) ;
  assign n2456 = n2454 | n2455 ;
  assign n2462 = n2424 & ~n2456 ;
  assign n2463 = n313 & ~n561 ;
  assign n2464 = ~n500 & n2463 ;
  assign n2465 = ( n828 & ~n2025 ) | ( n828 & n2464 ) | ( ~n2025 & n2464 ) ;
  assign n2466 = ~n828 & n2465 ;
  assign n2467 = ( ~n261 & n290 ) | ( ~n261 & n2466 ) | ( n290 & n2466 ) ;
  assign n2468 = ~n290 & n2467 ;
  assign n2469 = ( n144 & ~n668 ) | ( n144 & n2468 ) | ( ~n668 & n2468 ) ;
  assign n2470 = ~n144 & n2469 ;
  assign n2471 = ( ~n208 & n310 ) | ( ~n208 & n2470 ) | ( n310 & n2470 ) ;
  assign n2472 = ~n310 & n2471 ;
  assign n2473 = ( n136 & ~n564 ) | ( n136 & n2472 ) | ( ~n564 & n2472 ) ;
  assign n2474 = ~n136 & n2473 ;
  assign n2684 = n2462 & n2474 ;
  assign n2696 = n2695 ^ n2684 ^ 1'b0 ;
  assign n2697 = n2422 & n2696 ;
  assign n2423 = ~x0 & n2420 ;
  assign n2475 = n2474 ^ n2462 ^ 1'b0 ;
  assign n2698 = n2423 & ~n2475 ;
  assign n2457 = n2456 ^ n2424 ^ 1'b0 ;
  assign n2459 = ~n25 & n2421 ;
  assign n2699 = n2457 & n2459 ;
  assign n2700 = ( ~n2697 & n2698 ) | ( ~n2697 & n2699 ) | ( n2698 & n2699 ) ;
  assign n2701 = n2697 | n2700 ;
  assign n2478 = x0 & n2421 ;
  assign n2406 = n2405 ^ n2389 ^ 1'b0 ;
  assign n2272 = n2271 ^ n2250 ^ n2245 ;
  assign n2242 = n2241 ^ n2230 ^ n2204 ;
  assign n2185 = n2184 ^ n2171 ^ n2155 ;
  assign n2059 = n2058 ^ n2037 ^ n2016 ;
  assign n2060 = n2015 ^ n2014 ^ n1988 ;
  assign n1928 = n1927 ^ n1896 ^ n1860 ;
  assign n1846 = n1845 ^ n1831 ^ n1794 ;
  assign n1751 = n1750 ^ n1714 ^ n1673 ;
  assign n1620 = n1619 ^ n1605 ^ n1558 ;
  assign n1622 = n1557 ^ n1489 ^ n344 ;
  assign n1621 = n1556 ^ n1519 ^ n1518 ;
  assign n1623 = n1555 ^ n1523 ^ 1'b0 ;
  assign n1624 = n1622 & ~n1623 ;
  assign n1625 = n1621 & ~n1624 ;
  assign n1759 = ( n1620 & ~n1622 ) | ( n1620 & n1625 ) | ( ~n1622 & n1625 ) ;
  assign n1853 = ( n1620 & n1751 ) | ( n1620 & n1759 ) | ( n1751 & n1759 ) ;
  assign n1935 = ( n1751 & n1846 ) | ( n1751 & n1853 ) | ( n1846 & n1853 ) ;
  assign n2061 = ( n1846 & n1928 ) | ( n1846 & n1935 ) | ( n1928 & n1935 ) ;
  assign n2062 = ( n1928 & ~n2060 ) | ( n1928 & n2061 ) | ( ~n2060 & n2061 ) ;
  assign n2154 = ( n2059 & ~n2060 ) | ( n2059 & n2062 ) | ( ~n2060 & n2062 ) ;
  assign n2277 = ( n2059 & n2154 ) | ( n2059 & n2185 ) | ( n2154 & n2185 ) ;
  assign n2278 = ( n2185 & n2242 ) | ( n2185 & n2277 ) | ( n2242 & n2277 ) ;
  assign n2412 = ( n2242 & ~n2272 ) | ( n2242 & n2278 ) | ( ~n2272 & n2278 ) ;
  assign n2479 = ( ~n2272 & n2406 ) | ( ~n2272 & n2412 ) | ( n2406 & n2412 ) ;
  assign n2480 = ( n2406 & n2457 ) | ( n2406 & n2479 ) | ( n2457 & n2479 ) ;
  assign n2702 = ( n2457 & ~n2475 ) | ( n2457 & n2480 ) | ( ~n2475 & n2480 ) ;
  assign n2703 = n2702 ^ n2696 ^ n2475 ;
  assign n2704 = ( n2478 & n2701 ) | ( n2478 & ~n2703 ) | ( n2701 & ~n2703 ) ;
  assign n2705 = n2703 ^ n2701 ^ 1'b0 ;
  assign n2706 = ( n2701 & n2704 ) | ( n2701 & ~n2705 ) | ( n2704 & ~n2705 ) ;
  assign n2707 = n2706 ^ n539 ^ n537 ;
  assign n2458 = n2423 & n2457 ;
  assign n2460 = n2406 & n2459 ;
  assign n2461 = n2458 | n2460 ;
  assign n2476 = ~n2461 & n2475 ;
  assign n2477 = ( n2422 & n2461 ) | ( n2422 & ~n2476 ) | ( n2461 & ~n2476 ) ;
  assign n2481 = n2480 ^ n2475 ^ n2457 ;
  assign n2482 = ( n2477 & n2478 ) | ( n2477 & ~n2481 ) | ( n2478 & ~n2481 ) ;
  assign n2483 = n2481 ^ n2477 ^ 1'b0 ;
  assign n2484 = ( n2477 & n2482 ) | ( n2477 & ~n2483 ) | ( n2482 & ~n2483 ) ;
  assign n2485 = n2484 ^ n539 ^ n537 ;
  assign n2486 = n2422 & n2457 ;
  assign n2487 = n2406 & n2423 ;
  assign n2488 = ~n2272 & n2459 ;
  assign n2489 = ( ~n2486 & n2487 ) | ( ~n2486 & n2488 ) | ( n2487 & n2488 ) ;
  assign n2490 = n2486 | n2489 ;
  assign n2491 = n2490 ^ n2478 ^ 1'b0 ;
  assign n2492 = n2479 ^ n2457 ^ n2406 ;
  assign n2493 = ( n2478 & ~n2491 ) | ( n2478 & n2492 ) | ( ~n2491 & n2492 ) ;
  assign n2494 = ( n2490 & n2491 ) | ( n2490 & n2493 ) | ( n2491 & n2493 ) ;
  assign n2495 = n2494 ^ n539 ^ n537 ;
  assign n2197 = n1040 ^ n541 ^ 1'b0 ;
  assign n2275 = n1038 & n2197 ;
  assign n2198 = n1038 & ~n2197 ;
  assign n2294 = n2185 & n2198 ;
  assign n2199 = n1040 ^ n856 ^ 1'b0 ;
  assign n2200 = ~n1038 & n2197 ;
  assign n2201 = ~n2199 & n2200 ;
  assign n2295 = ~n2060 & n2201 ;
  assign n2203 = ~n1038 & n2199 ;
  assign n2296 = n2059 & n2203 ;
  assign n2297 = ( ~n2294 & n2295 ) | ( ~n2294 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = n2294 | n2297 ;
  assign n2186 = n2185 ^ n2154 ^ n2059 ;
  assign n2299 = n2298 ^ n2275 ^ 1'b0 ;
  assign n2300 = ( n2186 & ~n2275 ) | ( n2186 & n2299 ) | ( ~n2275 & n2299 ) ;
  assign n2301 = ( n2275 & n2298 ) | ( n2275 & n2300 ) | ( n2298 & n2300 ) ;
  assign n2302 = n2301 ^ n536 ^ x5 ;
  assign n2303 = n2059 & n2198 ;
  assign n2304 = n1928 & n2201 ;
  assign n2305 = ~n2060 & n2203 ;
  assign n2306 = ( ~n2303 & n2304 ) | ( ~n2303 & n2305 ) | ( n2304 & n2305 ) ;
  assign n2307 = n2303 | n2306 ;
  assign n2063 = n2062 ^ n2060 ^ n2059 ;
  assign n2308 = n2063 & ~n2307 ;
  assign n2309 = ( n2275 & n2307 ) | ( n2275 & ~n2308 ) | ( n2307 & ~n2308 ) ;
  assign n2310 = n2309 ^ n536 ^ x5 ;
  assign n2311 = n1846 & n2201 ;
  assign n2312 = n1928 & n2203 ;
  assign n2313 = n2311 | n2312 ;
  assign n2314 = n2060 & ~n2313 ;
  assign n2315 = ( n2198 & n2313 ) | ( n2198 & ~n2314 ) | ( n2313 & ~n2314 ) ;
  assign n2077 = n2061 ^ n2060 ^ n1928 ;
  assign n2316 = n2077 & ~n2315 ;
  assign n2317 = ( n2275 & n2315 ) | ( n2275 & ~n2316 ) | ( n2315 & ~n2316 ) ;
  assign n2318 = n2317 ^ n536 ^ x5 ;
  assign n2319 = n1928 & n2198 ;
  assign n2320 = n1751 & n2201 ;
  assign n2321 = n1846 & n2203 ;
  assign n2322 = ( ~n2319 & n2320 ) | ( ~n2319 & n2321 ) | ( n2320 & n2321 ) ;
  assign n2323 = n2319 | n2322 ;
  assign n1936 = n1935 ^ n1928 ^ n1846 ;
  assign n2324 = n2323 ^ n2275 ^ 1'b0 ;
  assign n2325 = ( n1936 & ~n2275 ) | ( n1936 & n2324 ) | ( ~n2275 & n2324 ) ;
  assign n2326 = ( n2275 & n2323 ) | ( n2275 & n2325 ) | ( n2323 & n2325 ) ;
  assign n2327 = n2326 ^ n536 ^ x5 ;
  assign n2328 = n1846 & n2198 ;
  assign n2329 = n1620 & n2201 ;
  assign n2330 = n1751 & n2203 ;
  assign n2331 = ( ~n2328 & n2329 ) | ( ~n2328 & n2330 ) | ( n2329 & n2330 ) ;
  assign n2332 = n2328 | n2331 ;
  assign n1854 = n1853 ^ n1846 ^ n1751 ;
  assign n2333 = n2332 ^ n2275 ^ 1'b0 ;
  assign n2334 = ( n1854 & ~n2275 ) | ( n1854 & n2333 ) | ( ~n2275 & n2333 ) ;
  assign n2335 = ( n2275 & n2332 ) | ( n2275 & n2334 ) | ( n2332 & n2334 ) ;
  assign n2336 = n2335 ^ n536 ^ x5 ;
  assign n1653 = n1621 & ~n1623 ;
  assign n1654 = n1653 ^ n1622 ^ 1'b0 ;
  assign n1941 = n548 ^ n545 ^ 1'b0 ;
  assign n1942 = n544 ^ n541 ^ 1'b0 ;
  assign n1943 = n1941 & n1942 ;
  assign n2126 = ~n1654 & n1943 ;
  assign n2127 = n2126 ^ n548 ^ 1'b0 ;
  assign n2066 = ~n1941 & n1942 ;
  assign n2128 = ~n1622 & n2066 ;
  assign n2068 = n546 & ~n1942 ;
  assign n2129 = n1621 & n2068 ;
  assign n2070 = n1941 & ~n1942 ;
  assign n2071 = ~n546 & n2070 ;
  assign n2130 = n1623 & n2071 ;
  assign n2131 = ( ~n2128 & n2129 ) | ( ~n2128 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2132 = n2128 | n2131 ;
  assign n2133 = n2132 ^ n548 ^ 1'b0 ;
  assign n2134 = ( ~n548 & n2127 ) | ( ~n548 & n2133 ) | ( n2127 & n2133 ) ;
  assign n1644 = n1623 ^ n1621 ^ 1'b0 ;
  assign n2116 = n1644 & n1943 ;
  assign n2117 = n2116 ^ n548 ^ 1'b0 ;
  assign n2118 = n1623 & n2068 ;
  assign n2119 = n1621 & n2066 ;
  assign n2120 = n2118 | n2119 ;
  assign n2121 = n2120 ^ n548 ^ 1'b0 ;
  assign n2122 = ( ~n548 & n2117 ) | ( ~n548 & n2121 ) | ( n2117 & n2121 ) ;
  assign n2123 = n1623 & n1942 ;
  assign n2124 = n548 & ~n2123 ;
  assign n2125 = n2122 & n2124 ;
  assign n2337 = n2134 ^ n2125 ^ 1'b0 ;
  assign n2338 = n2124 ^ n2122 ^ 1'b0 ;
  assign n2339 = n1620 & n2203 ;
  assign n2340 = n1751 & n2198 ;
  assign n2341 = n2339 | n2340 ;
  assign n2342 = n1622 & ~n2341 ;
  assign n2343 = ( n2201 & n2341 ) | ( n2201 & ~n2342 ) | ( n2341 & ~n2342 ) ;
  assign n1760 = n1759 ^ n1751 ^ n1620 ;
  assign n2344 = n2343 ^ n2275 ^ 1'b0 ;
  assign n2345 = ( n1760 & ~n2275 ) | ( n1760 & n2344 ) | ( ~n2275 & n2344 ) ;
  assign n2346 = ( n2275 & n2343 ) | ( n2275 & n2345 ) | ( n2343 & n2345 ) ;
  assign n2347 = n2346 ^ n536 ^ x5 ;
  assign n2348 = n1038 & n1623 ;
  assign n2349 = n541 & ~n2348 ;
  assign n2350 = n1644 & n2275 ;
  assign n2351 = n1623 & n2203 ;
  assign n2352 = n1621 & n2198 ;
  assign n2353 = ( ~n2350 & n2351 ) | ( ~n2350 & n2352 ) | ( n2351 & n2352 ) ;
  assign n2354 = n2350 | n2353 ;
  assign n2355 = n2354 ^ n536 ^ x5 ;
  assign n2356 = n2349 & n2355 ;
  assign n2357 = n1623 & n2201 ;
  assign n2358 = n1621 & n2203 ;
  assign n2359 = n2357 | n2358 ;
  assign n2360 = n1622 & ~n2359 ;
  assign n2361 = ( n2198 & n2359 ) | ( n2198 & ~n2360 ) | ( n2359 & ~n2360 ) ;
  assign n2362 = n1654 & ~n2361 ;
  assign n2363 = ( n2275 & n2361 ) | ( n2275 & ~n2362 ) | ( n2361 & ~n2362 ) ;
  assign n2364 = n2363 ^ n536 ^ x5 ;
  assign n2365 = n2356 & n2364 ;
  assign n2366 = n1621 & n2201 ;
  assign n2367 = n1620 & n2198 ;
  assign n2368 = n2366 | n2367 ;
  assign n2369 = n1622 & ~n2368 ;
  assign n2370 = ( n2203 & n2368 ) | ( n2203 & ~n2369 ) | ( n2368 & ~n2369 ) ;
  assign n1626 = n1625 ^ n1622 ^ n1620 ;
  assign n2371 = n1626 & ~n2370 ;
  assign n2372 = ( n2275 & n2370 ) | ( n2275 & ~n2371 ) | ( n2370 & ~n2371 ) ;
  assign n2373 = n2372 ^ n536 ^ x5 ;
  assign n2374 = ( n2123 & n2365 ) | ( n2123 & n2373 ) | ( n2365 & n2373 ) ;
  assign n2375 = ( n2338 & n2347 ) | ( n2338 & n2374 ) | ( n2347 & n2374 ) ;
  assign n2376 = ( n2336 & n2337 ) | ( n2336 & n2375 ) | ( n2337 & n2375 ) ;
  assign n2136 = ~n1626 & n1943 ;
  assign n2137 = n2136 ^ n548 ^ 1'b0 ;
  assign n2138 = ~n1622 & n2068 ;
  assign n2139 = n1621 & n2071 ;
  assign n2140 = n1620 & n2066 ;
  assign n2141 = ( ~n2138 & n2139 ) | ( ~n2138 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = n2138 | n2141 ;
  assign n2143 = n2142 ^ n548 ^ 1'b0 ;
  assign n2144 = ( ~n548 & n2137 ) | ( ~n548 & n2143 ) | ( n2137 & n2143 ) ;
  assign n2135 = n2125 & n2134 ;
  assign n1668 = n548 ^ n222 ^ 1'b0 ;
  assign n1764 = n1623 & n1668 ;
  assign n2377 = n2144 ^ n2135 ^ n1764 ;
  assign n2378 = ( n2327 & n2376 ) | ( n2327 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2145 = ( n1764 & n2135 ) | ( n1764 & n2144 ) | ( n2135 & n2144 ) ;
  assign n2107 = n1760 & n1943 ;
  assign n2108 = n2107 ^ n548 ^ 1'b0 ;
  assign n2109 = ~n1622 & n2071 ;
  assign n2110 = n1620 & n2068 ;
  assign n2111 = n1751 & n2066 ;
  assign n2112 = ( ~n2109 & n2110 ) | ( ~n2109 & n2111 ) | ( n2110 & n2111 ) ;
  assign n2113 = n2109 | n2112 ;
  assign n2114 = n2113 ^ n548 ^ 1'b0 ;
  assign n2115 = ( ~n548 & n2108 ) | ( ~n548 & n2114 ) | ( n2108 & n2114 ) ;
  assign n1757 = n225 & n1668 ;
  assign n1766 = n1644 & n1757 ;
  assign n1672 = ~n225 & n1668 ;
  assign n1767 = n1621 & n1672 ;
  assign n1667 = n224 ^ n222 ^ 1'b0 ;
  assign n1753 = n1667 & ~n1668 ;
  assign n1768 = n1623 & n1753 ;
  assign n1769 = ( ~n1766 & n1767 ) | ( ~n1766 & n1768 ) | ( n1767 & n1768 ) ;
  assign n1770 = n1766 | n1769 ;
  assign n1771 = n1770 ^ n219 ^ x11 ;
  assign n1765 = n220 & ~n1764 ;
  assign n2106 = n1771 ^ n1765 ^ 1'b0 ;
  assign n2379 = n2145 ^ n2115 ^ n2106 ;
  assign n2380 = ( n2318 & n2378 ) | ( n2318 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2146 = ( n2106 & n2115 ) | ( n2106 & n2145 ) | ( n2115 & n2145 ) ;
  assign n1773 = ~n1622 & n1672 ;
  assign n1774 = n1621 & n1753 ;
  assign n1669 = n225 & ~n1668 ;
  assign n1670 = ~n1667 & n1669 ;
  assign n1775 = n1623 & n1670 ;
  assign n1776 = ( ~n1773 & n1774 ) | ( ~n1773 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1777 = n1773 | n1776 ;
  assign n1778 = ( ~n1654 & n1757 ) | ( ~n1654 & n1777 ) | ( n1757 & n1777 ) ;
  assign n1779 = n1777 ^ n1654 ^ 1'b0 ;
  assign n1780 = ( n1777 & n1778 ) | ( n1777 & ~n1779 ) | ( n1778 & ~n1779 ) ;
  assign n1781 = n1780 ^ n219 ^ x11 ;
  assign n1772 = n1765 & n1771 ;
  assign n2105 = n1781 ^ n1772 ^ 1'b0 ;
  assign n2096 = n1854 & n1943 ;
  assign n2097 = n2096 ^ n548 ^ 1'b0 ;
  assign n2098 = n1846 & n2066 ;
  assign n2099 = n1751 & n2068 ;
  assign n2100 = n1620 & n2071 ;
  assign n2101 = ( ~n2098 & n2099 ) | ( ~n2098 & n2100 ) | ( n2099 & n2100 ) ;
  assign n2102 = n2098 | n2101 ;
  assign n2103 = n2102 ^ n548 ^ 1'b0 ;
  assign n2104 = ( ~n548 & n2097 ) | ( ~n548 & n2103 ) | ( n2097 & n2103 ) ;
  assign n2381 = n2146 ^ n2105 ^ n2104 ;
  assign n2382 = ( n2310 & n2380 ) | ( n2310 & n2381 ) | ( n2380 & n2381 ) ;
  assign n1783 = ~n1622 & n1753 ;
  assign n1784 = n1620 & n1672 ;
  assign n1785 = n1621 & n1670 ;
  assign n1786 = ( ~n1783 & n1784 ) | ( ~n1783 & n1785 ) | ( n1784 & n1785 ) ;
  assign n1787 = n1783 | n1786 ;
  assign n1788 = ( ~n1626 & n1757 ) | ( ~n1626 & n1787 ) | ( n1757 & n1787 ) ;
  assign n1789 = n1787 ^ n1626 ^ 1'b0 ;
  assign n1790 = ( n1787 & n1788 ) | ( n1787 & ~n1789 ) | ( n1788 & ~n1789 ) ;
  assign n1791 = n1790 ^ n219 ^ x11 ;
  assign n1782 = n1772 & n1781 ;
  assign n228 = n227 ^ n220 ^ 1'b0 ;
  assign n1642 = n228 & n1623 ;
  assign n2148 = n1791 ^ n1782 ^ n1642 ;
  assign n2147 = ( n2104 & n2105 ) | ( n2104 & n2146 ) | ( n2105 & n2146 ) ;
  assign n2087 = n1936 & n1943 ;
  assign n2088 = n2087 ^ n548 ^ 1'b0 ;
  assign n2089 = n1928 & n2066 ;
  assign n2090 = n1846 & n2068 ;
  assign n2091 = n1751 & n2071 ;
  assign n2092 = ( ~n2089 & n2090 ) | ( ~n2089 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = n2089 | n2092 ;
  assign n2094 = n2093 ^ n548 ^ 1'b0 ;
  assign n2095 = ( ~n548 & n2088 ) | ( ~n548 & n2094 ) | ( n2088 & n2094 ) ;
  assign n2383 = n2148 ^ n2147 ^ n2095 ;
  assign n2384 = ( n2302 & n2382 ) | ( n2302 & n2383 ) | ( n2382 & n2383 ) ;
  assign n1792 = ( n1642 & n1782 ) | ( n1642 & n1791 ) | ( n1782 & n1791 ) ;
  assign n1671 = ~n1622 & n1670 ;
  assign n1752 = n1672 & n1751 ;
  assign n1754 = n1620 & n1753 ;
  assign n1755 = ( ~n1671 & n1752 ) | ( ~n1671 & n1754 ) | ( n1752 & n1754 ) ;
  assign n1756 = n1671 | n1755 ;
  assign n1758 = n1757 ^ n1756 ^ 1'b0 ;
  assign n1761 = ( n1757 & ~n1758 ) | ( n1757 & n1760 ) | ( ~n1758 & n1760 ) ;
  assign n1762 = ( n1756 & n1758 ) | ( n1756 & n1761 ) | ( n1758 & n1761 ) ;
  assign n1763 = n1762 ^ n219 ^ x11 ;
  assign n231 = n228 & n230 ;
  assign n1645 = n231 & n1644 ;
  assign n1646 = n1645 ^ n218 ^ 1'b0 ;
  assign n1635 = n228 & ~n230 ;
  assign n1647 = n1621 & n1635 ;
  assign n1629 = n229 ^ n227 ^ 1'b0 ;
  assign n1630 = ~n228 & n1629 ;
  assign n1648 = n1623 & n1630 ;
  assign n1649 = n1647 | n1648 ;
  assign n1650 = n1649 ^ n218 ^ 1'b0 ;
  assign n1651 = ( ~n218 & n1646 ) | ( ~n218 & n1650 ) | ( n1646 & n1650 ) ;
  assign n1643 = n218 & ~n1642 ;
  assign n1666 = n1651 ^ n1643 ^ 1'b0 ;
  assign n2150 = n1792 ^ n1763 ^ n1666 ;
  assign n2149 = ( n2095 & n2147 ) | ( n2095 & n2148 ) | ( n2147 & n2148 ) ;
  assign n2078 = n1943 & ~n2077 ;
  assign n2079 = n2078 ^ n548 ^ 1'b0 ;
  assign n2080 = ~n2060 & n2066 ;
  assign n2081 = n1928 & n2068 ;
  assign n2082 = n1846 & n2071 ;
  assign n2083 = ( ~n2080 & n2081 ) | ( ~n2080 & n2082 ) | ( n2081 & n2082 ) ;
  assign n2084 = n2080 | n2083 ;
  assign n2085 = n2084 ^ n548 ^ 1'b0 ;
  assign n2086 = ( ~n548 & n2079 ) | ( ~n548 & n2085 ) | ( n2079 & n2085 ) ;
  assign n2385 = n2150 ^ n2149 ^ n2086 ;
  assign n2284 = n2198 & n2242 ;
  assign n2285 = n2059 & n2201 ;
  assign n2286 = n2185 & n2203 ;
  assign n2287 = ( ~n2284 & n2285 ) | ( ~n2284 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = n2284 | n2287 ;
  assign n2289 = n2288 ^ n2275 ^ 1'b0 ;
  assign n2290 = n2277 ^ n2242 ^ n2185 ;
  assign n2291 = ( n2275 & ~n2289 ) | ( n2275 & n2290 ) | ( ~n2289 & n2290 ) ;
  assign n2292 = ( n2288 & n2289 ) | ( n2288 & n2291 ) | ( n2289 & n2291 ) ;
  assign n2293 = n2292 ^ n536 ^ x5 ;
  assign n2496 = n2385 ^ n2293 ^ 1'b0 ;
  assign n2497 = n2384 & n2496 ;
  assign n2498 = n2384 | n2496 ;
  assign n2499 = n540 & n2478 ;
  assign n2500 = ~n1654 & n2499 ;
  assign n2501 = n1623 & n2423 ;
  assign n2502 = n1621 & n2422 ;
  assign n2503 = ( n540 & n2501 ) | ( n540 & ~n2502 ) | ( n2501 & ~n2502 ) ;
  assign n2504 = ~n2501 & n2503 ;
  assign n2505 = ( n1644 & n2499 ) | ( n1644 & ~n2504 ) | ( n2499 & ~n2504 ) ;
  assign n2506 = n2505 ^ n2504 ^ 1'b0 ;
  assign n2507 = ( n2504 & ~n2505 ) | ( n2504 & n2506 ) | ( ~n2505 & n2506 ) ;
  assign n2508 = n1621 & n2423 ;
  assign n2509 = n1623 & n2459 ;
  assign n2510 = n2508 | n2509 ;
  assign n2511 = ~n1622 & n2422 ;
  assign n2512 = ( n540 & n2510 ) | ( n540 & n2511 ) | ( n2510 & n2511 ) ;
  assign n2513 = n2511 ^ n2510 ^ 1'b0 ;
  assign n2514 = ( n540 & n2512 ) | ( n540 & n2513 ) | ( n2512 & n2513 ) ;
  assign n2515 = ( n2500 & n2507 ) | ( n2500 & ~n2514 ) | ( n2507 & ~n2514 ) ;
  assign n2516 = ~n2500 & n2515 ;
  assign n2517 = ( x0 & n1623 ) | ( x0 & ~n2516 ) | ( n1623 & ~n2516 ) ;
  assign n2518 = n2517 ^ n2516 ^ 1'b0 ;
  assign n2519 = ( n2516 & ~n2517 ) | ( n2516 & n2518 ) | ( ~n2517 & n2518 ) ;
  assign n2520 = ~n1622 & n2423 ;
  assign n2521 = n1621 & n2459 ;
  assign n2522 = n1620 & n2422 ;
  assign n2523 = ( ~n2520 & n2521 ) | ( ~n2520 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2524 = n2520 | n2523 ;
  assign n2525 = ( ~n1626 & n2478 ) | ( ~n1626 & n2524 ) | ( n2478 & n2524 ) ;
  assign n2526 = n2524 ^ n1626 ^ 1'b0 ;
  assign n2527 = ( n2524 & n2525 ) | ( n2524 & ~n2526 ) | ( n2525 & ~n2526 ) ;
  assign n2528 = n2527 ^ n539 ^ n537 ;
  assign n2529 = ( n2348 & n2519 ) | ( n2348 & n2528 ) | ( n2519 & n2528 ) ;
  assign n2530 = n1751 & n2422 ;
  assign n2531 = ~n1622 & n2459 ;
  assign n2532 = n1620 & n2423 ;
  assign n2533 = ( ~n2530 & n2531 ) | ( ~n2530 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2534 = n2530 | n2533 ;
  assign n2535 = n540 & n2534 ;
  assign n2536 = n2355 ^ n2349 ^ 1'b0 ;
  assign n2537 = n2529 | n2536 ;
  assign n2538 = n1760 & n2499 ;
  assign n2539 = n2537 & ~n2538 ;
  assign n2540 = n1760 & n2478 ;
  assign n2541 = ( n540 & n2534 ) | ( n540 & ~n2540 ) | ( n2534 & ~n2540 ) ;
  assign n2542 = n2540 | n2541 ;
  assign n2543 = ( n2535 & n2539 ) | ( n2535 & n2542 ) | ( n2539 & n2542 ) ;
  assign n2544 = ~n2535 & n2543 ;
  assign n2545 = n2544 ^ n2529 ^ 1'b0 ;
  assign n2546 = ( ~n2529 & n2536 ) | ( ~n2529 & n2545 ) | ( n2536 & n2545 ) ;
  assign n2547 = ( n2529 & n2544 ) | ( n2529 & n2546 ) | ( n2544 & n2546 ) ;
  assign n2548 = n2356 | n2364 ;
  assign n2549 = n1846 & n2422 ;
  assign n2550 = n1751 & n2423 ;
  assign n2551 = n1620 & n2459 ;
  assign n2552 = ( ~n2549 & n2550 ) | ( ~n2549 & n2551 ) | ( n2550 & n2551 ) ;
  assign n2553 = n2549 | n2552 ;
  assign n2554 = n2553 ^ n1854 ^ 1'b0 ;
  assign n2555 = ( ~n1854 & n2478 ) | ( ~n1854 & n2554 ) | ( n2478 & n2554 ) ;
  assign n2556 = ( n1854 & n2553 ) | ( n1854 & n2555 ) | ( n2553 & n2555 ) ;
  assign n2557 = n2556 ^ n539 ^ n537 ;
  assign n2558 = n2547 | n2557 ;
  assign n2559 = ( n2365 & n2548 ) | ( n2365 & n2558 ) | ( n2548 & n2558 ) ;
  assign n2560 = ~n2365 & n2559 ;
  assign n2561 = n2560 ^ n2547 ^ 1'b0 ;
  assign n2562 = ( ~n2547 & n2557 ) | ( ~n2547 & n2561 ) | ( n2557 & n2561 ) ;
  assign n2563 = ( n2547 & n2560 ) | ( n2547 & n2562 ) | ( n2560 & n2562 ) ;
  assign n2564 = n1928 & n2422 ;
  assign n2565 = n1846 & n2423 ;
  assign n2566 = n1751 & n2459 ;
  assign n2567 = ( ~n2564 & n2565 ) | ( ~n2564 & n2566 ) | ( n2565 & n2566 ) ;
  assign n2568 = n2564 | n2567 ;
  assign n2569 = n540 & n2568 ;
  assign n2570 = n1936 & n2478 ;
  assign n2571 = ( n540 & n2568 ) | ( n540 & ~n2570 ) | ( n2568 & ~n2570 ) ;
  assign n2572 = n2570 | n2571 ;
  assign n2573 = n2373 ^ n2365 ^ n2123 ;
  assign n2574 = n2563 | n2573 ;
  assign n2575 = n1936 & n2499 ;
  assign n2576 = n2574 & ~n2575 ;
  assign n2577 = ( n2569 & n2572 ) | ( n2569 & n2576 ) | ( n2572 & n2576 ) ;
  assign n2578 = ~n2569 & n2577 ;
  assign n2579 = n2578 ^ n2563 ^ 1'b0 ;
  assign n2580 = ( ~n2563 & n2573 ) | ( ~n2563 & n2579 ) | ( n2573 & n2579 ) ;
  assign n2581 = ( n2563 & n2578 ) | ( n2563 & n2580 ) | ( n2578 & n2580 ) ;
  assign n2582 = n2347 ^ n2338 ^ 1'b0 ;
  assign n2583 = n2374 & n2582 ;
  assign n2584 = n2374 | n2582 ;
  assign n2585 = ~n2060 & n2422 ;
  assign n2586 = n1928 & n2423 ;
  assign n2587 = n1846 & n2459 ;
  assign n2588 = ( ~n2585 & n2586 ) | ( ~n2585 & n2587 ) | ( n2586 & n2587 ) ;
  assign n2589 = n2585 | n2588 ;
  assign n2590 = ( ~n2077 & n2478 ) | ( ~n2077 & n2589 ) | ( n2478 & n2589 ) ;
  assign n2591 = n2589 ^ n2077 ^ 1'b0 ;
  assign n2592 = ( n2589 & n2590 ) | ( n2589 & ~n2591 ) | ( n2590 & ~n2591 ) ;
  assign n2593 = n2592 ^ n539 ^ n537 ;
  assign n2594 = n2581 | n2593 ;
  assign n2595 = ( n2583 & n2584 ) | ( n2583 & n2594 ) | ( n2584 & n2594 ) ;
  assign n2596 = ~n2583 & n2595 ;
  assign n2597 = n2596 ^ n2581 ^ 1'b0 ;
  assign n2598 = ( ~n2581 & n2593 ) | ( ~n2581 & n2597 ) | ( n2593 & n2597 ) ;
  assign n2599 = ( n2581 & n2596 ) | ( n2581 & n2598 ) | ( n2596 & n2598 ) ;
  assign n2600 = n2059 & n2422 ;
  assign n2601 = ~n2060 & n2423 ;
  assign n2602 = n1928 & n2459 ;
  assign n2603 = ( ~n2600 & n2601 ) | ( ~n2600 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = n2600 | n2603 ;
  assign n2605 = n540 & n2604 ;
  assign n2606 = ~n2063 & n2478 ;
  assign n2607 = ( n540 & n2604 ) | ( n540 & ~n2606 ) | ( n2604 & ~n2606 ) ;
  assign n2608 = n2606 | n2607 ;
  assign n2609 = n2375 ^ n2337 ^ n2336 ;
  assign n2610 = n2599 | n2609 ;
  assign n2611 = ~n2063 & n2499 ;
  assign n2612 = n2610 & ~n2611 ;
  assign n2613 = ( n2605 & n2608 ) | ( n2605 & n2612 ) | ( n2608 & n2612 ) ;
  assign n2614 = ~n2605 & n2613 ;
  assign n2615 = n2614 ^ n2599 ^ 1'b0 ;
  assign n2616 = ( ~n2599 & n2609 ) | ( ~n2599 & n2615 ) | ( n2609 & n2615 ) ;
  assign n2617 = ( n2599 & n2614 ) | ( n2599 & n2616 ) | ( n2614 & n2616 ) ;
  assign n2618 = n2185 & n2422 ;
  assign n2619 = n2059 & n2423 ;
  assign n2620 = ~n2060 & n2459 ;
  assign n2621 = ( ~n2618 & n2619 ) | ( ~n2618 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2622 = n2618 | n2621 ;
  assign n2623 = n540 & n2622 ;
  assign n2624 = n2186 & n2478 ;
  assign n2625 = ( n540 & n2622 ) | ( n540 & ~n2624 ) | ( n2622 & ~n2624 ) ;
  assign n2626 = n2624 | n2625 ;
  assign n2627 = n2377 ^ n2376 ^ n2327 ;
  assign n2628 = n2617 | n2627 ;
  assign n2629 = n2186 & n2499 ;
  assign n2630 = n2628 & ~n2629 ;
  assign n2631 = ( n2623 & n2626 ) | ( n2623 & n2630 ) | ( n2626 & n2630 ) ;
  assign n2632 = ~n2623 & n2631 ;
  assign n2633 = n2632 ^ n2617 ^ 1'b0 ;
  assign n2634 = ( ~n2617 & n2627 ) | ( ~n2617 & n2633 ) | ( n2627 & n2633 ) ;
  assign n2635 = ( n2617 & n2632 ) | ( n2617 & n2634 ) | ( n2632 & n2634 ) ;
  assign n2636 = n2242 & n2422 ;
  assign n2637 = n2185 & n2423 ;
  assign n2638 = n2059 & n2459 ;
  assign n2639 = ( ~n2636 & n2637 ) | ( ~n2636 & n2638 ) | ( n2637 & n2638 ) ;
  assign n2640 = n2636 | n2639 ;
  assign n2641 = n540 & n2640 ;
  assign n2642 = n2290 & n2478 ;
  assign n2643 = ( n540 & n2640 ) | ( n540 & ~n2642 ) | ( n2640 & ~n2642 ) ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n2379 ^ n2378 ^ n2318 ;
  assign n2646 = n2635 | n2645 ;
  assign n2647 = n2290 & n2499 ;
  assign n2648 = n2646 & ~n2647 ;
  assign n2649 = ( n2641 & n2644 ) | ( n2641 & n2648 ) | ( n2644 & n2648 ) ;
  assign n2650 = ~n2641 & n2649 ;
  assign n2651 = n2650 ^ n2635 ^ 1'b0 ;
  assign n2652 = ( ~n2635 & n2645 ) | ( ~n2635 & n2651 ) | ( n2645 & n2651 ) ;
  assign n2653 = ( n2635 & n2650 ) | ( n2635 & n2652 ) | ( n2650 & n2652 ) ;
  assign n2654 = ~n2272 & n2422 ;
  assign n2655 = n2242 & n2423 ;
  assign n2656 = n2185 & n2459 ;
  assign n2657 = ( ~n2654 & n2655 ) | ( ~n2654 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = n2654 | n2657 ;
  assign n2276 = n2272 ^ n2242 ^ 1'b0 ;
  assign n2279 = n2278 ^ n2276 ^ 1'b0 ;
  assign n2659 = ( ~n2279 & n2478 ) | ( ~n2279 & n2658 ) | ( n2478 & n2658 ) ;
  assign n2660 = n2658 ^ n2279 ^ 1'b0 ;
  assign n2661 = ( n2658 & n2659 ) | ( n2658 & ~n2660 ) | ( n2659 & ~n2660 ) ;
  assign n2662 = n2661 ^ n539 ^ n537 ;
  assign n2663 = n2381 ^ n2380 ^ n2310 ;
  assign n2664 = ( n2653 & n2662 ) | ( n2653 & n2663 ) | ( n2662 & n2663 ) ;
  assign n2665 = n2406 & n2422 ;
  assign n2666 = ~n2272 & n2423 ;
  assign n2667 = n2242 & n2459 ;
  assign n2668 = ( ~n2665 & n2666 ) | ( ~n2665 & n2667 ) | ( n2666 & n2667 ) ;
  assign n2669 = n2665 | n2668 ;
  assign n2413 = n2412 ^ n2406 ^ n2272 ;
  assign n2670 = ( ~n2413 & n2478 ) | ( ~n2413 & n2669 ) | ( n2478 & n2669 ) ;
  assign n2671 = n2669 ^ n2413 ^ 1'b0 ;
  assign n2672 = ( n2669 & n2670 ) | ( n2669 & ~n2671 ) | ( n2670 & ~n2671 ) ;
  assign n2673 = n2672 ^ n539 ^ n537 ;
  assign n2674 = n2383 ^ n2382 ^ n2302 ;
  assign n2675 = ( n2664 & n2673 ) | ( n2664 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = n2495 | n2675 ;
  assign n2677 = ( n2497 & n2498 ) | ( n2497 & n2676 ) | ( n2498 & n2676 ) ;
  assign n2678 = ~n2497 & n2677 ;
  assign n2679 = n2678 ^ n2495 ^ 1'b0 ;
  assign n2680 = ( ~n2495 & n2675 ) | ( ~n2495 & n2679 ) | ( n2675 & n2679 ) ;
  assign n2681 = ( n2495 & n2678 ) | ( n2495 & n2680 ) | ( n2678 & n2680 ) ;
  assign n1655 = n231 & ~n1654 ;
  assign n1656 = n1655 ^ n218 ^ 1'b0 ;
  assign n1657 = ~n1622 & n1635 ;
  assign n1632 = ~n228 & n230 ;
  assign n1633 = ~n1629 & n1632 ;
  assign n1658 = n1623 & n1633 ;
  assign n1659 = n1621 & n1630 ;
  assign n1660 = ( ~n1657 & n1658 ) | ( ~n1657 & n1659 ) | ( n1658 & n1659 ) ;
  assign n1661 = n1657 | n1660 ;
  assign n1662 = n1661 ^ n218 ^ 1'b0 ;
  assign n1663 = ( ~n218 & n1656 ) | ( ~n218 & n1662 ) | ( n1656 & n1662 ) ;
  assign n1652 = n1643 & n1651 ;
  assign n1858 = n1663 ^ n1652 ^ 1'b0 ;
  assign n1847 = n1672 & n1846 ;
  assign n1848 = n1751 & n1753 ;
  assign n1849 = n1620 & n1670 ;
  assign n1850 = ( ~n1847 & n1848 ) | ( ~n1847 & n1849 ) | ( n1848 & n1849 ) ;
  assign n1851 = n1847 | n1850 ;
  assign n1852 = n1851 ^ n1757 ^ 1'b0 ;
  assign n1855 = ( n1757 & ~n1852 ) | ( n1757 & n1854 ) | ( ~n1852 & n1854 ) ;
  assign n1856 = ( n1851 & n1852 ) | ( n1851 & n1855 ) | ( n1852 & n1855 ) ;
  assign n1857 = n1856 ^ n219 ^ x11 ;
  assign n1793 = ( n1666 & n1763 ) | ( n1666 & n1792 ) | ( n1763 & n1792 ) ;
  assign n2152 = n1858 ^ n1857 ^ n1793 ;
  assign n2151 = ( n2086 & n2149 ) | ( n2086 & n2150 ) | ( n2149 & n2150 ) ;
  assign n2064 = n1943 & ~n2063 ;
  assign n2065 = n2064 ^ n548 ^ 1'b0 ;
  assign n2067 = n2059 & n2066 ;
  assign n2069 = ~n2060 & n2068 ;
  assign n2072 = n1928 & n2071 ;
  assign n2073 = ( ~n2067 & n2069 ) | ( ~n2067 & n2072 ) | ( n2069 & n2072 ) ;
  assign n2074 = n2067 | n2073 ;
  assign n2075 = n2074 ^ n548 ^ 1'b0 ;
  assign n2076 = ( ~n548 & n2065 ) | ( ~n548 & n2075 ) | ( n2065 & n2075 ) ;
  assign n2387 = n2152 ^ n2151 ^ n2076 ;
  assign n2386 = ( n2293 & n2384 ) | ( n2293 & n2385 ) | ( n2384 & n2385 ) ;
  assign n2202 = n2185 & n2201 ;
  assign n2243 = n2203 & n2242 ;
  assign n2244 = n2202 | n2243 ;
  assign n2273 = ~n2244 & n2272 ;
  assign n2274 = ( n2198 & n2244 ) | ( n2198 & ~n2273 ) | ( n2244 & ~n2273 ) ;
  assign n2280 = ( n2274 & n2275 ) | ( n2274 & ~n2279 ) | ( n2275 & ~n2279 ) ;
  assign n2281 = n2279 ^ n2274 ^ 1'b0 ;
  assign n2282 = ( n2274 & n2280 ) | ( n2274 & ~n2281 ) | ( n2280 & ~n2281 ) ;
  assign n2283 = n2282 ^ n536 ^ x5 ;
  assign n2682 = n2387 ^ n2386 ^ n2283 ;
  assign n2683 = ( n2485 & n2681 ) | ( n2485 & n2682 ) | ( n2681 & n2682 ) ;
  assign n2407 = n2198 & n2406 ;
  assign n2408 = n2203 & ~n2272 ;
  assign n2409 = n2201 & n2242 ;
  assign n2410 = ( ~n2407 & n2408 ) | ( ~n2407 & n2409 ) | ( n2408 & n2409 ) ;
  assign n2411 = n2407 | n2410 ;
  assign n2414 = ( n2275 & n2411 ) | ( n2275 & ~n2413 ) | ( n2411 & ~n2413 ) ;
  assign n2415 = n2414 ^ n2275 ^ 1'b0 ;
  assign n2416 = ( n2411 & n2414 ) | ( n2411 & ~n2415 ) | ( n2414 & ~n2415 ) ;
  assign n2417 = n2416 ^ n536 ^ x5 ;
  assign n2388 = ( n2283 & n2386 ) | ( n2283 & n2387 ) | ( n2386 & n2387 ) ;
  assign n2187 = n1943 & n2186 ;
  assign n2188 = n2187 ^ n548 ^ 1'b0 ;
  assign n2189 = n2066 & n2185 ;
  assign n2190 = n2059 & n2068 ;
  assign n2191 = ~n2060 & n2071 ;
  assign n2192 = ( ~n2189 & n2190 ) | ( ~n2189 & n2191 ) | ( n2190 & n2191 ) ;
  assign n2193 = n2189 | n2192 ;
  assign n2194 = n2193 ^ n548 ^ 1'b0 ;
  assign n2195 = ( ~n548 & n2188 ) | ( ~n548 & n2194 ) | ( n2188 & n2194 ) ;
  assign n2153 = ( n2076 & n2151 ) | ( n2076 & n2152 ) | ( n2151 & n2152 ) ;
  assign n1929 = n1672 & n1928 ;
  assign n1930 = n1753 & n1846 ;
  assign n1931 = n1670 & n1751 ;
  assign n1932 = ( ~n1929 & n1930 ) | ( ~n1929 & n1931 ) | ( n1930 & n1931 ) ;
  assign n1933 = n1929 | n1932 ;
  assign n1934 = n1933 ^ n1757 ^ 1'b0 ;
  assign n1937 = ( ~n1757 & n1934 ) | ( ~n1757 & n1936 ) | ( n1934 & n1936 ) ;
  assign n1938 = ( n1757 & n1933 ) | ( n1757 & n1937 ) | ( n1933 & n1937 ) ;
  assign n1939 = n1938 ^ n219 ^ x11 ;
  assign n1859 = ( n1793 & n1857 ) | ( n1793 & n1858 ) | ( n1857 & n1858 ) ;
  assign n1664 = n1652 & n1663 ;
  assign n1641 = n218 & n1623 ;
  assign n1627 = n231 & ~n1626 ;
  assign n1628 = n1627 ^ n218 ^ 1'b0 ;
  assign n1631 = ~n1622 & n1630 ;
  assign n1634 = n1621 & n1633 ;
  assign n1636 = n1620 & n1635 ;
  assign n1637 = ( ~n1631 & n1634 ) | ( ~n1631 & n1636 ) | ( n1634 & n1636 ) ;
  assign n1638 = n1631 | n1637 ;
  assign n1639 = n1638 ^ n218 ^ 1'b0 ;
  assign n1640 = ( ~n218 & n1628 ) | ( ~n218 & n1639 ) | ( n1628 & n1639 ) ;
  assign n1665 = n1664 ^ n1641 ^ n1640 ;
  assign n1940 = n1939 ^ n1859 ^ n1665 ;
  assign n2196 = n2195 ^ n2153 ^ n1940 ;
  assign n2418 = n2417 ^ n2388 ^ n2196 ;
  assign n2708 = n2707 ^ n2683 ^ n2418 ;
  assign n2709 = n2682 ^ n2485 ^ 1'b0 ;
  assign n2710 = n269 | n511 ;
  assign n2711 = ( n332 & n377 ) | ( n332 & ~n2710 ) | ( n377 & ~n2710 ) ;
  assign n2712 = n2710 | n2711 ;
  assign n2713 = n275 | n799 ;
  assign n2714 = n1919 | n2713 ;
  assign n2715 = ( n238 & n364 ) | ( n238 & ~n2714 ) | ( n364 & ~n2714 ) ;
  assign n2716 = n2714 | n2715 ;
  assign n2717 = ( n134 & n379 ) | ( n134 & ~n2716 ) | ( n379 & ~n2716 ) ;
  assign n2718 = n2716 | n2717 ;
  assign n2719 = n566 | n2259 ;
  assign n2720 = ( n193 & n243 ) | ( n193 & ~n2719 ) | ( n243 & ~n2719 ) ;
  assign n2721 = n2719 | n2720 ;
  assign n2722 = ( ~n2712 & n2718 ) | ( ~n2712 & n2721 ) | ( n2718 & n2721 ) ;
  assign n2723 = n2712 | n2722 ;
  assign n2724 = ( n319 & n1720 ) | ( n319 & ~n2723 ) | ( n1720 & ~n2723 ) ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = ( n102 & n303 ) | ( n102 & ~n2725 ) | ( n303 & ~n2725 ) ;
  assign n2727 = n2725 | n2726 ;
  assign n2728 = ( n316 & n349 ) | ( n316 & ~n2727 ) | ( n349 & ~n2727 ) ;
  assign n2729 = n2727 | n2728 ;
  assign n2730 = ( n370 & n445 ) | ( n370 & ~n2729 ) | ( n445 & ~n2729 ) ;
  assign n2731 = n2729 | n2730 ;
  assign n2732 = n2731 ^ n2709 ^ 1'b0 ;
  assign n2733 = ( n2681 & n2709 ) | ( n2681 & n2732 ) | ( n2709 & n2732 ) ;
  assign n2734 = n2733 ^ n2709 ^ 1'b0 ;
  assign n2735 = ( n215 & n2708 ) | ( n215 & n2734 ) | ( n2708 & n2734 ) ;
  assign n2736 = n122 | n258 ;
  assign n2737 = n137 | n2736 ;
  assign n2738 = n72 | n2737 ;
  assign n2739 = ( n163 & n328 ) | ( n163 & ~n2738 ) | ( n328 & ~n2738 ) ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n136 | n232 ;
  assign n2742 = n1961 | n2741 ;
  assign n2743 = n2740 | n2742 ;
  assign n2744 = ( n195 & n299 ) | ( n195 & ~n2743 ) | ( n299 & ~n2743 ) ;
  assign n2745 = n2743 | n2744 ;
  assign n2746 = ( n168 & n349 ) | ( n168 & ~n2745 ) | ( n349 & ~n2745 ) ;
  assign n2747 = n2745 | n2746 ;
  assign n2748 = ( n156 & n445 ) | ( n156 & ~n2747 ) | ( n445 & ~n2747 ) ;
  assign n2749 = n2747 | n2748 ;
  assign n2750 = ( n142 & n182 ) | ( n142 & ~n2749 ) | ( n182 & ~n2749 ) ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n234 | n2751 ;
  assign n2753 = n282 | n2752 ;
  assign n2754 = ( n310 & n426 ) | ( n310 & ~n2753 ) | ( n426 & ~n2753 ) ;
  assign n2755 = n2753 | n2754 ;
  assign n2756 = n350 | n2252 ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = n814 | n2432 ;
  assign n2759 = n477 | n2758 ;
  assign n2760 = ( n138 & n451 ) | ( n138 & ~n2759 ) | ( n451 & ~n2759 ) ;
  assign n2761 = n2759 | n2760 ;
  assign n2762 = ( n2429 & ~n2757 ) | ( n2429 & n2761 ) | ( ~n2757 & n2761 ) ;
  assign n2763 = n2757 | n2762 ;
  assign n2764 = ( n255 & n304 ) | ( n255 & ~n2763 ) | ( n304 & ~n2763 ) ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = ( n149 & n157 ) | ( n149 & ~n2765 ) | ( n157 & ~n2765 ) ;
  assign n2767 = n2765 | n2766 ;
  assign n2768 = ( n87 & n325 ) | ( n87 & ~n2767 ) | ( n325 & ~n2767 ) ;
  assign n2769 = n2767 | n2768 ;
  assign n2770 = ( n118 & n263 ) | ( n118 & ~n2769 ) | ( n263 & ~n2769 ) ;
  assign n2771 = n2769 | n2770 ;
  assign n2841 = ( n2418 & n2683 ) | ( n2418 & n2707 ) | ( n2683 & n2707 ) ;
  assign n2773 = n384 | n786 ;
  assign n2774 = n240 | n2773 ;
  assign n2775 = n792 | n2774 ;
  assign n2776 = ( n500 & n813 ) | ( n500 & ~n2775 ) | ( n813 & ~n2775 ) ;
  assign n2777 = n2775 | n2776 ;
  assign n2778 = ( n394 & n807 ) | ( n394 & ~n2777 ) | ( n807 & ~n2777 ) ;
  assign n2779 = n2777 | n2778 ;
  assign n2780 = ( n328 & n349 ) | ( n328 & ~n2779 ) | ( n349 & ~n2779 ) ;
  assign n2781 = n2779 | n2780 ;
  assign n2772 = n2684 & ~n2695 ;
  assign n2782 = n2781 ^ n2772 ^ 1'b0 ;
  assign n2783 = n2422 & n2782 ;
  assign n2784 = n2423 & n2696 ;
  assign n2785 = n2459 & ~n2475 ;
  assign n2786 = ( ~n2783 & n2784 ) | ( ~n2783 & n2785 ) | ( n2784 & n2785 ) ;
  assign n2787 = n2783 | n2786 ;
  assign n2788 = n2787 ^ n2478 ^ 1'b0 ;
  assign n2789 = ( ~n2475 & n2696 ) | ( ~n2475 & n2702 ) | ( n2696 & n2702 ) ;
  assign n2790 = n2789 ^ n2782 ^ n2696 ;
  assign n2791 = ( n2478 & ~n2788 ) | ( n2478 & n2790 ) | ( ~n2788 & n2790 ) ;
  assign n2792 = ( n2787 & n2788 ) | ( n2787 & n2791 ) | ( n2788 & n2791 ) ;
  assign n2793 = n2792 ^ n539 ^ n537 ;
  assign n2836 = ( n2196 & n2388 ) | ( n2196 & n2417 ) | ( n2388 & n2417 ) ;
  assign n2827 = n2198 & n2457 ;
  assign n2828 = n2203 & n2406 ;
  assign n2829 = n2201 & ~n2272 ;
  assign n2830 = ( ~n2827 & n2828 ) | ( ~n2827 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = n2827 | n2830 ;
  assign n2832 = n2831 ^ n2275 ^ 1'b0 ;
  assign n2833 = ( ~n2275 & n2492 ) | ( ~n2275 & n2832 ) | ( n2492 & n2832 ) ;
  assign n2834 = ( n2275 & n2831 ) | ( n2275 & n2833 ) | ( n2831 & n2833 ) ;
  assign n2835 = n2834 ^ n536 ^ x5 ;
  assign n2825 = ( n1940 & n2153 ) | ( n1940 & n2195 ) | ( n2153 & n2195 ) ;
  assign n2816 = n1943 & n2290 ;
  assign n2817 = n2816 ^ n548 ^ 1'b0 ;
  assign n2818 = n2066 & n2242 ;
  assign n2819 = n2068 & n2185 ;
  assign n2820 = n2059 & n2071 ;
  assign n2821 = ( ~n2818 & n2819 ) | ( ~n2818 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2822 = n2818 | n2821 ;
  assign n2823 = n2822 ^ n548 ^ 1'b0 ;
  assign n2824 = ( ~n548 & n2817 ) | ( ~n548 & n2823 ) | ( n2817 & n2823 ) ;
  assign n2814 = ( n1665 & n1859 ) | ( n1665 & n1939 ) | ( n1859 & n1939 ) ;
  assign n2806 = n1672 & ~n2060 ;
  assign n2807 = n1753 & n1928 ;
  assign n2808 = n1670 & n1846 ;
  assign n2809 = ( ~n2806 & n2807 ) | ( ~n2806 & n2808 ) | ( n2807 & n2808 ) ;
  assign n2810 = n2806 | n2809 ;
  assign n2811 = n2077 & ~n2810 ;
  assign n2812 = ( n1757 & n2810 ) | ( n1757 & ~n2811 ) | ( n2810 & ~n2811 ) ;
  assign n2813 = n2812 ^ n219 ^ x11 ;
  assign n2804 = ( n1640 & n1641 ) | ( n1640 & n1664 ) | ( n1641 & n1664 ) ;
  assign n2795 = ~n1622 & n1633 ;
  assign n2796 = n1635 & n1751 ;
  assign n2797 = n1620 & n1630 ;
  assign n2798 = ( ~n2795 & n2796 ) | ( ~n2795 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2799 = n2795 | n2798 ;
  assign n2800 = n2799 ^ n231 ^ 1'b0 ;
  assign n2801 = ( ~n231 & n1760 ) | ( ~n231 & n2800 ) | ( n1760 & n2800 ) ;
  assign n2802 = ( n231 & n2799 ) | ( n231 & n2801 ) | ( n2799 & n2801 ) ;
  assign n2794 = n218 & n1621 ;
  assign n2803 = n2802 ^ n2794 ^ n218 ;
  assign n2805 = n2804 ^ n2803 ^ 1'b0 ;
  assign n2815 = n2814 ^ n2813 ^ n2805 ;
  assign n2826 = n2825 ^ n2824 ^ n2815 ;
  assign n2837 = n2836 ^ n2835 ^ n2826 ;
  assign n2838 = n2793 & n2837 ;
  assign n2839 = n2793 | n2837 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2842 = n2841 ^ n2840 ^ 1'b0 ;
  assign n2935 = ( n2735 & n2771 ) | ( n2735 & n2842 ) | ( n2771 & n2842 ) ;
  assign n2898 = n2423 & n2782 ;
  assign n2899 = n2459 & n2696 ;
  assign n2900 = n2898 | n2899 ;
  assign n2922 = n2772 & ~n2781 ;
  assign n2901 = n438 | n2741 ;
  assign n2902 = ( n157 & n580 ) | ( n157 & ~n2901 ) | ( n580 & ~n2901 ) ;
  assign n2903 = n2901 | n2902 ;
  assign n2904 = ( n105 & n305 ) | ( n105 & ~n2903 ) | ( n305 & ~n2903 ) ;
  assign n2905 = n2903 | n2904 ;
  assign n2906 = ( n178 & n266 ) | ( n178 & ~n2905 ) | ( n266 & ~n2905 ) ;
  assign n2907 = n2905 | n2906 ;
  assign n2908 = n399 | n2263 ;
  assign n2909 = n278 | n485 ;
  assign n2910 = ( n889 & n2908 ) | ( n889 & ~n2909 ) | ( n2908 & ~n2909 ) ;
  assign n2911 = ~n2908 & n2910 ;
  assign n2912 = ( n261 & ~n2907 ) | ( n261 & n2911 ) | ( ~n2907 & n2911 ) ;
  assign n2913 = ~n261 & n2912 ;
  assign n2914 = ( n195 & ~n303 ) | ( n195 & n2913 ) | ( ~n303 & n2913 ) ;
  assign n2915 = ~n195 & n2914 ;
  assign n2916 = ( n321 & ~n445 ) | ( n321 & n2915 ) | ( ~n445 & n2915 ) ;
  assign n2917 = ~n321 & n2916 ;
  assign n2918 = ( ~n131 & n426 ) | ( ~n131 & n2917 ) | ( n426 & n2917 ) ;
  assign n2919 = ~n426 & n2918 ;
  assign n2920 = ( ~n163 & n253 ) | ( ~n163 & n2919 ) | ( n253 & n2919 ) ;
  assign n2921 = ~n253 & n2920 ;
  assign n2923 = n2922 ^ n2921 ^ 1'b0 ;
  assign n2924 = ~n2900 & n2923 ;
  assign n2925 = ( n2422 & n2900 ) | ( n2422 & ~n2924 ) | ( n2900 & ~n2924 ) ;
  assign n2927 = ( n2696 & n2782 ) | ( n2696 & n2789 ) | ( n2782 & n2789 ) ;
  assign n2926 = n2923 ^ n2782 ^ 1'b0 ;
  assign n2928 = n2927 ^ n2926 ^ 1'b0 ;
  assign n2929 = ( n2478 & n2925 ) | ( n2478 & ~n2928 ) | ( n2925 & ~n2928 ) ;
  assign n2930 = n2928 ^ n2925 ^ 1'b0 ;
  assign n2931 = ( n2925 & n2929 ) | ( n2925 & ~n2930 ) | ( n2929 & ~n2930 ) ;
  assign n2932 = n2931 ^ n539 ^ n537 ;
  assign n2896 = ( n2826 & n2835 ) | ( n2826 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2888 = n2203 & n2457 ;
  assign n2889 = n2201 & n2406 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = n2475 & ~n2890 ;
  assign n2892 = ( n2198 & n2890 ) | ( n2198 & ~n2891 ) | ( n2890 & ~n2891 ) ;
  assign n2893 = n2481 & ~n2892 ;
  assign n2894 = ( n2275 & n2892 ) | ( n2275 & ~n2893 ) | ( n2892 & ~n2893 ) ;
  assign n2895 = n2894 ^ n536 ^ x5 ;
  assign n2878 = n1943 & ~n2279 ;
  assign n2879 = n2878 ^ n548 ^ 1'b0 ;
  assign n2880 = n2066 & ~n2272 ;
  assign n2881 = n2068 & n2242 ;
  assign n2882 = n2071 & n2185 ;
  assign n2883 = ( ~n2880 & n2881 ) | ( ~n2880 & n2882 ) | ( n2881 & n2882 ) ;
  assign n2884 = n2880 | n2883 ;
  assign n2885 = n2884 ^ n548 ^ 1'b0 ;
  assign n2886 = ( ~n548 & n2879 ) | ( ~n548 & n2885 ) | ( n2879 & n2885 ) ;
  assign n2877 = ( n2815 & n2824 ) | ( n2815 & n2825 ) | ( n2824 & n2825 ) ;
  assign n2875 = ( n2805 & n2813 ) | ( n2805 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2865 = n1635 & n1846 ;
  assign n2866 = n1620 & n1633 ;
  assign n2867 = n1630 & n1751 ;
  assign n2868 = ( ~n2865 & n2866 ) | ( ~n2865 & n2867 ) | ( n2866 & n2867 ) ;
  assign n2869 = n2865 | n2868 ;
  assign n2870 = n2869 ^ n231 ^ 1'b0 ;
  assign n2871 = ( ~n231 & n1854 ) | ( ~n231 & n2870 ) | ( n1854 & n2870 ) ;
  assign n2872 = ( n231 & n2869 ) | ( n231 & n2871 ) | ( n2869 & n2871 ) ;
  assign n2864 = n218 & n1622 ;
  assign n2873 = n2872 ^ n2864 ^ 1'b0 ;
  assign n2863 = ( n2794 & n2804 ) | ( n2794 & ~n2805 ) | ( n2804 & ~n2805 ) ;
  assign n2874 = n2873 ^ n2863 ^ 1'b0 ;
  assign n2855 = n1672 & n2059 ;
  assign n2856 = n1753 & ~n2060 ;
  assign n2857 = n1670 & n1928 ;
  assign n2858 = ( ~n2855 & n2856 ) | ( ~n2855 & n2857 ) | ( n2856 & n2857 ) ;
  assign n2859 = n2855 | n2858 ;
  assign n2860 = n2063 & ~n2859 ;
  assign n2861 = ( n1757 & n2859 ) | ( n1757 & ~n2860 ) | ( n2859 & ~n2860 ) ;
  assign n2862 = n2861 ^ n219 ^ x11 ;
  assign n2876 = n2875 ^ n2874 ^ n2862 ;
  assign n2887 = n2886 ^ n2877 ^ n2876 ;
  assign n2897 = n2896 ^ n2895 ^ n2887 ;
  assign n2933 = n2932 ^ n2897 ^ 1'b0 ;
  assign n2854 = ( n2793 & n2837 ) | ( n2793 & n2841 ) | ( n2837 & n2841 ) ;
  assign n2934 = n2933 ^ n2854 ^ 1'b0 ;
  assign n2844 = n912 | n2741 ;
  assign n2845 = n73 | n2844 ;
  assign n2846 = ( n975 & n1904 ) | ( n975 & ~n2845 ) | ( n1904 & ~n2845 ) ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = ( n372 & n401 ) | ( n372 & ~n2847 ) | ( n401 & ~n2847 ) ;
  assign n2849 = n2847 | n2848 ;
  assign n2850 = ( n174 & n2429 ) | ( n174 & ~n2849 ) | ( n2429 & ~n2849 ) ;
  assign n2851 = n2849 | n2850 ;
  assign n2852 = ( n240 & n288 ) | ( n240 & ~n2851 ) | ( n288 & ~n2851 ) ;
  assign n2853 = n2851 | n2852 ;
  assign n2936 = n2935 ^ n2934 ^ n2853 ;
  assign n2843 = n2842 ^ n2771 ^ n2735 ;
  assign n2937 = n2936 ^ n2843 ^ 1'b0 ;
  assign n3039 = n2843 & n2936 ;
  assign n3037 = ( n2853 & n2934 ) | ( n2853 & n2935 ) | ( n2934 & n2935 ) ;
  assign n3004 = n2423 & ~n2923 ;
  assign n3005 = n2459 & n2782 ;
  assign n3006 = n3004 | n3005 ;
  assign n3008 = n332 | n1961 ;
  assign n3009 = ( n509 & n604 ) | ( n509 & ~n3008 ) | ( n604 & ~n3008 ) ;
  assign n3010 = n3008 | n3009 ;
  assign n3011 = ( n325 & n404 ) | ( n325 & ~n3010 ) | ( n404 & ~n3010 ) ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = ( n138 & n475 ) | ( n138 & ~n3012 ) | ( n475 & ~n3012 ) ;
  assign n3014 = n3012 | n3013 ;
  assign n3015 = n302 | n458 ;
  assign n3016 = ( n568 & n991 ) | ( n568 & ~n3015 ) | ( n991 & ~n3015 ) ;
  assign n3017 = ~n568 & n3016 ;
  assign n3018 = ~n3014 & n3017 ;
  assign n3019 = ( ~n298 & n668 ) | ( ~n298 & n3018 ) | ( n668 & n3018 ) ;
  assign n3020 = ~n668 & n3019 ;
  assign n3021 = ( ~n175 & n212 ) | ( ~n175 & n3020 ) | ( n212 & n3020 ) ;
  assign n3022 = ~n212 & n3021 ;
  assign n3023 = ( ~n146 & n399 ) | ( ~n146 & n3022 ) | ( n399 & n3022 ) ;
  assign n3024 = ~n399 & n3023 ;
  assign n3007 = n2921 & ~n2922 ;
  assign n3025 = n3024 ^ n3007 ^ n2921 ;
  assign n3026 = ~n3006 & n3025 ;
  assign n3027 = ( n2422 & n3006 ) | ( n2422 & ~n3026 ) | ( n3006 & ~n3026 ) ;
  assign n3028 = n3027 ^ n2478 ^ 1'b0 ;
  assign n3030 = ( n2782 & ~n2923 ) | ( n2782 & n2927 ) | ( ~n2923 & n2927 ) ;
  assign n3029 = n3025 ^ n2923 ^ 1'b0 ;
  assign n3031 = n3030 ^ n3029 ^ 1'b0 ;
  assign n3032 = ( n2478 & ~n3028 ) | ( n2478 & n3031 ) | ( ~n3028 & n3031 ) ;
  assign n3033 = ( n3027 & n3028 ) | ( n3027 & n3032 ) | ( n3028 & n3032 ) ;
  assign n3034 = n3033 ^ n539 ^ n537 ;
  assign n3002 = ( n2887 & n2895 ) | ( n2887 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2994 = n2198 & n2696 ;
  assign n2995 = n2203 & ~n2475 ;
  assign n2996 = n2201 & n2457 ;
  assign n2997 = ( ~n2994 & n2995 ) | ( ~n2994 & n2996 ) | ( n2995 & n2996 ) ;
  assign n2998 = n2994 | n2997 ;
  assign n2999 = n2703 & ~n2998 ;
  assign n3000 = ( n2275 & n2998 ) | ( n2275 & ~n2999 ) | ( n2998 & ~n2999 ) ;
  assign n3001 = n3000 ^ n536 ^ x5 ;
  assign n2984 = n1943 & ~n2413 ;
  assign n2985 = n2984 ^ n548 ^ 1'b0 ;
  assign n2986 = n2066 & n2406 ;
  assign n2987 = n2068 & ~n2272 ;
  assign n2988 = n2071 & n2242 ;
  assign n2989 = ( ~n2986 & n2987 ) | ( ~n2986 & n2988 ) | ( n2987 & n2988 ) ;
  assign n2990 = n2986 | n2989 ;
  assign n2991 = n2990 ^ n548 ^ 1'b0 ;
  assign n2992 = ( ~n548 & n2985 ) | ( ~n548 & n2991 ) | ( n2985 & n2991 ) ;
  assign n2983 = ( n2876 & n2877 ) | ( n2876 & n2886 ) | ( n2877 & n2886 ) ;
  assign n2981 = ( n2862 & n2874 ) | ( n2862 & n2875 ) | ( n2874 & n2875 ) ;
  assign n2976 = n2863 & n2873 ;
  assign n2977 = n218 & ~n1622 ;
  assign n2978 = n2872 | n2977 ;
  assign n2979 = ( ~n2872 & n2976 ) | ( ~n2872 & n2978 ) | ( n2976 & n2978 ) ;
  assign n2967 = n1635 & n1928 ;
  assign n2968 = n1633 & n1751 ;
  assign n2969 = n1630 & n1846 ;
  assign n2970 = ( ~n2967 & n2968 ) | ( ~n2967 & n2969 ) | ( n2968 & n2969 ) ;
  assign n2971 = n2967 | n2970 ;
  assign n2972 = n2971 ^ n231 ^ 1'b0 ;
  assign n2973 = ( ~n231 & n1936 ) | ( ~n231 & n2972 ) | ( n1936 & n2972 ) ;
  assign n2974 = ( n231 & n2971 ) | ( n231 & n2973 ) | ( n2971 & n2973 ) ;
  assign n2966 = n218 & ~n1620 ;
  assign n2975 = n2974 ^ n2966 ^ 1'b0 ;
  assign n2980 = n2979 ^ n2975 ^ 1'b0 ;
  assign n2957 = n1672 & n2185 ;
  assign n2958 = n1753 & n2059 ;
  assign n2959 = n1670 & ~n2060 ;
  assign n2960 = ( ~n2957 & n2958 ) | ( ~n2957 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2961 = n2957 | n2960 ;
  assign n2962 = n2961 ^ n1757 ^ 1'b0 ;
  assign n2963 = ( ~n1757 & n2186 ) | ( ~n1757 & n2962 ) | ( n2186 & n2962 ) ;
  assign n2964 = ( n1757 & n2961 ) | ( n1757 & n2963 ) | ( n2961 & n2963 ) ;
  assign n2965 = n2964 ^ n219 ^ x11 ;
  assign n2982 = n2981 ^ n2980 ^ n2965 ;
  assign n2993 = n2992 ^ n2983 ^ n2982 ;
  assign n3003 = n3002 ^ n3001 ^ n2993 ;
  assign n3035 = n3034 ^ n3003 ^ 1'b0 ;
  assign n2956 = ( n2854 & n2897 ) | ( n2854 & n2932 ) | ( n2897 & n2932 ) ;
  assign n3036 = n3035 ^ n2956 ^ 1'b0 ;
  assign n2940 = n362 | n1832 ;
  assign n2941 = ( n1960 & n2751 ) | ( n1960 & ~n2940 ) | ( n2751 & ~n2940 ) ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n124 | n381 ;
  assign n2944 = ( n284 & n564 ) | ( n284 & ~n2943 ) | ( n564 & ~n2943 ) ;
  assign n2945 = n2943 | n2944 ;
  assign n2946 = ( n604 & ~n2942 ) | ( n604 & n2945 ) | ( ~n2942 & n2945 ) ;
  assign n2947 = n2942 | n2946 ;
  assign n2948 = ( n2429 & n2434 ) | ( n2429 & ~n2947 ) | ( n2434 & ~n2947 ) ;
  assign n2949 = n2947 | n2948 ;
  assign n2950 = ( n158 & n243 ) | ( n158 & ~n2949 ) | ( n243 & ~n2949 ) ;
  assign n2951 = n2949 | n2950 ;
  assign n2952 = ( n199 & n423 ) | ( n199 & ~n2951 ) | ( n423 & ~n2951 ) ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = ( n178 & n325 ) | ( n178 & ~n2953 ) | ( n325 & ~n2953 ) ;
  assign n2955 = n2953 | n2954 ;
  assign n3038 = n3037 ^ n3036 ^ n2955 ;
  assign n3040 = n3039 ^ n3038 ^ 1'b0 ;
  assign n2938 = x23 ^ x22 ^ 1'b0 ;
  assign n2939 = n2937 & n2938 ;
  assign n3041 = n3040 ^ n2939 ^ 1'b0 ;
  assign n3123 = n3038 & n3039 ;
  assign n3121 = ( n2955 & n3036 ) | ( n2955 & n3037 ) | ( n3036 & n3037 ) ;
  assign n3105 = n194 | n2253 ;
  assign n3106 = ( n258 & n304 ) | ( n258 & ~n3105 ) | ( n304 & ~n3105 ) ;
  assign n3107 = n3105 | n3106 ;
  assign n3108 = ( n116 & n253 ) | ( n116 & ~n3107 ) | ( n253 & ~n3107 ) ;
  assign n3109 = n3107 | n3108 ;
  assign n3110 = n320 | n420 ;
  assign n3111 = n586 | n3110 ;
  assign n3112 = n3109 | n3111 ;
  assign n3113 = ( n105 & n2718 ) | ( n105 & ~n3112 ) | ( n2718 & ~n3112 ) ;
  assign n3114 = n3112 | n3113 ;
  assign n3115 = ( n144 & n161 ) | ( n144 & ~n3114 ) | ( n161 & ~n3114 ) ;
  assign n3116 = n3114 | n3115 ;
  assign n3117 = ( n188 & n203 ) | ( n188 & ~n3116 ) | ( n203 & ~n3116 ) ;
  assign n3118 = n3116 | n3117 ;
  assign n3119 = ( n84 & n399 ) | ( n84 & ~n3118 ) | ( n399 & ~n3118 ) ;
  assign n3120 = n3118 | n3119 ;
  assign n3103 = ( n2956 & n3003 ) | ( n2956 & n3034 ) | ( n3003 & n3034 ) ;
  assign n3091 = n3029 & n3030 ;
  assign n3092 = n2923 & ~n3091 ;
  assign n3093 = n3025 | n3092 ;
  assign n3094 = n3025 & ~n3091 ;
  assign n3095 = n3093 & ~n3094 ;
  assign n3096 = n2478 & n3095 ;
  assign n3097 = n2423 & ~n3025 ;
  assign n3098 = n2459 & ~n2923 ;
  assign n3099 = ( ~n3096 & n3097 ) | ( ~n3096 & n3098 ) | ( n3097 & n3098 ) ;
  assign n3100 = n3096 | n3099 ;
  assign n3101 = n3100 ^ n539 ^ n537 ;
  assign n3089 = ( n2993 & n3001 ) | ( n2993 & n3002 ) | ( n3001 & n3002 ) ;
  assign n3080 = n2198 & n2782 ;
  assign n3081 = n2201 & ~n2475 ;
  assign n3082 = n2203 & n2696 ;
  assign n3083 = ( ~n3080 & n3081 ) | ( ~n3080 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = n3080 | n3083 ;
  assign n3085 = n3084 ^ n2275 ^ 1'b0 ;
  assign n3086 = ( ~n2275 & n2790 ) | ( ~n2275 & n3085 ) | ( n2790 & n3085 ) ;
  assign n3087 = ( n2275 & n3084 ) | ( n2275 & n3086 ) | ( n3084 & n3086 ) ;
  assign n3088 = n3087 ^ n536 ^ x5 ;
  assign n3070 = n1943 & n2492 ;
  assign n3071 = n3070 ^ n548 ^ 1'b0 ;
  assign n3072 = n2066 & n2457 ;
  assign n3073 = n2068 & n2406 ;
  assign n3074 = n2071 & ~n2272 ;
  assign n3075 = ( ~n3072 & n3073 ) | ( ~n3072 & n3074 ) | ( n3073 & n3074 ) ;
  assign n3076 = n3072 | n3075 ;
  assign n3077 = n3076 ^ n548 ^ 1'b0 ;
  assign n3078 = ( ~n548 & n3071 ) | ( ~n548 & n3077 ) | ( n3071 & n3077 ) ;
  assign n3069 = ( n2982 & n2983 ) | ( n2982 & n2992 ) | ( n2983 & n2992 ) ;
  assign n3067 = ( n2965 & n2980 ) | ( n2965 & n2981 ) | ( n2980 & n2981 ) ;
  assign n3062 = n2975 & n2979 ;
  assign n3063 = n218 & ~n2974 ;
  assign n3064 = n1620 & n3063 ;
  assign n3065 = n3062 | n3064 ;
  assign n3054 = n1635 & ~n2060 ;
  assign n3055 = n1633 & n1846 ;
  assign n3056 = n1630 & n1928 ;
  assign n3057 = ( ~n3054 & n3055 ) | ( ~n3054 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3058 = n3054 | n3057 ;
  assign n3059 = n2077 & ~n3058 ;
  assign n3060 = ( n231 & n3058 ) | ( n231 & ~n3059 ) | ( n3058 & ~n3059 ) ;
  assign n3053 = n218 & ~n1751 ;
  assign n3061 = n3060 ^ n3053 ^ 1'b0 ;
  assign n3066 = n3065 ^ n3061 ^ 1'b0 ;
  assign n3044 = n1672 & n2242 ;
  assign n3045 = n1753 & n2185 ;
  assign n3046 = n1670 & n2059 ;
  assign n3047 = ( ~n3044 & n3045 ) | ( ~n3044 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3048 = n3044 | n3047 ;
  assign n3049 = n3048 ^ n1757 ^ 1'b0 ;
  assign n3050 = ( ~n1757 & n2290 ) | ( ~n1757 & n3049 ) | ( n2290 & n3049 ) ;
  assign n3051 = ( n1757 & n3048 ) | ( n1757 & n3050 ) | ( n3048 & n3050 ) ;
  assign n3052 = n3051 ^ n219 ^ x11 ;
  assign n3068 = n3067 ^ n3066 ^ n3052 ;
  assign n3079 = n3078 ^ n3069 ^ n3068 ;
  assign n3090 = n3089 ^ n3088 ^ n3079 ;
  assign n3102 = n3101 ^ n3090 ^ 1'b0 ;
  assign n3104 = n3103 ^ n3102 ^ 1'b0 ;
  assign n3122 = n3121 ^ n3120 ^ n3104 ;
  assign n3124 = n3123 ^ n3122 ^ 1'b0 ;
  assign n3042 = n2937 | n3040 ;
  assign n3043 = n2938 & n3042 ;
  assign n3125 = n3124 ^ n3043 ^ 1'b0 ;
  assign n3197 = n3122 & n3123 ;
  assign n3183 = n96 | n1832 ;
  assign n3184 = ( n750 & n799 ) | ( n750 & ~n3183 ) | ( n799 & ~n3183 ) ;
  assign n3185 = n3183 | n3184 ;
  assign n3186 = ( n983 & n1949 ) | ( n983 & ~n3185 ) | ( n1949 & ~n3185 ) ;
  assign n3187 = n3185 | n3186 ;
  assign n3188 = ( n487 & n629 ) | ( n487 & ~n3187 ) | ( n629 & ~n3187 ) ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = ( n158 & n303 ) | ( n158 & ~n3189 ) | ( n303 & ~n3189 ) ;
  assign n3191 = n3189 | n3190 ;
  assign n3192 = ( n148 & n263 ) | ( n148 & ~n3191 ) | ( n263 & ~n3191 ) ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = ( n232 & n564 ) | ( n232 & ~n3193 ) | ( n564 & ~n3193 ) ;
  assign n3195 = n3193 | n3194 ;
  assign n3181 = ( n3090 & n3101 ) | ( n3090 & n3103 ) | ( n3101 & n3103 ) ;
  assign n3129 = ( n3079 & n3088 ) | ( n3079 & n3089 ) | ( n3088 & n3089 ) ;
  assign n3173 = n2478 & ~n3093 ;
  assign n3174 = n2459 & ~n3025 ;
  assign n3175 = n3173 | n3174 ;
  assign n3176 = n3175 ^ n539 ^ n537 ;
  assign n3165 = n2203 & n2782 ;
  assign n3166 = n2201 & n2696 ;
  assign n3167 = n3165 | n3166 ;
  assign n3168 = n2923 & ~n3167 ;
  assign n3169 = ( n2198 & n3167 ) | ( n2198 & ~n3168 ) | ( n3167 & ~n3168 ) ;
  assign n3170 = n2928 & ~n3169 ;
  assign n3171 = ( n2275 & n3169 ) | ( n2275 & ~n3170 ) | ( n3169 & ~n3170 ) ;
  assign n3172 = n3171 ^ n536 ^ x5 ;
  assign n3155 = n1943 & ~n2481 ;
  assign n3156 = n3155 ^ n548 ^ 1'b0 ;
  assign n3157 = n2068 & n2457 ;
  assign n3158 = n2071 & n2406 ;
  assign n3159 = n3157 | n3158 ;
  assign n3160 = n2475 & ~n3159 ;
  assign n3161 = ( n2066 & n3159 ) | ( n2066 & ~n3160 ) | ( n3159 & ~n3160 ) ;
  assign n3162 = n3161 ^ n548 ^ 1'b0 ;
  assign n3163 = ( ~n548 & n3156 ) | ( ~n548 & n3162 ) | ( n3156 & n3162 ) ;
  assign n3154 = ( n3068 & n3069 ) | ( n3068 & n3078 ) | ( n3069 & n3078 ) ;
  assign n3152 = ( n3052 & n3066 ) | ( n3052 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3147 = n3061 & n3065 ;
  assign n3148 = n218 & ~n3060 ;
  assign n3149 = n1751 & n3148 ;
  assign n3150 = n3147 | n3149 ;
  assign n3139 = n1635 & n2059 ;
  assign n3140 = n1633 & n1928 ;
  assign n3141 = n1630 & ~n2060 ;
  assign n3142 = ( ~n3139 & n3140 ) | ( ~n3139 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3143 = n3139 | n3142 ;
  assign n3144 = n2063 & ~n3143 ;
  assign n3145 = ( n231 & n3143 ) | ( n231 & ~n3144 ) | ( n3143 & ~n3144 ) ;
  assign n3138 = n218 & ~n1846 ;
  assign n3146 = n3145 ^ n3138 ^ 1'b0 ;
  assign n3151 = n3150 ^ n3146 ^ 1'b0 ;
  assign n3130 = n1672 & ~n2272 ;
  assign n3131 = n1753 & n2242 ;
  assign n3132 = n1670 & n2185 ;
  assign n3133 = ( ~n3130 & n3131 ) | ( ~n3130 & n3132 ) | ( n3131 & n3132 ) ;
  assign n3134 = n3130 | n3133 ;
  assign n3135 = n2279 & ~n3134 ;
  assign n3136 = ( n1757 & n3134 ) | ( n1757 & ~n3135 ) | ( n3134 & ~n3135 ) ;
  assign n3137 = n3136 ^ n219 ^ x11 ;
  assign n3153 = n3152 ^ n3151 ^ n3137 ;
  assign n3164 = n3163 ^ n3154 ^ n3153 ;
  assign n3177 = n3176 ^ n3172 ^ n3164 ;
  assign n3178 = n3129 & n3177 ;
  assign n3179 = n3129 | n3177 ;
  assign n3180 = ~n3178 & n3179 ;
  assign n3182 = n3181 ^ n3180 ^ 1'b0 ;
  assign n3128 = ( n3104 & n3120 ) | ( n3104 & ~n3122 ) | ( n3120 & ~n3122 ) ;
  assign n3196 = n3195 ^ n3182 ^ n3128 ;
  assign n3198 = n3197 ^ n3196 ^ 1'b0 ;
  assign n3126 = n3042 | n3124 ;
  assign n3127 = n2938 & n3126 ;
  assign n3199 = n3198 ^ n3127 ^ 1'b0 ;
  assign n3268 = n3196 & n3197 ;
  assign n3266 = ( n3128 & n3182 ) | ( n3128 & n3195 ) | ( n3182 & n3195 ) ;
  assign n3256 = n753 | n2253 ;
  assign n3257 = n560 | n3256 ;
  assign n3258 = ( n704 & n1508 ) | ( n704 & ~n3257 ) | ( n1508 & ~n3257 ) ;
  assign n3259 = n3257 | n3258 ;
  assign n3260 = ( n361 & n645 ) | ( n361 & ~n3259 ) | ( n645 & ~n3259 ) ;
  assign n3261 = n3259 | n3260 ;
  assign n3262 = ( n261 & n347 ) | ( n261 & ~n3261 ) | ( n347 & ~n3261 ) ;
  assign n3263 = n3261 | n3262 ;
  assign n3264 = ( n389 & n437 ) | ( n389 & ~n3263 ) | ( n437 & ~n3263 ) ;
  assign n3265 = n3263 | n3264 ;
  assign n3254 = ( n3129 & n3177 ) | ( n3129 & n3181 ) | ( n3177 & n3181 ) ;
  assign n3202 = ( n3164 & n3172 ) | ( n3164 & n3176 ) | ( n3172 & n3176 ) ;
  assign n3249 = ( n3153 & n3154 ) | ( n3153 & n3163 ) | ( n3154 & n3163 ) ;
  assign n3240 = n2203 & ~n2923 ;
  assign n3241 = n2201 & n2782 ;
  assign n3242 = n3240 | n3241 ;
  assign n3243 = n3025 & ~n3242 ;
  assign n3244 = ( n2198 & n3242 ) | ( n2198 & ~n3243 ) | ( n3242 & ~n3243 ) ;
  assign n3245 = n3244 ^ n2275 ^ 1'b0 ;
  assign n3246 = ( ~n2275 & n3031 ) | ( ~n2275 & n3245 ) | ( n3031 & n3245 ) ;
  assign n3247 = ( n2275 & n3244 ) | ( n2275 & n3246 ) | ( n3244 & n3246 ) ;
  assign n3248 = n3247 ^ n536 ^ x5 ;
  assign n3238 = ( n3137 & n3151 ) | ( n3137 & n3152 ) | ( n3151 & n3152 ) ;
  assign n3229 = n1943 & ~n2703 ;
  assign n3230 = n3229 ^ n548 ^ 1'b0 ;
  assign n3231 = n2066 & n2696 ;
  assign n3232 = n2068 & ~n2475 ;
  assign n3233 = n2071 & n2457 ;
  assign n3234 = ( ~n3231 & n3232 ) | ( ~n3231 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3235 = n3231 | n3234 ;
  assign n3236 = n3235 ^ n548 ^ 1'b0 ;
  assign n3237 = ( ~n548 & n3230 ) | ( ~n548 & n3236 ) | ( n3230 & n3236 ) ;
  assign n3218 = n231 & n2186 ;
  assign n3219 = n3218 ^ n218 ^ 1'b0 ;
  assign n3220 = n1635 & n2185 ;
  assign n3221 = n1633 & ~n2060 ;
  assign n3222 = n1630 & n2059 ;
  assign n3223 = ( ~n3220 & n3221 ) | ( ~n3220 & n3222 ) | ( n3221 & n3222 ) ;
  assign n3224 = n3220 | n3223 ;
  assign n3225 = n3224 ^ n218 ^ 1'b0 ;
  assign n3226 = ( ~n218 & n3219 ) | ( ~n218 & n3225 ) | ( n3219 & n3225 ) ;
  assign n3216 = n218 & n1928 ;
  assign n3217 = n3216 ^ n540 ^ 1'b0 ;
  assign n3227 = n3226 ^ n3217 ^ 1'b0 ;
  assign n3212 = n218 & n1846 ;
  assign n3213 = ~n3145 & n3212 ;
  assign n3214 = n3146 & n3150 ;
  assign n3215 = n3213 | n3214 ;
  assign n3203 = n1672 & n2406 ;
  assign n3204 = n1753 & ~n2272 ;
  assign n3205 = n1670 & n2242 ;
  assign n3206 = ( ~n3203 & n3204 ) | ( ~n3203 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3207 = n3203 | n3206 ;
  assign n3208 = ( n1757 & ~n2413 ) | ( n1757 & n3207 ) | ( ~n2413 & n3207 ) ;
  assign n3209 = n3207 ^ n2413 ^ 1'b0 ;
  assign n3210 = ( n3207 & n3208 ) | ( n3207 & ~n3209 ) | ( n3208 & ~n3209 ) ;
  assign n3211 = n3210 ^ n219 ^ x11 ;
  assign n3228 = n3227 ^ n3215 ^ n3211 ;
  assign n3239 = n3238 ^ n3237 ^ n3228 ;
  assign n3250 = n3249 ^ n3248 ^ n3239 ;
  assign n3251 = n3202 & n3250 ;
  assign n3252 = n3202 | n3250 ;
  assign n3253 = ~n3251 & n3252 ;
  assign n3255 = n3254 ^ n3253 ^ 1'b0 ;
  assign n3267 = n3266 ^ n3265 ^ n3255 ;
  assign n3269 = n3268 ^ n3267 ^ 1'b0 ;
  assign n3200 = n3126 | n3198 ;
  assign n3201 = n2938 & n3200 ;
  assign n3270 = n3269 ^ n3201 ^ 1'b0 ;
  assign n3340 = n3267 & n3268 ;
  assign n3338 = ( n3255 & n3265 ) | ( n3255 & n3266 ) | ( n3265 & n3266 ) ;
  assign n3324 = n113 | n303 ;
  assign n3325 = n296 | n3324 ;
  assign n3326 = n159 | n814 ;
  assign n3327 = n3325 | n3326 ;
  assign n3328 = ( n300 & n1910 ) | ( n300 & ~n3327 ) | ( n1910 & ~n3327 ) ;
  assign n3329 = n3327 | n3328 ;
  assign n3330 = ( n2446 & n3014 ) | ( n2446 & ~n3329 ) | ( n3014 & ~n3329 ) ;
  assign n3331 = n3329 | n3330 ;
  assign n3332 = ( n151 & n2945 ) | ( n151 & ~n3331 ) | ( n2945 & ~n3331 ) ;
  assign n3333 = n3331 | n3332 ;
  assign n3334 = ( n187 & n347 ) | ( n187 & ~n3333 ) | ( n347 & ~n3333 ) ;
  assign n3335 = n3333 | n3334 ;
  assign n3336 = ( n68 & n136 ) | ( n68 & ~n3335 ) | ( n136 & ~n3335 ) ;
  assign n3337 = n3335 | n3336 ;
  assign n3322 = ( n3202 & n3250 ) | ( n3202 & n3254 ) | ( n3250 & n3254 ) ;
  assign n3273 = ( n3239 & n3248 ) | ( n3239 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3317 = ( n3228 & n3237 ) | ( n3228 & n3238 ) | ( n3237 & n3238 ) ;
  assign n3315 = ( n3211 & n3215 ) | ( n3211 & n3227 ) | ( n3215 & n3227 ) ;
  assign n3309 = n218 & n540 ;
  assign n3310 = n1928 & n3309 ;
  assign n3311 = n3217 & n3226 ;
  assign n3312 = n3310 | n3311 ;
  assign n3307 = n218 | n2060 ;
  assign n3308 = n3307 ^ n2060 ^ n540 ;
  assign n3313 = n3312 ^ n3308 ^ 1'b0 ;
  assign n3298 = n231 & n2290 ;
  assign n3299 = n3298 ^ n218 ^ 1'b0 ;
  assign n3300 = n1635 & n2242 ;
  assign n3301 = n1633 & n2059 ;
  assign n3302 = n1630 & n2185 ;
  assign n3303 = ( ~n3300 & n3301 ) | ( ~n3300 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3304 = n3300 | n3303 ;
  assign n3305 = n3304 ^ n218 ^ 1'b0 ;
  assign n3306 = ( ~n218 & n3299 ) | ( ~n218 & n3305 ) | ( n3299 & n3305 ) ;
  assign n3289 = n1672 & n2457 ;
  assign n3290 = n1753 & n2406 ;
  assign n3291 = n1670 & ~n2272 ;
  assign n3292 = ( ~n3289 & n3290 ) | ( ~n3289 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3293 = n3289 | n3292 ;
  assign n3294 = n3293 ^ n1757 ^ 1'b0 ;
  assign n3295 = ( ~n1757 & n2492 ) | ( ~n1757 & n3294 ) | ( n2492 & n3294 ) ;
  assign n3296 = ( n1757 & n3293 ) | ( n1757 & n3295 ) | ( n3293 & n3295 ) ;
  assign n3297 = n3296 ^ n219 ^ x11 ;
  assign n3314 = n3313 ^ n3306 ^ n3297 ;
  assign n3280 = n1943 & n2790 ;
  assign n3281 = n3280 ^ n548 ^ 1'b0 ;
  assign n3282 = n2066 & n2782 ;
  assign n3283 = n2071 & ~n2475 ;
  assign n3284 = n2068 & n2696 ;
  assign n3285 = ( ~n3282 & n3283 ) | ( ~n3282 & n3284 ) | ( n3283 & n3284 ) ;
  assign n3286 = n3282 | n3285 ;
  assign n3287 = n3286 ^ n548 ^ 1'b0 ;
  assign n3288 = ( ~n548 & n3281 ) | ( ~n548 & n3287 ) | ( n3281 & n3287 ) ;
  assign n3316 = n3315 ^ n3314 ^ n3288 ;
  assign n3274 = n2275 & n3095 ;
  assign n3275 = n2203 & ~n3025 ;
  assign n3276 = n2201 & ~n2923 ;
  assign n3277 = ( ~n3274 & n3275 ) | ( ~n3274 & n3276 ) | ( n3275 & n3276 ) ;
  assign n3278 = n3274 | n3277 ;
  assign n3279 = n3278 ^ n536 ^ x5 ;
  assign n3318 = n3317 ^ n3316 ^ n3279 ;
  assign n3319 = n3273 & n3318 ;
  assign n3320 = n3273 | n3318 ;
  assign n3321 = ~n3319 & n3320 ;
  assign n3323 = n3322 ^ n3321 ^ 1'b0 ;
  assign n3339 = n3338 ^ n3337 ^ n3323 ;
  assign n3341 = n3340 ^ n3339 ^ 1'b0 ;
  assign n3271 = n3200 | n3269 ;
  assign n3272 = n2938 & n3271 ;
  assign n3342 = n3341 ^ n3272 ^ 1'b0 ;
  assign n3412 = n3339 & n3340 ;
  assign n3410 = ( n3323 & n3337 ) | ( n3323 & n3338 ) | ( n3337 & n3338 ) ;
  assign n3392 = n126 | n302 ;
  assign n3393 = n434 | n3392 ;
  assign n3394 = ( n265 & n1832 ) | ( n265 & ~n3393 ) | ( n1832 & ~n3393 ) ;
  assign n3395 = n3393 | n3394 ;
  assign n3396 = ( n151 & n244 ) | ( n151 & ~n3395 ) | ( n244 & ~n3395 ) ;
  assign n3397 = n3395 | n3396 ;
  assign n3398 = ( n283 & n668 ) | ( n283 & ~n3397 ) | ( n668 & ~n3397 ) ;
  assign n3399 = n3397 | n3398 ;
  assign n3400 = n267 | n2755 ;
  assign n3401 = ( n1502 & n2693 ) | ( n1502 & ~n3400 ) | ( n2693 & ~n3400 ) ;
  assign n3402 = n3400 | n3401 ;
  assign n3403 = n3399 | n3402 ;
  assign n3404 = ( n102 & n315 ) | ( n102 & ~n3403 ) | ( n315 & ~n3403 ) ;
  assign n3405 = n3403 | n3404 ;
  assign n3406 = ( n404 & n414 ) | ( n404 & ~n3405 ) | ( n414 & ~n3405 ) ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = ( n240 & n273 ) | ( n240 & ~n3407 ) | ( n273 & ~n3407 ) ;
  assign n3409 = n3407 | n3408 ;
  assign n3390 = ( n3273 & n3318 ) | ( n3273 & n3322 ) | ( n3318 & n3322 ) ;
  assign n3345 = ( n3279 & n3316 ) | ( n3279 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3385 = ( n3288 & n3314 ) | ( n3288 & n3315 ) | ( n3314 & n3315 ) ;
  assign n3381 = n2275 & ~n3093 ;
  assign n3382 = n2201 & ~n3025 ;
  assign n3383 = n3381 | n3382 ;
  assign n3384 = n3383 ^ n536 ^ x5 ;
  assign n3371 = n1943 & ~n2928 ;
  assign n3372 = n3371 ^ n548 ^ 1'b0 ;
  assign n3373 = n2068 & n2782 ;
  assign n3374 = n2071 & n2696 ;
  assign n3375 = n3373 | n3374 ;
  assign n3376 = n2923 & ~n3375 ;
  assign n3377 = ( n2066 & n3375 ) | ( n2066 & ~n3376 ) | ( n3375 & ~n3376 ) ;
  assign n3378 = n3377 ^ n548 ^ 1'b0 ;
  assign n3379 = ( ~n548 & n3372 ) | ( ~n548 & n3378 ) | ( n3372 & n3378 ) ;
  assign n3370 = ( n3297 & n3306 ) | ( n3297 & n3313 ) | ( n3306 & n3313 ) ;
  assign n3365 = ~n2060 & n3309 ;
  assign n3366 = n3308 & n3312 ;
  assign n3367 = n3365 | n3366 ;
  assign n3363 = n218 & n2059 ;
  assign n3364 = n3363 ^ n540 ^ 1'b0 ;
  assign n3368 = n3367 ^ n3364 ^ 1'b0 ;
  assign n3354 = n231 & ~n2279 ;
  assign n3355 = n3354 ^ n218 ^ 1'b0 ;
  assign n3356 = n1635 & ~n2272 ;
  assign n3357 = n1633 & n2185 ;
  assign n3358 = n1630 & n2242 ;
  assign n3359 = ( ~n3356 & n3357 ) | ( ~n3356 & n3358 ) | ( n3357 & n3358 ) ;
  assign n3360 = n3356 | n3359 ;
  assign n3361 = n3360 ^ n218 ^ 1'b0 ;
  assign n3362 = ( ~n218 & n3355 ) | ( ~n218 & n3361 ) | ( n3355 & n3361 ) ;
  assign n3346 = n1753 & n2457 ;
  assign n3347 = n1670 & n2406 ;
  assign n3348 = n3346 | n3347 ;
  assign n3349 = n2475 & ~n3348 ;
  assign n3350 = ( n1672 & n3348 ) | ( n1672 & ~n3349 ) | ( n3348 & ~n3349 ) ;
  assign n3351 = n2481 & ~n3350 ;
  assign n3352 = ( n1757 & n3350 ) | ( n1757 & ~n3351 ) | ( n3350 & ~n3351 ) ;
  assign n3353 = n3352 ^ n219 ^ x11 ;
  assign n3369 = n3368 ^ n3362 ^ n3353 ;
  assign n3380 = n3379 ^ n3370 ^ n3369 ;
  assign n3386 = n3385 ^ n3384 ^ n3380 ;
  assign n3387 = n3345 & n3386 ;
  assign n3388 = n3345 | n3386 ;
  assign n3389 = ~n3387 & n3388 ;
  assign n3391 = n3390 ^ n3389 ^ 1'b0 ;
  assign n3411 = n3410 ^ n3409 ^ n3391 ;
  assign n3413 = n3412 ^ n3411 ^ 1'b0 ;
  assign n3343 = n3271 | n3341 ;
  assign n3344 = n2938 & n3343 ;
  assign n3414 = n3413 ^ n3344 ^ 1'b0 ;
  assign n3470 = n3411 & n3412 ;
  assign n3468 = ( n3391 & n3409 ) | ( n3391 & n3410 ) | ( n3409 & n3410 ) ;
  assign n3465 = ( n3380 & n3384 ) | ( n3380 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3463 = ( n3369 & n3370 ) | ( n3369 & n3379 ) | ( n3370 & n3379 ) ;
  assign n3454 = n1943 & n3031 ;
  assign n3455 = n3454 ^ n548 ^ 1'b0 ;
  assign n3456 = n2068 & ~n2923 ;
  assign n3457 = n2071 & n2782 ;
  assign n3458 = n3456 | n3457 ;
  assign n3459 = n3025 & ~n3458 ;
  assign n3460 = ( n2066 & n3458 ) | ( n2066 & ~n3459 ) | ( n3458 & ~n3459 ) ;
  assign n3461 = n3460 ^ n548 ^ 1'b0 ;
  assign n3462 = ( ~n548 & n3455 ) | ( ~n548 & n3461 ) | ( n3455 & n3461 ) ;
  assign n3452 = ( n3353 & n3362 ) | ( n3353 & n3368 ) | ( n3362 & n3368 ) ;
  assign n3444 = n1672 & n2696 ;
  assign n3445 = n1753 & ~n2475 ;
  assign n3446 = n1670 & n2457 ;
  assign n3447 = ( ~n3444 & n3445 ) | ( ~n3444 & n3446 ) | ( n3445 & n3446 ) ;
  assign n3448 = n3444 | n3447 ;
  assign n3449 = n2703 & ~n3448 ;
  assign n3450 = ( n1757 & n3448 ) | ( n1757 & ~n3449 ) | ( n3448 & ~n3449 ) ;
  assign n3451 = n3450 ^ n219 ^ x11 ;
  assign n3440 = n2059 & n3309 ;
  assign n3441 = n3364 & n3367 ;
  assign n3442 = n3440 | n3441 ;
  assign n3431 = n231 & ~n2413 ;
  assign n3432 = n3431 ^ n218 ^ 1'b0 ;
  assign n3433 = n1635 & n2406 ;
  assign n3434 = n1633 & n2242 ;
  assign n3435 = n1630 & ~n2272 ;
  assign n3436 = ( ~n3433 & n3434 ) | ( ~n3433 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3437 = n3433 | n3436 ;
  assign n3438 = n3437 ^ n218 ^ 1'b0 ;
  assign n3439 = ( ~n218 & n3432 ) | ( ~n218 & n3438 ) | ( n3432 & n3438 ) ;
  assign n3429 = n218 & n2185 ;
  assign n3430 = n3429 ^ n542 ^ 1'b0 ;
  assign n3443 = n3442 ^ n3439 ^ n3430 ;
  assign n3453 = n3452 ^ n3451 ^ n3443 ;
  assign n3464 = n3463 ^ n3462 ^ n3453 ;
  assign n3466 = n3465 ^ n3464 ^ 1'b0 ;
  assign n3428 = ( n3345 & n3386 ) | ( n3345 & n3390 ) | ( n3386 & n3390 ) ;
  assign n3467 = n3466 ^ n3428 ^ 1'b0 ;
  assign n3417 = n735 | n1977 ;
  assign n3418 = ( n561 & n3325 ) | ( n561 & ~n3417 ) | ( n3325 & ~n3417 ) ;
  assign n3419 = n3417 | n3418 ;
  assign n3420 = ( n304 & n3399 ) | ( n304 & ~n3419 ) | ( n3399 & ~n3419 ) ;
  assign n3421 = n3419 | n3420 ;
  assign n3422 = ( n193 & n389 ) | ( n193 & ~n3421 ) | ( n389 & ~n3421 ) ;
  assign n3423 = n3421 | n3422 ;
  assign n3424 = ( n445 & n907 ) | ( n445 & ~n3423 ) | ( n907 & ~n3423 ) ;
  assign n3425 = n3423 | n3424 ;
  assign n3426 = ( n178 & n475 ) | ( n178 & ~n3425 ) | ( n475 & ~n3425 ) ;
  assign n3427 = n3425 | n3426 ;
  assign n3469 = n3468 ^ n3467 ^ n3427 ;
  assign n3471 = n3470 ^ n3469 ^ 1'b0 ;
  assign n3415 = n3343 | n3413 ;
  assign n3416 = n2938 & n3415 ;
  assign n3472 = n3471 ^ n3416 ^ 1'b0 ;
  assign n3536 = n3469 & n3470 ;
  assign n3534 = ( n3427 & n3467 ) | ( n3427 & n3468 ) | ( n3467 & n3468 ) ;
  assign n3514 = n691 | n1833 ;
  assign n3515 = ( n190 & n671 ) | ( n190 & ~n3514 ) | ( n671 & ~n3514 ) ;
  assign n3516 = n3514 | n3515 ;
  assign n3517 = n382 | n1545 ;
  assign n3518 = ( n255 & n299 ) | ( n255 & ~n3517 ) | ( n299 & ~n3517 ) ;
  assign n3519 = n3517 | n3518 ;
  assign n3520 = ( n349 & n451 ) | ( n349 & ~n3519 ) | ( n451 & ~n3519 ) ;
  assign n3521 = n3519 | n3520 ;
  assign n3522 = ( n72 & n205 ) | ( n72 & ~n3521 ) | ( n205 & ~n3521 ) ;
  assign n3523 = n3521 | n3522 ;
  assign n3524 = ( n263 & n426 ) | ( n263 & ~n3523 ) | ( n426 & ~n3523 ) ;
  assign n3525 = n3523 | n3524 ;
  assign n3526 = ( n194 & ~n3516 ) | ( n194 & n3525 ) | ( ~n3516 & n3525 ) ;
  assign n3527 = n3516 | n3526 ;
  assign n3528 = ( n235 & n305 ) | ( n235 & ~n3527 ) | ( n305 & ~n3527 ) ;
  assign n3529 = n3527 | n3528 ;
  assign n3530 = ( n284 & n328 ) | ( n284 & ~n3529 ) | ( n328 & ~n3529 ) ;
  assign n3531 = n3529 | n3530 ;
  assign n3532 = ( n266 & n399 ) | ( n266 & ~n3531 ) | ( n399 & ~n3531 ) ;
  assign n3533 = n3531 | n3532 ;
  assign n3512 = ( n3428 & n3464 ) | ( n3428 & n3465 ) | ( n3464 & n3465 ) ;
  assign n3475 = ( n3453 & n3462 ) | ( n3453 & n3463 ) | ( n3462 & n3463 ) ;
  assign n3501 = n1943 & n3095 ;
  assign n3502 = n3501 ^ n548 ^ 1'b0 ;
  assign n3503 = n2068 & ~n3025 ;
  assign n3504 = n2071 & ~n2923 ;
  assign n3505 = n3503 | n3504 ;
  assign n3506 = n3505 ^ n548 ^ 1'b0 ;
  assign n3507 = ( ~n548 & n3502 ) | ( ~n548 & n3506 ) | ( n3502 & n3506 ) ;
  assign n3500 = ( n3443 & n3451 ) | ( n3443 & n3452 ) | ( n3451 & n3452 ) ;
  assign n3498 = ( n3430 & n3439 ) | ( n3430 & n3442 ) | ( n3439 & n3442 ) ;
  assign n3495 = n218 & n2242 ;
  assign n3494 = ( n540 & n541 ) | ( n540 & ~n3429 ) | ( n541 & ~n3429 ) ;
  assign n3496 = n3495 ^ n3494 ^ 1'b0 ;
  assign n3485 = n231 & n2492 ;
  assign n3486 = n3485 ^ n218 ^ 1'b0 ;
  assign n3487 = n1635 & n2457 ;
  assign n3488 = n1633 & ~n2272 ;
  assign n3489 = n1630 & n2406 ;
  assign n3490 = ( ~n3487 & n3488 ) | ( ~n3487 & n3489 ) | ( n3488 & n3489 ) ;
  assign n3491 = n3487 | n3490 ;
  assign n3492 = n3491 ^ n218 ^ 1'b0 ;
  assign n3493 = ( ~n218 & n3486 ) | ( ~n218 & n3492 ) | ( n3486 & n3492 ) ;
  assign n3497 = n3496 ^ n3493 ^ 1'b0 ;
  assign n3476 = n1672 & n2782 ;
  assign n3477 = n1670 & ~n2475 ;
  assign n3478 = n1753 & n2696 ;
  assign n3479 = ( ~n3476 & n3477 ) | ( ~n3476 & n3478 ) | ( n3477 & n3478 ) ;
  assign n3480 = n3476 | n3479 ;
  assign n3481 = n3480 ^ n1757 ^ 1'b0 ;
  assign n3482 = ( ~n1757 & n2790 ) | ( ~n1757 & n3481 ) | ( n2790 & n3481 ) ;
  assign n3483 = ( n1757 & n3480 ) | ( n1757 & n3482 ) | ( n3480 & n3482 ) ;
  assign n3484 = n3483 ^ n219 ^ x11 ;
  assign n3499 = n3498 ^ n3497 ^ n3484 ;
  assign n3508 = n3507 ^ n3500 ^ n3499 ;
  assign n3509 = n3475 & n3508 ;
  assign n3510 = n3475 | n3508 ;
  assign n3511 = ~n3509 & n3510 ;
  assign n3513 = n3512 ^ n3511 ^ 1'b0 ;
  assign n3535 = n3534 ^ n3533 ^ n3513 ;
  assign n3537 = n3536 ^ n3535 ^ 1'b0 ;
  assign n3473 = n3415 | n3471 ;
  assign n3474 = n2938 & n3473 ;
  assign n3538 = n3537 ^ n3474 ^ 1'b0 ;
  assign n3587 = n3535 & n3536 ;
  assign n3585 = ( n3513 & n3533 ) | ( n3513 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3573 = n561 | n598 ;
  assign n3574 = n2761 | n3573 ;
  assign n3575 = ( n298 & n2434 ) | ( n298 & ~n3574 ) | ( n2434 & ~n3574 ) ;
  assign n3576 = n3574 | n3575 ;
  assign n3577 = ( n315 & n2693 ) | ( n315 & ~n3576 ) | ( n2693 & ~n3576 ) ;
  assign n3578 = n3576 | n3577 ;
  assign n3579 = ( n72 & n199 ) | ( n72 & ~n3578 ) | ( n199 & ~n3578 ) ;
  assign n3580 = n3578 | n3579 ;
  assign n3581 = ( n111 & n462 ) | ( n111 & ~n3580 ) | ( n462 & ~n3580 ) ;
  assign n3582 = n3580 | n3581 ;
  assign n3583 = ( n142 & n379 ) | ( n142 & ~n3582 ) | ( n379 & ~n3582 ) ;
  assign n3584 = n3582 | n3583 ;
  assign n3570 = ( n3499 & n3500 ) | ( n3499 & n3507 ) | ( n3500 & n3507 ) ;
  assign n3568 = ( n3484 & n3497 ) | ( n3484 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3563 = n2071 & ~n3025 ;
  assign n3564 = n3563 ^ n548 ^ 1'b0 ;
  assign n3565 = n1943 & ~n3093 ;
  assign n3566 = n3565 ^ n548 ^ 1'b0 ;
  assign n3567 = ( ~n548 & n3564 ) | ( ~n548 & n3566 ) | ( n3564 & n3566 ) ;
  assign n3561 = ( ~n3493 & n3494 ) | ( ~n3493 & n3495 ) | ( n3494 & n3495 ) ;
  assign n3551 = n231 & ~n2481 ;
  assign n3552 = n3551 ^ n218 ^ 1'b0 ;
  assign n3553 = n1630 & n2457 ;
  assign n3554 = n1633 & n2406 ;
  assign n3555 = n3553 | n3554 ;
  assign n3556 = n2475 & ~n3555 ;
  assign n3557 = ( n1635 & n3555 ) | ( n1635 & ~n3556 ) | ( n3555 & ~n3556 ) ;
  assign n3558 = n3557 ^ n218 ^ 1'b0 ;
  assign n3559 = ( ~n218 & n3552 ) | ( ~n218 & n3558 ) | ( n3552 & n3558 ) ;
  assign n3550 = n218 & ~n2276 ;
  assign n3560 = n3559 ^ n3550 ^ 1'b0 ;
  assign n3542 = n1753 & n2782 ;
  assign n3543 = n1670 & n2696 ;
  assign n3544 = n3542 | n3543 ;
  assign n3545 = n2923 & ~n3544 ;
  assign n3546 = ( n1672 & n3544 ) | ( n1672 & ~n3545 ) | ( n3544 & ~n3545 ) ;
  assign n3547 = n2928 & ~n3546 ;
  assign n3548 = ( n1757 & n3546 ) | ( n1757 & ~n3547 ) | ( n3546 & ~n3547 ) ;
  assign n3549 = n3548 ^ n219 ^ x11 ;
  assign n3562 = n3561 ^ n3560 ^ n3549 ;
  assign n3569 = n3568 ^ n3567 ^ n3562 ;
  assign n3571 = n3570 ^ n3569 ^ 1'b0 ;
  assign n3541 = ( n3475 & n3508 ) | ( n3475 & n3512 ) | ( n3508 & n3512 ) ;
  assign n3572 = n3571 ^ n3541 ^ 1'b0 ;
  assign n3586 = n3585 ^ n3584 ^ n3572 ;
  assign n3588 = n3587 ^ n3586 ^ 1'b0 ;
  assign n3539 = n3473 | n3537 ;
  assign n3540 = n2938 & n3539 ;
  assign n3589 = n3588 ^ n3540 ^ 1'b0 ;
  assign n3635 = n3586 & n3587 ;
  assign n3633 = ( n3572 & n3584 ) | ( n3572 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3622 = n358 | n2252 ;
  assign n3623 = ( n145 & n492 ) | ( n145 & ~n3622 ) | ( n492 & ~n3622 ) ;
  assign n3624 = n3622 | n3623 ;
  assign n3625 = ( n120 & n2429 ) | ( n120 & ~n3624 ) | ( n2429 & ~n3624 ) ;
  assign n3626 = n3624 | n3625 ;
  assign n3627 = ( n920 & n2693 ) | ( n920 & ~n3626 ) | ( n2693 & ~n3626 ) ;
  assign n3628 = n3626 | n3627 ;
  assign n3629 = ( n309 & n669 ) | ( n309 & ~n3628 ) | ( n669 & ~n3628 ) ;
  assign n3630 = n3628 | n3629 ;
  assign n3631 = ( n301 & n484 ) | ( n301 & ~n3630 ) | ( n484 & ~n3630 ) ;
  assign n3632 = n3630 | n3631 ;
  assign n3620 = ( n3541 & n3569 ) | ( n3541 & n3570 ) | ( n3569 & n3570 ) ;
  assign n3618 = ( n3562 & n3567 ) | ( n3562 & n3568 ) | ( n3567 & n3568 ) ;
  assign n3613 = n2272 | n3495 ;
  assign n3614 = n218 & ~n3613 ;
  assign n3615 = n3550 & ~n3614 ;
  assign n3616 = ( n3559 & n3614 ) | ( n3559 & ~n3615 ) | ( n3614 & ~n3615 ) ;
  assign n3611 = n218 & n2406 ;
  assign n3612 = n3611 ^ n3495 ^ n548 ;
  assign n3602 = n231 & ~n2703 ;
  assign n3603 = n3602 ^ n218 ^ 1'b0 ;
  assign n3604 = n1635 & n2696 ;
  assign n3605 = n1630 & ~n2475 ;
  assign n3606 = n1633 & n2457 ;
  assign n3607 = ( ~n3604 & n3605 ) | ( ~n3604 & n3606 ) | ( n3605 & n3606 ) ;
  assign n3608 = n3604 | n3607 ;
  assign n3609 = n3608 ^ n218 ^ 1'b0 ;
  assign n3610 = ( ~n218 & n3603 ) | ( ~n218 & n3609 ) | ( n3603 & n3609 ) ;
  assign n3617 = n3616 ^ n3612 ^ n3610 ;
  assign n3600 = ( ~n3549 & n3560 ) | ( ~n3549 & n3561 ) | ( n3560 & n3561 ) ;
  assign n3592 = n1753 & ~n2923 ;
  assign n3593 = n1670 & n2782 ;
  assign n3594 = n3592 | n3593 ;
  assign n3595 = n3025 & ~n3594 ;
  assign n3596 = ( n1672 & n3594 ) | ( n1672 & ~n3595 ) | ( n3594 & ~n3595 ) ;
  assign n3597 = n3596 ^ n1757 ^ 1'b0 ;
  assign n3598 = ( ~n1757 & n3031 ) | ( ~n1757 & n3597 ) | ( n3031 & n3597 ) ;
  assign n3599 = ( n1757 & n3596 ) | ( n1757 & n3598 ) | ( n3596 & n3598 ) ;
  assign n3601 = n3600 ^ n3599 ^ n220 ;
  assign n3619 = n3618 ^ n3617 ^ n3601 ;
  assign n3621 = n3620 ^ n3619 ^ 1'b0 ;
  assign n3634 = n3633 ^ n3632 ^ n3621 ;
  assign n3636 = n3635 ^ n3634 ^ 1'b0 ;
  assign n3590 = n3539 | n3588 ;
  assign n3591 = n2938 & n3590 ;
  assign n3637 = n3636 ^ n3591 ^ 1'b0 ;
  assign n3675 = n3634 & n3635 ;
  assign n3673 = ( n3621 & n3632 ) | ( n3621 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3667 = n699 | n717 ;
  assign n3668 = n783 | n3667 ;
  assign n3669 = ( n428 & n2907 ) | ( n428 & ~n3668 ) | ( n2907 & ~n3668 ) ;
  assign n3670 = n3668 | n3669 ;
  assign n3671 = ( n125 & n520 ) | ( n125 & ~n3670 ) | ( n520 & ~n3670 ) ;
  assign n3672 = n3670 | n3671 ;
  assign n3664 = n3617 ^ n3601 ^ 1'b0 ;
  assign n3665 = ( n3618 & n3620 ) | ( n3618 & n3664 ) | ( n3620 & n3664 ) ;
  assign n3661 = n3599 ^ n219 ^ x11 ;
  assign n3662 = ( n3600 & n3617 ) | ( n3600 & ~n3661 ) | ( n3617 & ~n3661 ) ;
  assign n3659 = ( n3610 & ~n3612 ) | ( n3610 & n3616 ) | ( ~n3612 & n3616 ) ;
  assign n3656 = n218 & n2457 ;
  assign n3655 = ( n3495 & n3611 ) | ( n3495 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3657 = n3656 ^ n3655 ^ 1'b0 ;
  assign n3646 = n231 & n2790 ;
  assign n3647 = n3646 ^ n218 ^ 1'b0 ;
  assign n3648 = n1635 & n2782 ;
  assign n3649 = n1633 & ~n2475 ;
  assign n3650 = n1630 & n2696 ;
  assign n3651 = ( ~n3648 & n3649 ) | ( ~n3648 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = n3648 | n3651 ;
  assign n3653 = n3652 ^ n218 ^ 1'b0 ;
  assign n3654 = ( ~n218 & n3647 ) | ( ~n218 & n3653 ) | ( n3647 & n3653 ) ;
  assign n3658 = n3657 ^ n3654 ^ 1'b0 ;
  assign n3640 = n1757 & n3095 ;
  assign n3641 = n1753 & ~n3025 ;
  assign n3642 = n1670 & ~n2923 ;
  assign n3643 = ( ~n3640 & n3641 ) | ( ~n3640 & n3642 ) | ( n3641 & n3642 ) ;
  assign n3644 = n3640 | n3643 ;
  assign n3645 = n3644 ^ n219 ^ x11 ;
  assign n3660 = n3659 ^ n3658 ^ n3645 ;
  assign n3663 = n3662 ^ n3660 ^ 1'b0 ;
  assign n3666 = n3665 ^ n3663 ^ 1'b0 ;
  assign n3674 = n3673 ^ n3672 ^ n3666 ;
  assign n3676 = n3675 ^ n3674 ^ 1'b0 ;
  assign n3638 = n3590 | n3636 ;
  assign n3639 = n2938 & n3638 ;
  assign n3677 = n3676 ^ n3639 ^ 1'b0 ;
  assign n3715 = n3674 & n3675 ;
  assign n3713 = ( n3666 & n3672 ) | ( n3666 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3701 = n107 | n321 ;
  assign n3702 = n305 | n3701 ;
  assign n3703 = ( n209 & n462 ) | ( n209 & ~n3702 ) | ( n462 & ~n3702 ) ;
  assign n3704 = n3702 | n3703 ;
  assign n3705 = n1733 | n3704 ;
  assign n3706 = n750 | n3705 ;
  assign n3707 = ( n2031 & n3109 ) | ( n2031 & ~n3706 ) | ( n3109 & ~n3706 ) ;
  assign n3708 = n3706 | n3707 ;
  assign n3709 = ( n100 & n1727 ) | ( n100 & ~n3708 ) | ( n1727 & ~n3708 ) ;
  assign n3710 = n3708 | n3709 ;
  assign n3711 = ( n250 & n426 ) | ( n250 & ~n3710 ) | ( n426 & ~n3710 ) ;
  assign n3712 = n3710 | n3711 ;
  assign n3699 = ( n3660 & n3662 ) | ( n3660 & ~n3665 ) | ( n3662 & ~n3665 ) ;
  assign n3697 = ( n3645 & ~n3658 ) | ( n3645 & n3659 ) | ( ~n3658 & n3659 ) ;
  assign n3692 = n1757 & ~n3093 ;
  assign n3693 = n1670 & ~n3025 ;
  assign n3694 = n3692 | n3693 ;
  assign n3695 = n3694 ^ n219 ^ x11 ;
  assign n3683 = n231 & ~n2928 ;
  assign n3684 = n3683 ^ n218 ^ 1'b0 ;
  assign n3685 = n1630 & n2782 ;
  assign n3686 = n1633 & n2696 ;
  assign n3687 = n3685 | n3686 ;
  assign n3688 = n2923 & ~n3687 ;
  assign n3689 = ( n1635 & n3687 ) | ( n1635 & ~n3688 ) | ( n3687 & ~n3688 ) ;
  assign n3690 = n3689 ^ n218 ^ 1'b0 ;
  assign n3691 = ( ~n218 & n3684 ) | ( ~n218 & n3690 ) | ( n3684 & n3690 ) ;
  assign n3681 = n218 & ~n2475 ;
  assign n3680 = ( n3654 & n3655 ) | ( n3654 & ~n3656 ) | ( n3655 & ~n3656 ) ;
  assign n3682 = n3681 ^ n3680 ^ n3656 ;
  assign n3696 = n3695 ^ n3691 ^ n3682 ;
  assign n3698 = n3697 ^ n3696 ^ 1'b0 ;
  assign n3700 = n3699 ^ n3698 ^ 1'b0 ;
  assign n3714 = n3713 ^ n3712 ^ n3700 ;
  assign n3716 = n3715 ^ n3714 ^ 1'b0 ;
  assign n3678 = n3638 | n3676 ;
  assign n3679 = n2938 & n3678 ;
  assign n3717 = n3716 ^ n3679 ^ 1'b0 ;
  assign n3756 = n3714 & n3715 ;
  assign n3754 = ( n3700 & n3712 ) | ( n3700 & n3713 ) | ( n3712 & n3713 ) ;
  assign n3737 = n169 | n389 ;
  assign n3738 = n174 | n3737 ;
  assign n3739 = ( n233 & n325 ) | ( n233 & ~n3738 ) | ( n325 & ~n3738 ) ;
  assign n3740 = n3738 | n3739 ;
  assign n3741 = n244 | n3740 ;
  assign n3742 = ( n928 & n2945 ) | ( n928 & ~n3741 ) | ( n2945 & ~n3741 ) ;
  assign n3743 = n3741 | n3742 ;
  assign n3744 = ( n196 & n2220 ) | ( n196 & ~n3743 ) | ( n2220 & ~n3743 ) ;
  assign n3745 = n3743 | n3744 ;
  assign n3746 = ( n367 & n2718 ) | ( n367 & ~n3745 ) | ( n2718 & ~n3745 ) ;
  assign n3747 = n3745 | n3746 ;
  assign n3748 = ( n235 & n376 ) | ( n235 & ~n3747 ) | ( n376 & ~n3747 ) ;
  assign n3749 = n3747 | n3748 ;
  assign n3750 = ( n116 & n404 ) | ( n116 & ~n3749 ) | ( n404 & ~n3749 ) ;
  assign n3751 = n3749 | n3750 ;
  assign n3752 = ( n212 & n331 ) | ( n212 & ~n3751 ) | ( n331 & ~n3751 ) ;
  assign n3753 = n3751 | n3752 ;
  assign n3735 = ( n3696 & ~n3697 ) | ( n3696 & n3699 ) | ( ~n3697 & n3699 ) ;
  assign n3733 = ( ~n3682 & n3691 ) | ( ~n3682 & n3695 ) | ( n3691 & n3695 ) ;
  assign n3731 = ( n3656 & n3680 ) | ( n3656 & ~n3681 ) | ( n3680 & ~n3681 ) ;
  assign n3722 = n231 & n3031 ;
  assign n3723 = n3722 ^ n218 ^ 1'b0 ;
  assign n3724 = n1630 & ~n2923 ;
  assign n3725 = n1633 & n2782 ;
  assign n3726 = n3724 | n3725 ;
  assign n3727 = n3025 & ~n3726 ;
  assign n3728 = ( n1635 & n3726 ) | ( n1635 & ~n3727 ) | ( n3726 & ~n3727 ) ;
  assign n3729 = n3728 ^ n218 ^ 1'b0 ;
  assign n3730 = ( ~n218 & n3723 ) | ( ~n218 & n3729 ) | ( n3723 & n3729 ) ;
  assign n3720 = n218 & n2696 ;
  assign n3721 = n3720 ^ n3681 ^ n220 ;
  assign n3732 = n3731 ^ n3730 ^ n3721 ;
  assign n3734 = n3733 ^ n3732 ^ 1'b0 ;
  assign n3736 = n3735 ^ n3734 ^ 1'b0 ;
  assign n3755 = n3754 ^ n3753 ^ n3736 ;
  assign n3757 = n3756 ^ n3755 ^ 1'b0 ;
  assign n3718 = n3678 | n3716 ;
  assign n3719 = n2938 & n3718 ;
  assign n3758 = n3757 ^ n3719 ^ 1'b0 ;
  assign n3791 = n3755 & n3756 ;
  assign n3776 = n332 | n1733 ;
  assign n3777 = n323 | n3776 ;
  assign n3778 = ( n697 & n1549 ) | ( n697 & ~n3777 ) | ( n1549 & ~n3777 ) ;
  assign n3779 = n3777 | n3778 ;
  assign n3780 = ( n260 & n972 ) | ( n260 & ~n3779 ) | ( n972 & ~n3779 ) ;
  assign n3781 = n3779 | n3780 ;
  assign n3782 = ( n236 & n2693 ) | ( n236 & ~n3781 ) | ( n2693 & ~n3781 ) ;
  assign n3783 = n3781 | n3782 ;
  assign n3784 = ( n149 & n363 ) | ( n149 & ~n3783 ) | ( n363 & ~n3783 ) ;
  assign n3785 = n3783 | n3784 ;
  assign n3786 = ( n148 & n376 ) | ( n148 & ~n3785 ) | ( n376 & ~n3785 ) ;
  assign n3787 = n3785 | n3786 ;
  assign n3788 = ( n84 & n125 ) | ( n84 & ~n3787 ) | ( n125 & ~n3787 ) ;
  assign n3789 = n3787 | n3788 ;
  assign n3774 = ( n3732 & ~n3733 ) | ( n3732 & n3735 ) | ( ~n3733 & n3735 ) ;
  assign n3773 = ( ~n3721 & n3730 ) | ( ~n3721 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3770 = n218 & n2782 ;
  assign n3769 = ( ~n220 & n3681 ) | ( ~n220 & n3720 ) | ( n3681 & n3720 ) ;
  assign n3771 = n3770 ^ n3769 ^ 1'b0 ;
  assign n3762 = n231 & n3095 ;
  assign n3763 = n3762 ^ n218 ^ 1'b0 ;
  assign n3764 = n1630 & ~n3025 ;
  assign n3765 = n1633 & ~n2923 ;
  assign n3766 = n3764 | n3765 ;
  assign n3767 = n3766 ^ n218 ^ 1'b0 ;
  assign n3768 = ( ~n218 & n3763 ) | ( ~n218 & n3767 ) | ( n3763 & n3767 ) ;
  assign n3772 = n3771 ^ n3768 ^ 1'b0 ;
  assign n3775 = n3774 ^ n3773 ^ n3772 ;
  assign n3761 = ( n3736 & n3753 ) | ( n3736 & ~n3755 ) | ( n3753 & ~n3755 ) ;
  assign n3790 = n3789 ^ n3775 ^ n3761 ;
  assign n3792 = n3791 ^ n3790 ^ 1'b0 ;
  assign n3759 = n3718 | n3757 ;
  assign n3760 = n2938 & n3759 ;
  assign n3793 = n3792 ^ n3760 ^ 1'b0 ;
  assign n3823 = n3790 & n3791 ;
  assign n3821 = ( n3761 & n3775 ) | ( n3761 & n3789 ) | ( n3775 & n3789 ) ;
  assign n3807 = n315 | n872 ;
  assign n3808 = ( n200 & n256 ) | ( n200 & ~n3807 ) | ( n256 & ~n3807 ) ;
  assign n3809 = n3807 | n3808 ;
  assign n3810 = n267 | n3809 ;
  assign n3811 = ( n377 & n3704 ) | ( n377 & ~n3810 ) | ( n3704 & ~n3810 ) ;
  assign n3812 = n3810 | n3811 ;
  assign n3813 = ( n935 & n1741 ) | ( n935 & ~n3812 ) | ( n1741 & ~n3812 ) ;
  assign n3814 = n3812 | n3813 ;
  assign n3815 = ( n137 & n149 ) | ( n137 & ~n3814 ) | ( n149 & ~n3814 ) ;
  assign n3816 = n3814 | n3815 ;
  assign n3817 = ( n156 & n379 ) | ( n156 & ~n3816 ) | ( n379 & ~n3816 ) ;
  assign n3818 = n3816 | n3817 ;
  assign n3819 = ( n78 & n84 ) | ( n78 & ~n3818 ) | ( n84 & ~n3818 ) ;
  assign n3820 = n3818 | n3819 ;
  assign n3799 = n1633 & ~n3025 ;
  assign n3800 = n3799 ^ n218 ^ 1'b0 ;
  assign n3801 = n231 & ~n3093 ;
  assign n3802 = n3801 ^ n218 ^ 1'b0 ;
  assign n3803 = ( ~n218 & n3800 ) | ( ~n218 & n3802 ) | ( n3800 & n3802 ) ;
  assign n3798 = n218 & ~n2926 ;
  assign n3804 = n3803 ^ n3798 ^ 1'b0 ;
  assign n3797 = ( n3768 & n3769 ) | ( n3768 & ~n3770 ) | ( n3769 & ~n3770 ) ;
  assign n3805 = n3804 ^ n3797 ^ 1'b0 ;
  assign n3796 = ( n3772 & ~n3773 ) | ( n3772 & n3774 ) | ( ~n3773 & n3774 ) ;
  assign n3806 = n3805 ^ n3796 ^ 1'b0 ;
  assign n3822 = n3821 ^ n3820 ^ n3806 ;
  assign n3824 = n3823 ^ n3822 ^ 1'b0 ;
  assign n3794 = n3759 | n3792 ;
  assign n3795 = n2938 & n3794 ;
  assign n3825 = n3824 ^ n3795 ^ 1'b0 ;
  assign n3853 = n3822 & n3823 ;
  assign n3848 = n3806 & n3820 ;
  assign n3849 = n3806 | n3820 ;
  assign n3850 = n3821 & n3849 ;
  assign n3851 = n3848 | n3850 ;
  assign n3828 = n365 | n1906 ;
  assign n3829 = ( n1951 & n3740 ) | ( n1951 & ~n3828 ) | ( n3740 & ~n3828 ) ;
  assign n3830 = n3828 | n3829 ;
  assign n3831 = ( n491 & n2740 ) | ( n491 & ~n3830 ) | ( n2740 & ~n3830 ) ;
  assign n3832 = n3830 | n3831 ;
  assign n3833 = ( n405 & n2721 ) | ( n405 & ~n3832 ) | ( n2721 & ~n3832 ) ;
  assign n3834 = n3832 | n3833 ;
  assign n3835 = ( n134 & n273 ) | ( n134 & ~n3834 ) | ( n273 & ~n3834 ) ;
  assign n3836 = n3834 | n3835 ;
  assign n3843 = ( n3796 & ~n3797 ) | ( n3796 & n3804 ) | ( ~n3797 & n3804 ) ;
  assign n3839 = n2923 | n3770 ;
  assign n3840 = n218 & ~n3839 ;
  assign n3841 = n3798 & ~n3840 ;
  assign n3842 = ( n3803 & n3840 ) | ( n3803 & ~n3841 ) | ( n3840 & ~n3841 ) ;
  assign n3837 = n3770 ^ n3025 ^ 1'b0 ;
  assign n3838 = n218 & n3837 ;
  assign n3844 = n3843 ^ n3842 ^ n3838 ;
  assign n3845 = n3836 | n3844 ;
  assign n3846 = n3836 & n3844 ;
  assign n3847 = n3845 & ~n3846 ;
  assign n3852 = n3851 ^ n3847 ^ 1'b0 ;
  assign n3854 = n3853 ^ n3852 ^ 1'b0 ;
  assign n3826 = n3794 | n3824 ;
  assign n3827 = n2938 & n3826 ;
  assign n3855 = n3854 ^ n3827 ^ 1'b0 ;
  assign n3871 = n3852 & n3853 ;
  assign n3869 = ( n3836 & n3844 ) | ( n3836 & n3851 ) | ( n3844 & n3851 ) ;
  assign n3858 = n246 | n617 ;
  assign n3859 = ( n711 & n2252 ) | ( n711 & ~n3858 ) | ( n2252 & ~n3858 ) ;
  assign n3860 = n3858 | n3859 ;
  assign n3861 = ( n481 & n2446 ) | ( n481 & ~n3860 ) | ( n2446 & ~n3860 ) ;
  assign n3862 = n3860 | n3861 ;
  assign n3863 = ( n100 & n196 ) | ( n100 & ~n3862 ) | ( n196 & ~n3862 ) ;
  assign n3864 = n3862 | n3863 ;
  assign n3865 = ( n208 & n305 ) | ( n208 & ~n3864 ) | ( n305 & ~n3864 ) ;
  assign n3866 = n3864 | n3865 ;
  assign n3867 = ( n150 & n182 ) | ( n150 & ~n3866 ) | ( n182 & ~n3866 ) ;
  assign n3868 = n3866 | n3867 ;
  assign n3870 = n3869 ^ n3868 ^ 1'b0 ;
  assign n3872 = n3871 ^ n3870 ^ 1'b0 ;
  assign n3856 = n3826 | n3854 ;
  assign n3857 = n2938 & n3856 ;
  assign n3873 = n3872 ^ n3857 ^ 1'b0 ;
  assign n3890 = n3856 | n3872 ;
  assign n3891 = n2938 & n3890 ;
  assign n3875 = n3868 & n3869 ;
  assign n3876 = n436 | n2212 ;
  assign n3877 = ( n420 & n879 ) | ( n420 & ~n3876 ) | ( n879 & ~n3876 ) ;
  assign n3878 = n3876 | n3877 ;
  assign n3879 = ( n674 & n862 ) | ( n674 & ~n3878 ) | ( n862 & ~n3878 ) ;
  assign n3880 = n3878 | n3879 ;
  assign n3881 = ( n185 & n363 ) | ( n185 & ~n3880 ) | ( n363 & ~n3880 ) ;
  assign n3882 = n3880 | n3881 ;
  assign n3883 = ( n122 & n305 ) | ( n122 & ~n3882 ) | ( n305 & ~n3882 ) ;
  assign n3884 = n3882 | n3883 ;
  assign n3885 = ( n232 & n283 ) | ( n232 & ~n3884 ) | ( n283 & ~n3884 ) ;
  assign n3886 = n3884 | n3885 ;
  assign n3888 = n3875 | n3886 ;
  assign n3887 = n3875 & n3886 ;
  assign n3874 = n3870 & n3871 ;
  assign n3889 = n3888 ^ n3887 ^ n3874 ;
  assign n3892 = n3891 ^ n3889 ^ 1'b0 ;
  assign n3907 = n3874 & n3888 ;
  assign n3895 = n3325 | n3809 ;
  assign n3896 = ( n272 & n2397 ) | ( n272 & ~n3895 ) | ( n2397 & ~n3895 ) ;
  assign n3897 = n3895 | n3896 ;
  assign n3898 = ( n238 & n742 ) | ( n238 & ~n3897 ) | ( n742 & ~n3897 ) ;
  assign n3899 = n3897 | n3898 ;
  assign n3900 = ( n123 & n405 ) | ( n123 & ~n3899 ) | ( n405 & ~n3899 ) ;
  assign n3901 = n3899 | n3900 ;
  assign n3902 = ( n124 & n205 ) | ( n124 & ~n3901 ) | ( n205 & ~n3901 ) ;
  assign n3903 = n3901 | n3902 ;
  assign n3904 = ( n188 & n559 ) | ( n188 & ~n3903 ) | ( n559 & ~n3903 ) ;
  assign n3905 = n3903 | n3904 ;
  assign n3906 = n3905 ^ n3887 ^ 1'b0 ;
  assign n3908 = n3907 ^ n3906 ^ 1'b0 ;
  assign n3893 = n3889 | n3890 ;
  assign n3894 = n2938 & n3893 ;
  assign n3909 = n3908 ^ n3894 ^ 1'b0 ;
  assign n3927 = n3893 | n3908 ;
  assign n3928 = n2938 & n3927 ;
  assign n3911 = n3887 & n3905 ;
  assign n3912 = n162 | n814 ;
  assign n3913 = n687 | n3912 ;
  assign n3914 = ( n786 & n3525 ) | ( n786 & ~n3913 ) | ( n3525 & ~n3913 ) ;
  assign n3915 = n3913 | n3914 ;
  assign n3916 = ( n151 & n389 ) | ( n151 & ~n3915 ) | ( n389 & ~n3915 ) ;
  assign n3917 = n3915 | n3916 ;
  assign n3918 = ( n122 & n309 ) | ( n122 & ~n3917 ) | ( n309 & ~n3917 ) ;
  assign n3919 = n3917 | n3918 ;
  assign n3920 = ( n282 & n445 ) | ( n282 & ~n3919 ) | ( n445 & ~n3919 ) ;
  assign n3921 = n3919 | n3920 ;
  assign n3922 = ( n131 & n310 ) | ( n131 & ~n3921 ) | ( n310 & ~n3921 ) ;
  assign n3923 = n3921 | n3922 ;
  assign n3925 = n3911 | n3923 ;
  assign n3924 = n3911 & n3923 ;
  assign n3910 = n3906 & n3907 ;
  assign n3926 = n3925 ^ n3924 ^ n3910 ;
  assign n3929 = n3928 ^ n3926 ^ 1'b0 ;
  assign n3937 = n3910 & n3925 ;
  assign n3932 = n504 | n2774 ;
  assign n3933 = n840 | n3932 ;
  assign n3934 = ( n233 & n376 ) | ( n233 & ~n3933 ) | ( n376 & ~n3933 ) ;
  assign n3935 = n3933 | n3934 ;
  assign n3936 = n3935 ^ n3924 ^ 1'b0 ;
  assign n3938 = n3937 ^ n3936 ^ 1'b0 ;
  assign n3930 = n3926 | n3927 ;
  assign n3931 = n2938 & n3930 ;
  assign n3939 = n3938 ^ n3931 ^ 1'b0 ;
  assign n3946 = n3930 | n3938 ;
  assign n3947 = n2938 & n3946 ;
  assign n3941 = n3924 & n3935 ;
  assign n3942 = n795 | n840 ;
  assign n3944 = n3941 | n3942 ;
  assign n3943 = n3941 & n3942 ;
  assign n3940 = n3936 & n3937 ;
  assign n3945 = n3944 ^ n3943 ^ n3940 ;
  assign n3948 = n3947 ^ n3945 ^ 1'b0 ;
  assign n3951 = n3940 & n3944 ;
  assign n3949 = n3945 | n3946 ;
  assign n3950 = n2938 & n3949 ;
  assign n3952 = n3951 ^ n3950 ^ n3943 ;
  assign n3953 = x21 | n48 ;
  assign n3954 = ( x22 & ~n3952 ) | ( x22 & n3953 ) | ( ~n3952 & n3953 ) ;
  assign n3955 = ~n3952 & n3954 ;
  assign n3956 = ( ~n3943 & n3949 ) | ( ~n3943 & n3951 ) | ( n3949 & n3951 ) ;
  assign n3957 = n3956 ^ n3943 ^ 1'b0 ;
  assign n3958 = x22 | n3953 ;
  assign n3959 = n2938 & ~n3958 ;
  assign n3960 = ( n2938 & n3957 ) | ( n2938 & n3959 ) | ( n3957 & n3959 ) ;
  assign y0 = n2937 ;
  assign y1 = n3041 ;
  assign y2 = n3125 ;
  assign y3 = n3199 ;
  assign y4 = n3270 ;
  assign y5 = n3342 ;
  assign y6 = n3414 ;
  assign y7 = n3472 ;
  assign y8 = n3538 ;
  assign y9 = n3589 ;
  assign y10 = n3637 ;
  assign y11 = n3677 ;
  assign y12 = n3717 ;
  assign y13 = n3758 ;
  assign y14 = n3793 ;
  assign y15 = n3825 ;
  assign y16 = n3855 ;
  assign y17 = n3873 ;
  assign y18 = n3892 ;
  assign y19 = n3909 ;
  assign y20 = n3929 ;
  assign y21 = n3939 ;
  assign y22 = n3948 ;
  assign y23 = ~n3955 ;
  assign y24 = n3960 ;
endmodule
