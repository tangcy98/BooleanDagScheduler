module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 ;
  assign n300 = x9 | x10 ;
  assign n390 = x11 & n300 ;
  assign n391 = x12 | n390 ;
  assign n64 = x12 & n390 ;
  assign n301 = ~n64 ;
  assign n65 = n391 & n301 ;
  assign n66 = x13 | n391 ;
  assign n69 = x14 & n66 ;
  assign n302 = ~x14 ;
  assign n67 = n302 & n66 ;
  assign n120 = n69 ^ n67 ^ x14 ;
  assign n68 = n67 ^ n66 ^ x15 ;
  assign n70 = x15 & n69 ;
  assign n71 = x16 & n70 ;
  assign n72 = x16 | n70 ;
  assign n303 = ~n71 ;
  assign n73 = n303 & n72 ;
  assign n74 = x17 & n72 ;
  assign n75 = x18 & n74 ;
  assign n76 = x18 | n74 ;
  assign n304 = ~n75 ;
  assign n77 = n304 & n76 ;
  assign n78 = x19 & n76 ;
  assign n79 = x20 & n78 ;
  assign n80 = x21 | n79 ;
  assign n104 = x21 & n79 ;
  assign n305 = ~n104 ;
  assign n105 = n80 & n305 ;
  assign n106 = n105 ^ n104 ^ x22 ;
  assign n81 = x22 | n80 ;
  assign n306 = ~x23 ;
  assign n82 = n306 & n81 ;
  assign n83 = n82 ^ n81 ^ x24 ;
  assign n84 = x23 & n81 ;
  assign n307 = ~x24 ;
  assign n85 = n307 & n84 ;
  assign n86 = n85 ^ n84 ^ x25 ;
  assign n87 = x24 & n84 ;
  assign n88 = x25 & n87 ;
  assign n89 = x26 & n88 ;
  assign n90 = x26 | n88 ;
  assign n308 = ~n89 ;
  assign n91 = n308 & n90 ;
  assign n309 = ~x27 ;
  assign n92 = n309 & n90 ;
  assign n93 = n92 ^ n90 ^ x28 ;
  assign n94 = x27 & n90 ;
  assign n310 = ~x28 ;
  assign n95 = n310 & n94 ;
  assign n96 = n95 ^ n94 ^ x29 ;
  assign n97 = ( x9 & n93 ) | ( x9 & n96 ) | ( n93 & n96 ) ;
  assign n311 = ~x9 ;
  assign n98 = n311 & n97 ;
  assign n99 = n94 ^ n92 ^ x27 ;
  assign n100 = ( n91 & n98 ) | ( n91 & n99 ) | ( n98 & n99 ) ;
  assign n312 = ~n91 ;
  assign n101 = n312 & n100 ;
  assign n313 = ~n83 ;
  assign n102 = ( n313 & n86 ) | ( n313 & n101 ) | ( n86 & n101 ) ;
  assign n103 = n83 & n102 ;
  assign n107 = n84 ^ n82 ^ x23 ;
  assign n108 = ( n103 & n106 ) | ( n103 & n107 ) | ( n106 & n107 ) ;
  assign n314 = ~n106 ;
  assign n109 = n314 & n108 ;
  assign n315 = ~x19 ;
  assign n110 = n315 & n76 ;
  assign n111 = n110 ^ n76 ^ x20 ;
  assign n316 = ~n105 ;
  assign n112 = n316 & n111 ;
  assign n113 = n109 & n112 ;
  assign n114 = n110 ^ n78 ^ x19 ;
  assign n115 = ( n77 & n113 ) | ( n77 & n114 ) | ( n113 & n114 ) ;
  assign n317 = ~n77 ;
  assign n116 = n317 & n115 ;
  assign n117 = n73 ^ n71 ^ x17 ;
  assign n118 = ( n73 & n116 ) | ( n73 & n117 ) | ( n116 & n117 ) ;
  assign n318 = ~n73 ;
  assign n119 = n318 & n118 ;
  assign n319 = ~n120 ;
  assign n121 = ( n68 & n119 ) | ( n68 & n319 ) | ( n119 & n319 ) ;
  assign n122 = n120 & n121 ;
  assign n123 = n65 ^ n64 ^ x13 ;
  assign n320 = ~n123 ;
  assign n124 = ( n65 & n122 ) | ( n65 & n320 ) | ( n122 & n320 ) ;
  assign n321 = ~n65 ;
  assign n125 = n321 & n124 ;
  assign n126 = n125 ^ n300 ^ 1'b0 ;
  assign n127 = ( x11 & n300 ) | ( x11 & n126 ) | ( n300 & n126 ) ;
  assign n128 = n127 ^ n300 ^ 1'b0 ;
  assign n322 = ~x10 ;
  assign n129 = x9 & n322 ;
  assign n130 = n129 ^ n300 ^ x9 ;
  assign n323 = ~n130 ;
  assign n131 = x8 & n323 ;
  assign n132 = n128 & n131 ;
  assign n324 = ~x6 ;
  assign n133 = ( n324 & x7 ) | ( n324 & n132 ) | ( x7 & n132 ) ;
  assign n134 = x6 & n133 ;
  assign n325 = ~x4 ;
  assign n135 = ( n325 & x5 ) | ( n325 & n134 ) | ( x5 & n134 ) ;
  assign n136 = x4 & n135 ;
  assign n326 = ~x2 ;
  assign n137 = ( n326 & x3 ) | ( n326 & n136 ) | ( x3 & n136 ) ;
  assign n138 = x2 & n137 ;
  assign n327 = ~x0 ;
  assign n139 = ( n327 & x1 ) | ( n327 & n138 ) | ( x1 & n138 ) ;
  assign n140 = x0 & n139 ;
  assign n141 = x28 & n94 ;
  assign n142 = n140 ^ x29 ^ 1'b0 ;
  assign n328 = ~x29 ;
  assign n143 = ( n328 & n141 ) | ( n328 & n142 ) | ( n141 & n142 ) ;
  assign n144 = ( x29 & n140 ) | ( x29 & n143 ) | ( n140 & n143 ) ;
  assign n145 = x1 | x2 ;
  assign n329 = ~n145 ;
  assign n146 = ( x3 & x4 ) | ( x3 & n329 ) | ( x4 & n329 ) ;
  assign n147 = n145 | n146 ;
  assign n330 = ~n147 ;
  assign n148 = ( x5 & x6 ) | ( x5 & n330 ) | ( x6 & n330 ) ;
  assign n149 = n147 | n148 ;
  assign n331 = ~n149 ;
  assign n150 = ( x7 & x8 ) | ( x7 & n331 ) | ( x8 & n331 ) ;
  assign n151 = n149 | n150 ;
  assign n152 = n129 ^ x11 ^ x10 ;
  assign n332 = ~n152 ;
  assign n153 = ( n130 & n151 ) | ( n130 & n332 ) | ( n151 & n332 ) ;
  assign n333 = ~n151 ;
  assign n154 = n333 & n153 ;
  assign n155 = ( n321 & n123 ) | ( n321 & n154 ) | ( n123 & n154 ) ;
  assign n156 = n65 & n155 ;
  assign n334 = ~n68 ;
  assign n157 = ( n334 & n120 ) | ( n334 & n156 ) | ( n120 & n156 ) ;
  assign n158 = n319 & n157 ;
  assign n335 = ~n117 ;
  assign n159 = n73 & n335 ;
  assign n160 = n158 & n159 ;
  assign n336 = ~n114 ;
  assign n161 = n77 & n336 ;
  assign n162 = n160 & n161 ;
  assign n163 = ( n105 & n111 ) | ( n105 & n162 ) | ( n111 & n162 ) ;
  assign n337 = ~n111 ;
  assign n164 = n337 & n163 ;
  assign n338 = ~n107 ;
  assign n165 = n106 & n338 ;
  assign n166 = n164 & n165 ;
  assign n339 = ~n86 ;
  assign n167 = ( n83 & n339 ) | ( n83 & n166 ) | ( n339 & n166 ) ;
  assign n168 = n313 & n167 ;
  assign n340 = ~n99 ;
  assign n169 = n91 & n340 ;
  assign n170 = n168 & n169 ;
  assign n341 = ~n93 ;
  assign n171 = x9 & n341 ;
  assign n172 = n170 & n171 ;
  assign n173 = ( x29 & n141 ) | ( x29 & n172 ) | ( n141 & n172 ) ;
  assign n342 = ~n172 ;
  assign n174 = n342 & n173 ;
  assign n343 = ~n174 ;
  assign n175 = n144 & n343 ;
  assign n176 = x39 | x40 ;
  assign n177 = x41 & n176 ;
  assign n178 = x42 | n177 ;
  assign n179 = x43 | n178 ;
  assign n344 = ~x44 ;
  assign n180 = n344 & n179 ;
  assign n181 = n180 ^ n179 ^ x45 ;
  assign n345 = ~n178 ;
  assign n182 = x43 & n345 ;
  assign n346 = ~x43 ;
  assign n183 = n346 & n178 ;
  assign n184 = n182 | n183 ;
  assign n185 = n183 ^ x44 ^ x43 ;
  assign n347 = ~n185 ;
  assign n186 = n184 & n347 ;
  assign n348 = ~n181 ;
  assign n187 = ( x45 & n348 ) | ( x45 & n186 ) | ( n348 & n186 ) ;
  assign n188 = x46 | n187 ;
  assign n189 = x47 & n188 ;
  assign n190 = x48 | n189 ;
  assign n191 = x49 & n190 ;
  assign n192 = x50 & n191 ;
  assign n193 = x51 | n192 ;
  assign n194 = x52 | n193 ;
  assign n195 = x53 & n194 ;
  assign n196 = x54 & n195 ;
  assign n197 = x55 & n196 ;
  assign n198 = x56 | n197 ;
  assign n199 = x57 & n198 ;
  assign n200 = x58 & n199 ;
  assign n201 = x59 & n200 ;
  assign n349 = ~n201 ;
  assign n202 = x0 & n349 ;
  assign n350 = ~x53 ;
  assign n203 = n350 & n194 ;
  assign n204 = n203 ^ n194 ^ x54 ;
  assign n351 = ~x54 ;
  assign n205 = n351 & n195 ;
  assign n206 = n205 ^ n195 ^ x55 ;
  assign n207 = x51 & n192 ;
  assign n352 = ~n207 ;
  assign n208 = n193 & n352 ;
  assign n353 = ~x49 ;
  assign n209 = n353 & n190 ;
  assign n236 = n209 ^ n191 ^ x49 ;
  assign n210 = n209 ^ n190 ^ x50 ;
  assign n213 = x46 & n187 ;
  assign n354 = ~n213 ;
  assign n214 = n188 & n354 ;
  assign n233 = n214 ^ n213 ^ x47 ;
  assign n211 = x48 & n189 ;
  assign n355 = ~n211 ;
  assign n212 = n190 & n355 ;
  assign n356 = ~x41 ;
  assign n215 = n356 & n176 ;
  assign n227 = n215 ^ n177 ^ x41 ;
  assign n216 = n215 ^ n176 ^ x42 ;
  assign n217 = x39 & x40 ;
  assign n357 = ~n217 ;
  assign n218 = n176 & n357 ;
  assign n219 = x31 | x32 ;
  assign n220 = x33 | n219 ;
  assign n358 = ~n220 ;
  assign n221 = ( x34 & x35 ) | ( x34 & n358 ) | ( x35 & n358 ) ;
  assign n222 = n220 | n221 ;
  assign n359 = ~n222 ;
  assign n223 = ( x36 & x37 ) | ( x36 & n359 ) | ( x37 & n359 ) ;
  assign n224 = n222 | n223 ;
  assign n360 = ~n224 ;
  assign n225 = ( x38 & n218 ) | ( x38 & n360 ) | ( n218 & n360 ) ;
  assign n361 = ~x38 ;
  assign n226 = n361 & n225 ;
  assign n228 = ( n216 & n226 ) | ( n216 & n227 ) | ( n226 & n227 ) ;
  assign n362 = ~n227 ;
  assign n229 = n362 & n228 ;
  assign n230 = n186 & n229 ;
  assign n231 = ( n181 & n214 ) | ( n181 & n230 ) | ( n214 & n230 ) ;
  assign n232 = n348 & n231 ;
  assign n234 = ( n212 & n232 ) | ( n212 & n233 ) | ( n232 & n233 ) ;
  assign n363 = ~n233 ;
  assign n235 = n363 & n234 ;
  assign n364 = ~n210 ;
  assign n237 = ( n364 & n235 ) | ( n364 & n236 ) | ( n235 & n236 ) ;
  assign n365 = ~n236 ;
  assign n238 = n365 & n237 ;
  assign n239 = n208 & n238 ;
  assign n240 = n208 ^ n207 ^ x52 ;
  assign n241 = n203 ^ n195 ^ x53 ;
  assign n366 = ~n241 ;
  assign n242 = n240 & n366 ;
  assign n243 = n239 & n242 ;
  assign n367 = ~n206 ;
  assign n244 = ( n204 & n367 ) | ( n204 & n243 ) | ( n367 & n243 ) ;
  assign n368 = ~n204 ;
  assign n245 = n368 & n244 ;
  assign n246 = x56 & n197 ;
  assign n369 = ~n246 ;
  assign n247 = n198 & n369 ;
  assign n370 = ~x57 ;
  assign n248 = n370 & n198 ;
  assign n249 = n248 ^ n199 ^ x57 ;
  assign n371 = ~n249 ;
  assign n250 = n247 & n371 ;
  assign n251 = n245 & n250 ;
  assign n252 = n248 ^ n198 ^ x58 ;
  assign n372 = ~n252 ;
  assign n253 = x39 & n372 ;
  assign n254 = n251 & n253 ;
  assign n255 = ( x59 & n200 ) | ( x59 & n254 ) | ( n200 & n254 ) ;
  assign n373 = ~n254 ;
  assign n256 = n373 & n255 ;
  assign n257 = x0 | x30 ;
  assign n258 = n201 & n257 ;
  assign n374 = ~x39 ;
  assign n259 = x30 & n374 ;
  assign n260 = x59 & n259 ;
  assign n261 = n252 & n260 ;
  assign n262 = ( n247 & n249 ) | ( n247 & n261 ) | ( n249 & n261 ) ;
  assign n375 = ~n247 ;
  assign n263 = n375 & n262 ;
  assign n264 = ( n368 & n206 ) | ( n368 & n263 ) | ( n206 & n263 ) ;
  assign n265 = n204 & n264 ;
  assign n266 = ( n240 & n241 ) | ( n240 & n265 ) | ( n241 & n265 ) ;
  assign n376 = ~n240 ;
  assign n267 = n376 & n266 ;
  assign n377 = ~n208 ;
  assign n268 = n377 & n210 ;
  assign n269 = n267 & n268 ;
  assign n270 = ( n212 & n236 ) | ( n212 & n269 ) | ( n236 & n269 ) ;
  assign n378 = ~n212 ;
  assign n271 = n378 & n270 ;
  assign n272 = ( n214 & n233 ) | ( n214 & n271 ) | ( n233 & n271 ) ;
  assign n379 = ~n214 ;
  assign n273 = n379 & n272 ;
  assign n274 = ( n181 & n347 ) | ( n181 & n273 ) | ( n347 & n273 ) ;
  assign n275 = n185 & n274 ;
  assign n380 = ~n184 ;
  assign n276 = ( n380 & n216 ) | ( n380 & n275 ) | ( n216 & n275 ) ;
  assign n381 = ~n216 ;
  assign n277 = n381 & n276 ;
  assign n278 = ( n218 & n227 ) | ( n218 & n277 ) | ( n227 & n277 ) ;
  assign n382 = ~n218 ;
  assign n279 = n382 & n278 ;
  assign n383 = ~x37 ;
  assign n280 = ( n383 & x38 ) | ( n383 & n279 ) | ( x38 & n279 ) ;
  assign n281 = x37 & n280 ;
  assign n384 = ~x35 ;
  assign n282 = ( n384 & x36 ) | ( n384 & n281 ) | ( x36 & n281 ) ;
  assign n283 = x35 & n282 ;
  assign n385 = ~x33 ;
  assign n284 = ( n385 & x34 ) | ( n385 & n283 ) | ( x34 & n283 ) ;
  assign n285 = x33 & n284 ;
  assign n386 = ~x31 ;
  assign n286 = ( n386 & x32 ) | ( n386 & n285 ) | ( x32 & n285 ) ;
  assign n287 = x31 & n286 ;
  assign n387 = ~n256 ;
  assign n288 = ( n387 & n258 ) | ( n387 & n287 ) | ( n258 & n287 ) ;
  assign n289 = n256 | n288 ;
  assign n290 = ( n144 & n202 ) | ( n144 & n289 ) | ( n202 & n289 ) ;
  assign n388 = ~n202 ;
  assign n291 = n388 & n290 ;
  assign n292 = x29 & n141 ;
  assign n293 = ( n342 & n291 ) | ( n342 & n292 ) | ( n291 & n292 ) ;
  assign n294 = n291 ^ n172 ^ 1'b0 ;
  assign n389 = ~n294 ;
  assign n295 = ( n291 & n293 ) | ( n291 & n389 ) | ( n293 & n389 ) ;
  assign n296 = x0 & n201 ;
  assign n297 = x30 & n296 ;
  assign n298 = n256 | n297 ;
  assign n299 = ( n144 & n174 ) | ( n144 & n298 ) | ( n174 & n298 ) ;
  assign n63 = n343 & n299 ;
  assign n61 = ~n175 ;
  assign n62 = ~n295 ;
  assign y0 = n61 ;
  assign y1 = n62 ;
  assign y2 = n63 ;
endmodule
