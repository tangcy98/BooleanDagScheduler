module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 ;
  assign n1205 = x38 | x100 ;
  assign n1206 = x39 | x87 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = ~x224 & x833 ;
  assign n1209 = x332 | x929 ;
  assign n1210 = n1208 & ~n1209 ;
  assign n1211 = x265 & ~x332 ;
  assign n1212 = x224 & ~n1211 ;
  assign n1213 = x222 | n1212 ;
  assign n1214 = n1213 ^ n1210 ^ 1'b0 ;
  assign n1215 = ( n1210 & n1213 ) | ( n1210 & n1214 ) | ( n1213 & n1214 ) ;
  assign n1216 = ( x223 & ~n1210 ) | ( x223 & n1215 ) | ( ~n1210 & n1215 ) ;
  assign n1217 = x332 | x1144 ;
  assign n1218 = n1217 ^ n1216 ^ 1'b0 ;
  assign n1219 = x222 & ~n1208 ;
  assign n1220 = x223 | n1219 ;
  assign n1221 = ( n1217 & n1218 ) | ( n1217 & ~n1220 ) | ( n1218 & ~n1220 ) ;
  assign n1222 = ( n1216 & ~n1218 ) | ( n1216 & n1221 ) | ( ~n1218 & n1221 ) ;
  assign n1223 = x234 & ~x332 ;
  assign n1224 = x95 & ~x479 ;
  assign n1225 = x58 | x90 ;
  assign n1226 = x88 | x98 ;
  assign n1227 = x77 | n1226 ;
  assign n1228 = x50 | n1227 ;
  assign n1229 = x102 | n1228 ;
  assign n1230 = x63 | x107 ;
  assign n1231 = x65 | x71 ;
  assign n1232 = x83 | x103 ;
  assign n1233 = x67 | x69 ;
  assign n1234 = x66 | x73 ;
  assign n1235 = x61 | x76 ;
  assign n1236 = x85 | x106 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = x48 | n1237 ;
  assign n1239 = x89 | n1238 ;
  assign n1240 = x49 | n1239 ;
  assign n1241 = x104 | n1240 ;
  assign n1242 = x45 | n1241 ;
  assign n1243 = x68 | x84 ;
  assign n1244 = x82 | x111 ;
  assign n1245 = x36 | n1244 ;
  assign n1246 = n1243 | n1245 ;
  assign n1247 = n1242 | n1246 ;
  assign n1248 = n1234 | n1247 ;
  assign n1249 = n1233 | n1248 ;
  assign n1250 = n1232 | n1249 ;
  assign n1251 = n1231 | n1250 ;
  assign n1252 = n1230 | n1251 ;
  assign n1253 = x64 | n1252 ;
  assign n1254 = x81 | n1253 ;
  assign n1255 = n1229 | n1254 ;
  assign n1256 = x47 | x91 ;
  assign n1257 = x109 | x110 ;
  assign n1258 = x97 | x108 ;
  assign n1259 = x94 | n1258 ;
  assign n1260 = x53 | x60 ;
  assign n1261 = x86 | n1260 ;
  assign n1262 = x46 | n1261 ;
  assign n1263 = n1259 | n1262 ;
  assign n1264 = n1257 | n1263 ;
  assign n1265 = n1256 | n1264 ;
  assign n1266 = n1255 | n1265 ;
  assign n1267 = n1225 | n1266 ;
  assign n1268 = x35 | x93 ;
  assign n1269 = n1267 | n1268 ;
  assign n1270 = x72 | x96 ;
  assign n1271 = x51 | x70 ;
  assign n1272 = n1270 | n1271 ;
  assign n1273 = n1269 | n1272 ;
  assign n1274 = x32 | x40 ;
  assign n1275 = n1273 | n1274 ;
  assign n1276 = x95 | n1275 ;
  assign n1277 = ~n1224 & n1276 ;
  assign n1278 = ~x137 & x198 ;
  assign n1279 = ~x95 & n1278 ;
  assign n1280 = n1277 | n1279 ;
  assign n1281 = n1223 & n1280 ;
  assign n1282 = x144 | x174 ;
  assign n1283 = x189 | n1282 ;
  assign n1284 = x223 | n1283 ;
  assign n1285 = x234 | x332 ;
  assign n1286 = x70 | n1269 ;
  assign n1287 = x51 | x96 ;
  assign n1288 = x40 | x72 ;
  assign n1289 = x32 | x95 ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = n1287 | n1290 ;
  assign n1292 = n1286 | n1291 ;
  assign n1293 = n1278 | n1292 ;
  assign n1294 = ~n1285 & n1293 ;
  assign n1295 = ( ~n1281 & n1284 ) | ( ~n1281 & n1294 ) | ( n1284 & n1294 ) ;
  assign n1296 = n1281 | n1295 ;
  assign n1297 = ~x223 & n1283 ;
  assign n1298 = n1292 ^ x234 ^ 1'b0 ;
  assign n1299 = ( n1277 & n1292 ) | ( n1277 & n1298 ) | ( n1292 & n1298 ) ;
  assign n1300 = x142 & ~x198 ;
  assign n1301 = x137 | n1300 ;
  assign n1302 = n1301 ^ n1299 ^ 1'b0 ;
  assign n1303 = ( n1299 & n1301 ) | ( n1299 & n1302 ) | ( n1301 & n1302 ) ;
  assign n1304 = ( x332 & n1224 ) | ( x332 & n1285 ) | ( n1224 & n1285 ) ;
  assign n1305 = ( ~n1299 & n1303 ) | ( ~n1299 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1306 = ( ~n1296 & n1297 ) | ( ~n1296 & n1305 ) | ( n1297 & n1305 ) ;
  assign n1307 = n1306 ^ n1296 ^ 1'b0 ;
  assign n1308 = ( n1296 & ~n1306 ) | ( n1296 & n1307 ) | ( ~n1306 & n1307 ) ;
  assign n1309 = ( x222 & x224 ) | ( x222 & ~n1308 ) | ( x224 & ~n1308 ) ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = n1310 ^ n1222 ^ 1'b0 ;
  assign n1312 = ( n1222 & n1310 ) | ( n1222 & n1311 ) | ( n1310 & n1311 ) ;
  assign n1313 = ( x299 & ~n1222 ) | ( x299 & n1312 ) | ( ~n1222 & n1312 ) ;
  assign n1314 = x215 & ~n1217 ;
  assign n1315 = ~x216 & x833 ;
  assign n1316 = x1144 & ~n1315 ;
  assign n1317 = x929 & n1315 ;
  assign n1318 = ( x332 & ~n1316 ) | ( x332 & n1317 ) | ( ~n1316 & n1317 ) ;
  assign n1319 = n1316 | n1318 ;
  assign n1320 = x221 & n1319 ;
  assign n1321 = x216 & ~n1211 ;
  assign n1322 = x153 & ~x332 ;
  assign n1323 = x105 & x228 ;
  assign n1324 = n1322 & ~n1323 ;
  assign n1325 = x216 | n1324 ;
  assign n1326 = x95 & x234 ;
  assign n1327 = x137 | n1326 ;
  assign n1328 = x152 | x161 ;
  assign n1329 = x166 | n1328 ;
  assign n1330 = ~x146 & n1329 ;
  assign n1331 = x210 | n1330 ;
  assign n1332 = n1331 ^ n1327 ^ 1'b0 ;
  assign n1333 = ( n1327 & n1331 ) | ( n1327 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ( n1299 & ~n1327 ) | ( n1299 & n1333 ) | ( ~n1327 & n1333 ) ;
  assign n1335 = n1334 ^ x332 ^ 1'b0 ;
  assign n1336 = ( x105 & x332 ) | ( x105 & ~n1334 ) | ( x332 & ~n1334 ) ;
  assign n1337 = ( x105 & ~n1335 ) | ( x105 & n1336 ) | ( ~n1335 & n1336 ) ;
  assign n1338 = x105 | n1322 ;
  assign n1339 = ( x228 & n1337 ) | ( x228 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1340 = ~n1337 & n1339 ;
  assign n1341 = n1325 | n1340 ;
  assign n1342 = ~n1321 & n1341 ;
  assign n1343 = x221 | n1342 ;
  assign n1344 = ( x215 & ~n1320 ) | ( x215 & n1343 ) | ( ~n1320 & n1343 ) ;
  assign n1345 = ~x215 & n1344 ;
  assign n1346 = ( x299 & n1314 ) | ( x299 & ~n1345 ) | ( n1314 & ~n1345 ) ;
  assign n1347 = ~n1314 & n1346 ;
  assign n1348 = ( n1207 & n1313 ) | ( n1207 & ~n1347 ) | ( n1313 & ~n1347 ) ;
  assign n1349 = ~n1207 & n1348 ;
  assign n1350 = n1217 ^ x215 ^ 1'b0 ;
  assign n1351 = n1319 ^ x221 ^ 1'b0 ;
  assign n1352 = ~n1304 & n1323 ;
  assign n1353 = ( ~n1321 & n1325 ) | ( ~n1321 & n1352 ) | ( n1325 & n1352 ) ;
  assign n1354 = ~n1321 & n1353 ;
  assign n1355 = ( ~n1319 & n1351 ) | ( ~n1319 & n1354 ) | ( n1351 & n1354 ) ;
  assign n1356 = ( ~n1217 & n1350 ) | ( ~n1217 & n1355 ) | ( n1350 & n1355 ) ;
  assign n1357 = x299 & n1356 ;
  assign n1358 = x299 | n1222 ;
  assign n1359 = x222 | x224 ;
  assign n1360 = x223 | n1359 ;
  assign n1361 = n1304 & ~n1360 ;
  assign n1362 = n1358 | n1361 ;
  assign n1363 = ~n1357 & n1362 ;
  assign n1364 = n1207 & ~n1363 ;
  assign n1365 = ( x75 & n1349 ) | ( x75 & ~n1364 ) | ( n1349 & ~n1364 ) ;
  assign n1366 = ~n1349 & n1365 ;
  assign n1367 = x215 & n1217 ;
  assign n1368 = x299 & ~n1367 ;
  assign n1369 = n1255 | n1263 ;
  assign n1370 = x58 | x91 ;
  assign n1371 = x47 | n1370 ;
  assign n1372 = n1257 | n1371 ;
  assign n1373 = n1369 | n1372 ;
  assign n1374 = x90 | x93 ;
  assign n1375 = x70 | x96 ;
  assign n1376 = x35 | x51 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = n1374 | n1377 ;
  assign n1379 = n1373 | n1378 ;
  assign n1380 = n1288 | n1379 ;
  assign n1381 = x32 & n1380 ;
  assign n1382 = ( x32 & x225 ) | ( x32 & n1381 ) | ( x225 & n1381 ) ;
  assign n1383 = n1382 ^ n1381 ^ x32 ;
  assign n1384 = x95 | n1383 ;
  assign n1385 = x60 & ~n1255 ;
  assign n1386 = x53 | n1385 ;
  assign n1387 = x86 | x94 ;
  assign n1388 = x60 | n1255 ;
  assign n1389 = x53 & n1388 ;
  assign n1390 = n1387 | n1389 ;
  assign n1391 = n1386 & ~n1390 ;
  assign n1392 = x46 | n1257 ;
  assign n1393 = n1256 | n1258 ;
  assign n1394 = n1392 | n1393 ;
  assign n1395 = x58 | n1394 ;
  assign n1396 = n1374 | n1395 ;
  assign n1397 = n1391 & ~n1396 ;
  assign n1398 = x35 | n1397 ;
  assign n1399 = x93 | n1267 ;
  assign n1400 = x35 & n1399 ;
  assign n1401 = x35 & ~n1399 ;
  assign n1402 = ~x225 & n1401 ;
  assign n1403 = x70 | n1402 ;
  assign n1404 = x51 | n1403 ;
  assign n1405 = n1400 | n1404 ;
  assign n1406 = n1398 & ~n1405 ;
  assign n1407 = x96 | n1406 ;
  assign n1408 = x47 | n1264 ;
  assign n1409 = n1255 | n1408 ;
  assign n1410 = x35 | x70 ;
  assign n1411 = x51 | n1410 ;
  assign n1412 = x93 | n1225 ;
  assign n1413 = x91 | n1412 ;
  assign n1414 = n1411 | n1413 ;
  assign n1415 = n1409 | n1414 ;
  assign n1416 = x96 & n1415 ;
  assign n1417 = n1288 | n1416 ;
  assign n1418 = n1407 & ~n1417 ;
  assign n1419 = x32 | n1418 ;
  assign n1420 = ~n1384 & n1419 ;
  assign n1421 = n1224 | n1420 ;
  assign n1422 = x95 & n1275 ;
  assign n1423 = x137 | n1422 ;
  assign n1424 = n1421 & ~n1423 ;
  assign n1425 = x210 & x234 ;
  assign n1426 = x137 & ~n1422 ;
  assign n1427 = x96 & ~n1415 ;
  assign n1428 = x51 | x72 ;
  assign n1429 = x40 | n1428 ;
  assign n1430 = n1269 | n1429 ;
  assign n1431 = n1427 & ~n1430 ;
  assign n1432 = x72 & n1379 ;
  assign n1433 = x40 | n1432 ;
  assign n1434 = x51 & n1286 ;
  assign n1435 = x96 | n1434 ;
  assign n1436 = ~x51 & x70 ;
  assign n1437 = n1435 | n1436 ;
  assign n1438 = n1400 | n1402 ;
  assign n1439 = x58 & n1266 ;
  assign n1440 = x90 & n1373 ;
  assign n1441 = x93 | n1440 ;
  assign n1442 = n1439 | n1441 ;
  assign n1443 = x91 & ~n1409 ;
  assign n1444 = n1225 | n1443 ;
  assign n1445 = x109 | n1369 ;
  assign n1446 = x110 & n1445 ;
  assign n1447 = x47 & ~n1255 ;
  assign n1448 = ~n1264 & n1447 ;
  assign n1449 = x47 & ~n1448 ;
  assign n1450 = x91 | n1449 ;
  assign n1451 = n1446 | n1450 ;
  assign n1452 = x47 | x110 ;
  assign n1453 = x109 & ~n1369 ;
  assign n1454 = x102 | n1254 ;
  assign n1455 = n1226 | n1454 ;
  assign n1456 = x50 | n1260 ;
  assign n1457 = x77 | n1456 ;
  assign n1458 = n1387 | n1457 ;
  assign n1459 = n1455 | n1458 ;
  assign n1460 = x97 | n1459 ;
  assign n1461 = x108 & n1460 ;
  assign n1462 = x97 & n1459 ;
  assign n1463 = n1227 | n1454 ;
  assign n1464 = n1456 | n1463 ;
  assign n1465 = ~x86 & x94 ;
  assign n1466 = ~n1464 & n1465 ;
  assign n1467 = x97 | n1466 ;
  assign n1564 = ( x94 & n1387 ) | ( x94 & n1464 ) | ( n1387 & n1464 ) ;
  assign n1468 = x50 & n1463 ;
  assign n1469 = x60 | n1468 ;
  assign n1470 = x77 & ~n1455 ;
  assign n1471 = x50 | n1470 ;
  assign n1472 = x98 | n1454 ;
  assign n1473 = x88 & n1472 ;
  assign n1474 = x81 & n1253 ;
  assign n1475 = x102 & n1254 ;
  assign n1476 = n1474 | n1475 ;
  assign n1477 = x64 & n1252 ;
  assign n1478 = x63 & ~x107 ;
  assign n1479 = ~n1251 & n1478 ;
  assign n1480 = x64 | n1479 ;
  assign n1537 = ( x65 & n1231 ) | ( x65 & n1250 ) | ( n1231 & n1250 ) ;
  assign n1481 = x67 | n1248 ;
  assign n1482 = x69 & n1481 ;
  assign n1483 = ( x103 & n1232 ) | ( x103 & n1249 ) | ( n1232 & n1249 ) ;
  assign n1484 = n1482 | n1483 ;
  assign n1485 = x69 | x83 ;
  assign n1486 = x67 & n1248 ;
  assign n1487 = n1234 | n1242 ;
  assign n1488 = x84 | n1487 ;
  assign n1489 = x68 & n1488 ;
  assign n1490 = x68 | x111 ;
  assign n1491 = x84 & n1487 ;
  assign n1492 = ( x66 & x73 ) | ( x66 & n1242 ) | ( x73 & n1242 ) ;
  assign n1493 = x104 & n1240 ;
  assign n1494 = x45 | n1493 ;
  assign n1495 = x89 & n1238 ;
  assign n1496 = x49 | n1495 ;
  assign n1497 = x85 & x106 ;
  assign n1498 = n1235 | n1497 ;
  assign n1499 = x61 & x76 ;
  assign n1500 = ( n1236 & n1498 ) | ( n1236 & n1499 ) | ( n1498 & n1499 ) ;
  assign n1501 = n1498 & n1500 ;
  assign n1502 = ( x48 & n1237 ) | ( x48 & n1501 ) | ( n1237 & n1501 ) ;
  assign n1503 = n1237 & n1502 ;
  assign n1504 = ( n1239 & n1496 ) | ( n1239 & n1503 ) | ( n1496 & n1503 ) ;
  assign n1505 = n1503 ^ n1496 ^ 1'b0 ;
  assign n1506 = ( n1239 & n1504 ) | ( n1239 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1507 = ( n1241 & n1494 ) | ( n1241 & n1506 ) | ( n1494 & n1506 ) ;
  assign n1508 = n1506 ^ n1494 ^ 1'b0 ;
  assign n1509 = ( n1241 & n1507 ) | ( n1241 & n1508 ) | ( n1507 & n1508 ) ;
  assign n1510 = ( x45 & n1241 ) | ( x45 & ~n1509 ) | ( n1241 & ~n1509 ) ;
  assign n1511 = ~n1509 & n1510 ;
  assign n1512 = n1234 | n1511 ;
  assign n1513 = ~n1492 & n1512 ;
  assign n1514 = x84 | n1513 ;
  assign n1515 = n1514 ^ n1491 ^ 1'b0 ;
  assign n1516 = ( n1491 & n1514 ) | ( n1491 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = ( n1490 & ~n1491 ) | ( n1490 & n1516 ) | ( ~n1491 & n1516 ) ;
  assign n1518 = x68 | n1488 ;
  assign n1519 = ( x82 & n1244 ) | ( x82 & n1518 ) | ( n1244 & n1518 ) ;
  assign n1520 = ( n1489 & n1517 ) | ( n1489 & ~n1519 ) | ( n1517 & ~n1519 ) ;
  assign n1521 = ~n1489 & n1520 ;
  assign n1522 = x36 | x67 ;
  assign n1523 = x82 & ~n1490 ;
  assign n1524 = ~n1488 & n1523 ;
  assign n1525 = ( ~n1521 & n1522 ) | ( ~n1521 & n1524 ) | ( n1522 & n1524 ) ;
  assign n1526 = n1521 | n1525 ;
  assign n1527 = n1244 | n1518 ;
  assign n1528 = x36 & n1527 ;
  assign n1529 = ( n1486 & n1526 ) | ( n1486 & ~n1528 ) | ( n1526 & ~n1528 ) ;
  assign n1530 = ~n1486 & n1529 ;
  assign n1531 = ( ~n1484 & n1485 ) | ( ~n1484 & n1530 ) | ( n1485 & n1530 ) ;
  assign n1532 = ~n1484 & n1531 ;
  assign n1533 = x103 & ~n1485 ;
  assign n1534 = ~n1481 & n1533 ;
  assign n1535 = ( x71 & ~n1532 ) | ( x71 & n1534 ) | ( ~n1532 & n1534 ) ;
  assign n1536 = n1532 | n1535 ;
  assign n1538 = n1537 ^ n1536 ^ 1'b0 ;
  assign n1539 = ( n1536 & n1537 ) | ( n1536 & n1538 ) | ( n1537 & n1538 ) ;
  assign n1540 = ( x107 & ~n1537 ) | ( x107 & n1539 ) | ( ~n1537 & n1539 ) ;
  assign n1541 = ( x63 & n1230 ) | ( x63 & n1251 ) | ( n1230 & n1251 ) ;
  assign n1542 = n1540 & ~n1541 ;
  assign n1543 = ( ~n1477 & n1480 ) | ( ~n1477 & n1542 ) | ( n1480 & n1542 ) ;
  assign n1544 = ~n1477 & n1543 ;
  assign n1545 = x65 & ~x71 ;
  assign n1546 = ~n1250 & n1545 ;
  assign n1547 = ( ~n1541 & n1542 ) | ( ~n1541 & n1546 ) | ( n1542 & n1546 ) ;
  assign n1548 = n1547 ^ x64 ^ 1'b0 ;
  assign n1549 = ( ~n1252 & n1547 ) | ( ~n1252 & n1548 ) | ( n1547 & n1548 ) ;
  assign n1550 = ( x81 & x102 ) | ( x81 & ~n1549 ) | ( x102 & ~n1549 ) ;
  assign n1551 = n1549 | n1550 ;
  assign n1552 = ~n1476 & n1551 ;
  assign n1553 = ( ~n1476 & n1544 ) | ( ~n1476 & n1552 ) | ( n1544 & n1552 ) ;
  assign n1554 = n1226 | n1553 ;
  assign n1555 = x98 & n1454 ;
  assign n1556 = x77 | n1555 ;
  assign n1557 = ( n1473 & n1554 ) | ( n1473 & ~n1556 ) | ( n1554 & ~n1556 ) ;
  assign n1558 = ~n1473 & n1557 ;
  assign n1559 = n1471 | n1558 ;
  assign n1560 = ~n1469 & n1559 ;
  assign n1561 = n1386 | n1560 ;
  assign n1562 = ~n1389 & n1561 ;
  assign n1563 = x86 | n1562 ;
  assign n1565 = n1563 | n1564 ;
  assign n1566 = ( n1467 & ~n1564 ) | ( n1467 & n1565 ) | ( ~n1564 & n1565 ) ;
  assign n1567 = n1566 ^ n1462 ^ 1'b0 ;
  assign n1568 = ( n1462 & n1566 ) | ( n1462 & n1567 ) | ( n1566 & n1567 ) ;
  assign n1569 = ( x108 & ~n1462 ) | ( x108 & n1568 ) | ( ~n1462 & n1568 ) ;
  assign n1570 = ( x46 & ~n1461 ) | ( x46 & n1569 ) | ( ~n1461 & n1569 ) ;
  assign n1571 = ~x46 & n1570 ;
  assign n1572 = ~x109 & n1571 ;
  assign n1573 = n1453 | n1572 ;
  assign n1574 = n1452 | n1573 ;
  assign n1575 = ~n1451 & n1574 ;
  assign n1576 = n1444 | n1575 ;
  assign n1577 = ~n1442 & n1576 ;
  assign n1578 = x93 & ~n1267 ;
  assign n1579 = ( x35 & ~n1577 ) | ( x35 & n1578 ) | ( ~n1577 & n1578 ) ;
  assign n1580 = n1577 | n1579 ;
  assign n1581 = ~n1438 & n1580 ;
  assign n1582 = x51 | n1581 ;
  assign n1583 = ~n1437 & n1582 ;
  assign n1584 = x72 | n1583 ;
  assign n1585 = ~n1433 & n1584 ;
  assign n1586 = x40 & ~n1273 ;
  assign n1587 = ( x32 & ~n1585 ) | ( x32 & n1586 ) | ( ~n1585 & n1586 ) ;
  assign n1588 = n1585 | n1587 ;
  assign n1589 = n1431 | n1588 ;
  assign n1590 = ( x95 & ~n1383 ) | ( x95 & n1589 ) | ( ~n1383 & n1589 ) ;
  assign n1591 = n1426 & n1590 ;
  assign n1592 = ( n1424 & n1425 ) | ( n1424 & ~n1591 ) | ( n1425 & ~n1591 ) ;
  assign n1593 = ~n1424 & n1592 ;
  assign n1594 = x841 & ~n1267 ;
  assign n1595 = ~x93 & n1594 ;
  assign n1596 = ~n1428 & n1595 ;
  assign n1597 = x35 | x40 ;
  assign n1598 = ( x225 & n1375 ) | ( x225 & ~n1597 ) | ( n1375 & ~n1597 ) ;
  assign n1599 = ~n1375 & n1598 ;
  assign n1600 = x32 & ~n1599 ;
  assign n1601 = ( x32 & ~n1596 ) | ( x32 & n1600 ) | ( ~n1596 & n1600 ) ;
  assign n1602 = ( x95 & n1589 ) | ( x95 & ~n1601 ) | ( n1589 & ~n1601 ) ;
  assign n1603 = n1602 ^ n1422 ^ 1'b0 ;
  assign n1604 = ( x137 & n1422 ) | ( x137 & ~n1602 ) | ( n1422 & ~n1602 ) ;
  assign n1605 = ( x137 & ~n1603 ) | ( x137 & n1604 ) | ( ~n1603 & n1604 ) ;
  assign n1606 = n1419 & ~n1601 ;
  assign n1607 = x95 | n1606 ;
  assign n1608 = ( ~x95 & n1224 ) | ( ~x95 & n1607 ) | ( n1224 & n1607 ) ;
  assign n1609 = ~n1422 & n1608 ;
  assign n1610 = x829 & x950 ;
  assign n1611 = x1092 & x1093 ;
  assign n1612 = n1610 & n1611 ;
  assign n1613 = n1608 & ~n1612 ;
  assign n1614 = ~x833 & x957 ;
  assign n1615 = x1091 & ~n1614 ;
  assign n1616 = ~n1330 & n1615 ;
  assign n1617 = ~n1613 & n1616 ;
  assign n1618 = n1609 & ~n1617 ;
  assign n1619 = ~n1422 & n1616 ;
  assign n1620 = x95 & x479 ;
  assign n1621 = x97 | n1391 ;
  assign n1622 = x108 | n1462 ;
  assign n1623 = x110 | n1622 ;
  assign n1624 = x46 | x109 ;
  assign n1625 = n1256 | n1624 ;
  assign n1626 = n1412 | n1625 ;
  assign n1627 = n1623 | n1626 ;
  assign n1628 = ( x35 & n1621 ) | ( x35 & ~n1627 ) | ( n1621 & ~n1627 ) ;
  assign n1629 = n1628 ^ n1621 ^ 1'b0 ;
  assign n1630 = ( x35 & n1628 ) | ( x35 & ~n1629 ) | ( n1628 & ~n1629 ) ;
  assign n1631 = ~n1405 & n1630 ;
  assign n1632 = x96 | n1631 ;
  assign n1633 = ~n1417 & n1632 ;
  assign n1634 = x32 | n1633 ;
  assign n1635 = n1634 ^ n1601 ^ 1'b0 ;
  assign n1636 = ( n1601 & n1634 ) | ( n1601 & n1635 ) | ( n1634 & n1635 ) ;
  assign n1637 = ( x95 & ~n1601 ) | ( x95 & n1636 ) | ( ~n1601 & n1636 ) ;
  assign n1638 = ( n1612 & n1620 ) | ( n1612 & n1637 ) | ( n1620 & n1637 ) ;
  assign n1639 = ~n1620 & n1638 ;
  assign n1640 = x137 | n1639 ;
  assign n1641 = ( x137 & n1619 ) | ( x137 & n1640 ) | ( n1619 & n1640 ) ;
  assign n1642 = ( ~n1605 & n1618 ) | ( ~n1605 & n1641 ) | ( n1618 & n1641 ) ;
  assign n1643 = ~n1605 & n1642 ;
  assign n1644 = ( x210 & x234 ) | ( x210 & n1643 ) | ( x234 & n1643 ) ;
  assign n1645 = x234 & n1644 ;
  assign n1648 = n1224 | n1422 ;
  assign n1646 = ~n1383 & n1588 ;
  assign n1647 = x95 | n1646 ;
  assign n1649 = n1648 ^ n1647 ^ 1'b0 ;
  assign n1650 = ( x137 & ~n1647 ) | ( x137 & n1648 ) | ( ~n1647 & n1648 ) ;
  assign n1651 = ( x137 & ~n1649 ) | ( x137 & n1650 ) | ( ~n1649 & n1650 ) ;
  assign n1652 = x40 | n1270 ;
  assign n1653 = n1406 & ~n1652 ;
  assign n1654 = x32 | n1653 ;
  assign n1655 = ~n1384 & n1654 ;
  assign n1656 = x137 | n1655 ;
  assign n1657 = ( x210 & n1651 ) | ( x210 & n1656 ) | ( n1651 & n1656 ) ;
  assign n1658 = ~n1651 & n1657 ;
  assign n1659 = n1588 & ~n1601 ;
  assign n1660 = x95 | n1659 ;
  assign n1661 = n1660 ^ n1648 ^ 1'b0 ;
  assign n1662 = ( x137 & n1648 ) | ( x137 & ~n1660 ) | ( n1648 & ~n1660 ) ;
  assign n1663 = ( x137 & ~n1661 ) | ( x137 & n1662 ) | ( ~n1661 & n1662 ) ;
  assign n1664 = x210 | x234 ;
  assign n1665 = x95 | n1601 ;
  assign n1666 = n1654 & ~n1665 ;
  assign n1667 = x137 | n1666 ;
  assign n1668 = n1330 & ~n1667 ;
  assign n1669 = n1664 | n1668 ;
  assign n1670 = n1612 & n1615 ;
  assign n1671 = n1630 & n1670 ;
  assign n1672 = n1398 & ~n1670 ;
  assign n1673 = n1671 | n1672 ;
  assign n1674 = n1405 | n1652 ;
  assign n1675 = ( x32 & n1673 ) | ( x32 & ~n1674 ) | ( n1673 & ~n1674 ) ;
  assign n1676 = n1675 ^ n1673 ^ 1'b0 ;
  assign n1677 = ( x32 & n1675 ) | ( x32 & ~n1676 ) | ( n1675 & ~n1676 ) ;
  assign n1678 = n1677 ^ n1665 ^ 1'b0 ;
  assign n1679 = ( n1665 & n1677 ) | ( n1665 & n1678 ) | ( n1677 & n1678 ) ;
  assign n1680 = ( x137 & ~n1665 ) | ( x137 & n1679 ) | ( ~n1665 & n1679 ) ;
  assign n1681 = ( n1330 & ~n1669 ) | ( n1330 & n1680 ) | ( ~n1669 & n1680 ) ;
  assign n1682 = ~n1669 & n1681 ;
  assign n1683 = ( n1658 & ~n1663 ) | ( n1658 & n1682 ) | ( ~n1663 & n1682 ) ;
  assign n1684 = n1663 ^ n1658 ^ 1'b0 ;
  assign n1685 = ( n1658 & n1683 ) | ( n1658 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1686 = ( ~n1593 & n1645 ) | ( ~n1593 & n1685 ) | ( n1645 & n1685 ) ;
  assign n1687 = ~n1593 & n1686 ;
  assign n1688 = ( x153 & x332 ) | ( x153 & ~n1687 ) | ( x332 & ~n1687 ) ;
  assign n1689 = ~x332 & n1688 ;
  assign n1690 = x225 & x841 ;
  assign n1691 = ( x32 & n1381 ) | ( x32 & n1690 ) | ( n1381 & n1690 ) ;
  assign n1692 = x95 | n1691 ;
  assign n1693 = x70 & n1269 ;
  assign n1694 = n1287 | n1693 ;
  assign n1695 = n1288 | n1694 ;
  assign n1696 = n1403 & ~n1695 ;
  assign n1697 = x32 | n1696 ;
  assign n1698 = ~n1692 & n1697 ;
  assign n1699 = x137 & ~n1698 ;
  assign n1700 = x32 | n1586 ;
  assign n1701 = x93 & n1267 ;
  assign n1702 = n1439 | n1440 ;
  assign n1703 = x109 & n1369 ;
  assign n1704 = x46 | n1461 ;
  assign n1705 = ~x53 & n1560 ;
  assign n1706 = x86 | n1705 ;
  assign n1707 = n1564 | n1706 ;
  assign n1708 = ( n1467 & ~n1564 ) | ( n1467 & n1707 ) | ( ~n1564 & n1707 ) ;
  assign n1709 = ~n1462 & n1708 ;
  assign n1710 = x108 | n1709 ;
  assign n1711 = ~n1704 & n1710 ;
  assign n1712 = x109 | n1711 ;
  assign n1713 = ~n1703 & n1712 ;
  assign n1714 = n1452 | n1713 ;
  assign n1715 = ~n1451 & n1714 ;
  assign n1716 = ( n1225 & n1443 ) | ( n1225 & ~n1715 ) | ( n1443 & ~n1715 ) ;
  assign n1717 = n1715 | n1716 ;
  assign n1718 = n1717 ^ n1702 ^ 1'b0 ;
  assign n1719 = ( n1702 & n1717 ) | ( n1702 & n1718 ) | ( n1717 & n1718 ) ;
  assign n1720 = ( x93 & ~n1702 ) | ( x93 & n1719 ) | ( ~n1702 & n1719 ) ;
  assign n1721 = ( x35 & ~n1701 ) | ( x35 & n1720 ) | ( ~n1701 & n1720 ) ;
  assign n1722 = ~x35 & n1721 ;
  assign n1723 = n1404 | n1722 ;
  assign n1724 = n1435 | n1693 ;
  assign n1725 = n1723 & ~n1724 ;
  assign n1726 = x72 | n1725 ;
  assign n1727 = ~n1433 & n1726 ;
  assign n1728 = n1700 | n1727 ;
  assign n1729 = n1670 | n1728 ;
  assign n1730 = n1670 & ~n1700 ;
  assign n1731 = ~x97 & n1708 ;
  assign n1732 = x108 | n1731 ;
  assign n1733 = ( x109 & ~n1704 ) | ( x109 & n1732 ) | ( ~n1704 & n1732 ) ;
  assign n1734 = ~x109 & n1733 ;
  assign n1735 = n1369 & ~n1734 ;
  assign n1736 = ( x109 & n1734 ) | ( x109 & ~n1735 ) | ( n1734 & ~n1735 ) ;
  assign n1737 = n1452 | n1736 ;
  assign n1738 = ~n1451 & n1737 ;
  assign n1739 = ( n1225 & n1443 ) | ( n1225 & ~n1738 ) | ( n1443 & ~n1738 ) ;
  assign n1740 = n1738 | n1739 ;
  assign n1741 = n1740 ^ n1702 ^ 1'b0 ;
  assign n1742 = ( n1702 & n1740 ) | ( n1702 & n1741 ) | ( n1740 & n1741 ) ;
  assign n1743 = ( x93 & ~n1702 ) | ( x93 & n1742 ) | ( ~n1702 & n1742 ) ;
  assign n1744 = ( x35 & ~n1701 ) | ( x35 & n1743 ) | ( ~n1701 & n1743 ) ;
  assign n1745 = ~x35 & n1744 ;
  assign n1746 = n1404 | n1745 ;
  assign n1747 = ~n1724 & n1746 ;
  assign n1748 = x72 | n1747 ;
  assign n1749 = ~n1433 & n1748 ;
  assign n1750 = ( n1691 & n1730 ) | ( n1691 & ~n1749 ) | ( n1730 & ~n1749 ) ;
  assign n1751 = n1750 ^ n1730 ^ 1'b0 ;
  assign n1752 = ( n1691 & n1750 ) | ( n1691 & ~n1751 ) | ( n1750 & ~n1751 ) ;
  assign n1753 = ( x95 & n1729 ) | ( x95 & ~n1752 ) | ( n1729 & ~n1752 ) ;
  assign n1754 = n1753 ^ n1729 ^ 1'b0 ;
  assign n1755 = ( x95 & n1753 ) | ( x95 & ~n1754 ) | ( n1753 & ~n1754 ) ;
  assign n1756 = n1755 ^ n1648 ^ 1'b0 ;
  assign n1757 = ( n1648 & n1755 ) | ( n1648 & n1756 ) | ( n1755 & n1756 ) ;
  assign n1758 = ( x137 & ~n1648 ) | ( x137 & n1757 ) | ( ~n1648 & n1757 ) ;
  assign n1759 = n1758 ^ n1699 ^ 1'b0 ;
  assign n1760 = ( n1699 & n1758 ) | ( n1699 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1761 = ( x210 & ~n1699 ) | ( x210 & n1760 ) | ( ~n1699 & n1760 ) ;
  assign n1762 = ~n1382 & n1728 ;
  assign n1763 = x95 | n1762 ;
  assign n1764 = ( x137 & ~n1648 ) | ( x137 & n1763 ) | ( ~n1648 & n1763 ) ;
  assign n1765 = ~x137 & n1764 ;
  assign n1766 = x95 | n1382 ;
  assign n1767 = ~x137 & x210 ;
  assign n1768 = ( x210 & n1766 ) | ( x210 & n1767 ) | ( n1766 & n1767 ) ;
  assign n1769 = ( x210 & ~n1697 ) | ( x210 & n1768 ) | ( ~n1697 & n1768 ) ;
  assign n1770 = n1223 & ~n1769 ;
  assign n1771 = ( n1223 & n1765 ) | ( n1223 & n1770 ) | ( n1765 & n1770 ) ;
  assign n1772 = n1761 & n1771 ;
  assign n1773 = x72 | n1427 ;
  assign n1774 = n1725 | n1773 ;
  assign n1775 = ~n1433 & n1774 ;
  assign n1776 = n1700 | n1775 ;
  assign n1777 = n1670 | n1776 ;
  assign n1778 = n1747 | n1773 ;
  assign n1779 = ~n1433 & n1778 ;
  assign n1780 = ( n1691 & n1730 ) | ( n1691 & ~n1779 ) | ( n1730 & ~n1779 ) ;
  assign n1781 = n1780 ^ n1730 ^ 1'b0 ;
  assign n1782 = ( n1691 & n1780 ) | ( n1691 & ~n1781 ) | ( n1780 & ~n1781 ) ;
  assign n1783 = ( x95 & n1777 ) | ( x95 & ~n1782 ) | ( n1777 & ~n1782 ) ;
  assign n1784 = ~x95 & n1783 ;
  assign n1785 = x95 & ~n1275 ;
  assign n1786 = ( x137 & ~n1784 ) | ( x137 & n1785 ) | ( ~n1784 & n1785 ) ;
  assign n1787 = n1784 | n1786 ;
  assign n1788 = n1224 & ~n1275 ;
  assign n1789 = x137 & ~n1788 ;
  assign n1790 = x72 | n1274 ;
  assign n1791 = n1427 & ~n1790 ;
  assign n1792 = n1697 | n1791 ;
  assign n1793 = ~n1692 & n1792 ;
  assign n1794 = n1789 & ~n1793 ;
  assign n1795 = ( x210 & n1787 ) | ( x210 & ~n1794 ) | ( n1787 & ~n1794 ) ;
  assign n1796 = n1795 ^ n1787 ^ 1'b0 ;
  assign n1797 = ( x210 & n1795 ) | ( x210 & ~n1796 ) | ( n1795 & ~n1796 ) ;
  assign n1798 = ~n1766 & n1792 ;
  assign n1799 = n1788 | n1798 ;
  assign n1800 = ( x137 & ~x210 ) | ( x137 & n1799 ) | ( ~x210 & n1799 ) ;
  assign n1801 = x210 ^ x137 ^ 1'b0 ;
  assign n1802 = ( x210 & ~n1800 ) | ( x210 & n1801 ) | ( ~n1800 & n1801 ) ;
  assign n1803 = n1802 ^ n1423 ^ 1'b0 ;
  assign n1804 = ~n1382 & n1776 ;
  assign n1805 = x95 | n1804 ;
  assign n1806 = ( n1423 & n1803 ) | ( n1423 & ~n1805 ) | ( n1803 & ~n1805 ) ;
  assign n1807 = ( n1802 & ~n1803 ) | ( n1802 & n1806 ) | ( ~n1803 & n1806 ) ;
  assign n1808 = ( x234 & x332 ) | ( x234 & ~n1807 ) | ( x332 & ~n1807 ) ;
  assign n1809 = n1807 | n1808 ;
  assign n1810 = n1797 & ~n1809 ;
  assign n1811 = ( n1329 & ~n1772 ) | ( n1329 & n1810 ) | ( ~n1772 & n1810 ) ;
  assign n1812 = n1772 | n1811 ;
  assign n1813 = x146 & ~n1761 ;
  assign n1814 = n1698 ^ x137 ^ 1'b0 ;
  assign n1815 = ~n1691 & n1728 ;
  assign n1816 = x95 | n1815 ;
  assign n1817 = ~n1648 & n1816 ;
  assign n1818 = ( n1698 & ~n1814 ) | ( n1698 & n1817 ) | ( ~n1814 & n1817 ) ;
  assign n1819 = ( x146 & x210 ) | ( x146 & ~n1818 ) | ( x210 & ~n1818 ) ;
  assign n1820 = n1818 | n1819 ;
  assign n1821 = ( n1771 & n1813 ) | ( n1771 & n1820 ) | ( n1813 & n1820 ) ;
  assign n1822 = ~n1813 & n1821 ;
  assign n1823 = x146 & ~n1797 ;
  assign n1824 = ~n1691 & n1776 ;
  assign n1825 = x95 | n1824 ;
  assign n1826 = ~n1422 & n1825 ;
  assign n1827 = x137 | n1826 ;
  assign n1828 = ~n1794 & n1827 ;
  assign n1829 = ( x146 & x210 ) | ( x146 & ~n1828 ) | ( x210 & ~n1828 ) ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = ( ~n1809 & n1823 ) | ( ~n1809 & n1830 ) | ( n1823 & n1830 ) ;
  assign n1832 = ~n1823 & n1831 ;
  assign n1833 = ( n1329 & n1822 ) | ( n1329 & ~n1832 ) | ( n1822 & ~n1832 ) ;
  assign n1834 = ~n1822 & n1833 ;
  assign n1835 = ( x153 & n1812 ) | ( x153 & ~n1834 ) | ( n1812 & ~n1834 ) ;
  assign n1836 = ~x153 & n1835 ;
  assign n1837 = ( x228 & ~n1689 ) | ( x228 & n1836 ) | ( ~n1689 & n1836 ) ;
  assign n1838 = n1689 | n1837 ;
  assign n1839 = x46 & ~n1258 ;
  assign n1840 = ~n1459 & n1839 ;
  assign n1841 = x109 | n1840 ;
  assign n1842 = n1571 | n1841 ;
  assign n1843 = ~n1703 & n1842 ;
  assign n1844 = n1452 | n1843 ;
  assign n1845 = ~n1451 & n1844 ;
  assign n1846 = ( n1225 & n1443 ) | ( n1225 & ~n1845 ) | ( n1443 & ~n1845 ) ;
  assign n1847 = n1845 | n1846 ;
  assign n1848 = ( n1439 & ~n1441 ) | ( n1439 & n1847 ) | ( ~n1441 & n1847 ) ;
  assign n1849 = ~n1439 & n1848 ;
  assign n1850 = ( x35 & n1578 ) | ( x35 & ~n1849 ) | ( n1578 & ~n1849 ) ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = n1851 ^ n1438 ^ 1'b0 ;
  assign n1853 = ( n1438 & n1851 ) | ( n1438 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = ( x51 & ~n1438 ) | ( x51 & n1853 ) | ( ~n1438 & n1853 ) ;
  assign n1855 = ( n1435 & ~n1436 ) | ( n1435 & n1854 ) | ( ~n1436 & n1854 ) ;
  assign n1856 = ~n1435 & n1855 ;
  assign n1857 = x72 | n1856 ;
  assign n1858 = ~n1433 & n1857 ;
  assign n1859 = n1700 | n1858 ;
  assign n1860 = ~n1383 & n1859 ;
  assign n1861 = x95 | n1860 ;
  assign n1862 = n1861 ^ n1648 ^ 1'b0 ;
  assign n1863 = ( x137 & n1648 ) | ( x137 & ~n1861 ) | ( n1648 & ~n1861 ) ;
  assign n1864 = ( x137 & ~n1862 ) | ( x137 & n1863 ) | ( ~n1862 & n1863 ) ;
  assign n1865 = ( x137 & n1655 ) | ( x137 & ~n1864 ) | ( n1655 & ~n1864 ) ;
  assign n1866 = ~n1864 & n1865 ;
  assign n1867 = ~n1601 & n1859 ;
  assign n1868 = x95 | n1867 ;
  assign n1869 = n1868 ^ n1648 ^ 1'b0 ;
  assign n1870 = ( x137 & n1648 ) | ( x137 & ~n1868 ) | ( n1648 & ~n1868 ) ;
  assign n1871 = ( x137 & ~n1869 ) | ( x137 & n1870 ) | ( ~n1869 & n1870 ) ;
  assign n1872 = n1680 & ~n1871 ;
  assign n1873 = n1866 ^ x210 ^ 1'b0 ;
  assign n1874 = ( n1866 & n1872 ) | ( n1866 & ~n1873 ) | ( n1872 & ~n1873 ) ;
  assign n1875 = x146 & n1874 ;
  assign n1876 = n1667 & ~n1871 ;
  assign n1877 = x210 | n1876 ;
  assign n1878 = x210 & ~n1866 ;
  assign n1879 = ( x146 & n1877 ) | ( x146 & ~n1878 ) | ( n1877 & ~n1878 ) ;
  assign n1880 = ~x146 & n1879 ;
  assign n1881 = ( n1285 & ~n1875 ) | ( n1285 & n1880 ) | ( ~n1875 & n1880 ) ;
  assign n1882 = n1875 | n1881 ;
  assign n1883 = n1421 ^ x137 ^ 1'b0 ;
  assign n1884 = x479 & n1422 ;
  assign n1885 = n1431 | n1859 ;
  assign n1886 = ~n1383 & n1885 ;
  assign n1887 = ~x95 & n1886 ;
  assign n1888 = ( x95 & ~n1884 ) | ( x95 & n1887 ) | ( ~n1884 & n1887 ) ;
  assign n1889 = ( n1421 & n1883 ) | ( n1421 & n1888 ) | ( n1883 & n1888 ) ;
  assign n1890 = x210 & ~n1889 ;
  assign n1891 = x146 | n1890 ;
  assign n1892 = ~n1601 & n1885 ;
  assign n1893 = ~x95 & n1892 ;
  assign n1894 = ( x95 & ~n1884 ) | ( x95 & n1893 ) | ( ~n1884 & n1893 ) ;
  assign n1895 = x137 & ~n1894 ;
  assign n1896 = x137 | n1608 ;
  assign n1897 = ~n1895 & n1896 ;
  assign n1898 = x210 | n1897 ;
  assign n1899 = n1223 & ~n1898 ;
  assign n1900 = ( n1223 & n1891 ) | ( n1223 & n1899 ) | ( n1891 & n1899 ) ;
  assign n1901 = n1613 | n1640 ;
  assign n1902 = n1615 & ~n1895 ;
  assign n1903 = n1901 & n1902 ;
  assign n1904 = ( ~n1615 & n1897 ) | ( ~n1615 & n1903 ) | ( n1897 & n1903 ) ;
  assign n1905 = n1903 ^ n1615 ^ 1'b0 ;
  assign n1906 = ( n1903 & n1904 ) | ( n1903 & ~n1905 ) | ( n1904 & ~n1905 ) ;
  assign n1907 = x210 | n1906 ;
  assign n1908 = ~n1890 & n1907 ;
  assign n1909 = ( x146 & ~n1900 ) | ( x146 & n1908 ) | ( ~n1900 & n1908 ) ;
  assign n1910 = n1909 ^ n1900 ^ 1'b0 ;
  assign n1911 = ( n1900 & ~n1909 ) | ( n1900 & n1910 ) | ( ~n1909 & n1910 ) ;
  assign n1912 = n1329 & ~n1911 ;
  assign n1913 = n1882 & n1912 ;
  assign n1914 = ~x234 & n1874 ;
  assign n1915 = x332 | n1914 ;
  assign n1916 = x234 & n1908 ;
  assign n1917 = ( ~n1329 & n1915 ) | ( ~n1329 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = ~n1329 & n1917 ;
  assign n1919 = ( x105 & n1913 ) | ( x105 & ~n1918 ) | ( n1913 & ~n1918 ) ;
  assign n1920 = ~n1913 & n1919 ;
  assign n1921 = ~x105 & n1322 ;
  assign n1922 = ( x228 & n1920 ) | ( x228 & ~n1921 ) | ( n1920 & ~n1921 ) ;
  assign n1923 = ~n1920 & n1922 ;
  assign n1924 = ( x216 & n1838 ) | ( x216 & ~n1923 ) | ( n1838 & ~n1923 ) ;
  assign n1925 = n1924 ^ n1838 ^ 1'b0 ;
  assign n1926 = ( x216 & n1924 ) | ( x216 & ~n1925 ) | ( n1924 & ~n1925 ) ;
  assign n1927 = n1926 ^ n1321 ^ 1'b0 ;
  assign n1928 = ( n1321 & n1926 ) | ( n1321 & n1927 ) | ( n1926 & n1927 ) ;
  assign n1929 = ( x221 & ~n1321 ) | ( x221 & n1928 ) | ( ~n1321 & n1928 ) ;
  assign n1930 = n1929 ^ n1320 ^ 1'b0 ;
  assign n1931 = ( n1320 & n1929 ) | ( n1320 & n1930 ) | ( n1929 & n1930 ) ;
  assign n1932 = ( x215 & ~n1320 ) | ( x215 & n1931 ) | ( ~n1320 & n1931 ) ;
  assign n1933 = n1368 & n1932 ;
  assign n1934 = x198 & ~n1889 ;
  assign n1935 = x198 | n1906 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = x234 & n1936 ;
  assign n1938 = x198 & ~n1866 ;
  assign n1939 = x198 | n1872 ;
  assign n1940 = ~n1938 & n1939 ;
  assign n1941 = ~x234 & n1940 ;
  assign n1942 = ( x332 & ~n1937 ) | ( x332 & n1941 ) | ( ~n1937 & n1941 ) ;
  assign n1943 = n1937 | n1942 ;
  assign n1944 = ( x223 & ~n1283 ) | ( x223 & n1943 ) | ( ~n1283 & n1943 ) ;
  assign n1945 = ~x223 & n1944 ;
  assign n1946 = x142 | n1934 ;
  assign n1947 = x198 | n1897 ;
  assign n1948 = n1223 & ~n1947 ;
  assign n1949 = ( n1223 & n1946 ) | ( n1223 & n1948 ) | ( n1946 & n1948 ) ;
  assign n1950 = ( x142 & n1936 ) | ( x142 & ~n1949 ) | ( n1936 & ~n1949 ) ;
  assign n1951 = n1950 ^ n1949 ^ 1'b0 ;
  assign n1952 = ( n1949 & ~n1950 ) | ( n1949 & n1951 ) | ( ~n1950 & n1951 ) ;
  assign n1953 = x142 & n1940 ;
  assign n1954 = x198 | n1876 ;
  assign n1955 = x142 | n1938 ;
  assign n1956 = n1954 & ~n1955 ;
  assign n1957 = ( n1285 & ~n1953 ) | ( n1285 & n1956 ) | ( ~n1953 & n1956 ) ;
  assign n1958 = n1953 | n1957 ;
  assign n1959 = ( x223 & n1283 ) | ( x223 & n1958 ) | ( n1283 & n1958 ) ;
  assign n1960 = ~x223 & n1959 ;
  assign n1961 = ( n1945 & ~n1952 ) | ( n1945 & n1960 ) | ( ~n1952 & n1960 ) ;
  assign n1962 = n1952 ^ n1945 ^ 1'b0 ;
  assign n1963 = ( n1945 & n1961 ) | ( n1945 & ~n1962 ) | ( n1961 & ~n1962 ) ;
  assign n1964 = ( x222 & ~x224 ) | ( x222 & n1963 ) | ( ~x224 & n1963 ) ;
  assign n1965 = ~x222 & n1964 ;
  assign n1966 = ( x299 & n1222 ) | ( x299 & ~n1965 ) | ( n1222 & ~n1965 ) ;
  assign n1967 = n1965 | n1966 ;
  assign n1968 = ( x39 & ~n1933 ) | ( x39 & n1967 ) | ( ~n1933 & n1967 ) ;
  assign n1969 = ~x39 & n1968 ;
  assign n1970 = x137 & ~n1299 ;
  assign n1971 = n1304 | n1970 ;
  assign n1972 = ~n1360 & n1971 ;
  assign n1973 = ( x299 & n1222 ) | ( x299 & ~n1972 ) | ( n1222 & ~n1972 ) ;
  assign n1974 = n1972 | n1973 ;
  assign n1975 = n1211 ^ x216 ^ 1'b0 ;
  assign n1976 = x332 | n1276 ;
  assign n1977 = x137 | x153 ;
  assign n1978 = n1976 | n1977 ;
  assign n1979 = x137 & ~n1292 ;
  assign n1980 = n1322 & ~n1979 ;
  assign n1981 = x228 | n1980 ;
  assign n1982 = n1978 & ~n1981 ;
  assign n1983 = ( n1338 & n1921 ) | ( n1338 & ~n1971 ) | ( n1921 & ~n1971 ) ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = ( x228 & n1982 ) | ( x228 & ~n1984 ) | ( n1982 & ~n1984 ) ;
  assign n1986 = ( ~n1211 & n1975 ) | ( ~n1211 & n1985 ) | ( n1975 & n1985 ) ;
  assign n1987 = ( n1319 & ~n1351 ) | ( n1319 & n1986 ) | ( ~n1351 & n1986 ) ;
  assign n1988 = ( n1217 & ~n1350 ) | ( n1217 & n1987 ) | ( ~n1350 & n1987 ) ;
  assign n1989 = x299 & ~n1988 ;
  assign n1990 = n1974 & ~n1989 ;
  assign n1991 = x39 & n1990 ;
  assign n1992 = ( x38 & ~n1969 ) | ( x38 & n1991 ) | ( ~n1969 & n1991 ) ;
  assign n1993 = n1969 | n1992 ;
  assign n1994 = x38 | x39 ;
  assign n1995 = x210 & ~x252 ;
  assign n1996 = n1330 | n1995 ;
  assign n1997 = ~n1978 & n1996 ;
  assign n1998 = n1330 & n1979 ;
  assign n1999 = x252 | n1767 ;
  assign n2000 = ( n1330 & n1976 ) | ( n1330 & ~n1999 ) | ( n1976 & ~n1999 ) ;
  assign n2001 = n1999 | n2000 ;
  assign n2002 = ( n1322 & n1998 ) | ( n1322 & n2001 ) | ( n1998 & n2001 ) ;
  assign n2003 = ~n1998 & n2002 ;
  assign n2004 = ( ~x228 & n1997 ) | ( ~x228 & n2003 ) | ( n1997 & n2003 ) ;
  assign n2005 = ~x228 & n2004 ;
  assign n2006 = ( x216 & n1340 ) | ( x216 & ~n2005 ) | ( n1340 & ~n2005 ) ;
  assign n2007 = n2005 | n2006 ;
  assign n2008 = n2007 ^ n1321 ^ 1'b0 ;
  assign n2009 = ( n1321 & n2007 ) | ( n1321 & n2008 ) | ( n2007 & n2008 ) ;
  assign n2010 = ( x221 & ~n1321 ) | ( x221 & n2009 ) | ( ~n1321 & n2009 ) ;
  assign n2011 = ( x215 & ~n1320 ) | ( x215 & n2010 ) | ( ~n1320 & n2010 ) ;
  assign n2012 = ~x215 & n2011 ;
  assign n2013 = ( x299 & n1314 ) | ( x299 & ~n2012 ) | ( n1314 & ~n2012 ) ;
  assign n2014 = ~n1314 & n2013 ;
  assign n2015 = ( n1313 & n1994 ) | ( n1313 & ~n2014 ) | ( n1994 & ~n2014 ) ;
  assign n2016 = ~n1994 & n2015 ;
  assign n2017 = ~n1363 & n1994 ;
  assign n2018 = x100 & ~n2017 ;
  assign n2019 = n2018 ^ n2016 ^ 1'b0 ;
  assign n2020 = ( n2016 & n2018 ) | ( n2016 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2021 = ( x87 & ~n2016 ) | ( x87 & n2020 ) | ( ~n2016 & n2020 ) ;
  assign n2022 = x215 | x221 ;
  assign n2023 = n1325 | n2022 ;
  assign n2024 = n1971 & ~n2023 ;
  assign n2025 = n1356 & ~n2024 ;
  assign n2026 = x299 & n2025 ;
  assign n2027 = ( x39 & n1974 ) | ( x39 & ~n2026 ) | ( n1974 & ~n2026 ) ;
  assign n2028 = ~x39 & n2027 ;
  assign n2029 = x39 & n1363 ;
  assign n2030 = x38 & ~n2029 ;
  assign n2031 = n2030 ^ n2028 ^ 1'b0 ;
  assign n2032 = ( n2028 & n2030 ) | ( n2028 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = ( x100 & ~n2028 ) | ( x100 & n2032 ) | ( ~n2028 & n2032 ) ;
  assign n2034 = ~n2021 & n2033 ;
  assign n2035 = ( n1993 & n2021 ) | ( n1993 & ~n2034 ) | ( n2021 & ~n2034 ) ;
  assign n2036 = x39 | n1205 ;
  assign n2037 = n2036 ^ n1990 ^ 1'b0 ;
  assign n2038 = ( n1363 & n1990 ) | ( n1363 & n2037 ) | ( n1990 & n2037 ) ;
  assign n2039 = x87 & ~n2038 ;
  assign n2040 = ( x75 & n2035 ) | ( x75 & ~n2039 ) | ( n2035 & ~n2039 ) ;
  assign n2041 = ~x75 & n2040 ;
  assign n2042 = ( ~x92 & n1366 ) | ( ~x92 & n2041 ) | ( n1366 & n2041 ) ;
  assign n2043 = ~x92 & n2042 ;
  assign n2044 = x75 | x87 ;
  assign n2045 = n2038 | n2044 ;
  assign n2046 = x92 & ~n2044 ;
  assign n2047 = ( x92 & n1363 ) | ( x92 & n2046 ) | ( n1363 & n2046 ) ;
  assign n2048 = n2045 & n2047 ;
  assign n2049 = ( x54 & ~n2043 ) | ( x54 & n2048 ) | ( ~n2043 & n2048 ) ;
  assign n2050 = n2043 | n2049 ;
  assign n2051 = x87 | x100 ;
  assign n2052 = x38 | n2051 ;
  assign n2053 = x75 | x92 ;
  assign n2054 = n2052 | n2053 ;
  assign n2055 = n2028 & ~n2054 ;
  assign n2056 = n1207 | n2053 ;
  assign n2057 = n1363 & n2056 ;
  assign n2058 = n2055 | n2057 ;
  assign n2059 = x54 & ~n2058 ;
  assign n2060 = ( x74 & n2050 ) | ( x74 & ~n2059 ) | ( n2050 & ~n2059 ) ;
  assign n2061 = ~x74 & n2060 ;
  assign n2062 = x54 & ~n1363 ;
  assign n2063 = x74 & ~n2062 ;
  assign n2064 = ( n2058 & n2059 ) | ( n2058 & n2063 ) | ( n2059 & n2063 ) ;
  assign n2065 = ( ~x55 & n2061 ) | ( ~x55 & n2064 ) | ( n2061 & n2064 ) ;
  assign n2066 = ~x55 & n2065 ;
  assign n2067 = x54 | x74 ;
  assign n2068 = n2053 | n2067 ;
  assign n2069 = n2051 | n2068 ;
  assign n2070 = n1994 | n2069 ;
  assign n2071 = n1356 & n2070 ;
  assign n2072 = x228 & n1338 ;
  assign n2073 = ~x228 & n1322 ;
  assign n2074 = n1292 & n2073 ;
  assign n2075 = x216 | n2074 ;
  assign n2076 = ~x332 & n1299 ;
  assign n2077 = x105 & ~n2076 ;
  assign n2078 = ~n2075 & n2077 ;
  assign n2079 = ( n2072 & n2075 ) | ( n2072 & ~n2078 ) | ( n2075 & ~n2078 ) ;
  assign n2080 = n2079 ^ n1321 ^ 1'b0 ;
  assign n2081 = ( n1321 & n2079 ) | ( n1321 & n2080 ) | ( n2079 & n2080 ) ;
  assign n2082 = ( x221 & ~n1321 ) | ( x221 & n2081 ) | ( ~n1321 & n2081 ) ;
  assign n2083 = n2082 ^ n1320 ^ 1'b0 ;
  assign n2084 = ( n1320 & n2082 ) | ( n1320 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2085 = ( x215 & ~n1320 ) | ( x215 & n2084 ) | ( ~n1320 & n2084 ) ;
  assign n2086 = ( ~n1367 & n2070 ) | ( ~n1367 & n2085 ) | ( n2070 & n2085 ) ;
  assign n2087 = ~n2070 & n2086 ;
  assign n2088 = ( x55 & n2071 ) | ( x55 & ~n2087 ) | ( n2071 & ~n2087 ) ;
  assign n2089 = ~n2071 & n2088 ;
  assign n2090 = ( x56 & ~n2066 ) | ( x56 & n2089 ) | ( ~n2066 & n2089 ) ;
  assign n2091 = n2066 | n2090 ;
  assign n2092 = x56 & n1356 ;
  assign n2093 = x62 & ~n2092 ;
  assign n2094 = n2093 ^ x59 ^ 1'b0 ;
  assign n2095 = x100 | n1994 ;
  assign n2096 = x92 | n2044 ;
  assign n2097 = n2067 | n2096 ;
  assign n2098 = x55 | n2097 ;
  assign n2099 = n2095 | n2098 ;
  assign n2100 = n2099 ^ n1988 ^ 1'b0 ;
  assign n2101 = ( ~n1356 & n1988 ) | ( ~n1356 & n2100 ) | ( n1988 & n2100 ) ;
  assign n2102 = x56 | n2101 ;
  assign n2103 = ( n2093 & ~n2094 ) | ( n2093 & n2102 ) | ( ~n2094 & n2102 ) ;
  assign n2104 = ( x59 & n2094 ) | ( x59 & n2103 ) | ( n2094 & n2103 ) ;
  assign n2105 = x56 & ~n2101 ;
  assign n2106 = x62 | n2105 ;
  assign n2107 = ~n2104 & n2106 ;
  assign n2108 = ( n2091 & n2104 ) | ( n2091 & ~n2107 ) | ( n2104 & ~n2107 ) ;
  assign n2109 = x56 | x62 ;
  assign n2110 = n2099 | n2109 ;
  assign n2111 = n2024 & ~n2110 ;
  assign n2112 = ~x59 & n2111 ;
  assign n2113 = x57 & ~n1356 ;
  assign n2114 = ( x57 & n2112 ) | ( x57 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2115 = x59 & n1356 ;
  assign n2116 = ~n2111 & n2115 ;
  assign n2117 = x57 | n2116 ;
  assign n2118 = ~n2114 & n2117 ;
  assign n2119 = ( n2108 & n2114 ) | ( n2108 & ~n2118 ) | ( n2114 & ~n2118 ) ;
  assign n2120 = x57 | x59 ;
  assign n2121 = ~x939 & n1315 ;
  assign n2122 = x1146 | n1315 ;
  assign n2123 = ( x221 & n2121 ) | ( x221 & n2122 ) | ( n2121 & n2122 ) ;
  assign n2124 = ~n2121 & n2123 ;
  assign n2125 = x216 & ~x221 ;
  assign n2126 = x276 & n2125 ;
  assign n2127 = x216 | n1323 ;
  assign n2128 = ~n2126 & n2127 ;
  assign n2129 = x221 | n2128 ;
  assign n2130 = ( x215 & ~n2124 ) | ( x215 & n2129 ) | ( ~n2124 & n2129 ) ;
  assign n2131 = ~x215 & n2130 ;
  assign n2132 = x1146 & ~n2131 ;
  assign n2133 = ( x215 & n2131 ) | ( x215 & ~n2132 ) | ( n2131 & ~n2132 ) ;
  assign n2134 = x1146 ^ x215 ^ 1'b0 ;
  assign n2135 = n2124 | n2126 ;
  assign n2136 = ( x1146 & ~n2134 ) | ( x1146 & n2135 ) | ( ~n2134 & n2135 ) ;
  assign n2137 = n2133 ^ x154 ^ 1'b0 ;
  assign n2138 = ( n2133 & ~n2136 ) | ( n2133 & n2137 ) | ( ~n2136 & n2137 ) ;
  assign n2139 = n2120 & n2138 ;
  assign n2140 = x215 & x1146 ;
  assign n2141 = n2124 | n2140 ;
  assign n2142 = x228 | n1292 ;
  assign n2143 = x216 | n2142 ;
  assign n2144 = n2141 | n2143 ;
  assign n2145 = x154 & n2136 ;
  assign n2146 = n2144 | n2145 ;
  assign n2147 = x55 | n2070 ;
  assign n2148 = n2138 | n2147 ;
  assign n2149 = n2146 & ~n2148 ;
  assign n2150 = x56 | n2098 ;
  assign n2151 = n2095 | n2150 ;
  assign n2152 = ~n2138 & n2151 ;
  assign n2153 = n2149 | n2152 ;
  assign n2154 = x62 & n2153 ;
  assign n2155 = n2099 & ~n2138 ;
  assign n2156 = x56 & ~n2155 ;
  assign n2157 = n2156 ^ n2149 ^ 1'b0 ;
  assign n2158 = ( n2149 & n2156 ) | ( n2149 & n2157 ) | ( n2156 & n2157 ) ;
  assign n2159 = ( x62 & ~n2149 ) | ( x62 & n2158 ) | ( ~n2149 & n2158 ) ;
  assign n2160 = x223 & ~x1146 ;
  assign n2161 = ~x222 & x224 ;
  assign n2162 = ~x939 & n1208 ;
  assign n2163 = x1146 | n1208 ;
  assign n2164 = ( x222 & n2162 ) | ( x222 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = ~n2162 & n2164 ;
  assign n2166 = x223 | n2165 ;
  assign n2167 = x224 & ~x276 ;
  assign n2168 = x222 | n2167 ;
  assign n2169 = ~n2166 & n2168 ;
  assign n2170 = x222 | x223 ;
  assign n2171 = ( n2161 & ~n2169 ) | ( n2161 & n2170 ) | ( ~n2169 & n2170 ) ;
  assign n2172 = ( x299 & ~n2160 ) | ( x299 & n2171 ) | ( ~n2160 & n2171 ) ;
  assign n2173 = ~x299 & n2172 ;
  assign n2174 = x299 & ~n2138 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = n2067 & ~n2175 ;
  assign n2177 = n2044 | n2095 ;
  assign n2178 = ~n2175 & n2177 ;
  assign n2179 = x299 & ~n2133 ;
  assign n2180 = n2144 & n2179 ;
  assign n2181 = ( ~x154 & n2173 ) | ( ~x154 & n2180 ) | ( n2173 & n2180 ) ;
  assign n2182 = ~x154 & n2181 ;
  assign n2183 = x299 & ~n2136 ;
  assign n2184 = n2183 ^ n2173 ^ x299 ;
  assign n2185 = x154 & n2184 ;
  assign n2186 = ( n2036 & ~n2182 ) | ( n2036 & n2185 ) | ( ~n2182 & n2185 ) ;
  assign n2187 = n2182 | n2186 ;
  assign n2188 = n2044 | n2187 ;
  assign n2189 = ( x92 & n2178 ) | ( x92 & n2188 ) | ( n2178 & n2188 ) ;
  assign n2190 = ~n2178 & n2189 ;
  assign n2191 = x75 & ~n2175 ;
  assign n2192 = n2036 & ~n2175 ;
  assign n2193 = x87 & ~n2187 ;
  assign n2194 = ( x87 & n2192 ) | ( x87 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = x252 | n1292 ;
  assign n2196 = n1292 ^ x146 ^ 1'b0 ;
  assign n2197 = ( n1292 & n2195 ) | ( n1292 & n2196 ) | ( n2195 & n2196 ) ;
  assign n2198 = x152 & n2197 ;
  assign n2199 = x161 | x166 ;
  assign n2200 = n2195 | n2199 ;
  assign n2201 = ~n2197 & n2199 ;
  assign n2202 = ( x152 & n2200 ) | ( x152 & ~n2201 ) | ( n2200 & ~n2201 ) ;
  assign n2203 = ~x152 & n2202 ;
  assign n2204 = x38 | x216 ;
  assign n2205 = x228 | n2204 ;
  assign n2206 = ~x154 & x299 ;
  assign n2207 = ~x39 & n2206 ;
  assign n2208 = ( n2141 & ~n2205 ) | ( n2141 & n2207 ) | ( ~n2205 & n2207 ) ;
  assign n2209 = ~n2141 & n2208 ;
  assign n2210 = ( n2198 & ~n2203 ) | ( n2198 & n2209 ) | ( ~n2203 & n2209 ) ;
  assign n2211 = ~n2198 & n2210 ;
  assign n2212 = x100 & n2175 ;
  assign n2213 = ~n2211 & n2212 ;
  assign n2214 = x38 & ~n2175 ;
  assign n2215 = x216 | x228 ;
  assign n2216 = n2141 | n2215 ;
  assign n2217 = x39 & n1292 ;
  assign n2218 = x40 & n1273 ;
  assign n2219 = n1381 | n2218 ;
  assign n2220 = n1400 | n1693 ;
  assign n2221 = x70 | n1580 ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2223 = x51 | n2222 ;
  assign n2224 = ~n1435 & n2223 ;
  assign n2225 = n1773 | n2224 ;
  assign n2226 = ~n1432 & n2225 ;
  assign n2227 = ( n1274 & ~n2219 ) | ( n1274 & n2226 ) | ( ~n2219 & n2226 ) ;
  assign n2228 = ~n2219 & n2227 ;
  assign n2229 = x95 | n2228 ;
  assign n2230 = ~n1422 & n2229 ;
  assign n2231 = x39 | n2230 ;
  assign n2232 = ~n2217 & n2231 ;
  assign n2233 = n2179 & ~n2232 ;
  assign n2234 = ( n2179 & n2216 ) | ( n2179 & n2233 ) | ( n2216 & n2233 ) ;
  assign n2235 = ( ~x154 & n2173 ) | ( ~x154 & n2234 ) | ( n2173 & n2234 ) ;
  assign n2236 = ~x154 & n2235 ;
  assign n2237 = ( x38 & n2185 ) | ( x38 & ~n2236 ) | ( n2185 & ~n2236 ) ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = ( x100 & ~n2214 ) | ( x100 & n2238 ) | ( ~n2214 & n2238 ) ;
  assign n2240 = ~x100 & n2239 ;
  assign n2241 = ( x87 & ~n2213 ) | ( x87 & n2240 ) | ( ~n2213 & n2240 ) ;
  assign n2242 = n2213 | n2241 ;
  assign n2243 = n2242 ^ n2194 ^ 1'b0 ;
  assign n2244 = ( n2194 & n2242 ) | ( n2194 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = ( x75 & ~n2194 ) | ( x75 & n2244 ) | ( ~n2194 & n2244 ) ;
  assign n2246 = ( x92 & ~n2191 ) | ( x92 & n2245 ) | ( ~n2191 & n2245 ) ;
  assign n2247 = ~x92 & n2246 ;
  assign n2248 = ( n2067 & ~n2190 ) | ( n2067 & n2247 ) | ( ~n2190 & n2247 ) ;
  assign n2249 = n2190 | n2248 ;
  assign n2250 = ( x55 & ~n2176 ) | ( x55 & n2249 ) | ( ~n2176 & n2249 ) ;
  assign n2251 = ~x55 & n2250 ;
  assign n2252 = x55 & ~n2138 ;
  assign n2253 = n2252 ^ x56 ^ 1'b0 ;
  assign n2254 = n2070 | n2146 ;
  assign n2255 = ( n2252 & ~n2253 ) | ( n2252 & n2254 ) | ( ~n2253 & n2254 ) ;
  assign n2256 = ( x56 & n2253 ) | ( x56 & n2255 ) | ( n2253 & n2255 ) ;
  assign n2257 = ( ~n2159 & n2251 ) | ( ~n2159 & n2256 ) | ( n2251 & n2256 ) ;
  assign n2258 = ~n2159 & n2257 ;
  assign n2259 = ( n2120 & ~n2154 ) | ( n2120 & n2258 ) | ( ~n2154 & n2258 ) ;
  assign n2260 = n2154 | n2259 ;
  assign n2261 = ( x239 & ~n2139 ) | ( x239 & n2260 ) | ( ~n2139 & n2260 ) ;
  assign n2262 = ~x239 & n2261 ;
  assign n2263 = x216 | x221 ;
  assign n2264 = x215 | n2263 ;
  assign n2265 = n1224 & n1323 ;
  assign n2266 = ~n2264 & n2265 ;
  assign n2267 = n2136 | n2266 ;
  assign n2268 = x154 & n2267 ;
  assign n2269 = ~x215 & n2267 ;
  assign n2270 = x154 | n2133 ;
  assign n2271 = ( n2268 & ~n2269 ) | ( n2268 & n2270 ) | ( ~n2269 & n2270 ) ;
  assign n2272 = ~n2268 & n2271 ;
  assign n2273 = n2120 & n2272 ;
  assign n2274 = x239 & ~n2273 ;
  assign n2275 = n2274 ^ n2262 ^ 1'b0 ;
  assign n2276 = n2144 | n2268 ;
  assign n2277 = ~n2272 & n2276 ;
  assign n2278 = ~n2147 & n2277 ;
  assign n2279 = ~x56 & n2278 ;
  assign n2280 = n2151 & ~n2272 ;
  assign n2281 = ( x62 & n2279 ) | ( x62 & n2280 ) | ( n2279 & n2280 ) ;
  assign n2282 = n2280 ^ n2279 ^ 1'b0 ;
  assign n2283 = ( x62 & n2281 ) | ( x62 & n2282 ) | ( n2281 & n2282 ) ;
  assign n2284 = n2099 & ~n2272 ;
  assign n2285 = x56 & ~n2284 ;
  assign n2286 = n2285 ^ n2278 ^ 1'b0 ;
  assign n2287 = ( n2278 & n2285 ) | ( n2278 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = ( x62 & ~n2278 ) | ( x62 & n2287 ) | ( ~n2278 & n2287 ) ;
  assign n2289 = x299 & ~n2272 ;
  assign n2290 = x223 | x299 ;
  assign n2291 = n1359 | n2290 ;
  assign n2292 = n1224 & ~n2291 ;
  assign n2293 = n2173 | n2292 ;
  assign n2294 = n2289 | n2293 ;
  assign n2295 = n2067 & ~n2294 ;
  assign n2296 = x92 & n2294 ;
  assign n2297 = x299 & ~n2277 ;
  assign n2298 = ~n2177 & n2297 ;
  assign n2299 = n2296 & ~n2298 ;
  assign n2300 = x75 & ~n2294 ;
  assign n2301 = x87 & n2294 ;
  assign n2302 = ~n2036 & n2297 ;
  assign n2303 = n2301 & ~n2302 ;
  assign n2304 = n2294 & ~n2297 ;
  assign n2305 = x39 & ~n2304 ;
  assign n2306 = x72 | n2224 ;
  assign n2307 = ~n1432 & n2306 ;
  assign n2308 = n1274 | n2307 ;
  assign n2309 = ~n2219 & n2308 ;
  assign n2310 = x95 | n2309 ;
  assign n2311 = ~n1648 & n2310 ;
  assign n2312 = ~x228 & n2311 ;
  assign n2313 = ~n1290 & n1427 ;
  assign n2314 = n1224 | n2313 ;
  assign n2315 = n1323 & ~n2314 ;
  assign n2316 = n2312 | n2315 ;
  assign n2317 = ~x154 & n2316 ;
  assign n2318 = x105 & n2314 ;
  assign n2319 = ~n1422 & n2314 ;
  assign n2320 = n2318 ^ x228 ^ 1'b0 ;
  assign n2321 = ( n2318 & n2319 ) | ( n2318 & ~n2320 ) | ( n2319 & ~n2320 ) ;
  assign n2322 = x154 & ~n2321 ;
  assign n2323 = ( n2264 & ~n2317 ) | ( n2264 & n2322 ) | ( ~n2317 & n2322 ) ;
  assign n2324 = n2317 | n2323 ;
  assign n2325 = n2183 & n2324 ;
  assign n2326 = x224 | n2314 ;
  assign n2327 = ( n2166 & ~n2169 ) | ( n2166 & n2326 ) | ( ~n2169 & n2326 ) ;
  assign n2328 = n2327 ^ n2160 ^ 1'b0 ;
  assign n2329 = ( n2160 & n2327 ) | ( n2160 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = ( x299 & ~n2160 ) | ( x299 & n2329 ) | ( ~n2160 & n2329 ) ;
  assign n2331 = n2330 ^ n2325 ^ 1'b0 ;
  assign n2332 = ( n2325 & n2330 ) | ( n2325 & n2331 ) | ( n2330 & n2331 ) ;
  assign n2333 = ( x39 & ~n2325 ) | ( x39 & n2332 ) | ( ~n2325 & n2332 ) ;
  assign n2334 = ( n1205 & ~n2305 ) | ( n1205 & n2333 ) | ( ~n2305 & n2333 ) ;
  assign n2335 = ~n1205 & n2334 ;
  assign n2336 = n1205 & n2294 ;
  assign n2337 = x100 & n2211 ;
  assign n2338 = n2336 & ~n2337 ;
  assign n2339 = ( ~x87 & n2335 ) | ( ~x87 & n2338 ) | ( n2335 & n2338 ) ;
  assign n2340 = ~x87 & n2339 ;
  assign n2341 = ( x75 & ~n2303 ) | ( x75 & n2340 ) | ( ~n2303 & n2340 ) ;
  assign n2342 = n2303 | n2341 ;
  assign n2343 = ( x92 & ~n2300 ) | ( x92 & n2342 ) | ( ~n2300 & n2342 ) ;
  assign n2344 = ~x92 & n2343 ;
  assign n2345 = ( n2067 & ~n2299 ) | ( n2067 & n2344 ) | ( ~n2299 & n2344 ) ;
  assign n2346 = n2299 | n2345 ;
  assign n2347 = ( x55 & ~n2295 ) | ( x55 & n2346 ) | ( ~n2295 & n2346 ) ;
  assign n2348 = ~x55 & n2347 ;
  assign n2349 = x55 & ~n2272 ;
  assign n2350 = n2349 ^ x56 ^ 1'b0 ;
  assign n2351 = n2070 | n2276 ;
  assign n2352 = ( n2349 & ~n2350 ) | ( n2349 & n2351 ) | ( ~n2350 & n2351 ) ;
  assign n2353 = ( x56 & n2350 ) | ( x56 & n2352 ) | ( n2350 & n2352 ) ;
  assign n2354 = ( ~n2288 & n2348 ) | ( ~n2288 & n2353 ) | ( n2348 & n2353 ) ;
  assign n2355 = ~n2288 & n2354 ;
  assign n2356 = ( n2120 & ~n2283 ) | ( n2120 & n2355 ) | ( ~n2283 & n2355 ) ;
  assign n2357 = n2283 | n2356 ;
  assign n2358 = ( n2274 & ~n2275 ) | ( n2274 & n2357 ) | ( ~n2275 & n2357 ) ;
  assign n2359 = ( n2262 & n2275 ) | ( n2262 & n2358 ) | ( n2275 & n2358 ) ;
  assign n2360 = x1145 ^ x215 ^ 1'b0 ;
  assign n2361 = ~x927 & n1315 ;
  assign n2362 = x1145 | n1315 ;
  assign n2363 = ( x221 & n2361 ) | ( x221 & n2362 ) | ( n2361 & n2362 ) ;
  assign n2364 = ~n2361 & n2363 ;
  assign n2365 = x216 & x274 ;
  assign n2366 = x221 | n2365 ;
  assign n2367 = x151 & ~n1323 ;
  assign n2368 = ( ~x216 & n1323 ) | ( ~x216 & n2367 ) | ( n1323 & n2367 ) ;
  assign n2369 = ( ~n2364 & n2366 ) | ( ~n2364 & n2368 ) | ( n2366 & n2368 ) ;
  assign n2370 = ~n2364 & n2369 ;
  assign n2371 = ( ~x1145 & n2360 ) | ( ~x1145 & n2370 ) | ( n2360 & n2370 ) ;
  assign n2372 = ~n2022 & n2265 ;
  assign n2373 = ~n2365 & n2372 ;
  assign n2374 = n2371 & ~n2373 ;
  assign n2375 = n2151 & n2374 ;
  assign n2376 = ~n1224 & n1323 ;
  assign n2377 = n2367 | n2376 ;
  assign n2378 = x151 | n2142 ;
  assign n2379 = n2378 ^ n2377 ^ 1'b0 ;
  assign n2380 = ( n2377 & n2378 ) | ( n2377 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = ( x216 & ~n2377 ) | ( x216 & n2380 ) | ( ~n2377 & n2380 ) ;
  assign n2382 = ~n2366 & n2381 ;
  assign n2383 = n2364 | n2382 ;
  assign n2384 = ( x1145 & ~n2360 ) | ( x1145 & n2383 ) | ( ~n2360 & n2383 ) ;
  assign n2385 = n2151 | n2384 ;
  assign n2386 = ( x62 & n2375 ) | ( x62 & n2385 ) | ( n2375 & n2385 ) ;
  assign n2387 = ~n2375 & n2386 ;
  assign n2388 = x235 & ~n2120 ;
  assign n2389 = x223 & ~x1145 ;
  assign n2390 = x224 & x274 ;
  assign n2391 = n2161 & ~n2390 ;
  assign n2392 = x1145 | n1208 ;
  assign n2393 = ( x222 & x927 ) | ( x222 & n1219 ) | ( x927 & n1219 ) ;
  assign n2394 = n2392 & n2393 ;
  assign n2395 = ( x223 & ~n2391 ) | ( x223 & n2394 ) | ( ~n2391 & n2394 ) ;
  assign n2396 = n2391 | n2395 ;
  assign n2397 = ( x299 & ~n2389 ) | ( x299 & n2396 ) | ( ~n2389 & n2396 ) ;
  assign n2398 = ~x299 & n2397 ;
  assign n2399 = n2292 | n2398 ;
  assign n2400 = x299 & ~n2374 ;
  assign n2401 = n2399 | n2400 ;
  assign n2402 = n1994 & ~n2401 ;
  assign n2403 = x215 & x1145 ;
  assign n2404 = n2198 | n2203 ;
  assign n2405 = x228 | n2404 ;
  assign n2406 = ~n2376 & n2405 ;
  assign n2407 = ~x151 & n2406 ;
  assign n2408 = ( ~n2366 & n2381 ) | ( ~n2366 & n2407 ) | ( n2381 & n2407 ) ;
  assign n2409 = ~n2366 & n2408 ;
  assign n2410 = ( ~x215 & n2364 ) | ( ~x215 & n2409 ) | ( n2364 & n2409 ) ;
  assign n2411 = ~x215 & n2410 ;
  assign n2412 = ( x299 & n2403 ) | ( x299 & n2411 ) | ( n2403 & n2411 ) ;
  assign n2413 = n2411 ^ n2403 ^ 1'b0 ;
  assign n2414 = ( x299 & n2412 ) | ( x299 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2415 = ( n1994 & n2399 ) | ( n1994 & ~n2414 ) | ( n2399 & ~n2414 ) ;
  assign n2416 = n2414 | n2415 ;
  assign n2417 = ( x100 & n2402 ) | ( x100 & n2416 ) | ( n2402 & n2416 ) ;
  assign n2418 = ~n2402 & n2417 ;
  assign n2419 = x299 & ~n2403 ;
  assign n2420 = x151 & n2321 ;
  assign n2421 = x216 | n2420 ;
  assign n2422 = ( x151 & n2316 ) | ( x151 & ~n2421 ) | ( n2316 & ~n2421 ) ;
  assign n2423 = ~n2421 & n2422 ;
  assign n2424 = ( x221 & n2365 ) | ( x221 & ~n2423 ) | ( n2365 & ~n2423 ) ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = n2425 ^ n2364 ^ 1'b0 ;
  assign n2427 = ( n2364 & n2425 ) | ( n2364 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2428 = ( x215 & ~n2364 ) | ( x215 & n2427 ) | ( ~n2364 & n2427 ) ;
  assign n2429 = n2419 & n2428 ;
  assign n2430 = x223 & x1145 ;
  assign n2431 = x222 | n2390 ;
  assign n2432 = n2326 & ~n2431 ;
  assign n2433 = ( ~x223 & n2394 ) | ( ~x223 & n2432 ) | ( n2394 & n2432 ) ;
  assign n2434 = ~x223 & n2433 ;
  assign n2435 = ( x299 & ~n2430 ) | ( x299 & n2434 ) | ( ~n2430 & n2434 ) ;
  assign n2436 = n2430 | n2435 ;
  assign n2437 = ( x39 & ~n2429 ) | ( x39 & n2436 ) | ( ~n2429 & n2436 ) ;
  assign n2438 = ~x39 & n2437 ;
  assign n2439 = x299 & n2384 ;
  assign n2440 = n2399 | n2439 ;
  assign n2441 = x39 & n2440 ;
  assign n2442 = ( x38 & ~n2438 ) | ( x38 & n2441 ) | ( ~n2438 & n2441 ) ;
  assign n2443 = n2438 | n2442 ;
  assign n2444 = x38 & ~n2401 ;
  assign n2445 = ( x100 & n2443 ) | ( x100 & ~n2444 ) | ( n2443 & ~n2444 ) ;
  assign n2446 = ~x100 & n2445 ;
  assign n2447 = ( ~x87 & n2418 ) | ( ~x87 & n2446 ) | ( n2418 & n2446 ) ;
  assign n2448 = ~x87 & n2447 ;
  assign n2449 = n2440 ^ n2036 ^ 1'b0 ;
  assign n2450 = ( n2401 & n2440 ) | ( n2401 & n2449 ) | ( n2440 & n2449 ) ;
  assign n2451 = x87 & n2450 ;
  assign n2452 = ( x75 & ~n2448 ) | ( x75 & n2451 ) | ( ~n2448 & n2451 ) ;
  assign n2453 = n2448 | n2452 ;
  assign n2454 = ( x92 & n2046 ) | ( x92 & n2401 ) | ( n2046 & n2401 ) ;
  assign n2455 = n2454 ^ n2067 ^ 1'b0 ;
  assign n2456 = n2044 | n2450 ;
  assign n2457 = ( n2454 & ~n2455 ) | ( n2454 & n2456 ) | ( ~n2455 & n2456 ) ;
  assign n2458 = ( n2067 & n2455 ) | ( n2067 & n2457 ) | ( n2455 & n2457 ) ;
  assign n2459 = x75 & ~n2401 ;
  assign n2460 = x92 | n2459 ;
  assign n2461 = ~n2458 & n2460 ;
  assign n2462 = ( n2453 & n2458 ) | ( n2453 & ~n2461 ) | ( n2458 & ~n2461 ) ;
  assign n2463 = n2070 & n2374 ;
  assign n2464 = x55 & ~n2463 ;
  assign n2465 = n2464 ^ x56 ^ 1'b0 ;
  assign n2466 = n2070 | n2384 ;
  assign n2467 = ( n2464 & ~n2465 ) | ( n2464 & n2466 ) | ( ~n2465 & n2466 ) ;
  assign n2468 = ( x56 & n2465 ) | ( x56 & n2467 ) | ( n2465 & n2467 ) ;
  assign n2469 = n2067 & ~n2401 ;
  assign n2470 = x55 | n2469 ;
  assign n2471 = ~n2468 & n2470 ;
  assign n2472 = ( n2462 & n2468 ) | ( n2462 & ~n2471 ) | ( n2468 & ~n2471 ) ;
  assign n2473 = ~n2099 & n2384 ;
  assign n2474 = n2099 & ~n2374 ;
  assign n2475 = ( x56 & n2473 ) | ( x56 & ~n2474 ) | ( n2473 & ~n2474 ) ;
  assign n2476 = ~n2473 & n2475 ;
  assign n2477 = ( x62 & n2472 ) | ( x62 & ~n2476 ) | ( n2472 & ~n2476 ) ;
  assign n2478 = ~x62 & n2477 ;
  assign n2479 = ( n2387 & n2388 ) | ( n2387 & ~n2478 ) | ( n2388 & ~n2478 ) ;
  assign n2480 = ~n2387 & n2479 ;
  assign n2481 = x235 & n2373 ;
  assign n2482 = ( n2120 & n2371 ) | ( n2120 & n2481 ) | ( n2371 & n2481 ) ;
  assign n2483 = ~n2481 & n2482 ;
  assign n2484 = x235 | n2120 ;
  assign n2485 = n2364 | n2403 ;
  assign n2486 = n2143 | n2485 ;
  assign n2487 = n2099 | n2486 ;
  assign n2488 = ~n2371 & n2487 ;
  assign n2489 = x56 & ~n2488 ;
  assign n2490 = x55 & ~n2371 ;
  assign n2491 = n2070 | n2486 ;
  assign n2492 = n2490 & n2491 ;
  assign n2493 = x299 & ~n2371 ;
  assign n2494 = n2398 | n2493 ;
  assign n2495 = n2067 & ~n2494 ;
  assign n2496 = n2177 & ~n2494 ;
  assign n2497 = x92 & ~n2496 ;
  assign n2498 = n2486 & n2493 ;
  assign n2499 = n2095 | n2398 ;
  assign n2500 = n2498 | n2499 ;
  assign n2501 = n2044 | n2500 ;
  assign n2502 = n2497 & n2501 ;
  assign n2503 = x75 & ~n2494 ;
  assign n2504 = n2036 & ~n2494 ;
  assign n2505 = x87 & ~n2500 ;
  assign n2506 = ( x87 & n2504 ) | ( x87 & n2505 ) | ( n2504 & n2505 ) ;
  assign n2507 = n2205 | n2485 ;
  assign n2508 = ~x100 & n2232 ;
  assign n2509 = ~x39 & x100 ;
  assign n2510 = ~n2404 & n2509 ;
  assign n2511 = n2508 | n2510 ;
  assign n2512 = n2493 & ~n2511 ;
  assign n2513 = ( n2493 & n2507 ) | ( n2493 & n2512 ) | ( n2507 & n2512 ) ;
  assign n2514 = ( x87 & n2398 ) | ( x87 & ~n2513 ) | ( n2398 & ~n2513 ) ;
  assign n2515 = n2513 | n2514 ;
  assign n2516 = n2515 ^ n2506 ^ 1'b0 ;
  assign n2517 = ( n2506 & n2515 ) | ( n2506 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = ( x75 & ~n2506 ) | ( x75 & n2517 ) | ( ~n2506 & n2517 ) ;
  assign n2519 = ( x92 & ~n2503 ) | ( x92 & n2518 ) | ( ~n2503 & n2518 ) ;
  assign n2520 = ~x92 & n2519 ;
  assign n2521 = ( n2067 & ~n2502 ) | ( n2067 & n2520 ) | ( ~n2502 & n2520 ) ;
  assign n2522 = n2502 | n2521 ;
  assign n2523 = ( x55 & ~n2495 ) | ( x55 & n2522 ) | ( ~n2495 & n2522 ) ;
  assign n2524 = ~x55 & n2523 ;
  assign n2525 = ( x56 & ~n2492 ) | ( x56 & n2524 ) | ( ~n2492 & n2524 ) ;
  assign n2526 = n2492 | n2525 ;
  assign n2527 = ( x62 & ~n2489 ) | ( x62 & n2526 ) | ( ~n2489 & n2526 ) ;
  assign n2528 = ~x62 & n2527 ;
  assign n2529 = x62 & ~n2371 ;
  assign n2530 = x56 | n2487 ;
  assign n2531 = n2529 & n2530 ;
  assign n2532 = ( ~n2484 & n2528 ) | ( ~n2484 & n2531 ) | ( n2528 & n2531 ) ;
  assign n2533 = n2484 | n2532 ;
  assign n2534 = ( n2480 & ~n2483 ) | ( n2480 & n2533 ) | ( ~n2483 & n2533 ) ;
  assign n2535 = ~n2480 & n2534 ;
  assign n2536 = x1143 ^ x215 ^ 1'b0 ;
  assign n2537 = ~x944 & n1315 ;
  assign n2538 = x1143 | n1315 ;
  assign n2539 = ( x221 & n2537 ) | ( x221 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2540 = ~n2537 & n2539 ;
  assign n2541 = x216 & x264 ;
  assign n2542 = x221 | n2541 ;
  assign n2543 = ~x105 & x146 ;
  assign n2544 = x284 & ~n1224 ;
  assign n2545 = x105 & ~n2544 ;
  assign n2546 = ( x228 & n2543 ) | ( x228 & ~n2545 ) | ( n2543 & ~n2545 ) ;
  assign n2547 = ~n2543 & n2546 ;
  assign n2548 = n2265 | n2547 ;
  assign n2549 = x146 | x228 ;
  assign n2550 = ~n2548 & n2549 ;
  assign n2551 = x216 | n2550 ;
  assign n2552 = n2551 ^ n2542 ^ 1'b0 ;
  assign n2553 = ( n2542 & n2551 ) | ( n2542 & n2552 ) | ( n2551 & n2552 ) ;
  assign n2554 = ( n2540 & ~n2542 ) | ( n2540 & n2553 ) | ( ~n2542 & n2553 ) ;
  assign n2555 = ( x1143 & ~n2536 ) | ( x1143 & n2554 ) | ( ~n2536 & n2554 ) ;
  assign n2556 = n2372 & ~n2541 ;
  assign n2557 = x238 & n2556 ;
  assign n2558 = ( n2120 & n2555 ) | ( n2120 & ~n2557 ) | ( n2555 & ~n2557 ) ;
  assign n2559 = ~n2555 & n2558 ;
  assign n2560 = n2555 | n2556 ;
  assign n2561 = n2151 & ~n2560 ;
  assign n2562 = x215 & x1143 ;
  assign n2563 = ( ~x146 & x284 ) | ( ~x146 & n2196 ) | ( x284 & n2196 ) ;
  assign n2564 = ~x228 & n2563 ;
  assign n2565 = n2547 | n2564 ;
  assign n2566 = ~x216 & n2565 ;
  assign n2567 = ( ~n2540 & n2542 ) | ( ~n2540 & n2566 ) | ( n2542 & n2566 ) ;
  assign n2568 = ~n2540 & n2567 ;
  assign n2569 = x215 | n2568 ;
  assign n2570 = ~n2562 & n2569 ;
  assign n2571 = ~n2151 & n2570 ;
  assign n2572 = ( x62 & n2561 ) | ( x62 & ~n2571 ) | ( n2561 & ~n2571 ) ;
  assign n2573 = ~n2561 & n2572 ;
  assign n2574 = x238 & ~n2120 ;
  assign n2575 = n2099 & n2560 ;
  assign n2576 = n2099 | n2570 ;
  assign n2577 = ( x56 & n2575 ) | ( x56 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2578 = ~n2575 & n2577 ;
  assign n2579 = ~n2070 & n2570 ;
  assign n2580 = n2070 & ~n2555 ;
  assign n2581 = x55 & ~n2580 ;
  assign n2582 = ( x55 & n2556 ) | ( x55 & n2581 ) | ( n2556 & n2581 ) ;
  assign n2583 = n2582 ^ n2579 ^ 1'b0 ;
  assign n2584 = ( n2579 & n2582 ) | ( n2579 & n2583 ) | ( n2582 & n2583 ) ;
  assign n2585 = ( x56 & ~n2579 ) | ( x56 & n2584 ) | ( ~n2579 & n2584 ) ;
  assign n2586 = x223 & x1143 ;
  assign n2587 = ~x944 & n1208 ;
  assign n2588 = x1143 | n1208 ;
  assign n2589 = ( x222 & n2587 ) | ( x222 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2590 = ~n2587 & n2589 ;
  assign n2591 = ~x224 & n2544 ;
  assign n2592 = ( x222 & x264 ) | ( x222 & n1359 ) | ( x264 & n1359 ) ;
  assign n2593 = ( ~n2590 & n2591 ) | ( ~n2590 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2594 = ~n2590 & n2593 ;
  assign n2595 = x223 | n2594 ;
  assign n2596 = n2595 ^ n2586 ^ 1'b0 ;
  assign n2597 = ( n2586 & n2595 ) | ( n2586 & n2596 ) | ( n2595 & n2596 ) ;
  assign n2598 = ( x299 & ~n2586 ) | ( x299 & n2597 ) | ( ~n2586 & n2597 ) ;
  assign n2599 = x299 & n2560 ;
  assign n2600 = n2598 & ~n2599 ;
  assign n2601 = n2044 & n2600 ;
  assign n2602 = x299 & ~n2570 ;
  assign n2603 = n2598 & ~n2602 ;
  assign n2604 = n2603 ^ n2036 ^ 1'b0 ;
  assign n2605 = ( n2600 & n2603 ) | ( n2600 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = ~n2044 & n2605 ;
  assign n2607 = ( x92 & n2601 ) | ( x92 & ~n2606 ) | ( n2601 & ~n2606 ) ;
  assign n2608 = ~n2601 & n2607 ;
  assign n2609 = x75 & n2600 ;
  assign n2610 = x87 & ~n2605 ;
  assign n2611 = x252 & ~n1329 ;
  assign n2612 = x284 | n2611 ;
  assign n2613 = ~x228 & n1292 ;
  assign n2614 = ( ~x228 & n2612 ) | ( ~x228 & n2613 ) | ( n2612 & n2613 ) ;
  assign n2615 = ( x146 & n2195 ) | ( x146 & ~n2614 ) | ( n2195 & ~n2614 ) ;
  assign n2616 = n2615 ^ n2614 ^ 1'b0 ;
  assign n2617 = ( n2614 & ~n2615 ) | ( n2614 & n2616 ) | ( ~n2615 & n2616 ) ;
  assign n2618 = n2547 | n2617 ;
  assign n2619 = x216 | n2618 ;
  assign n2620 = ( ~x216 & n2542 ) | ( ~x216 & n2619 ) | ( n2542 & n2619 ) ;
  assign n2621 = n2620 ^ n2540 ^ 1'b0 ;
  assign n2622 = ( n2540 & n2620 ) | ( n2540 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2623 = ( x215 & ~n2540 ) | ( x215 & n2622 ) | ( ~n2540 & n2622 ) ;
  assign n2624 = n2623 ^ n2562 ^ 1'b0 ;
  assign n2625 = ( x299 & n2562 ) | ( x299 & ~n2623 ) | ( n2562 & ~n2623 ) ;
  assign n2626 = ( x299 & ~n2624 ) | ( x299 & n2625 ) | ( ~n2624 & n2625 ) ;
  assign n2627 = ( n1994 & n2598 ) | ( n1994 & ~n2626 ) | ( n2598 & ~n2626 ) ;
  assign n2628 = ~n1994 & n2627 ;
  assign n2629 = n1994 & n2600 ;
  assign n2630 = ( x100 & n2628 ) | ( x100 & ~n2629 ) | ( n2628 & ~n2629 ) ;
  assign n2631 = ~n2628 & n2630 ;
  assign n2632 = x38 & n2600 ;
  assign n2633 = x39 & ~n2603 ;
  assign n2634 = ~n2318 & n2547 ;
  assign n2635 = ~x146 & n2319 ;
  assign n2636 = x146 & ~n2311 ;
  assign n2637 = ( x284 & n2635 ) | ( x284 & ~n2636 ) | ( n2635 & ~n2636 ) ;
  assign n2638 = ~n2635 & n2637 ;
  assign n2639 = x146 | x284 ;
  assign n2640 = n2230 | n2639 ;
  assign n2641 = n2640 ^ n2638 ^ 1'b0 ;
  assign n2642 = ( n2638 & n2640 ) | ( n2638 & n2641 ) | ( n2640 & n2641 ) ;
  assign n2643 = ( x228 & ~n2638 ) | ( x228 & n2642 ) | ( ~n2638 & n2642 ) ;
  assign n2644 = n2643 ^ n2634 ^ 1'b0 ;
  assign n2645 = ( n2634 & n2643 ) | ( n2634 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2646 = ( x216 & ~n2634 ) | ( x216 & n2645 ) | ( ~n2634 & n2645 ) ;
  assign n2647 = ( x221 & ~n2541 ) | ( x221 & n2646 ) | ( ~n2541 & n2646 ) ;
  assign n2648 = ~x221 & n2647 ;
  assign n2649 = ( ~x215 & n2540 ) | ( ~x215 & n2648 ) | ( n2540 & n2648 ) ;
  assign n2650 = ~x215 & n2649 ;
  assign n2651 = ( x299 & n2562 ) | ( x299 & ~n2650 ) | ( n2562 & ~n2650 ) ;
  assign n2652 = ~n2562 & n2651 ;
  assign n2653 = x299 | n2586 ;
  assign n2654 = ( ~x224 & n2314 ) | ( ~x224 & n2591 ) | ( n2314 & n2591 ) ;
  assign n2655 = ( ~n2590 & n2592 ) | ( ~n2590 & n2654 ) | ( n2592 & n2654 ) ;
  assign n2656 = ~n2590 & n2655 ;
  assign n2657 = n2314 & ~n2592 ;
  assign n2658 = n2656 & ~n2657 ;
  assign n2659 = x223 | n2658 ;
  assign n2660 = ~n2653 & n2659 ;
  assign n2661 = ( x39 & ~n2652 ) | ( x39 & n2660 ) | ( ~n2652 & n2660 ) ;
  assign n2662 = n2652 | n2661 ;
  assign n2663 = ( x38 & ~n2633 ) | ( x38 & n2662 ) | ( ~n2633 & n2662 ) ;
  assign n2664 = ~x38 & n2663 ;
  assign n2665 = ( x100 & ~n2632 ) | ( x100 & n2664 ) | ( ~n2632 & n2664 ) ;
  assign n2666 = n2632 | n2665 ;
  assign n2667 = n2666 ^ n2631 ^ 1'b0 ;
  assign n2668 = ( n2631 & n2666 ) | ( n2631 & n2667 ) | ( n2666 & n2667 ) ;
  assign n2669 = ( x87 & ~n2631 ) | ( x87 & n2668 ) | ( ~n2631 & n2668 ) ;
  assign n2670 = ( x75 & ~n2610 ) | ( x75 & n2669 ) | ( ~n2610 & n2669 ) ;
  assign n2671 = ~x75 & n2670 ;
  assign n2672 = ( x92 & ~n2609 ) | ( x92 & n2671 ) | ( ~n2609 & n2671 ) ;
  assign n2673 = n2609 | n2672 ;
  assign n2674 = ( n2067 & ~n2608 ) | ( n2067 & n2673 ) | ( ~n2608 & n2673 ) ;
  assign n2675 = ~n2067 & n2674 ;
  assign n2676 = n2067 & n2600 ;
  assign n2677 = x55 | n2676 ;
  assign n2678 = ( ~n2585 & n2675 ) | ( ~n2585 & n2677 ) | ( n2675 & n2677 ) ;
  assign n2679 = ~n2585 & n2678 ;
  assign n2680 = ( x62 & ~n2578 ) | ( x62 & n2679 ) | ( ~n2578 & n2679 ) ;
  assign n2681 = n2578 | n2680 ;
  assign n2682 = ( n2573 & n2574 ) | ( n2573 & n2681 ) | ( n2574 & n2681 ) ;
  assign n2683 = ~n2573 & n2682 ;
  assign n2684 = n2151 & ~n2555 ;
  assign n2685 = n2548 | n2564 ;
  assign n2686 = ~x216 & n2685 ;
  assign n2687 = ( ~n2540 & n2542 ) | ( ~n2540 & n2686 ) | ( n2542 & n2686 ) ;
  assign n2688 = ~n2540 & n2687 ;
  assign n2689 = ( ~x1143 & n2536 ) | ( ~x1143 & n2688 ) | ( n2536 & n2688 ) ;
  assign n2690 = ~n2151 & n2689 ;
  assign n2691 = ( x62 & n2684 ) | ( x62 & ~n2690 ) | ( n2684 & ~n2690 ) ;
  assign n2692 = ~n2684 & n2691 ;
  assign n2693 = ( x238 & n2120 ) | ( x238 & ~n2692 ) | ( n2120 & ~n2692 ) ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = ~n2070 & n2689 ;
  assign n2696 = n2695 ^ n2581 ^ 1'b0 ;
  assign n2697 = ( n2581 & n2695 ) | ( n2581 & n2696 ) | ( n2695 & n2696 ) ;
  assign n2698 = ( x56 & ~n2695 ) | ( x56 & n2697 ) | ( ~n2695 & n2697 ) ;
  assign n2699 = n1224 & ~n1360 ;
  assign n2700 = n2598 | n2699 ;
  assign n2701 = x299 & n2555 ;
  assign n2702 = n2700 & ~n2701 ;
  assign n2703 = n2044 & n2702 ;
  assign n2704 = x299 & ~n2689 ;
  assign n2705 = n2700 & ~n2704 ;
  assign n2706 = n2705 ^ n2036 ^ 1'b0 ;
  assign n2707 = ( n2702 & n2705 ) | ( n2702 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2708 = ~n2044 & n2707 ;
  assign n2709 = ( x92 & n2703 ) | ( x92 & ~n2708 ) | ( n2703 & ~n2708 ) ;
  assign n2710 = ~n2703 & n2709 ;
  assign n2711 = x75 & n2702 ;
  assign n2712 = x87 & ~n2707 ;
  assign n2713 = n2548 | n2617 ;
  assign n2714 = x216 | n2713 ;
  assign n2715 = ( ~x216 & n2542 ) | ( ~x216 & n2714 ) | ( n2542 & n2714 ) ;
  assign n2716 = n2715 ^ n2540 ^ 1'b0 ;
  assign n2717 = ( n2540 & n2715 ) | ( n2540 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2718 = ( x215 & ~n2540 ) | ( x215 & n2717 ) | ( ~n2540 & n2717 ) ;
  assign n2719 = n2718 ^ n2562 ^ 1'b0 ;
  assign n2720 = ( x299 & n2562 ) | ( x299 & ~n2718 ) | ( n2562 & ~n2718 ) ;
  assign n2721 = ( x299 & ~n2719 ) | ( x299 & n2720 ) | ( ~n2719 & n2720 ) ;
  assign n2722 = ( n1994 & n2700 ) | ( n1994 & ~n2721 ) | ( n2700 & ~n2721 ) ;
  assign n2723 = ~n1994 & n2722 ;
  assign n2724 = n1994 & n2702 ;
  assign n2725 = ( x100 & n2723 ) | ( x100 & ~n2724 ) | ( n2723 & ~n2724 ) ;
  assign n2726 = ~n2723 & n2725 ;
  assign n2727 = x38 & n2702 ;
  assign n2728 = x39 & ~n2705 ;
  assign n2729 = ~n2653 & n2656 ;
  assign n2730 = n2659 ^ n2653 ^ 1'b0 ;
  assign n2731 = ( n2653 & n2659 ) | ( n2653 & n2730 ) | ( n2659 & n2730 ) ;
  assign n2732 = ( x39 & ~n2653 ) | ( x39 & n2731 ) | ( ~n2653 & n2731 ) ;
  assign n2733 = x146 | n2311 ;
  assign n2734 = x146 & x284 ;
  assign n2735 = ~n2230 & n2734 ;
  assign n2736 = x146 & n2319 ;
  assign n2737 = ( x284 & ~n2735 ) | ( x284 & n2736 ) | ( ~n2735 & n2736 ) ;
  assign n2738 = ~n2735 & n2737 ;
  assign n2739 = ( x228 & n2733 ) | ( x228 & ~n2738 ) | ( n2733 & ~n2738 ) ;
  assign n2740 = n2739 ^ n2733 ^ 1'b0 ;
  assign n2741 = ( x228 & n2739 ) | ( x228 & ~n2740 ) | ( n2739 & ~n2740 ) ;
  assign n2742 = n1323 & n2314 ;
  assign n2743 = ( n2547 & n2741 ) | ( n2547 & ~n2742 ) | ( n2741 & ~n2742 ) ;
  assign n2744 = ~n2547 & n2743 ;
  assign n2745 = x216 | n2744 ;
  assign n2746 = ~n2542 & n2745 ;
  assign n2747 = ( ~x215 & n2540 ) | ( ~x215 & n2746 ) | ( n2540 & n2746 ) ;
  assign n2748 = ~x215 & n2747 ;
  assign n2749 = ( x299 & n2562 ) | ( x299 & ~n2748 ) | ( n2562 & ~n2748 ) ;
  assign n2750 = ~n2562 & n2749 ;
  assign n2751 = ( ~n2729 & n2732 ) | ( ~n2729 & n2750 ) | ( n2732 & n2750 ) ;
  assign n2752 = n2729 | n2751 ;
  assign n2753 = ( x38 & ~n2728 ) | ( x38 & n2752 ) | ( ~n2728 & n2752 ) ;
  assign n2754 = ~x38 & n2753 ;
  assign n2755 = ( x100 & ~n2727 ) | ( x100 & n2754 ) | ( ~n2727 & n2754 ) ;
  assign n2756 = n2727 | n2755 ;
  assign n2757 = n2756 ^ n2726 ^ 1'b0 ;
  assign n2758 = ( n2726 & n2756 ) | ( n2726 & n2757 ) | ( n2756 & n2757 ) ;
  assign n2759 = ( x87 & ~n2726 ) | ( x87 & n2758 ) | ( ~n2726 & n2758 ) ;
  assign n2760 = ( x75 & ~n2712 ) | ( x75 & n2759 ) | ( ~n2712 & n2759 ) ;
  assign n2761 = ~x75 & n2760 ;
  assign n2762 = ( x92 & ~n2711 ) | ( x92 & n2761 ) | ( ~n2711 & n2761 ) ;
  assign n2763 = n2711 | n2762 ;
  assign n2764 = ( n2067 & ~n2710 ) | ( n2067 & n2763 ) | ( ~n2710 & n2763 ) ;
  assign n2765 = ~n2067 & n2764 ;
  assign n2766 = n2067 & n2702 ;
  assign n2767 = x55 | n2766 ;
  assign n2768 = ( ~n2698 & n2765 ) | ( ~n2698 & n2767 ) | ( n2765 & n2767 ) ;
  assign n2769 = ~n2698 & n2768 ;
  assign n2770 = n2099 | n2689 ;
  assign n2771 = n2770 ^ x62 ^ 1'b0 ;
  assign n2772 = n2099 & n2555 ;
  assign n2773 = x56 & ~n2772 ;
  assign n2774 = ( n2770 & ~n2771 ) | ( n2770 & n2773 ) | ( ~n2771 & n2773 ) ;
  assign n2775 = ( x62 & n2771 ) | ( x62 & n2774 ) | ( n2771 & n2774 ) ;
  assign n2776 = ( ~n2694 & n2769 ) | ( ~n2694 & n2775 ) | ( n2769 & n2775 ) ;
  assign n2777 = ~n2694 & n2776 ;
  assign n2778 = ( ~n2559 & n2683 ) | ( ~n2559 & n2777 ) | ( n2683 & n2777 ) ;
  assign n2779 = n2559 | n2778 ;
  assign n2780 = x172 & ~x228 ;
  assign n2781 = n2142 & ~n2780 ;
  assign n2782 = x262 | n1292 ;
  assign n2783 = ~n2781 & n2782 ;
  assign n2784 = x215 & x1142 ;
  assign n2785 = ~x932 & n1315 ;
  assign n2786 = x1142 | n1315 ;
  assign n2787 = ( x221 & n2785 ) | ( x221 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2788 = ~n2785 & n2787 ;
  assign n2789 = x216 & x277 ;
  assign n2790 = x221 | n2789 ;
  assign n2791 = x262 & ~n1224 ;
  assign n2792 = x105 & n2791 ;
  assign n2793 = ~x105 & x172 ;
  assign n2794 = ( x228 & n2792 ) | ( x228 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2795 = ( ~x216 & n2780 ) | ( ~x216 & n2794 ) | ( n2780 & n2794 ) ;
  assign n2796 = ( ~n2788 & n2790 ) | ( ~n2788 & n2795 ) | ( n2790 & n2795 ) ;
  assign n2797 = ~n2788 & n2796 ;
  assign n2798 = x215 | n2797 ;
  assign n2799 = ~n2784 & n2798 ;
  assign n2800 = n2265 | n2794 ;
  assign n2801 = n2783 | n2800 ;
  assign n2802 = ~x216 & n2801 ;
  assign n2803 = ( ~n2788 & n2790 ) | ( ~n2788 & n2802 ) | ( n2790 & n2802 ) ;
  assign n2804 = ~n2788 & n2803 ;
  assign n2805 = x215 | n2804 ;
  assign n2806 = ~n2784 & n2805 ;
  assign n2807 = ( n2783 & n2799 ) | ( n2783 & n2806 ) | ( n2799 & n2806 ) ;
  assign n2808 = ~n2151 & n2807 ;
  assign n2809 = n2151 & n2799 ;
  assign n2810 = ( x62 & n2808 ) | ( x62 & ~n2809 ) | ( n2808 & ~n2809 ) ;
  assign n2811 = ~n2808 & n2810 ;
  assign n2812 = n2099 & ~n2799 ;
  assign n2813 = n2099 | n2807 ;
  assign n2814 = ( x56 & n2812 ) | ( x56 & n2813 ) | ( n2812 & n2813 ) ;
  assign n2815 = ~n2812 & n2814 ;
  assign n2816 = ~n2070 & n2807 ;
  assign n2817 = n2070 & n2799 ;
  assign n2818 = x55 & ~n2817 ;
  assign n2819 = n2818 ^ n2816 ^ 1'b0 ;
  assign n2820 = ( n2816 & n2818 ) | ( n2816 & n2819 ) | ( n2818 & n2819 ) ;
  assign n2821 = ( x56 & ~n2816 ) | ( x56 & n2820 ) | ( ~n2816 & n2820 ) ;
  assign n2822 = x223 & x1142 ;
  assign n2823 = ~x932 & n1208 ;
  assign n2824 = x1142 | n1208 ;
  assign n2825 = ( x222 & n2823 ) | ( x222 & n2824 ) | ( n2823 & n2824 ) ;
  assign n2826 = ~n2823 & n2825 ;
  assign n2827 = ~x224 & n2791 ;
  assign n2828 = ( x222 & x277 ) | ( x222 & n1359 ) | ( x277 & n1359 ) ;
  assign n2829 = ( ~n2826 & n2827 ) | ( ~n2826 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2830 = ~n2826 & n2829 ;
  assign n2831 = x223 | n2830 ;
  assign n2832 = n2831 ^ n2822 ^ 1'b0 ;
  assign n2833 = ( n2822 & n2831 ) | ( n2822 & n2832 ) | ( n2831 & n2832 ) ;
  assign n2834 = ( x299 & ~n2822 ) | ( x299 & n2833 ) | ( ~n2822 & n2833 ) ;
  assign n2835 = x299 & ~n2807 ;
  assign n2836 = n2834 & ~n2835 ;
  assign n2837 = x299 & ~n2799 ;
  assign n2838 = n2834 & ~n2837 ;
  assign n2839 = n2836 ^ n2036 ^ 1'b0 ;
  assign n2840 = ( n2836 & n2838 ) | ( n2836 & n2839 ) | ( n2838 & n2839 ) ;
  assign n2841 = ~n2044 & n2840 ;
  assign n2842 = n2044 & n2838 ;
  assign n2843 = ( x92 & n2841 ) | ( x92 & ~n2842 ) | ( n2841 & ~n2842 ) ;
  assign n2844 = ~n2841 & n2843 ;
  assign n2845 = x75 & n2838 ;
  assign n2846 = x87 & ~n2840 ;
  assign n2847 = x299 | n2822 ;
  assign n2848 = ( ~x224 & n2314 ) | ( ~x224 & n2827 ) | ( n2314 & n2827 ) ;
  assign n2849 = ( ~n2826 & n2828 ) | ( ~n2826 & n2848 ) | ( n2828 & n2848 ) ;
  assign n2850 = ~n2826 & n2849 ;
  assign n2851 = n2314 & ~n2828 ;
  assign n2852 = n2850 & ~n2851 ;
  assign n2853 = x223 | n2852 ;
  assign n2854 = n2853 ^ n2847 ^ 1'b0 ;
  assign n2855 = ( n2847 & n2853 ) | ( n2847 & n2854 ) | ( n2853 & n2854 ) ;
  assign n2856 = ( x39 & ~n2847 ) | ( x39 & n2855 ) | ( ~n2847 & n2855 ) ;
  assign n2857 = x299 & ~n2784 ;
  assign n2858 = n2857 ^ n2856 ^ 1'b0 ;
  assign n2859 = ~n2313 & n2792 ;
  assign n2860 = x228 & ~n2793 ;
  assign n2861 = ~n2859 & n2860 ;
  assign n2862 = x262 & n2311 ;
  assign n2863 = x172 | n2862 ;
  assign n2864 = x172 & ~x262 ;
  assign n2865 = ( x172 & n2319 ) | ( x172 & n2864 ) | ( n2319 & n2864 ) ;
  assign n2866 = x262 | n2230 ;
  assign n2867 = n2865 & n2866 ;
  assign n2868 = ( x228 & n2863 ) | ( x228 & ~n2867 ) | ( n2863 & ~n2867 ) ;
  assign n2869 = n2868 ^ n2863 ^ 1'b0 ;
  assign n2870 = ( x228 & n2868 ) | ( x228 & ~n2869 ) | ( n2868 & ~n2869 ) ;
  assign n2871 = ( x216 & ~n2861 ) | ( x216 & n2870 ) | ( ~n2861 & n2870 ) ;
  assign n2872 = ~x216 & n2871 ;
  assign n2873 = ( x221 & n2789 ) | ( x221 & ~n2872 ) | ( n2789 & ~n2872 ) ;
  assign n2874 = n2872 | n2873 ;
  assign n2875 = n2874 ^ n2788 ^ 1'b0 ;
  assign n2876 = ( n2788 & n2874 ) | ( n2788 & n2875 ) | ( n2874 & n2875 ) ;
  assign n2877 = ( x215 & ~n2788 ) | ( x215 & n2876 ) | ( ~n2788 & n2876 ) ;
  assign n2878 = ( n2857 & ~n2858 ) | ( n2857 & n2877 ) | ( ~n2858 & n2877 ) ;
  assign n2879 = ( n2856 & n2858 ) | ( n2856 & n2878 ) | ( n2858 & n2878 ) ;
  assign n2880 = x39 & ~n2836 ;
  assign n2881 = ( x38 & n2879 ) | ( x38 & ~n2880 ) | ( n2879 & ~n2880 ) ;
  assign n2882 = ~x38 & n2881 ;
  assign n2883 = x38 & n2838 ;
  assign n2884 = ( x100 & ~n2882 ) | ( x100 & n2883 ) | ( ~n2882 & n2883 ) ;
  assign n2885 = n2882 | n2884 ;
  assign n2886 = x215 & ~x1142 ;
  assign n2887 = n2405 & ~n2780 ;
  assign n2888 = x262 | n2404 ;
  assign n2889 = ~n2887 & n2888 ;
  assign n2890 = n2794 | n2889 ;
  assign n2891 = x216 | n2890 ;
  assign n2892 = ( ~x216 & n2790 ) | ( ~x216 & n2891 ) | ( n2790 & n2891 ) ;
  assign n2893 = ( x215 & ~n2788 ) | ( x215 & n2892 ) | ( ~n2788 & n2892 ) ;
  assign n2894 = ~x215 & n2893 ;
  assign n2895 = ( x299 & n2886 ) | ( x299 & ~n2894 ) | ( n2886 & ~n2894 ) ;
  assign n2896 = ~n2886 & n2895 ;
  assign n2897 = ( n1994 & n2834 ) | ( n1994 & ~n2896 ) | ( n2834 & ~n2896 ) ;
  assign n2898 = ~n1994 & n2897 ;
  assign n2899 = n1994 & n2838 ;
  assign n2900 = ( x100 & n2898 ) | ( x100 & ~n2899 ) | ( n2898 & ~n2899 ) ;
  assign n2901 = ~n2898 & n2900 ;
  assign n2902 = ( x87 & n2885 ) | ( x87 & ~n2901 ) | ( n2885 & ~n2901 ) ;
  assign n2903 = n2902 ^ n2885 ^ 1'b0 ;
  assign n2904 = ( x87 & n2902 ) | ( x87 & ~n2903 ) | ( n2902 & ~n2903 ) ;
  assign n2905 = ( x75 & ~n2846 ) | ( x75 & n2904 ) | ( ~n2846 & n2904 ) ;
  assign n2906 = ~x75 & n2905 ;
  assign n2907 = ( x92 & ~n2845 ) | ( x92 & n2906 ) | ( ~n2845 & n2906 ) ;
  assign n2908 = n2845 | n2907 ;
  assign n2909 = ( n2067 & ~n2844 ) | ( n2067 & n2908 ) | ( ~n2844 & n2908 ) ;
  assign n2910 = ~n2067 & n2909 ;
  assign n2911 = n2067 & n2838 ;
  assign n2912 = x55 | n2911 ;
  assign n2913 = ( ~n2821 & n2910 ) | ( ~n2821 & n2912 ) | ( n2910 & n2912 ) ;
  assign n2914 = ~n2821 & n2913 ;
  assign n2915 = ( x62 & ~n2815 ) | ( x62 & n2914 ) | ( ~n2815 & n2914 ) ;
  assign n2916 = n2815 | n2915 ;
  assign n2917 = ( n2120 & ~n2811 ) | ( n2120 & n2916 ) | ( ~n2811 & n2916 ) ;
  assign n2918 = ~n2120 & n2917 ;
  assign n2919 = n2120 & n2799 ;
  assign n2920 = ( x249 & n2918 ) | ( x249 & ~n2919 ) | ( n2918 & ~n2919 ) ;
  assign n2921 = ~n2918 & n2920 ;
  assign n2922 = ~n2151 & n2806 ;
  assign n2923 = n2266 | n2799 ;
  assign n2924 = n2151 & n2923 ;
  assign n2925 = ( x62 & n2922 ) | ( x62 & ~n2924 ) | ( n2922 & ~n2924 ) ;
  assign n2926 = ~n2922 & n2925 ;
  assign n2927 = n2099 & ~n2923 ;
  assign n2928 = n2099 | n2806 ;
  assign n2929 = ( x56 & n2927 ) | ( x56 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2930 = ~n2927 & n2929 ;
  assign n2931 = ~n2070 & n2806 ;
  assign n2932 = n2070 & n2923 ;
  assign n2933 = x55 & ~n2932 ;
  assign n2934 = n2933 ^ n2931 ^ 1'b0 ;
  assign n2935 = ( n2931 & n2933 ) | ( n2931 & n2934 ) | ( n2933 & n2934 ) ;
  assign n2936 = ( x56 & ~n2931 ) | ( x56 & n2935 ) | ( ~n2931 & n2935 ) ;
  assign n2937 = n2699 | n2834 ;
  assign n2938 = x299 & ~n2806 ;
  assign n2939 = n2937 & ~n2938 ;
  assign n2940 = x299 & ~n2923 ;
  assign n2941 = n2937 & ~n2940 ;
  assign n2942 = n2939 ^ n2036 ^ 1'b0 ;
  assign n2943 = ( n2939 & n2941 ) | ( n2939 & n2942 ) | ( n2941 & n2942 ) ;
  assign n2944 = ~n2044 & n2943 ;
  assign n2945 = n2044 & n2941 ;
  assign n2946 = ( x92 & n2944 ) | ( x92 & ~n2945 ) | ( n2944 & ~n2945 ) ;
  assign n2947 = ~n2944 & n2946 ;
  assign n2948 = x75 & n2941 ;
  assign n2949 = x87 & ~n2943 ;
  assign n2950 = n2800 | n2889 ;
  assign n2951 = x216 | n2950 ;
  assign n2952 = ( ~x216 & n2790 ) | ( ~x216 & n2951 ) | ( n2790 & n2951 ) ;
  assign n2953 = ( x215 & ~n2788 ) | ( x215 & n2952 ) | ( ~n2788 & n2952 ) ;
  assign n2954 = ~x215 & n2953 ;
  assign n2955 = ( x299 & n2886 ) | ( x299 & ~n2954 ) | ( n2886 & ~n2954 ) ;
  assign n2956 = ~n2886 & n2955 ;
  assign n2957 = ( n1994 & n2937 ) | ( n1994 & ~n2956 ) | ( n2937 & ~n2956 ) ;
  assign n2958 = ~n1994 & n2957 ;
  assign n2959 = n1994 & n2941 ;
  assign n2960 = ( x100 & n2958 ) | ( x100 & ~n2959 ) | ( n2958 & ~n2959 ) ;
  assign n2961 = ~n2958 & n2960 ;
  assign n2962 = x38 & n2941 ;
  assign n2963 = x39 & ~n2939 ;
  assign n2964 = ~n2318 & n2861 ;
  assign n2965 = x262 & n2230 ;
  assign n2966 = n2311 & n2864 ;
  assign n2967 = ~x262 & n2319 ;
  assign n2968 = ( x172 & ~n2966 ) | ( x172 & n2967 ) | ( ~n2966 & n2967 ) ;
  assign n2969 = ~n2966 & n2968 ;
  assign n2970 = ( x228 & ~n2965 ) | ( x228 & n2969 ) | ( ~n2965 & n2969 ) ;
  assign n2971 = n2965 | n2970 ;
  assign n2972 = ( x216 & ~n2964 ) | ( x216 & n2971 ) | ( ~n2964 & n2971 ) ;
  assign n2973 = ~x216 & n2972 ;
  assign n2974 = ( x221 & n2789 ) | ( x221 & ~n2973 ) | ( n2789 & ~n2973 ) ;
  assign n2975 = n2973 | n2974 ;
  assign n2976 = n2975 ^ n2788 ^ 1'b0 ;
  assign n2977 = ( n2788 & n2975 ) | ( n2788 & n2976 ) | ( n2975 & n2976 ) ;
  assign n2978 = ( x215 & ~n2788 ) | ( x215 & n2977 ) | ( ~n2788 & n2977 ) ;
  assign n2979 = n2857 & n2978 ;
  assign n2980 = ~n2847 & n2850 ;
  assign n2981 = ( ~n2856 & n2979 ) | ( ~n2856 & n2980 ) | ( n2979 & n2980 ) ;
  assign n2982 = n2856 | n2981 ;
  assign n2983 = ( x38 & ~n2963 ) | ( x38 & n2982 ) | ( ~n2963 & n2982 ) ;
  assign n2984 = ~x38 & n2983 ;
  assign n2985 = ( x100 & ~n2962 ) | ( x100 & n2984 ) | ( ~n2962 & n2984 ) ;
  assign n2986 = n2962 | n2985 ;
  assign n2987 = n2986 ^ n2961 ^ 1'b0 ;
  assign n2988 = ( n2961 & n2986 ) | ( n2961 & n2987 ) | ( n2986 & n2987 ) ;
  assign n2989 = ( x87 & ~n2961 ) | ( x87 & n2988 ) | ( ~n2961 & n2988 ) ;
  assign n2990 = ( x75 & ~n2949 ) | ( x75 & n2989 ) | ( ~n2949 & n2989 ) ;
  assign n2991 = ~x75 & n2990 ;
  assign n2992 = ( x92 & ~n2948 ) | ( x92 & n2991 ) | ( ~n2948 & n2991 ) ;
  assign n2993 = n2948 | n2992 ;
  assign n2994 = ( n2067 & ~n2947 ) | ( n2067 & n2993 ) | ( ~n2947 & n2993 ) ;
  assign n2995 = ~n2067 & n2994 ;
  assign n2996 = n2067 & n2941 ;
  assign n2997 = x55 | n2996 ;
  assign n2998 = ( ~n2936 & n2995 ) | ( ~n2936 & n2997 ) | ( n2995 & n2997 ) ;
  assign n2999 = ~n2936 & n2998 ;
  assign n3000 = ( x62 & ~n2930 ) | ( x62 & n2999 ) | ( ~n2930 & n2999 ) ;
  assign n3001 = n2930 | n3000 ;
  assign n3002 = ( n2120 & ~n2926 ) | ( n2120 & n3001 ) | ( ~n2926 & n3001 ) ;
  assign n3003 = ~n2120 & n3002 ;
  assign n3004 = n2120 & n2923 ;
  assign n3005 = x249 | n3004 ;
  assign n3006 = ( ~n2921 & n3003 ) | ( ~n2921 & n3005 ) | ( n3003 & n3005 ) ;
  assign n3007 = ~n2921 & n3006 ;
  assign n3008 = x216 & x270 ;
  assign n3009 = n2372 & ~n3008 ;
  assign n3010 = x241 & n3009 ;
  assign n3011 = x215 & x1141 ;
  assign n3012 = ~x935 & n1315 ;
  assign n3013 = x1141 | n1315 ;
  assign n3014 = ( x221 & n3012 ) | ( x221 & n3013 ) | ( n3012 & n3013 ) ;
  assign n3015 = ~n3012 & n3014 ;
  assign n3016 = x221 | n3008 ;
  assign n3017 = ~x105 & x171 ;
  assign n3018 = x861 & ~n1224 ;
  assign n3019 = x105 & ~n3018 ;
  assign n3020 = ( x228 & n3017 ) | ( x228 & ~n3019 ) | ( n3017 & ~n3019 ) ;
  assign n3021 = ~n3017 & n3020 ;
  assign n3022 = x216 | n3021 ;
  assign n3023 = x171 | x228 ;
  assign n3024 = ~n3022 & n3023 ;
  assign n3025 = ( ~n3015 & n3016 ) | ( ~n3015 & n3024 ) | ( n3016 & n3024 ) ;
  assign n3026 = ~n3015 & n3025 ;
  assign n3027 = x215 | n3026 ;
  assign n3028 = ~n3011 & n3027 ;
  assign n3029 = ( n2120 & n3010 ) | ( n2120 & n3028 ) | ( n3010 & n3028 ) ;
  assign n3030 = ~n3010 & n3029 ;
  assign n3031 = x223 & ~x1141 ;
  assign n3032 = x224 | n3018 ;
  assign n3033 = ( x222 & x270 ) | ( x222 & n1359 ) | ( x270 & n1359 ) ;
  assign n3034 = n3032 & ~n3033 ;
  assign n3035 = ~x935 & n1208 ;
  assign n3036 = x1141 | n1208 ;
  assign n3037 = ( x222 & n3035 ) | ( x222 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3038 = ~n3035 & n3037 ;
  assign n3039 = ( x223 & ~n3034 ) | ( x223 & n3038 ) | ( ~n3034 & n3038 ) ;
  assign n3040 = n3034 | n3039 ;
  assign n3041 = ( x299 & ~n3031 ) | ( x299 & n3040 ) | ( ~n3031 & n3040 ) ;
  assign n3042 = ~x299 & n3041 ;
  assign n3043 = x299 & ~n3028 ;
  assign n3044 = n3042 | n3043 ;
  assign n3045 = n1994 & ~n3044 ;
  assign n3046 = x100 & ~n3045 ;
  assign n3047 = x861 | n2404 ;
  assign n3048 = x171 & n2404 ;
  assign n3049 = ( x228 & n3047 ) | ( x228 & ~n3048 ) | ( n3047 & ~n3048 ) ;
  assign n3050 = ~x228 & n3049 ;
  assign n3051 = n3022 | n3050 ;
  assign n3052 = ~n3016 & n3051 ;
  assign n3053 = ( ~x215 & n3015 ) | ( ~x215 & n3052 ) | ( n3015 & n3052 ) ;
  assign n3054 = ~x215 & n3053 ;
  assign n3055 = ( x299 & n3011 ) | ( x299 & n3054 ) | ( n3011 & n3054 ) ;
  assign n3056 = n3054 ^ n3011 ^ 1'b0 ;
  assign n3057 = ( x299 & n3055 ) | ( x299 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3058 = ( n1994 & n3042 ) | ( n1994 & ~n3057 ) | ( n3042 & ~n3057 ) ;
  assign n3059 = n3057 | n3058 ;
  assign n3060 = n3046 & n3059 ;
  assign n3061 = x299 & ~n3011 ;
  assign n3062 = ~n2318 & n3021 ;
  assign n3063 = x171 & n2311 ;
  assign n3064 = x861 & n2319 ;
  assign n3065 = x171 | n3064 ;
  assign n3066 = x861 & ~n3065 ;
  assign n3067 = ( x861 & n3063 ) | ( x861 & n3066 ) | ( n3063 & n3066 ) ;
  assign n3068 = n2230 | n3065 ;
  assign n3069 = n3068 ^ n3067 ^ 1'b0 ;
  assign n3070 = ( n3067 & n3068 ) | ( n3067 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3071 = ( x228 & ~n3067 ) | ( x228 & n3070 ) | ( ~n3067 & n3070 ) ;
  assign n3072 = ( x216 & ~n3062 ) | ( x216 & n3071 ) | ( ~n3062 & n3071 ) ;
  assign n3073 = ~x216 & n3072 ;
  assign n3074 = ( x221 & n3008 ) | ( x221 & ~n3073 ) | ( n3008 & ~n3073 ) ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = n3075 ^ n3015 ^ 1'b0 ;
  assign n3077 = ( n3015 & n3075 ) | ( n3015 & n3076 ) | ( n3075 & n3076 ) ;
  assign n3078 = ( x215 & ~n3015 ) | ( x215 & n3077 ) | ( ~n3015 & n3077 ) ;
  assign n3079 = n3061 & n3078 ;
  assign n3080 = x223 & x1141 ;
  assign n3081 = x299 | n3080 ;
  assign n3082 = x861 & ~n2314 ;
  assign n3083 = x224 | n3082 ;
  assign n3084 = ~n3033 & n3083 ;
  assign n3085 = n3038 | n3084 ;
  assign n3086 = n3081 | n3085 ;
  assign n3087 = n2314 & ~n3033 ;
  assign n3088 = ( ~x223 & n3085 ) | ( ~x223 & n3087 ) | ( n3085 & n3087 ) ;
  assign n3089 = ~x223 & n3088 ;
  assign n3090 = ( ~x39 & n3081 ) | ( ~x39 & n3089 ) | ( n3081 & n3089 ) ;
  assign n3091 = ~x39 & n3090 ;
  assign n3092 = ( n3079 & n3086 ) | ( n3079 & n3091 ) | ( n3086 & n3091 ) ;
  assign n3093 = ~n3079 & n3092 ;
  assign n3094 = x171 & n1292 ;
  assign n3095 = ( ~x228 & x861 ) | ( ~x228 & n2613 ) | ( x861 & n2613 ) ;
  assign n3096 = ~n3094 & n3095 ;
  assign n3097 = n3022 | n3096 ;
  assign n3098 = ~n3016 & n3097 ;
  assign n3099 = n3015 | n3098 ;
  assign n3100 = x215 | n3099 ;
  assign n3101 = ( ~x215 & n3011 ) | ( ~x215 & n3100 ) | ( n3011 & n3100 ) ;
  assign n3102 = x299 & n3101 ;
  assign n3103 = n3042 | n3102 ;
  assign n3104 = x39 & n3103 ;
  assign n3105 = ( x38 & ~n3093 ) | ( x38 & n3104 ) | ( ~n3093 & n3104 ) ;
  assign n3106 = n3093 | n3105 ;
  assign n3107 = x38 & ~n3044 ;
  assign n3108 = ( x100 & n3106 ) | ( x100 & ~n3107 ) | ( n3106 & ~n3107 ) ;
  assign n3109 = ~x100 & n3108 ;
  assign n3110 = ( ~x87 & n3060 ) | ( ~x87 & n3109 ) | ( n3060 & n3109 ) ;
  assign n3111 = ~x87 & n3110 ;
  assign n3112 = n3103 ^ n2036 ^ 1'b0 ;
  assign n3113 = ( n3044 & n3103 ) | ( n3044 & n3112 ) | ( n3103 & n3112 ) ;
  assign n3114 = x87 & n3113 ;
  assign n3115 = ( x75 & ~n3111 ) | ( x75 & n3114 ) | ( ~n3111 & n3114 ) ;
  assign n3116 = n3111 | n3115 ;
  assign n3117 = ( x92 & n2046 ) | ( x92 & n3044 ) | ( n2046 & n3044 ) ;
  assign n3118 = n3117 ^ n2067 ^ 1'b0 ;
  assign n3119 = n2044 | n3113 ;
  assign n3120 = ( n3117 & ~n3118 ) | ( n3117 & n3119 ) | ( ~n3118 & n3119 ) ;
  assign n3121 = ( n2067 & n3118 ) | ( n2067 & n3120 ) | ( n3118 & n3120 ) ;
  assign n3122 = x75 & ~n3044 ;
  assign n3123 = x92 | n3122 ;
  assign n3124 = ~n3121 & n3123 ;
  assign n3125 = ( n3116 & n3121 ) | ( n3116 & ~n3124 ) | ( n3121 & ~n3124 ) ;
  assign n3126 = n2070 | n3101 ;
  assign n3127 = n3126 ^ x56 ^ 1'b0 ;
  assign n3128 = n2070 & n3028 ;
  assign n3129 = x55 & ~n3128 ;
  assign n3130 = ( n3126 & ~n3127 ) | ( n3126 & n3129 ) | ( ~n3127 & n3129 ) ;
  assign n3131 = ( x56 & n3127 ) | ( x56 & n3130 ) | ( n3127 & n3130 ) ;
  assign n3132 = n2067 & ~n3044 ;
  assign n3133 = x55 | n3132 ;
  assign n3134 = ~n3131 & n3133 ;
  assign n3135 = ( n3125 & n3131 ) | ( n3125 & ~n3134 ) | ( n3131 & ~n3134 ) ;
  assign n3136 = n2151 & n3028 ;
  assign n3137 = x62 & ~n3136 ;
  assign n3138 = n2151 | n3101 ;
  assign n3139 = n3137 & n3138 ;
  assign n3140 = ( x241 & n2120 ) | ( x241 & ~n3139 ) | ( n2120 & ~n3139 ) ;
  assign n3141 = n3139 | n3140 ;
  assign n3142 = n2099 & ~n3028 ;
  assign n3143 = x56 & ~n3142 ;
  assign n3144 = ~n2099 & n3101 ;
  assign n3145 = ( x62 & n3143 ) | ( x62 & ~n3144 ) | ( n3143 & ~n3144 ) ;
  assign n3146 = n3145 ^ n3143 ^ 1'b0 ;
  assign n3147 = ( x62 & n3145 ) | ( x62 & ~n3146 ) | ( n3145 & ~n3146 ) ;
  assign n3148 = ~n3141 & n3147 ;
  assign n3149 = ( n3135 & n3141 ) | ( n3135 & ~n3148 ) | ( n3141 & ~n3148 ) ;
  assign n3150 = ~n3009 & n3028 ;
  assign n3151 = n2099 & ~n3150 ;
  assign n3152 = x56 & ~n3151 ;
  assign n3153 = n2265 | n3022 ;
  assign n3154 = n3096 | n3153 ;
  assign n3155 = ~n3016 & n3154 ;
  assign n3156 = n3015 | n3155 ;
  assign n3157 = x215 | n3156 ;
  assign n3158 = ( ~x215 & n3011 ) | ( ~x215 & n3157 ) | ( n3011 & n3157 ) ;
  assign n3159 = ~n2099 & n3158 ;
  assign n3160 = ( x62 & n3152 ) | ( x62 & ~n3159 ) | ( n3152 & ~n3159 ) ;
  assign n3161 = n3160 ^ n3152 ^ 1'b0 ;
  assign n3162 = ( x62 & n3160 ) | ( x62 & ~n3161 ) | ( n3160 & ~n3161 ) ;
  assign n3163 = n2292 | n3042 ;
  assign n3164 = x299 & ~n3150 ;
  assign n3165 = n3163 | n3164 ;
  assign n3166 = n2067 & ~n3165 ;
  assign n3167 = n2044 & ~n3165 ;
  assign n3168 = x299 & n3158 ;
  assign n3169 = n3163 | n3168 ;
  assign n3170 = n3169 ^ n2036 ^ 1'b0 ;
  assign n3171 = ( n3165 & n3169 ) | ( n3165 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3172 = n2044 | n3171 ;
  assign n3173 = ( x92 & n3167 ) | ( x92 & n3172 ) | ( n3167 & n3172 ) ;
  assign n3174 = ~n3167 & n3173 ;
  assign n3175 = x75 & ~n3165 ;
  assign n3176 = x87 & n3171 ;
  assign n3177 = x38 & ~n3165 ;
  assign n3178 = x39 & n3169 ;
  assign n3179 = ~x861 & n2311 ;
  assign n3180 = x171 | n3179 ;
  assign n3181 = x861 & ~n2230 ;
  assign n3182 = x861 | n2319 ;
  assign n3183 = ( x171 & n3181 ) | ( x171 & n3182 ) | ( n3181 & n3182 ) ;
  assign n3184 = ~n3181 & n3183 ;
  assign n3185 = ( x228 & n3180 ) | ( x228 & ~n3184 ) | ( n3180 & ~n3184 ) ;
  assign n3186 = n3185 ^ n3180 ^ 1'b0 ;
  assign n3187 = ( x228 & n3185 ) | ( x228 & ~n3186 ) | ( n3185 & ~n3186 ) ;
  assign n3188 = ( n2742 & ~n3022 ) | ( n2742 & n3187 ) | ( ~n3022 & n3187 ) ;
  assign n3189 = ~n2742 & n3188 ;
  assign n3190 = ( x221 & n3008 ) | ( x221 & ~n3189 ) | ( n3008 & ~n3189 ) ;
  assign n3191 = n3189 | n3190 ;
  assign n3192 = n3191 ^ n3015 ^ 1'b0 ;
  assign n3193 = ( n3015 & n3191 ) | ( n3015 & n3192 ) | ( n3191 & n3192 ) ;
  assign n3194 = ( x215 & ~n3015 ) | ( x215 & n3193 ) | ( ~n3015 & n3193 ) ;
  assign n3195 = ( n3061 & ~n3091 ) | ( n3061 & n3194 ) | ( ~n3091 & n3194 ) ;
  assign n3196 = n3091 ^ n3061 ^ 1'b0 ;
  assign n3197 = ( n3091 & ~n3195 ) | ( n3091 & n3196 ) | ( ~n3195 & n3196 ) ;
  assign n3198 = ( x38 & ~n3178 ) | ( x38 & n3197 ) | ( ~n3178 & n3197 ) ;
  assign n3199 = n3178 | n3198 ;
  assign n3200 = ( x100 & ~n3177 ) | ( x100 & n3199 ) | ( ~n3177 & n3199 ) ;
  assign n3201 = ~x100 & n3200 ;
  assign n3202 = n1994 & ~n3165 ;
  assign n3203 = x100 & ~n3202 ;
  assign n3204 = n3050 | n3153 ;
  assign n3205 = ~n3016 & n3204 ;
  assign n3206 = ( ~x215 & n3015 ) | ( ~x215 & n3205 ) | ( n3015 & n3205 ) ;
  assign n3207 = ~x215 & n3206 ;
  assign n3208 = ( x299 & n3011 ) | ( x299 & n3207 ) | ( n3011 & n3207 ) ;
  assign n3209 = n3207 ^ n3011 ^ 1'b0 ;
  assign n3210 = ( x299 & n3208 ) | ( x299 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = ( n1994 & n3163 ) | ( n1994 & ~n3210 ) | ( n3163 & ~n3210 ) ;
  assign n3212 = n3210 | n3211 ;
  assign n3213 = n3203 & n3212 ;
  assign n3214 = ( ~x87 & n3201 ) | ( ~x87 & n3213 ) | ( n3201 & n3213 ) ;
  assign n3215 = ~x87 & n3214 ;
  assign n3216 = ( x75 & ~n3176 ) | ( x75 & n3215 ) | ( ~n3176 & n3215 ) ;
  assign n3217 = n3176 | n3216 ;
  assign n3218 = ( x92 & ~n3175 ) | ( x92 & n3217 ) | ( ~n3175 & n3217 ) ;
  assign n3219 = ~x92 & n3218 ;
  assign n3220 = ( n2067 & ~n3174 ) | ( n2067 & n3219 ) | ( ~n3174 & n3219 ) ;
  assign n3221 = n3174 | n3220 ;
  assign n3222 = ( x55 & ~n3166 ) | ( x55 & n3221 ) | ( ~n3166 & n3221 ) ;
  assign n3223 = ~x55 & n3222 ;
  assign n3224 = n2070 | n3158 ;
  assign n3225 = n3224 ^ x56 ^ 1'b0 ;
  assign n3226 = ( x55 & n3009 ) | ( x55 & n3129 ) | ( n3009 & n3129 ) ;
  assign n3227 = ( n3224 & ~n3225 ) | ( n3224 & n3226 ) | ( ~n3225 & n3226 ) ;
  assign n3228 = ( x56 & n3225 ) | ( x56 & n3227 ) | ( n3225 & n3227 ) ;
  assign n3229 = ( ~n3162 & n3223 ) | ( ~n3162 & n3228 ) | ( n3223 & n3228 ) ;
  assign n3230 = ~n3162 & n3229 ;
  assign n3231 = x241 & ~n2120 ;
  assign n3232 = n2151 & n3150 ;
  assign n3233 = n2151 | n3158 ;
  assign n3234 = ( x62 & n3232 ) | ( x62 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3235 = ~n3232 & n3234 ;
  assign n3236 = ( n3230 & n3231 ) | ( n3230 & ~n3235 ) | ( n3231 & ~n3235 ) ;
  assign n3237 = ~n3230 & n3236 ;
  assign n3238 = ( n3030 & n3149 ) | ( n3030 & ~n3237 ) | ( n3149 & ~n3237 ) ;
  assign n3239 = ~n3030 & n3238 ;
  assign n3240 = x216 & x282 ;
  assign n3241 = n2372 & ~n3240 ;
  assign n3242 = x248 & n3241 ;
  assign n3243 = x215 & x1140 ;
  assign n3244 = ~x921 & n1315 ;
  assign n3245 = x1140 | n1315 ;
  assign n3246 = ( x221 & n3244 ) | ( x221 & n3245 ) | ( n3244 & n3245 ) ;
  assign n3247 = ~n3244 & n3246 ;
  assign n3248 = x221 | n3240 ;
  assign n3249 = ~x105 & x170 ;
  assign n3250 = x869 & ~n1224 ;
  assign n3251 = x105 & ~n3250 ;
  assign n3252 = ( x228 & n3249 ) | ( x228 & ~n3251 ) | ( n3249 & ~n3251 ) ;
  assign n3253 = ~n3249 & n3252 ;
  assign n3254 = x216 | n3253 ;
  assign n3255 = x170 | x228 ;
  assign n3256 = ~n3254 & n3255 ;
  assign n3257 = ( ~n3247 & n3248 ) | ( ~n3247 & n3256 ) | ( n3248 & n3256 ) ;
  assign n3258 = ~n3247 & n3257 ;
  assign n3259 = x215 | n3258 ;
  assign n3260 = ~n3243 & n3259 ;
  assign n3261 = ( n2120 & n3242 ) | ( n2120 & n3260 ) | ( n3242 & n3260 ) ;
  assign n3262 = ~n3242 & n3261 ;
  assign n3263 = x223 & ~x1140 ;
  assign n3264 = x224 | n3250 ;
  assign n3265 = ( x222 & x282 ) | ( x222 & n1359 ) | ( x282 & n1359 ) ;
  assign n3266 = n3264 & ~n3265 ;
  assign n3267 = ~x921 & n1208 ;
  assign n3268 = x1140 | n1208 ;
  assign n3269 = ( x222 & n3267 ) | ( x222 & n3268 ) | ( n3267 & n3268 ) ;
  assign n3270 = ~n3267 & n3269 ;
  assign n3271 = ( x223 & ~n3266 ) | ( x223 & n3270 ) | ( ~n3266 & n3270 ) ;
  assign n3272 = n3266 | n3271 ;
  assign n3273 = ( x299 & ~n3263 ) | ( x299 & n3272 ) | ( ~n3263 & n3272 ) ;
  assign n3274 = ~x299 & n3273 ;
  assign n3275 = x299 & ~n3260 ;
  assign n3276 = n3274 | n3275 ;
  assign n3277 = n1994 & ~n3276 ;
  assign n3278 = x100 & ~n3277 ;
  assign n3279 = x869 | n2404 ;
  assign n3280 = x170 & n2404 ;
  assign n3281 = ( x228 & n3279 ) | ( x228 & ~n3280 ) | ( n3279 & ~n3280 ) ;
  assign n3282 = ~x228 & n3281 ;
  assign n3283 = n3254 | n3282 ;
  assign n3284 = ~n3248 & n3283 ;
  assign n3285 = ( ~x215 & n3247 ) | ( ~x215 & n3284 ) | ( n3247 & n3284 ) ;
  assign n3286 = ~x215 & n3285 ;
  assign n3287 = ( x299 & n3243 ) | ( x299 & n3286 ) | ( n3243 & n3286 ) ;
  assign n3288 = n3286 ^ n3243 ^ 1'b0 ;
  assign n3289 = ( x299 & n3287 ) | ( x299 & n3288 ) | ( n3287 & n3288 ) ;
  assign n3290 = ( n1994 & n3274 ) | ( n1994 & ~n3289 ) | ( n3274 & ~n3289 ) ;
  assign n3291 = n3289 | n3290 ;
  assign n3292 = n3278 & n3291 ;
  assign n3293 = x299 & ~n3243 ;
  assign n3294 = ~n2318 & n3253 ;
  assign n3295 = x170 & n2311 ;
  assign n3296 = x869 & n2319 ;
  assign n3297 = x170 | n3296 ;
  assign n3298 = x869 & ~n3297 ;
  assign n3299 = ( x869 & n3295 ) | ( x869 & n3298 ) | ( n3295 & n3298 ) ;
  assign n3300 = n2230 | n3297 ;
  assign n3301 = n3300 ^ n3299 ^ 1'b0 ;
  assign n3302 = ( n3299 & n3300 ) | ( n3299 & n3301 ) | ( n3300 & n3301 ) ;
  assign n3303 = ( x228 & ~n3299 ) | ( x228 & n3302 ) | ( ~n3299 & n3302 ) ;
  assign n3304 = ( x216 & ~n3294 ) | ( x216 & n3303 ) | ( ~n3294 & n3303 ) ;
  assign n3305 = ~x216 & n3304 ;
  assign n3306 = ( x221 & n3240 ) | ( x221 & ~n3305 ) | ( n3240 & ~n3305 ) ;
  assign n3307 = n3305 | n3306 ;
  assign n3308 = n3307 ^ n3247 ^ 1'b0 ;
  assign n3309 = ( n3247 & n3307 ) | ( n3247 & n3308 ) | ( n3307 & n3308 ) ;
  assign n3310 = ( x215 & ~n3247 ) | ( x215 & n3309 ) | ( ~n3247 & n3309 ) ;
  assign n3311 = n3293 & n3310 ;
  assign n3312 = x223 & x1140 ;
  assign n3313 = x299 | n3312 ;
  assign n3314 = x869 & ~n2314 ;
  assign n3315 = x224 | n3314 ;
  assign n3316 = ~n3265 & n3315 ;
  assign n3317 = n3270 | n3316 ;
  assign n3318 = n3313 | n3317 ;
  assign n3319 = n2314 & ~n3265 ;
  assign n3320 = ( ~x223 & n3317 ) | ( ~x223 & n3319 ) | ( n3317 & n3319 ) ;
  assign n3321 = ~x223 & n3320 ;
  assign n3322 = ( ~x39 & n3313 ) | ( ~x39 & n3321 ) | ( n3313 & n3321 ) ;
  assign n3323 = ~x39 & n3322 ;
  assign n3324 = ( n3311 & n3318 ) | ( n3311 & n3323 ) | ( n3318 & n3323 ) ;
  assign n3325 = ~n3311 & n3324 ;
  assign n3326 = x170 & n1292 ;
  assign n3327 = ( ~x228 & x869 ) | ( ~x228 & n2613 ) | ( x869 & n2613 ) ;
  assign n3328 = ~n3326 & n3327 ;
  assign n3329 = n3254 | n3328 ;
  assign n3330 = ~n3248 & n3329 ;
  assign n3331 = n3247 | n3330 ;
  assign n3332 = x215 | n3331 ;
  assign n3333 = ( ~x215 & n3243 ) | ( ~x215 & n3332 ) | ( n3243 & n3332 ) ;
  assign n3334 = x299 & n3333 ;
  assign n3335 = n3274 | n3334 ;
  assign n3336 = x39 & n3335 ;
  assign n3337 = ( x38 & ~n3325 ) | ( x38 & n3336 ) | ( ~n3325 & n3336 ) ;
  assign n3338 = n3325 | n3337 ;
  assign n3339 = x38 & ~n3276 ;
  assign n3340 = ( x100 & n3338 ) | ( x100 & ~n3339 ) | ( n3338 & ~n3339 ) ;
  assign n3341 = ~x100 & n3340 ;
  assign n3342 = ( ~x87 & n3292 ) | ( ~x87 & n3341 ) | ( n3292 & n3341 ) ;
  assign n3343 = ~x87 & n3342 ;
  assign n3344 = n3335 ^ n2036 ^ 1'b0 ;
  assign n3345 = ( n3276 & n3335 ) | ( n3276 & n3344 ) | ( n3335 & n3344 ) ;
  assign n3346 = x87 & n3345 ;
  assign n3347 = ( x75 & ~n3343 ) | ( x75 & n3346 ) | ( ~n3343 & n3346 ) ;
  assign n3348 = n3343 | n3347 ;
  assign n3349 = ( x92 & n2046 ) | ( x92 & n3276 ) | ( n2046 & n3276 ) ;
  assign n3350 = n3349 ^ n2067 ^ 1'b0 ;
  assign n3351 = n2044 | n3345 ;
  assign n3352 = ( n3349 & ~n3350 ) | ( n3349 & n3351 ) | ( ~n3350 & n3351 ) ;
  assign n3353 = ( n2067 & n3350 ) | ( n2067 & n3352 ) | ( n3350 & n3352 ) ;
  assign n3354 = x75 & ~n3276 ;
  assign n3355 = x92 | n3354 ;
  assign n3356 = ~n3353 & n3355 ;
  assign n3357 = ( n3348 & n3353 ) | ( n3348 & ~n3356 ) | ( n3353 & ~n3356 ) ;
  assign n3358 = n2070 | n3333 ;
  assign n3359 = n3358 ^ x56 ^ 1'b0 ;
  assign n3360 = n2070 & n3260 ;
  assign n3361 = x55 & ~n3360 ;
  assign n3362 = ( n3358 & ~n3359 ) | ( n3358 & n3361 ) | ( ~n3359 & n3361 ) ;
  assign n3363 = ( x56 & n3359 ) | ( x56 & n3362 ) | ( n3359 & n3362 ) ;
  assign n3364 = n2067 & ~n3276 ;
  assign n3365 = x55 | n3364 ;
  assign n3366 = ~n3363 & n3365 ;
  assign n3367 = ( n3357 & n3363 ) | ( n3357 & ~n3366 ) | ( n3363 & ~n3366 ) ;
  assign n3368 = n2151 & n3260 ;
  assign n3369 = x62 & ~n3368 ;
  assign n3370 = n2151 | n3333 ;
  assign n3371 = n3369 & n3370 ;
  assign n3372 = ( x248 & n2120 ) | ( x248 & ~n3371 ) | ( n2120 & ~n3371 ) ;
  assign n3373 = n3371 | n3372 ;
  assign n3374 = n2099 & ~n3260 ;
  assign n3375 = x56 & ~n3374 ;
  assign n3376 = ~n2099 & n3333 ;
  assign n3377 = ( x62 & n3375 ) | ( x62 & ~n3376 ) | ( n3375 & ~n3376 ) ;
  assign n3378 = n3377 ^ n3375 ^ 1'b0 ;
  assign n3379 = ( x62 & n3377 ) | ( x62 & ~n3378 ) | ( n3377 & ~n3378 ) ;
  assign n3380 = ~n3373 & n3379 ;
  assign n3381 = ( n3367 & n3373 ) | ( n3367 & ~n3380 ) | ( n3373 & ~n3380 ) ;
  assign n3382 = ~n3241 & n3260 ;
  assign n3383 = n2099 & ~n3382 ;
  assign n3384 = x56 & ~n3383 ;
  assign n3385 = n2265 | n3254 ;
  assign n3386 = n3328 | n3385 ;
  assign n3387 = ~n3248 & n3386 ;
  assign n3388 = n3247 | n3387 ;
  assign n3389 = x215 | n3388 ;
  assign n3390 = ( ~x215 & n3243 ) | ( ~x215 & n3389 ) | ( n3243 & n3389 ) ;
  assign n3391 = ~n2099 & n3390 ;
  assign n3392 = ( x62 & n3384 ) | ( x62 & ~n3391 ) | ( n3384 & ~n3391 ) ;
  assign n3393 = n3392 ^ n3384 ^ 1'b0 ;
  assign n3394 = ( x62 & n3392 ) | ( x62 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = n2292 | n3274 ;
  assign n3396 = x299 & ~n3382 ;
  assign n3397 = n3395 | n3396 ;
  assign n3398 = n2067 & ~n3397 ;
  assign n3399 = n2044 & ~n3397 ;
  assign n3400 = x299 & n3390 ;
  assign n3401 = n3395 | n3400 ;
  assign n3402 = n3401 ^ n2036 ^ 1'b0 ;
  assign n3403 = ( n3397 & n3401 ) | ( n3397 & n3402 ) | ( n3401 & n3402 ) ;
  assign n3404 = n2044 | n3403 ;
  assign n3405 = ( x92 & n3399 ) | ( x92 & n3404 ) | ( n3399 & n3404 ) ;
  assign n3406 = ~n3399 & n3405 ;
  assign n3407 = x75 & ~n3397 ;
  assign n3408 = x87 & n3403 ;
  assign n3409 = x38 & ~n3397 ;
  assign n3410 = x39 & n3401 ;
  assign n3411 = ~x869 & n2311 ;
  assign n3412 = x170 | n3411 ;
  assign n3413 = x869 & ~n2230 ;
  assign n3414 = x869 | n2319 ;
  assign n3415 = ( x170 & n3413 ) | ( x170 & n3414 ) | ( n3413 & n3414 ) ;
  assign n3416 = ~n3413 & n3415 ;
  assign n3417 = ( x228 & n3412 ) | ( x228 & ~n3416 ) | ( n3412 & ~n3416 ) ;
  assign n3418 = n3417 ^ n3412 ^ 1'b0 ;
  assign n3419 = ( x228 & n3417 ) | ( x228 & ~n3418 ) | ( n3417 & ~n3418 ) ;
  assign n3420 = ( n2742 & ~n3254 ) | ( n2742 & n3419 ) | ( ~n3254 & n3419 ) ;
  assign n3421 = ~n2742 & n3420 ;
  assign n3422 = ( x221 & n3240 ) | ( x221 & ~n3421 ) | ( n3240 & ~n3421 ) ;
  assign n3423 = n3421 | n3422 ;
  assign n3424 = n3423 ^ n3247 ^ 1'b0 ;
  assign n3425 = ( n3247 & n3423 ) | ( n3247 & n3424 ) | ( n3423 & n3424 ) ;
  assign n3426 = ( x215 & ~n3247 ) | ( x215 & n3425 ) | ( ~n3247 & n3425 ) ;
  assign n3427 = ( n3293 & ~n3323 ) | ( n3293 & n3426 ) | ( ~n3323 & n3426 ) ;
  assign n3428 = n3323 ^ n3293 ^ 1'b0 ;
  assign n3429 = ( n3323 & ~n3427 ) | ( n3323 & n3428 ) | ( ~n3427 & n3428 ) ;
  assign n3430 = ( x38 & ~n3410 ) | ( x38 & n3429 ) | ( ~n3410 & n3429 ) ;
  assign n3431 = n3410 | n3430 ;
  assign n3432 = ( x100 & ~n3409 ) | ( x100 & n3431 ) | ( ~n3409 & n3431 ) ;
  assign n3433 = ~x100 & n3432 ;
  assign n3434 = n1994 & ~n3397 ;
  assign n3435 = x100 & ~n3434 ;
  assign n3436 = n3282 | n3385 ;
  assign n3437 = ~n3248 & n3436 ;
  assign n3438 = ( ~x215 & n3247 ) | ( ~x215 & n3437 ) | ( n3247 & n3437 ) ;
  assign n3439 = ~x215 & n3438 ;
  assign n3440 = ( x299 & n3243 ) | ( x299 & n3439 ) | ( n3243 & n3439 ) ;
  assign n3441 = n3439 ^ n3243 ^ 1'b0 ;
  assign n3442 = ( x299 & n3440 ) | ( x299 & n3441 ) | ( n3440 & n3441 ) ;
  assign n3443 = ( n1994 & n3395 ) | ( n1994 & ~n3442 ) | ( n3395 & ~n3442 ) ;
  assign n3444 = n3442 | n3443 ;
  assign n3445 = n3435 & n3444 ;
  assign n3446 = ( ~x87 & n3433 ) | ( ~x87 & n3445 ) | ( n3433 & n3445 ) ;
  assign n3447 = ~x87 & n3446 ;
  assign n3448 = ( x75 & ~n3408 ) | ( x75 & n3447 ) | ( ~n3408 & n3447 ) ;
  assign n3449 = n3408 | n3448 ;
  assign n3450 = ( x92 & ~n3407 ) | ( x92 & n3449 ) | ( ~n3407 & n3449 ) ;
  assign n3451 = ~x92 & n3450 ;
  assign n3452 = ( n2067 & ~n3406 ) | ( n2067 & n3451 ) | ( ~n3406 & n3451 ) ;
  assign n3453 = n3406 | n3452 ;
  assign n3454 = ( x55 & ~n3398 ) | ( x55 & n3453 ) | ( ~n3398 & n3453 ) ;
  assign n3455 = ~x55 & n3454 ;
  assign n3456 = n2070 | n3390 ;
  assign n3457 = n3456 ^ x56 ^ 1'b0 ;
  assign n3458 = ( x55 & n3241 ) | ( x55 & n3361 ) | ( n3241 & n3361 ) ;
  assign n3459 = ( n3456 & ~n3457 ) | ( n3456 & n3458 ) | ( ~n3457 & n3458 ) ;
  assign n3460 = ( x56 & n3457 ) | ( x56 & n3459 ) | ( n3457 & n3459 ) ;
  assign n3461 = ( ~n3394 & n3455 ) | ( ~n3394 & n3460 ) | ( n3455 & n3460 ) ;
  assign n3462 = ~n3394 & n3461 ;
  assign n3463 = x248 & ~n2120 ;
  assign n3464 = n2151 & n3382 ;
  assign n3465 = n2151 | n3390 ;
  assign n3466 = ( x62 & n3464 ) | ( x62 & n3465 ) | ( n3464 & n3465 ) ;
  assign n3467 = ~n3464 & n3466 ;
  assign n3468 = ( n3462 & n3463 ) | ( n3462 & ~n3467 ) | ( n3463 & ~n3467 ) ;
  assign n3469 = ~n3462 & n3468 ;
  assign n3470 = ( n3262 & n3381 ) | ( n3262 & ~n3469 ) | ( n3381 & ~n3469 ) ;
  assign n3471 = ~n3262 & n3470 ;
  assign n3472 = x216 & ~x1139 ;
  assign n3473 = ~x833 & x1139 ;
  assign n3474 = x833 & x920 ;
  assign n3475 = x216 | n3474 ;
  assign n3476 = ( x221 & n3473 ) | ( x221 & n3475 ) | ( n3473 & n3475 ) ;
  assign n3477 = n3475 ^ n3473 ^ 1'b0 ;
  assign n3478 = ( x221 & n3476 ) | ( x221 & n3477 ) | ( n3476 & n3477 ) ;
  assign n3479 = ~n3472 & n3478 ;
  assign n3480 = x148 | x215 ;
  assign n3481 = x862 & ~n2321 ;
  assign n3482 = x216 | n3481 ;
  assign n3483 = n2230 ^ x228 ^ 1'b0 ;
  assign n3484 = ( x105 & n2230 ) | ( x105 & n3483 ) | ( n2230 & n3483 ) ;
  assign n3485 = ( x862 & ~n3482 ) | ( x862 & n3484 ) | ( ~n3482 & n3484 ) ;
  assign n3486 = ~n3482 & n3485 ;
  assign n3487 = x216 & x281 ;
  assign n3488 = ( x221 & ~n3486 ) | ( x221 & n3487 ) | ( ~n3486 & n3487 ) ;
  assign n3489 = n3486 | n3488 ;
  assign n3490 = n3479 | n3489 ;
  assign n3491 = ( ~n3479 & n3480 ) | ( ~n3479 & n3490 ) | ( n3480 & n3490 ) ;
  assign n3492 = x215 & x1139 ;
  assign n3493 = x299 & ~n3492 ;
  assign n3494 = x221 | n3487 ;
  assign n3495 = x216 | x862 ;
  assign n3496 = n2316 & ~n3495 ;
  assign n3497 = ( ~n3479 & n3494 ) | ( ~n3479 & n3496 ) | ( n3494 & n3496 ) ;
  assign n3498 = ~n3479 & n3497 ;
  assign n3499 = x148 & ~x215 ;
  assign n3500 = x216 | n3479 ;
  assign n3501 = n2316 | n3500 ;
  assign n3502 = n3499 & n3501 ;
  assign n3503 = ~n3498 & n3502 ;
  assign n3504 = n3493 & ~n3503 ;
  assign n3505 = n3491 & n3504 ;
  assign n3506 = x1139 | n1208 ;
  assign n3507 = ( x222 & x920 ) | ( x222 & n1219 ) | ( x920 & n1219 ) ;
  assign n3508 = n3506 & n3507 ;
  assign n3509 = x223 & x1139 ;
  assign n3510 = x224 | n3509 ;
  assign n3511 = n3508 | n3510 ;
  assign n3512 = x862 | n3511 ;
  assign n3513 = ( x222 & x281 ) | ( x222 & n1359 ) | ( x281 & n1359 ) ;
  assign n3514 = ( x223 & ~n3508 ) | ( x223 & n3513 ) | ( ~n3508 & n3513 ) ;
  assign n3515 = ~x223 & n3514 ;
  assign n3516 = x1139 & ~n3515 ;
  assign n3517 = ( x223 & n3515 ) | ( x223 & ~n3516 ) | ( n3515 & ~n3516 ) ;
  assign n3518 = n3512 & ~n3517 ;
  assign n3519 = n2314 & ~n3511 ;
  assign n3520 = ( x299 & n3518 ) | ( x299 & ~n3519 ) | ( n3518 & ~n3519 ) ;
  assign n3521 = n3520 ^ n3518 ^ 1'b0 ;
  assign n3522 = ( x299 & n3520 ) | ( x299 & ~n3521 ) | ( n3520 & ~n3521 ) ;
  assign n3523 = ( x39 & ~n3505 ) | ( x39 & n3522 ) | ( ~n3505 & n3522 ) ;
  assign n3524 = ~x39 & n3523 ;
  assign n3525 = n1224 & ~n3511 ;
  assign n3526 = x299 | n3517 ;
  assign n3527 = n3512 & ~n3526 ;
  assign n3528 = ~n3525 & n3527 ;
  assign n3529 = n2142 & ~n2376 ;
  assign n3530 = ~n3500 & n3529 ;
  assign n3531 = n3495 | n3529 ;
  assign n3532 = ~n3494 & n3531 ;
  assign n3533 = n3479 | n3532 ;
  assign n3534 = ( n3499 & n3530 ) | ( n3499 & n3533 ) | ( n3530 & n3533 ) ;
  assign n3535 = ~n3530 & n3534 ;
  assign n3536 = n3492 | n3535 ;
  assign n3537 = ~n1323 & n2142 ;
  assign n3538 = x862 & ~n2265 ;
  assign n3539 = ( x216 & ~n3537 ) | ( x216 & n3538 ) | ( ~n3537 & n3538 ) ;
  assign n3540 = n3537 | n3539 ;
  assign n3541 = n3540 ^ n3494 ^ 1'b0 ;
  assign n3542 = ( n3494 & n3540 ) | ( n3494 & n3541 ) | ( n3540 & n3541 ) ;
  assign n3543 = ( n3479 & ~n3494 ) | ( n3479 & n3542 ) | ( ~n3494 & n3542 ) ;
  assign n3544 = ~n3480 & n3543 ;
  assign n3545 = n3536 | n3544 ;
  assign n3546 = x299 & n3545 ;
  assign n3547 = n3528 | n3546 ;
  assign n3548 = x39 & n3547 ;
  assign n3549 = ( x38 & ~n3524 ) | ( x38 & n3548 ) | ( ~n3524 & n3548 ) ;
  assign n3550 = n3524 | n3549 ;
  assign n3551 = n2376 & ~n3495 ;
  assign n3552 = ( ~n3479 & n3494 ) | ( ~n3479 & n3551 ) | ( n3494 & n3551 ) ;
  assign n3553 = ~n3479 & n3552 ;
  assign n3554 = x148 & ~n1323 ;
  assign n3555 = ~n3500 & n3554 ;
  assign n3556 = x215 | n3555 ;
  assign n3557 = ( ~n3492 & n3553 ) | ( ~n3492 & n3556 ) | ( n3553 & n3556 ) ;
  assign n3558 = ~n3492 & n3557 ;
  assign n3559 = n2266 | n3558 ;
  assign n3560 = x299 & ~n3559 ;
  assign n3561 = n3528 | n3560 ;
  assign n3562 = x38 & ~n3561 ;
  assign n3563 = ( x100 & n3550 ) | ( x100 & ~n3562 ) | ( n3550 & ~n3562 ) ;
  assign n3564 = ~x100 & n3563 ;
  assign n3565 = n1994 & ~n3561 ;
  assign n3566 = ~n1323 & n2405 ;
  assign n3567 = ~n3494 & n3566 ;
  assign n3568 = n3543 | n3567 ;
  assign n3569 = ~n3480 & n3568 ;
  assign n3570 = n3492 | n3569 ;
  assign n3571 = n2406 & ~n3494 ;
  assign n3572 = n3533 | n3571 ;
  assign n3573 = n2406 & ~n3500 ;
  assign n3574 = n3499 & ~n3573 ;
  assign n3575 = n3572 & n3574 ;
  assign n3576 = ( x299 & n3570 ) | ( x299 & n3575 ) | ( n3570 & n3575 ) ;
  assign n3577 = n3575 ^ n3570 ^ 1'b0 ;
  assign n3578 = ( x299 & n3576 ) | ( x299 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3579 = ( n1994 & n3528 ) | ( n1994 & ~n3578 ) | ( n3528 & ~n3578 ) ;
  assign n3580 = n3578 | n3579 ;
  assign n3581 = ( x100 & n3565 ) | ( x100 & n3580 ) | ( n3565 & n3580 ) ;
  assign n3582 = ~n3565 & n3581 ;
  assign n3583 = ( ~x87 & n3564 ) | ( ~x87 & n3582 ) | ( n3564 & n3582 ) ;
  assign n3584 = ~x87 & n3583 ;
  assign n3585 = n3561 ^ n2036 ^ 1'b0 ;
  assign n3586 = ( n3547 & n3561 ) | ( n3547 & ~n3585 ) | ( n3561 & ~n3585 ) ;
  assign n3587 = x87 & n3586 ;
  assign n3588 = ( x75 & ~n3584 ) | ( x75 & n3587 ) | ( ~n3584 & n3587 ) ;
  assign n3589 = n3584 | n3588 ;
  assign n3590 = ( x92 & n2046 ) | ( x92 & n3561 ) | ( n2046 & n3561 ) ;
  assign n3591 = n3590 ^ n2067 ^ 1'b0 ;
  assign n3592 = n2044 | n3586 ;
  assign n3593 = ( n3590 & ~n3591 ) | ( n3590 & n3592 ) | ( ~n3591 & n3592 ) ;
  assign n3594 = ( n2067 & n3591 ) | ( n2067 & n3593 ) | ( n3591 & n3593 ) ;
  assign n3595 = x75 & ~n3561 ;
  assign n3596 = x92 | n3595 ;
  assign n3597 = ~n3594 & n3596 ;
  assign n3598 = ( n3589 & n3594 ) | ( n3589 & ~n3597 ) | ( n3594 & ~n3597 ) ;
  assign n3599 = n2070 & n3559 ;
  assign n3600 = x55 & ~n3599 ;
  assign n3601 = n3600 ^ x56 ^ 1'b0 ;
  assign n3602 = n2070 | n3545 ;
  assign n3603 = ( n3600 & ~n3601 ) | ( n3600 & n3602 ) | ( ~n3601 & n3602 ) ;
  assign n3604 = ( x56 & n3601 ) | ( x56 & n3603 ) | ( n3601 & n3603 ) ;
  assign n3605 = n2067 & ~n3561 ;
  assign n3606 = x55 | n3605 ;
  assign n3607 = ~n3604 & n3606 ;
  assign n3608 = ( n3598 & n3604 ) | ( n3598 & ~n3607 ) | ( n3604 & ~n3607 ) ;
  assign n3609 = n2151 & n3559 ;
  assign n3610 = x62 & ~n3609 ;
  assign n3611 = n3610 ^ n2120 ^ 1'b0 ;
  assign n3612 = n2151 | n3545 ;
  assign n3613 = ( n3610 & ~n3611 ) | ( n3610 & n3612 ) | ( ~n3611 & n3612 ) ;
  assign n3614 = ( n2120 & n3611 ) | ( n2120 & n3613 ) | ( n3611 & n3613 ) ;
  assign n3615 = ~n2099 & n3545 ;
  assign n3616 = n2099 & ~n3558 ;
  assign n3617 = x56 & ~n3616 ;
  assign n3618 = ( x56 & n2266 ) | ( x56 & n3617 ) | ( n2266 & n3617 ) ;
  assign n3619 = n3618 ^ n3615 ^ 1'b0 ;
  assign n3620 = ( n3615 & n3618 ) | ( n3615 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3621 = ( x62 & ~n3615 ) | ( x62 & n3620 ) | ( ~n3615 & n3620 ) ;
  assign n3622 = ~n3614 & n3621 ;
  assign n3623 = ( n3608 & n3614 ) | ( n3608 & ~n3622 ) | ( n3614 & ~n3622 ) ;
  assign n3624 = n2120 & n3558 ;
  assign n3627 = x862 & n3484 ;
  assign n3628 = ~x862 & n2321 ;
  assign n3629 = ( x216 & ~n3627 ) | ( x216 & n3628 ) | ( ~n3627 & n3628 ) ;
  assign n3630 = n3627 | n3629 ;
  assign n3631 = n3630 ^ n3494 ^ 1'b0 ;
  assign n3632 = ( n3494 & n3630 ) | ( n3494 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = ( n3479 & ~n3494 ) | ( n3479 & n3632 ) | ( ~n3494 & n3632 ) ;
  assign n3634 = n3499 & n3633 ;
  assign n3625 = n3480 | n3498 ;
  assign n3626 = ~n3492 & n3625 ;
  assign n3635 = n3634 ^ n3626 ^ 1'b0 ;
  assign n3636 = ( x299 & ~n3626 ) | ( x299 & n3634 ) | ( ~n3626 & n3634 ) ;
  assign n3637 = ( x299 & ~n3635 ) | ( x299 & n3636 ) | ( ~n3635 & n3636 ) ;
  assign n3638 = ( n2314 & ~n3526 ) | ( n2314 & n3527 ) | ( ~n3526 & n3527 ) ;
  assign n3639 = ( ~x39 & n3637 ) | ( ~x39 & n3638 ) | ( n3637 & n3638 ) ;
  assign n3640 = ~x39 & n3639 ;
  assign n3641 = n2292 | n3527 ;
  assign n3642 = n3533 & ~n3556 ;
  assign n3643 = n3536 | n3642 ;
  assign n3644 = x299 & n3643 ;
  assign n3645 = n3641 | n3644 ;
  assign n3646 = x39 & n3645 ;
  assign n3647 = ( x38 & ~n3640 ) | ( x38 & n3646 ) | ( ~n3640 & n3646 ) ;
  assign n3648 = n3640 | n3647 ;
  assign n3649 = x299 & ~n3558 ;
  assign n3650 = n3641 | n3649 ;
  assign n3651 = x38 & ~n3650 ;
  assign n3652 = ( x100 & n3648 ) | ( x100 & ~n3651 ) | ( n3648 & ~n3651 ) ;
  assign n3653 = ~x100 & n3652 ;
  assign n3654 = n1994 & ~n3650 ;
  assign n3655 = ~n3500 & n3566 ;
  assign n3656 = n3499 & n3533 ;
  assign n3657 = n3656 ^ n3655 ^ 1'b0 ;
  assign n3658 = ( n3655 & n3656 ) | ( n3655 & n3657 ) | ( n3656 & n3657 ) ;
  assign n3659 = ( n3492 & ~n3655 ) | ( n3492 & n3658 ) | ( ~n3655 & n3658 ) ;
  assign n3660 = ~n3480 & n3572 ;
  assign n3661 = ( x299 & n3659 ) | ( x299 & n3660 ) | ( n3659 & n3660 ) ;
  assign n3662 = n3660 ^ n3659 ^ 1'b0 ;
  assign n3663 = ( x299 & n3661 ) | ( x299 & n3662 ) | ( n3661 & n3662 ) ;
  assign n3664 = ( n1994 & n3641 ) | ( n1994 & ~n3663 ) | ( n3641 & ~n3663 ) ;
  assign n3665 = n3663 | n3664 ;
  assign n3666 = ( x100 & n3654 ) | ( x100 & n3665 ) | ( n3654 & n3665 ) ;
  assign n3667 = ~n3654 & n3666 ;
  assign n3668 = ( ~x87 & n3653 ) | ( ~x87 & n3667 ) | ( n3653 & n3667 ) ;
  assign n3669 = ~x87 & n3668 ;
  assign n3670 = n3650 ^ n2036 ^ 1'b0 ;
  assign n3671 = ( n3645 & n3650 ) | ( n3645 & ~n3670 ) | ( n3650 & ~n3670 ) ;
  assign n3672 = x87 & n3671 ;
  assign n3673 = ( x75 & ~n3669 ) | ( x75 & n3672 ) | ( ~n3669 & n3672 ) ;
  assign n3674 = n3669 | n3673 ;
  assign n3675 = x75 & ~n3650 ;
  assign n3676 = ( x92 & n3674 ) | ( x92 & ~n3675 ) | ( n3674 & ~n3675 ) ;
  assign n3677 = ~x92 & n3676 ;
  assign n3678 = n2044 & ~n3650 ;
  assign n3679 = n2044 | n3671 ;
  assign n3680 = ( x92 & n3678 ) | ( x92 & n3679 ) | ( n3678 & n3679 ) ;
  assign n3681 = ~n3678 & n3680 ;
  assign n3682 = ( n2067 & ~n3677 ) | ( n2067 & n3681 ) | ( ~n3677 & n3681 ) ;
  assign n3683 = n3677 | n3682 ;
  assign n3684 = n2070 & n3558 ;
  assign n3685 = x55 & ~n3684 ;
  assign n3686 = n3685 ^ x56 ^ 1'b0 ;
  assign n3687 = n2070 | n3643 ;
  assign n3688 = ( n3685 & ~n3686 ) | ( n3685 & n3687 ) | ( ~n3686 & n3687 ) ;
  assign n3689 = ( x56 & n3686 ) | ( x56 & n3688 ) | ( n3686 & n3688 ) ;
  assign n3690 = n2067 & ~n3650 ;
  assign n3691 = x55 | n3690 ;
  assign n3692 = ~n3689 & n3691 ;
  assign n3693 = ( n3683 & n3689 ) | ( n3683 & ~n3692 ) | ( n3689 & ~n3692 ) ;
  assign n3694 = n2151 & n3558 ;
  assign n3695 = x62 & ~n3694 ;
  assign n3696 = n3695 ^ n2120 ^ 1'b0 ;
  assign n3697 = n2151 | n3643 ;
  assign n3698 = ( n3695 & ~n3696 ) | ( n3695 & n3697 ) | ( ~n3696 & n3697 ) ;
  assign n3699 = ( n2120 & n3696 ) | ( n2120 & n3698 ) | ( n3696 & n3698 ) ;
  assign n3700 = ~n2099 & n3643 ;
  assign n3701 = n3700 ^ n3617 ^ 1'b0 ;
  assign n3702 = ( n3617 & n3700 ) | ( n3617 & n3701 ) | ( n3700 & n3701 ) ;
  assign n3703 = ( x62 & ~n3700 ) | ( x62 & n3702 ) | ( ~n3700 & n3702 ) ;
  assign n3704 = ~n3699 & n3703 ;
  assign n3705 = ( n3693 & n3699 ) | ( n3693 & ~n3704 ) | ( n3699 & ~n3704 ) ;
  assign n3706 = ( x247 & n3624 ) | ( x247 & n3705 ) | ( n3624 & n3705 ) ;
  assign n3707 = ~n3624 & n3706 ;
  assign n3708 = n2120 & n3559 ;
  assign n3709 = x247 | n3708 ;
  assign n3710 = ~n3707 & n3709 ;
  assign n3711 = ( n3623 & n3707 ) | ( n3623 & ~n3710 ) | ( n3707 & ~n3710 ) ;
  assign n3712 = x216 & x269 ;
  assign n3713 = n2372 & ~n3712 ;
  assign n3714 = x246 & n3713 ;
  assign n3715 = x215 & x1138 ;
  assign n3716 = ~x940 & n1315 ;
  assign n3717 = x1138 | n1315 ;
  assign n3718 = ( x221 & n3716 ) | ( x221 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3719 = ~n3716 & n3718 ;
  assign n3720 = x221 | n3712 ;
  assign n3721 = ~x105 & x169 ;
  assign n3722 = x877 & ~n1224 ;
  assign n3723 = x105 & ~n3722 ;
  assign n3724 = ( x228 & n3721 ) | ( x228 & ~n3723 ) | ( n3721 & ~n3723 ) ;
  assign n3725 = ~n3721 & n3724 ;
  assign n3726 = x216 | n3725 ;
  assign n3727 = x169 | x228 ;
  assign n3728 = ~n3726 & n3727 ;
  assign n3729 = ( ~n3719 & n3720 ) | ( ~n3719 & n3728 ) | ( n3720 & n3728 ) ;
  assign n3730 = ~n3719 & n3729 ;
  assign n3731 = x215 | n3730 ;
  assign n3732 = ~n3715 & n3731 ;
  assign n3733 = ( n2120 & n3714 ) | ( n2120 & n3732 ) | ( n3714 & n3732 ) ;
  assign n3734 = ~n3714 & n3733 ;
  assign n3735 = x223 & ~x1138 ;
  assign n3736 = x224 | n3722 ;
  assign n3737 = ( x222 & x269 ) | ( x222 & n1359 ) | ( x269 & n1359 ) ;
  assign n3738 = n3736 & ~n3737 ;
  assign n3739 = ~x940 & n1208 ;
  assign n3740 = x1138 | n1208 ;
  assign n3741 = ( x222 & n3739 ) | ( x222 & n3740 ) | ( n3739 & n3740 ) ;
  assign n3742 = ~n3739 & n3741 ;
  assign n3743 = ( x223 & ~n3738 ) | ( x223 & n3742 ) | ( ~n3738 & n3742 ) ;
  assign n3744 = n3738 | n3743 ;
  assign n3745 = ( x299 & ~n3735 ) | ( x299 & n3744 ) | ( ~n3735 & n3744 ) ;
  assign n3746 = ~x299 & n3745 ;
  assign n3747 = x299 & ~n3732 ;
  assign n3748 = n3746 | n3747 ;
  assign n3749 = n1994 & ~n3748 ;
  assign n3750 = x100 & ~n3749 ;
  assign n3751 = x877 | n2404 ;
  assign n3752 = x169 & n2404 ;
  assign n3753 = ( x228 & n3751 ) | ( x228 & ~n3752 ) | ( n3751 & ~n3752 ) ;
  assign n3754 = ~x228 & n3753 ;
  assign n3755 = n3726 | n3754 ;
  assign n3756 = ~n3720 & n3755 ;
  assign n3757 = ( ~x215 & n3719 ) | ( ~x215 & n3756 ) | ( n3719 & n3756 ) ;
  assign n3758 = ~x215 & n3757 ;
  assign n3759 = ( x299 & n3715 ) | ( x299 & n3758 ) | ( n3715 & n3758 ) ;
  assign n3760 = n3758 ^ n3715 ^ 1'b0 ;
  assign n3761 = ( x299 & n3759 ) | ( x299 & n3760 ) | ( n3759 & n3760 ) ;
  assign n3762 = ( n1994 & n3746 ) | ( n1994 & ~n3761 ) | ( n3746 & ~n3761 ) ;
  assign n3763 = n3761 | n3762 ;
  assign n3764 = n3750 & n3763 ;
  assign n3765 = x299 & ~n3715 ;
  assign n3766 = ~n2318 & n3725 ;
  assign n3767 = x169 & n2311 ;
  assign n3768 = x877 & n2319 ;
  assign n3769 = x169 | n3768 ;
  assign n3770 = x877 & ~n3769 ;
  assign n3771 = ( x877 & n3767 ) | ( x877 & n3770 ) | ( n3767 & n3770 ) ;
  assign n3772 = n2230 | n3769 ;
  assign n3773 = n3772 ^ n3771 ^ 1'b0 ;
  assign n3774 = ( n3771 & n3772 ) | ( n3771 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ( x228 & ~n3771 ) | ( x228 & n3774 ) | ( ~n3771 & n3774 ) ;
  assign n3776 = ( x216 & ~n3766 ) | ( x216 & n3775 ) | ( ~n3766 & n3775 ) ;
  assign n3777 = ~x216 & n3776 ;
  assign n3778 = ( x221 & n3712 ) | ( x221 & ~n3777 ) | ( n3712 & ~n3777 ) ;
  assign n3779 = n3777 | n3778 ;
  assign n3780 = n3779 ^ n3719 ^ 1'b0 ;
  assign n3781 = ( n3719 & n3779 ) | ( n3719 & n3780 ) | ( n3779 & n3780 ) ;
  assign n3782 = ( x215 & ~n3719 ) | ( x215 & n3781 ) | ( ~n3719 & n3781 ) ;
  assign n3783 = n3765 & n3782 ;
  assign n3784 = x223 & x1138 ;
  assign n3785 = x299 | n3784 ;
  assign n3786 = x877 & ~n2314 ;
  assign n3787 = x224 | n3786 ;
  assign n3788 = ~n3737 & n3787 ;
  assign n3789 = n3742 | n3788 ;
  assign n3790 = n3785 | n3789 ;
  assign n3791 = n2314 & ~n3737 ;
  assign n3792 = ( ~x223 & n3789 ) | ( ~x223 & n3791 ) | ( n3789 & n3791 ) ;
  assign n3793 = ~x223 & n3792 ;
  assign n3794 = ( ~x39 & n3785 ) | ( ~x39 & n3793 ) | ( n3785 & n3793 ) ;
  assign n3795 = ~x39 & n3794 ;
  assign n3796 = ( n3783 & n3790 ) | ( n3783 & n3795 ) | ( n3790 & n3795 ) ;
  assign n3797 = ~n3783 & n3796 ;
  assign n3798 = x877 | n1292 ;
  assign n3799 = x169 & n1292 ;
  assign n3800 = ( x228 & n3798 ) | ( x228 & ~n3799 ) | ( n3798 & ~n3799 ) ;
  assign n3801 = ~x228 & n3800 ;
  assign n3802 = n3726 | n3801 ;
  assign n3803 = ~n3720 & n3802 ;
  assign n3804 = n3719 | n3803 ;
  assign n3805 = x215 | n3804 ;
  assign n3806 = ( ~x215 & n3715 ) | ( ~x215 & n3805 ) | ( n3715 & n3805 ) ;
  assign n3807 = x299 & n3806 ;
  assign n3808 = n3746 | n3807 ;
  assign n3809 = x39 & n3808 ;
  assign n3810 = ( x38 & ~n3797 ) | ( x38 & n3809 ) | ( ~n3797 & n3809 ) ;
  assign n3811 = n3797 | n3810 ;
  assign n3812 = x38 & ~n3748 ;
  assign n3813 = ( x100 & n3811 ) | ( x100 & ~n3812 ) | ( n3811 & ~n3812 ) ;
  assign n3814 = ~x100 & n3813 ;
  assign n3815 = ( ~x87 & n3764 ) | ( ~x87 & n3814 ) | ( n3764 & n3814 ) ;
  assign n3816 = ~x87 & n3815 ;
  assign n3817 = n3808 ^ n2036 ^ 1'b0 ;
  assign n3818 = ( n3748 & n3808 ) | ( n3748 & n3817 ) | ( n3808 & n3817 ) ;
  assign n3819 = x87 & n3818 ;
  assign n3820 = ( x75 & ~n3816 ) | ( x75 & n3819 ) | ( ~n3816 & n3819 ) ;
  assign n3821 = n3816 | n3820 ;
  assign n3822 = ( x92 & n2046 ) | ( x92 & n3748 ) | ( n2046 & n3748 ) ;
  assign n3823 = n3822 ^ n2067 ^ 1'b0 ;
  assign n3824 = n2044 | n3818 ;
  assign n3825 = ( n3822 & ~n3823 ) | ( n3822 & n3824 ) | ( ~n3823 & n3824 ) ;
  assign n3826 = ( n2067 & n3823 ) | ( n2067 & n3825 ) | ( n3823 & n3825 ) ;
  assign n3827 = x75 & ~n3748 ;
  assign n3828 = x92 | n3827 ;
  assign n3829 = ~n3826 & n3828 ;
  assign n3830 = ( n3821 & n3826 ) | ( n3821 & ~n3829 ) | ( n3826 & ~n3829 ) ;
  assign n3831 = n2070 | n3806 ;
  assign n3832 = n3831 ^ x56 ^ 1'b0 ;
  assign n3833 = n2070 & n3732 ;
  assign n3834 = x55 & ~n3833 ;
  assign n3835 = ( n3831 & ~n3832 ) | ( n3831 & n3834 ) | ( ~n3832 & n3834 ) ;
  assign n3836 = ( x56 & n3832 ) | ( x56 & n3835 ) | ( n3832 & n3835 ) ;
  assign n3837 = n2067 & ~n3748 ;
  assign n3838 = x55 | n3837 ;
  assign n3839 = ~n3836 & n3838 ;
  assign n3840 = ( n3830 & n3836 ) | ( n3830 & ~n3839 ) | ( n3836 & ~n3839 ) ;
  assign n3841 = n2151 & n3732 ;
  assign n3842 = x62 & ~n3841 ;
  assign n3843 = n2151 | n3806 ;
  assign n3844 = n3842 & n3843 ;
  assign n3845 = ( x246 & n2120 ) | ( x246 & ~n3844 ) | ( n2120 & ~n3844 ) ;
  assign n3846 = n3844 | n3845 ;
  assign n3847 = n2099 & ~n3732 ;
  assign n3848 = x56 & ~n3847 ;
  assign n3849 = ~n2099 & n3806 ;
  assign n3850 = ( x62 & n3848 ) | ( x62 & ~n3849 ) | ( n3848 & ~n3849 ) ;
  assign n3851 = n3850 ^ n3848 ^ 1'b0 ;
  assign n3852 = ( x62 & n3850 ) | ( x62 & ~n3851 ) | ( n3850 & ~n3851 ) ;
  assign n3853 = ~n3846 & n3852 ;
  assign n3854 = ( n3840 & n3846 ) | ( n3840 & ~n3853 ) | ( n3846 & ~n3853 ) ;
  assign n3855 = ~n3713 & n3732 ;
  assign n3856 = n2099 & ~n3855 ;
  assign n3857 = x56 & ~n3856 ;
  assign n3858 = n2265 | n3726 ;
  assign n3859 = n3801 | n3858 ;
  assign n3860 = ~n3720 & n3859 ;
  assign n3861 = n3719 | n3860 ;
  assign n3862 = x215 | n3861 ;
  assign n3863 = ( ~x215 & n3715 ) | ( ~x215 & n3862 ) | ( n3715 & n3862 ) ;
  assign n3864 = ~n2099 & n3863 ;
  assign n3865 = ( x62 & n3857 ) | ( x62 & ~n3864 ) | ( n3857 & ~n3864 ) ;
  assign n3866 = n3865 ^ n3857 ^ 1'b0 ;
  assign n3867 = ( x62 & n3865 ) | ( x62 & ~n3866 ) | ( n3865 & ~n3866 ) ;
  assign n3868 = n2292 | n3746 ;
  assign n3869 = x299 & ~n3855 ;
  assign n3870 = n3868 | n3869 ;
  assign n3871 = n2067 & ~n3870 ;
  assign n3872 = n2044 & ~n3870 ;
  assign n3873 = x299 & n3863 ;
  assign n3874 = n3868 | n3873 ;
  assign n3875 = n3874 ^ n2036 ^ 1'b0 ;
  assign n3876 = ( n3870 & n3874 ) | ( n3870 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3877 = n2044 | n3876 ;
  assign n3878 = ( x92 & n3872 ) | ( x92 & n3877 ) | ( n3872 & n3877 ) ;
  assign n3879 = ~n3872 & n3878 ;
  assign n3880 = x75 & ~n3870 ;
  assign n3881 = x87 & n3876 ;
  assign n3882 = x38 & ~n3870 ;
  assign n3883 = x39 & n3874 ;
  assign n3884 = ~x877 & n2311 ;
  assign n3885 = x169 | n3884 ;
  assign n3886 = x877 & ~n2230 ;
  assign n3887 = x877 | n2319 ;
  assign n3888 = ( x169 & n3886 ) | ( x169 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ~n3886 & n3888 ;
  assign n3890 = ( x228 & n3885 ) | ( x228 & ~n3889 ) | ( n3885 & ~n3889 ) ;
  assign n3891 = n3890 ^ n3885 ^ 1'b0 ;
  assign n3892 = ( x228 & n3890 ) | ( x228 & ~n3891 ) | ( n3890 & ~n3891 ) ;
  assign n3893 = ( n2742 & ~n3726 ) | ( n2742 & n3892 ) | ( ~n3726 & n3892 ) ;
  assign n3894 = ~n2742 & n3893 ;
  assign n3895 = ( x221 & n3712 ) | ( x221 & ~n3894 ) | ( n3712 & ~n3894 ) ;
  assign n3896 = n3894 | n3895 ;
  assign n3897 = n3896 ^ n3719 ^ 1'b0 ;
  assign n3898 = ( n3719 & n3896 ) | ( n3719 & n3897 ) | ( n3896 & n3897 ) ;
  assign n3899 = ( x215 & ~n3719 ) | ( x215 & n3898 ) | ( ~n3719 & n3898 ) ;
  assign n3900 = ( n3765 & ~n3795 ) | ( n3765 & n3899 ) | ( ~n3795 & n3899 ) ;
  assign n3901 = n3795 ^ n3765 ^ 1'b0 ;
  assign n3902 = ( n3795 & ~n3900 ) | ( n3795 & n3901 ) | ( ~n3900 & n3901 ) ;
  assign n3903 = ( x38 & ~n3883 ) | ( x38 & n3902 ) | ( ~n3883 & n3902 ) ;
  assign n3904 = n3883 | n3903 ;
  assign n3905 = ( x100 & ~n3882 ) | ( x100 & n3904 ) | ( ~n3882 & n3904 ) ;
  assign n3906 = ~x100 & n3905 ;
  assign n3907 = n1994 & ~n3870 ;
  assign n3908 = x100 & ~n3907 ;
  assign n3909 = n3754 | n3858 ;
  assign n3910 = ~n3720 & n3909 ;
  assign n3911 = ( ~x215 & n3719 ) | ( ~x215 & n3910 ) | ( n3719 & n3910 ) ;
  assign n3912 = ~x215 & n3911 ;
  assign n3913 = ( x299 & n3715 ) | ( x299 & n3912 ) | ( n3715 & n3912 ) ;
  assign n3914 = n3912 ^ n3715 ^ 1'b0 ;
  assign n3915 = ( x299 & n3913 ) | ( x299 & n3914 ) | ( n3913 & n3914 ) ;
  assign n3916 = ( n1994 & n3868 ) | ( n1994 & ~n3915 ) | ( n3868 & ~n3915 ) ;
  assign n3917 = n3915 | n3916 ;
  assign n3918 = n3908 & n3917 ;
  assign n3919 = ( ~x87 & n3906 ) | ( ~x87 & n3918 ) | ( n3906 & n3918 ) ;
  assign n3920 = ~x87 & n3919 ;
  assign n3921 = ( x75 & ~n3881 ) | ( x75 & n3920 ) | ( ~n3881 & n3920 ) ;
  assign n3922 = n3881 | n3921 ;
  assign n3923 = ( x92 & ~n3880 ) | ( x92 & n3922 ) | ( ~n3880 & n3922 ) ;
  assign n3924 = ~x92 & n3923 ;
  assign n3925 = ( n2067 & ~n3879 ) | ( n2067 & n3924 ) | ( ~n3879 & n3924 ) ;
  assign n3926 = n3879 | n3925 ;
  assign n3927 = ( x55 & ~n3871 ) | ( x55 & n3926 ) | ( ~n3871 & n3926 ) ;
  assign n3928 = ~x55 & n3927 ;
  assign n3929 = n2070 | n3863 ;
  assign n3930 = n3929 ^ x56 ^ 1'b0 ;
  assign n3931 = ( x55 & n3713 ) | ( x55 & n3834 ) | ( n3713 & n3834 ) ;
  assign n3932 = ( n3929 & ~n3930 ) | ( n3929 & n3931 ) | ( ~n3930 & n3931 ) ;
  assign n3933 = ( x56 & n3930 ) | ( x56 & n3932 ) | ( n3930 & n3932 ) ;
  assign n3934 = ( ~n3867 & n3928 ) | ( ~n3867 & n3933 ) | ( n3928 & n3933 ) ;
  assign n3935 = ~n3867 & n3934 ;
  assign n3936 = x246 & ~n2120 ;
  assign n3937 = n2151 & n3855 ;
  assign n3938 = n2151 | n3863 ;
  assign n3939 = ( x62 & n3937 ) | ( x62 & n3938 ) | ( n3937 & n3938 ) ;
  assign n3940 = ~n3937 & n3939 ;
  assign n3941 = ( n3935 & n3936 ) | ( n3935 & ~n3940 ) | ( n3936 & ~n3940 ) ;
  assign n3942 = ~n3935 & n3941 ;
  assign n3943 = ( n3734 & n3854 ) | ( n3734 & ~n3942 ) | ( n3854 & ~n3942 ) ;
  assign n3944 = ~n3734 & n3943 ;
  assign n3945 = x216 & x280 ;
  assign n3946 = n2372 & ~n3945 ;
  assign n3947 = x240 & n3946 ;
  assign n3948 = x215 & x1137 ;
  assign n3949 = ~x933 & n1315 ;
  assign n3950 = x1137 | n1315 ;
  assign n3951 = ( x221 & n3949 ) | ( x221 & n3950 ) | ( n3949 & n3950 ) ;
  assign n3952 = ~n3949 & n3951 ;
  assign n3953 = x221 | n3945 ;
  assign n3954 = ~x105 & x168 ;
  assign n3955 = x878 & ~n1224 ;
  assign n3956 = x105 & ~n3955 ;
  assign n3957 = ( x228 & n3954 ) | ( x228 & ~n3956 ) | ( n3954 & ~n3956 ) ;
  assign n3958 = ~n3954 & n3957 ;
  assign n3959 = x216 | n3958 ;
  assign n3960 = x168 | x228 ;
  assign n3961 = ~n3959 & n3960 ;
  assign n3962 = ( ~n3952 & n3953 ) | ( ~n3952 & n3961 ) | ( n3953 & n3961 ) ;
  assign n3963 = ~n3952 & n3962 ;
  assign n3964 = x215 | n3963 ;
  assign n3965 = ~n3948 & n3964 ;
  assign n3966 = ( n2120 & n3947 ) | ( n2120 & n3965 ) | ( n3947 & n3965 ) ;
  assign n3967 = ~n3947 & n3966 ;
  assign n3968 = x223 & ~x1137 ;
  assign n3969 = x224 | n3955 ;
  assign n3970 = ( x222 & x280 ) | ( x222 & n1359 ) | ( x280 & n1359 ) ;
  assign n3971 = n3969 & ~n3970 ;
  assign n3972 = ~x933 & n1208 ;
  assign n3973 = x1137 | n1208 ;
  assign n3974 = ( x222 & n3972 ) | ( x222 & n3973 ) | ( n3972 & n3973 ) ;
  assign n3975 = ~n3972 & n3974 ;
  assign n3976 = ( x223 & ~n3971 ) | ( x223 & n3975 ) | ( ~n3971 & n3975 ) ;
  assign n3977 = n3971 | n3976 ;
  assign n3978 = ( x299 & ~n3968 ) | ( x299 & n3977 ) | ( ~n3968 & n3977 ) ;
  assign n3979 = ~x299 & n3978 ;
  assign n3980 = x299 & ~n3965 ;
  assign n3981 = n3979 | n3980 ;
  assign n3982 = n1994 & ~n3981 ;
  assign n3983 = x100 & ~n3982 ;
  assign n3984 = x878 | n2404 ;
  assign n3985 = x168 & n2404 ;
  assign n3986 = ( x228 & n3984 ) | ( x228 & ~n3985 ) | ( n3984 & ~n3985 ) ;
  assign n3987 = ~x228 & n3986 ;
  assign n3988 = n3959 | n3987 ;
  assign n3989 = ~n3953 & n3988 ;
  assign n3990 = ( ~x215 & n3952 ) | ( ~x215 & n3989 ) | ( n3952 & n3989 ) ;
  assign n3991 = ~x215 & n3990 ;
  assign n3992 = ( x299 & n3948 ) | ( x299 & n3991 ) | ( n3948 & n3991 ) ;
  assign n3993 = n3991 ^ n3948 ^ 1'b0 ;
  assign n3994 = ( x299 & n3992 ) | ( x299 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3995 = ( n1994 & n3979 ) | ( n1994 & ~n3994 ) | ( n3979 & ~n3994 ) ;
  assign n3996 = n3994 | n3995 ;
  assign n3997 = n3983 & n3996 ;
  assign n3998 = x299 & ~n3948 ;
  assign n3999 = ~n2318 & n3958 ;
  assign n4000 = x168 & n2311 ;
  assign n4001 = x878 & n2319 ;
  assign n4002 = x168 | n4001 ;
  assign n4003 = x878 & ~n4002 ;
  assign n4004 = ( x878 & n4000 ) | ( x878 & n4003 ) | ( n4000 & n4003 ) ;
  assign n4005 = n2230 | n4002 ;
  assign n4006 = n4005 ^ n4004 ^ 1'b0 ;
  assign n4007 = ( n4004 & n4005 ) | ( n4004 & n4006 ) | ( n4005 & n4006 ) ;
  assign n4008 = ( x228 & ~n4004 ) | ( x228 & n4007 ) | ( ~n4004 & n4007 ) ;
  assign n4009 = ( x216 & ~n3999 ) | ( x216 & n4008 ) | ( ~n3999 & n4008 ) ;
  assign n4010 = ~x216 & n4009 ;
  assign n4011 = ( x221 & n3945 ) | ( x221 & ~n4010 ) | ( n3945 & ~n4010 ) ;
  assign n4012 = n4010 | n4011 ;
  assign n4013 = n4012 ^ n3952 ^ 1'b0 ;
  assign n4014 = ( n3952 & n4012 ) | ( n3952 & n4013 ) | ( n4012 & n4013 ) ;
  assign n4015 = ( x215 & ~n3952 ) | ( x215 & n4014 ) | ( ~n3952 & n4014 ) ;
  assign n4016 = n3998 & n4015 ;
  assign n4017 = x223 & x1137 ;
  assign n4018 = x299 | n4017 ;
  assign n4019 = x878 & ~n2314 ;
  assign n4020 = x224 | n4019 ;
  assign n4021 = ~n3970 & n4020 ;
  assign n4022 = n3975 | n4021 ;
  assign n4023 = n4018 | n4022 ;
  assign n4024 = n2314 & ~n3970 ;
  assign n4025 = ( ~x223 & n4022 ) | ( ~x223 & n4024 ) | ( n4022 & n4024 ) ;
  assign n4026 = ~x223 & n4025 ;
  assign n4027 = ( ~x39 & n4018 ) | ( ~x39 & n4026 ) | ( n4018 & n4026 ) ;
  assign n4028 = ~x39 & n4027 ;
  assign n4029 = ( n4016 & n4023 ) | ( n4016 & n4028 ) | ( n4023 & n4028 ) ;
  assign n4030 = ~n4016 & n4029 ;
  assign n4031 = x878 | n1292 ;
  assign n4032 = x168 & n1292 ;
  assign n4033 = ( x228 & n4031 ) | ( x228 & ~n4032 ) | ( n4031 & ~n4032 ) ;
  assign n4034 = ~x228 & n4033 ;
  assign n4035 = n3959 | n4034 ;
  assign n4036 = ~n3953 & n4035 ;
  assign n4037 = n3952 | n4036 ;
  assign n4038 = x215 | n4037 ;
  assign n4039 = ( ~x215 & n3948 ) | ( ~x215 & n4038 ) | ( n3948 & n4038 ) ;
  assign n4040 = x299 & n4039 ;
  assign n4041 = n3979 | n4040 ;
  assign n4042 = x39 & n4041 ;
  assign n4043 = ( x38 & ~n4030 ) | ( x38 & n4042 ) | ( ~n4030 & n4042 ) ;
  assign n4044 = n4030 | n4043 ;
  assign n4045 = x38 & ~n3981 ;
  assign n4046 = ( x100 & n4044 ) | ( x100 & ~n4045 ) | ( n4044 & ~n4045 ) ;
  assign n4047 = ~x100 & n4046 ;
  assign n4048 = ( ~x87 & n3997 ) | ( ~x87 & n4047 ) | ( n3997 & n4047 ) ;
  assign n4049 = ~x87 & n4048 ;
  assign n4050 = n4041 ^ n2036 ^ 1'b0 ;
  assign n4051 = ( n3981 & n4041 ) | ( n3981 & n4050 ) | ( n4041 & n4050 ) ;
  assign n4052 = x87 & n4051 ;
  assign n4053 = ( x75 & ~n4049 ) | ( x75 & n4052 ) | ( ~n4049 & n4052 ) ;
  assign n4054 = n4049 | n4053 ;
  assign n4055 = ( x92 & n2046 ) | ( x92 & n3981 ) | ( n2046 & n3981 ) ;
  assign n4056 = n4055 ^ n2067 ^ 1'b0 ;
  assign n4057 = n2044 | n4051 ;
  assign n4058 = ( n4055 & ~n4056 ) | ( n4055 & n4057 ) | ( ~n4056 & n4057 ) ;
  assign n4059 = ( n2067 & n4056 ) | ( n2067 & n4058 ) | ( n4056 & n4058 ) ;
  assign n4060 = x75 & ~n3981 ;
  assign n4061 = x92 | n4060 ;
  assign n4062 = ~n4059 & n4061 ;
  assign n4063 = ( n4054 & n4059 ) | ( n4054 & ~n4062 ) | ( n4059 & ~n4062 ) ;
  assign n4064 = n2070 | n4039 ;
  assign n4065 = n4064 ^ x56 ^ 1'b0 ;
  assign n4066 = n2070 & n3965 ;
  assign n4067 = x55 & ~n4066 ;
  assign n4068 = ( n4064 & ~n4065 ) | ( n4064 & n4067 ) | ( ~n4065 & n4067 ) ;
  assign n4069 = ( x56 & n4065 ) | ( x56 & n4068 ) | ( n4065 & n4068 ) ;
  assign n4070 = n2067 & ~n3981 ;
  assign n4071 = x55 | n4070 ;
  assign n4072 = ~n4069 & n4071 ;
  assign n4073 = ( n4063 & n4069 ) | ( n4063 & ~n4072 ) | ( n4069 & ~n4072 ) ;
  assign n4074 = n2151 & n3965 ;
  assign n4075 = x62 & ~n4074 ;
  assign n4076 = n2151 | n4039 ;
  assign n4077 = n4075 & n4076 ;
  assign n4078 = ( x240 & n2120 ) | ( x240 & ~n4077 ) | ( n2120 & ~n4077 ) ;
  assign n4079 = n4077 | n4078 ;
  assign n4080 = n2099 & ~n3965 ;
  assign n4081 = x56 & ~n4080 ;
  assign n4082 = ~n2099 & n4039 ;
  assign n4083 = ( x62 & n4081 ) | ( x62 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  assign n4084 = n4083 ^ n4081 ^ 1'b0 ;
  assign n4085 = ( x62 & n4083 ) | ( x62 & ~n4084 ) | ( n4083 & ~n4084 ) ;
  assign n4086 = ~n4079 & n4085 ;
  assign n4087 = ( n4073 & n4079 ) | ( n4073 & ~n4086 ) | ( n4079 & ~n4086 ) ;
  assign n4088 = ~n3946 & n3965 ;
  assign n4089 = n2099 & ~n4088 ;
  assign n4090 = x56 & ~n4089 ;
  assign n4091 = n2265 | n3959 ;
  assign n4092 = n4034 | n4091 ;
  assign n4093 = ~n3953 & n4092 ;
  assign n4094 = n3952 | n4093 ;
  assign n4095 = x215 | n4094 ;
  assign n4096 = ( ~x215 & n3948 ) | ( ~x215 & n4095 ) | ( n3948 & n4095 ) ;
  assign n4097 = ~n2099 & n4096 ;
  assign n4098 = ( x62 & n4090 ) | ( x62 & ~n4097 ) | ( n4090 & ~n4097 ) ;
  assign n4099 = n4098 ^ n4090 ^ 1'b0 ;
  assign n4100 = ( x62 & n4098 ) | ( x62 & ~n4099 ) | ( n4098 & ~n4099 ) ;
  assign n4101 = n2292 | n3979 ;
  assign n4102 = x299 & ~n4088 ;
  assign n4103 = n4101 | n4102 ;
  assign n4104 = n2067 & ~n4103 ;
  assign n4105 = n2044 & ~n4103 ;
  assign n4106 = x299 & n4096 ;
  assign n4107 = n4101 | n4106 ;
  assign n4108 = n4107 ^ n2036 ^ 1'b0 ;
  assign n4109 = ( n4103 & n4107 ) | ( n4103 & n4108 ) | ( n4107 & n4108 ) ;
  assign n4110 = n2044 | n4109 ;
  assign n4111 = ( x92 & n4105 ) | ( x92 & n4110 ) | ( n4105 & n4110 ) ;
  assign n4112 = ~n4105 & n4111 ;
  assign n4113 = x75 & ~n4103 ;
  assign n4114 = x87 & n4109 ;
  assign n4115 = x38 & ~n4103 ;
  assign n4116 = x39 & n4107 ;
  assign n4117 = ~x878 & n2311 ;
  assign n4118 = x168 | n4117 ;
  assign n4119 = x878 & ~n2230 ;
  assign n4120 = x878 | n2319 ;
  assign n4121 = ( x168 & n4119 ) | ( x168 & n4120 ) | ( n4119 & n4120 ) ;
  assign n4122 = ~n4119 & n4121 ;
  assign n4123 = ( x228 & n4118 ) | ( x228 & ~n4122 ) | ( n4118 & ~n4122 ) ;
  assign n4124 = n4123 ^ n4118 ^ 1'b0 ;
  assign n4125 = ( x228 & n4123 ) | ( x228 & ~n4124 ) | ( n4123 & ~n4124 ) ;
  assign n4126 = ( n2742 & ~n3959 ) | ( n2742 & n4125 ) | ( ~n3959 & n4125 ) ;
  assign n4127 = ~n2742 & n4126 ;
  assign n4128 = ( x221 & n3945 ) | ( x221 & ~n4127 ) | ( n3945 & ~n4127 ) ;
  assign n4129 = n4127 | n4128 ;
  assign n4130 = n4129 ^ n3952 ^ 1'b0 ;
  assign n4131 = ( n3952 & n4129 ) | ( n3952 & n4130 ) | ( n4129 & n4130 ) ;
  assign n4132 = ( x215 & ~n3952 ) | ( x215 & n4131 ) | ( ~n3952 & n4131 ) ;
  assign n4133 = ( n3998 & ~n4028 ) | ( n3998 & n4132 ) | ( ~n4028 & n4132 ) ;
  assign n4134 = n4028 ^ n3998 ^ 1'b0 ;
  assign n4135 = ( n4028 & ~n4133 ) | ( n4028 & n4134 ) | ( ~n4133 & n4134 ) ;
  assign n4136 = ( x38 & ~n4116 ) | ( x38 & n4135 ) | ( ~n4116 & n4135 ) ;
  assign n4137 = n4116 | n4136 ;
  assign n4138 = ( x100 & ~n4115 ) | ( x100 & n4137 ) | ( ~n4115 & n4137 ) ;
  assign n4139 = ~x100 & n4138 ;
  assign n4140 = n1994 & ~n4103 ;
  assign n4141 = x100 & ~n4140 ;
  assign n4142 = n3987 | n4091 ;
  assign n4143 = ~n3953 & n4142 ;
  assign n4144 = ( ~x215 & n3952 ) | ( ~x215 & n4143 ) | ( n3952 & n4143 ) ;
  assign n4145 = ~x215 & n4144 ;
  assign n4146 = ( x299 & n3948 ) | ( x299 & n4145 ) | ( n3948 & n4145 ) ;
  assign n4147 = n4145 ^ n3948 ^ 1'b0 ;
  assign n4148 = ( x299 & n4146 ) | ( x299 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = ( n1994 & n4101 ) | ( n1994 & ~n4148 ) | ( n4101 & ~n4148 ) ;
  assign n4150 = n4148 | n4149 ;
  assign n4151 = n4141 & n4150 ;
  assign n4152 = ( ~x87 & n4139 ) | ( ~x87 & n4151 ) | ( n4139 & n4151 ) ;
  assign n4153 = ~x87 & n4152 ;
  assign n4154 = ( x75 & ~n4114 ) | ( x75 & n4153 ) | ( ~n4114 & n4153 ) ;
  assign n4155 = n4114 | n4154 ;
  assign n4156 = ( x92 & ~n4113 ) | ( x92 & n4155 ) | ( ~n4113 & n4155 ) ;
  assign n4157 = ~x92 & n4156 ;
  assign n4158 = ( n2067 & ~n4112 ) | ( n2067 & n4157 ) | ( ~n4112 & n4157 ) ;
  assign n4159 = n4112 | n4158 ;
  assign n4160 = ( x55 & ~n4104 ) | ( x55 & n4159 ) | ( ~n4104 & n4159 ) ;
  assign n4161 = ~x55 & n4160 ;
  assign n4162 = n2070 | n4096 ;
  assign n4163 = n4162 ^ x56 ^ 1'b0 ;
  assign n4164 = ( x55 & n3946 ) | ( x55 & n4067 ) | ( n3946 & n4067 ) ;
  assign n4165 = ( n4162 & ~n4163 ) | ( n4162 & n4164 ) | ( ~n4163 & n4164 ) ;
  assign n4166 = ( x56 & n4163 ) | ( x56 & n4165 ) | ( n4163 & n4165 ) ;
  assign n4167 = ( ~n4100 & n4161 ) | ( ~n4100 & n4166 ) | ( n4161 & n4166 ) ;
  assign n4168 = ~n4100 & n4167 ;
  assign n4169 = x240 & ~n2120 ;
  assign n4170 = n2151 & n4088 ;
  assign n4171 = n2151 | n4096 ;
  assign n4172 = ( x62 & n4170 ) | ( x62 & n4171 ) | ( n4170 & n4171 ) ;
  assign n4173 = ~n4170 & n4172 ;
  assign n4174 = ( n4168 & n4169 ) | ( n4168 & ~n4173 ) | ( n4169 & ~n4173 ) ;
  assign n4175 = ~n4168 & n4174 ;
  assign n4176 = ( n3967 & n4087 ) | ( n3967 & ~n4175 ) | ( n4087 & ~n4175 ) ;
  assign n4177 = ~n3967 & n4176 ;
  assign n4178 = x224 | x875 ;
  assign n4179 = n1224 | n4178 ;
  assign n4180 = x224 & ~x266 ;
  assign n4181 = ( x222 & n4179 ) | ( x222 & ~n4180 ) | ( n4179 & ~n4180 ) ;
  assign n4182 = ~x222 & n4181 ;
  assign n4183 = x1136 | n1208 ;
  assign n4184 = ( x222 & x928 ) | ( x222 & n1219 ) | ( x928 & n1219 ) ;
  assign n4185 = n4183 & n4184 ;
  assign n4186 = n4182 | n4185 ;
  assign n4187 = x1136 ^ x223 ^ 1'b0 ;
  assign n4188 = ( x1136 & n4186 ) | ( x1136 & ~n4187 ) | ( n4186 & ~n4187 ) ;
  assign n4189 = ~x299 & n4188 ;
  assign n4190 = x875 & ~n1224 ;
  assign n4191 = n1360 | n4190 ;
  assign n4192 = n4189 & n4191 ;
  assign n4193 = x215 & x1136 ;
  assign n4194 = ~x928 & n1315 ;
  assign n4195 = x1136 | n1315 ;
  assign n4196 = ( x221 & n4194 ) | ( x221 & n4195 ) | ( n4194 & n4195 ) ;
  assign n4197 = ~n4194 & n4196 ;
  assign n4198 = x266 ^ x216 ^ 1'b0 ;
  assign n4199 = x166 ^ x105 ^ 1'b0 ;
  assign n4200 = ( x166 & n4190 ) | ( x166 & n4199 ) | ( n4190 & n4199 ) ;
  assign n4201 = x228 ^ x166 ^ 1'b0 ;
  assign n4202 = ( x166 & n4200 ) | ( x166 & n4201 ) | ( n4200 & n4201 ) ;
  assign n4203 = ( x266 & ~n4198 ) | ( x266 & n4202 ) | ( ~n4198 & n4202 ) ;
  assign n4204 = x221 | n4203 ;
  assign n4205 = ( ~x221 & n4197 ) | ( ~x221 & n4204 ) | ( n4197 & n4204 ) ;
  assign n4206 = x215 | n4205 ;
  assign n4207 = ( ~x215 & n4193 ) | ( ~x215 & n4206 ) | ( n4193 & n4206 ) ;
  assign n4208 = x299 & n4207 ;
  assign n4209 = n4192 | n4208 ;
  assign n4210 = n1994 & ~n4209 ;
  assign n4211 = x100 & ~n4210 ;
  assign n4212 = x216 & x266 ;
  assign n4213 = x228 & n4200 ;
  assign n4214 = x875 | n2197 ;
  assign n4215 = x166 & n4214 ;
  assign n4216 = ~n1328 & n2195 ;
  assign n4217 = n1328 & n2197 ;
  assign n4218 = ( x875 & n4216 ) | ( x875 & ~n4217 ) | ( n4216 & ~n4217 ) ;
  assign n4219 = ~n4216 & n4218 ;
  assign n4220 = ( ~x228 & n4215 ) | ( ~x228 & n4219 ) | ( n4215 & n4219 ) ;
  assign n4221 = ~x228 & n4220 ;
  assign n4222 = ( ~x216 & n4213 ) | ( ~x216 & n4221 ) | ( n4213 & n4221 ) ;
  assign n4223 = ( ~x221 & n4212 ) | ( ~x221 & n4222 ) | ( n4212 & n4222 ) ;
  assign n4224 = ~x221 & n4223 ;
  assign n4225 = ( ~x215 & n4197 ) | ( ~x215 & n4224 ) | ( n4197 & n4224 ) ;
  assign n4226 = ~x215 & n4225 ;
  assign n4227 = ( x299 & n4193 ) | ( x299 & n4226 ) | ( n4193 & n4226 ) ;
  assign n4228 = n4226 ^ n4193 ^ 1'b0 ;
  assign n4229 = ( x299 & n4227 ) | ( x299 & n4228 ) | ( n4227 & n4228 ) ;
  assign n4230 = ( n1994 & n4192 ) | ( n1994 & ~n4229 ) | ( n4192 & ~n4229 ) ;
  assign n4231 = n4229 | n4230 ;
  assign n4232 = n4211 & n4231 ;
  assign n4233 = x228 & ~n2318 ;
  assign n4234 = ~n4200 & n4233 ;
  assign n4235 = x166 & n2319 ;
  assign n4236 = x166 | n2311 ;
  assign n4237 = ( x875 & n4235 ) | ( x875 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = x166 & ~x875 ;
  assign n4240 = ( ~n2230 & n4238 ) | ( ~n2230 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4241 = n4238 ^ n2230 ^ 1'b0 ;
  assign n4242 = ( n4238 & n4240 ) | ( n4238 & ~n4241 ) | ( n4240 & ~n4241 ) ;
  assign n4243 = ( ~n2318 & n2320 ) | ( ~n2318 & n4242 ) | ( n2320 & n4242 ) ;
  assign n4244 = ( x216 & ~n4234 ) | ( x216 & n4243 ) | ( ~n4234 & n4243 ) ;
  assign n4245 = ~x216 & n4244 ;
  assign n4246 = ( ~x221 & n4212 ) | ( ~x221 & n4245 ) | ( n4212 & n4245 ) ;
  assign n4247 = ~x221 & n4246 ;
  assign n4248 = ( ~x215 & n4197 ) | ( ~x215 & n4247 ) | ( n4197 & n4247 ) ;
  assign n4249 = ~x215 & n4248 ;
  assign n4250 = ( x299 & n4193 ) | ( x299 & ~n4249 ) | ( n4193 & ~n4249 ) ;
  assign n4251 = ~n4193 & n4250 ;
  assign n4252 = x223 & x1136 ;
  assign n4253 = x299 | n4252 ;
  assign n4254 = ~n1359 & n2314 ;
  assign n4255 = n4186 | n4254 ;
  assign n4256 = ~x223 & n4255 ;
  assign n4257 = ( ~x39 & n4253 ) | ( ~x39 & n4256 ) | ( n4253 & n4256 ) ;
  assign n4258 = ~x39 & n4257 ;
  assign n4259 = n4182 & ~n4254 ;
  assign n4260 = n4185 | n4253 ;
  assign n4261 = n4259 | n4260 ;
  assign n4262 = ( n4251 & n4258 ) | ( n4251 & n4261 ) | ( n4258 & n4261 ) ;
  assign n4263 = ~n4251 & n4262 ;
  assign n4264 = ~x166 & n1292 ;
  assign n4265 = x228 | n4264 ;
  assign n4266 = ( x875 & n1292 ) | ( x875 & ~n4265 ) | ( n1292 & ~n4265 ) ;
  assign n4267 = ~n4265 & n4266 ;
  assign n4268 = n4213 | n4267 ;
  assign n4269 = ( x266 & ~n4198 ) | ( x266 & n4268 ) | ( ~n4198 & n4268 ) ;
  assign n4270 = x221 | n4269 ;
  assign n4271 = ( ~x221 & n4197 ) | ( ~x221 & n4270 ) | ( n4197 & n4270 ) ;
  assign n4272 = x215 | n4271 ;
  assign n4273 = ( ~x215 & n4193 ) | ( ~x215 & n4272 ) | ( n4193 & n4272 ) ;
  assign n4274 = x299 & n4273 ;
  assign n4275 = n4192 | n4274 ;
  assign n4276 = x39 & n4275 ;
  assign n4277 = ( x38 & ~n4263 ) | ( x38 & n4276 ) | ( ~n4263 & n4276 ) ;
  assign n4278 = n4263 | n4277 ;
  assign n4279 = x38 & ~n4209 ;
  assign n4280 = ( x100 & n4278 ) | ( x100 & ~n4279 ) | ( n4278 & ~n4279 ) ;
  assign n4281 = ~x100 & n4280 ;
  assign n4282 = ( ~x87 & n4232 ) | ( ~x87 & n4281 ) | ( n4232 & n4281 ) ;
  assign n4283 = ~x87 & n4282 ;
  assign n4284 = n4275 ^ n2036 ^ 1'b0 ;
  assign n4285 = ( n4209 & n4275 ) | ( n4209 & n4284 ) | ( n4275 & n4284 ) ;
  assign n4286 = x87 & n4285 ;
  assign n4287 = ( x75 & ~n4283 ) | ( x75 & n4286 ) | ( ~n4283 & n4286 ) ;
  assign n4288 = n4283 | n4287 ;
  assign n4289 = x75 & ~n4209 ;
  assign n4290 = ( x92 & n4288 ) | ( x92 & ~n4289 ) | ( n4288 & ~n4289 ) ;
  assign n4291 = ~x92 & n4290 ;
  assign n4292 = n2044 & ~n4209 ;
  assign n4293 = n2044 | n4285 ;
  assign n4294 = ( x92 & n4292 ) | ( x92 & n4293 ) | ( n4292 & n4293 ) ;
  assign n4295 = ~n4292 & n4294 ;
  assign n4296 = ( n2067 & ~n4291 ) | ( n2067 & n4295 ) | ( ~n4291 & n4295 ) ;
  assign n4297 = n4291 | n4296 ;
  assign n4298 = n2070 | n4273 ;
  assign n4299 = n4298 ^ x56 ^ 1'b0 ;
  assign n4300 = n2070 & ~n4207 ;
  assign n4301 = x55 & ~n4300 ;
  assign n4302 = ( n4298 & ~n4299 ) | ( n4298 & n4301 ) | ( ~n4299 & n4301 ) ;
  assign n4303 = ( x56 & n4299 ) | ( x56 & n4302 ) | ( n4299 & n4302 ) ;
  assign n4304 = n2067 & ~n4209 ;
  assign n4305 = x55 | n4304 ;
  assign n4306 = ~n4303 & n4305 ;
  assign n4307 = ( n4297 & n4303 ) | ( n4297 & ~n4306 ) | ( n4303 & ~n4306 ) ;
  assign n4308 = n2099 & n4207 ;
  assign n4309 = ~n2099 & n4273 ;
  assign n4310 = ( x56 & n4308 ) | ( x56 & ~n4309 ) | ( n4308 & ~n4309 ) ;
  assign n4311 = ~n4308 & n4310 ;
  assign n4312 = ( x62 & n4307 ) | ( x62 & ~n4311 ) | ( n4307 & ~n4311 ) ;
  assign n4313 = ~x62 & n4312 ;
  assign n4314 = n2151 & ~n4207 ;
  assign n4315 = n2151 | n4273 ;
  assign n4316 = ( x62 & n4314 ) | ( x62 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4317 = ~n4314 & n4316 ;
  assign n4318 = ( n2120 & ~n4313 ) | ( n2120 & n4317 ) | ( ~n4313 & n4317 ) ;
  assign n4319 = n4313 | n4318 ;
  assign n4320 = n2266 | n4207 ;
  assign n4321 = n2120 & ~n4320 ;
  assign n4322 = x245 & ~n4321 ;
  assign n4323 = n2151 & ~n4320 ;
  assign n4324 = n2265 | n4213 ;
  assign n4325 = n4267 | n4324 ;
  assign n4326 = ( x266 & ~n4198 ) | ( x266 & n4325 ) | ( ~n4198 & n4325 ) ;
  assign n4327 = x221 | n4326 ;
  assign n4328 = ( ~x221 & n4197 ) | ( ~x221 & n4327 ) | ( n4197 & n4327 ) ;
  assign n4329 = x215 | n4328 ;
  assign n4330 = ( ~x215 & n4193 ) | ( ~x215 & n4329 ) | ( n4193 & n4329 ) ;
  assign n4331 = n2151 | n4330 ;
  assign n4332 = ( x62 & n4323 ) | ( x62 & n4331 ) | ( n4323 & n4331 ) ;
  assign n4333 = ~n4323 & n4332 ;
  assign n4334 = n2099 & n4320 ;
  assign n4335 = x56 & ~n4334 ;
  assign n4336 = ~n2099 & n4330 ;
  assign n4337 = ( x62 & n4335 ) | ( x62 & ~n4336 ) | ( n4335 & ~n4336 ) ;
  assign n4338 = n4337 ^ n4335 ^ 1'b0 ;
  assign n4339 = ( x62 & n4337 ) | ( x62 & ~n4338 ) | ( n4337 & ~n4338 ) ;
  assign n4340 = n4188 ^ x299 ^ 1'b0 ;
  assign n4341 = ( n4188 & n4320 ) | ( n4188 & n4340 ) | ( n4320 & n4340 ) ;
  assign n4342 = n2067 & ~n4341 ;
  assign n4343 = n2044 & ~n4341 ;
  assign n4344 = ( n4188 & n4330 ) | ( n4188 & n4340 ) | ( n4330 & n4340 ) ;
  assign n4345 = n4344 ^ n2036 ^ 1'b0 ;
  assign n4346 = ( n4341 & n4344 ) | ( n4341 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4347 = n2044 | n4346 ;
  assign n4348 = ( x92 & n4343 ) | ( x92 & n4347 ) | ( n4343 & n4347 ) ;
  assign n4349 = ~n4343 & n4348 ;
  assign n4350 = x75 & ~n4341 ;
  assign n4351 = x87 & n4346 ;
  assign n4352 = x38 & ~n4341 ;
  assign n4353 = x39 & n4344 ;
  assign n4354 = x299 & ~n4193 ;
  assign n4355 = x166 & n2311 ;
  assign n4356 = x166 | n2319 ;
  assign n4357 = ( x875 & ~n4355 ) | ( x875 & n4356 ) | ( ~n4355 & n4356 ) ;
  assign n4358 = ~x875 & n4357 ;
  assign n4359 = x166 | n2230 ;
  assign n4360 = x875 & n4359 ;
  assign n4361 = ( x228 & ~n4358 ) | ( x228 & n4360 ) | ( ~n4358 & n4360 ) ;
  assign n4362 = n4358 | n4361 ;
  assign n4363 = ( x216 & ~n4234 ) | ( x216 & n4362 ) | ( ~n4234 & n4362 ) ;
  assign n4364 = ~x216 & n4363 ;
  assign n4365 = ( ~x221 & n4212 ) | ( ~x221 & n4364 ) | ( n4212 & n4364 ) ;
  assign n4366 = ~x221 & n4365 ;
  assign n4367 = ( ~x215 & n4197 ) | ( ~x215 & n4366 ) | ( n4197 & n4366 ) ;
  assign n4368 = ~x215 & n4367 ;
  assign n4369 = ( n4258 & ~n4354 ) | ( n4258 & n4368 ) | ( ~n4354 & n4368 ) ;
  assign n4370 = n4354 ^ n4258 ^ 1'b0 ;
  assign n4371 = ( n4258 & n4369 ) | ( n4258 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = ( x38 & ~n4353 ) | ( x38 & n4371 ) | ( ~n4353 & n4371 ) ;
  assign n4373 = n4353 | n4372 ;
  assign n4374 = ( x100 & ~n4352 ) | ( x100 & n4373 ) | ( ~n4352 & n4373 ) ;
  assign n4375 = ~x100 & n4374 ;
  assign n4376 = n1994 & ~n4341 ;
  assign n4377 = x100 & ~n4376 ;
  assign n4378 = n4221 | n4324 ;
  assign n4379 = ~x216 & n4378 ;
  assign n4380 = ( ~x221 & n4212 ) | ( ~x221 & n4379 ) | ( n4212 & n4379 ) ;
  assign n4381 = ~x221 & n4380 ;
  assign n4382 = ( ~x215 & n4197 ) | ( ~x215 & n4381 ) | ( n4197 & n4381 ) ;
  assign n4383 = ~x215 & n4382 ;
  assign n4384 = ( x299 & n4193 ) | ( x299 & n4383 ) | ( n4193 & n4383 ) ;
  assign n4385 = n4383 ^ n4193 ^ 1'b0 ;
  assign n4386 = ( x299 & n4384 ) | ( x299 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4387 = ( n1994 & n4189 ) | ( n1994 & ~n4386 ) | ( n4189 & ~n4386 ) ;
  assign n4388 = n4386 | n4387 ;
  assign n4389 = n4377 & n4388 ;
  assign n4390 = ( ~x87 & n4375 ) | ( ~x87 & n4389 ) | ( n4375 & n4389 ) ;
  assign n4391 = ~x87 & n4390 ;
  assign n4392 = ( x75 & ~n4351 ) | ( x75 & n4391 ) | ( ~n4351 & n4391 ) ;
  assign n4393 = n4351 | n4392 ;
  assign n4394 = ( x92 & ~n4350 ) | ( x92 & n4393 ) | ( ~n4350 & n4393 ) ;
  assign n4395 = ~x92 & n4394 ;
  assign n4396 = ( n2067 & ~n4349 ) | ( n2067 & n4395 ) | ( ~n4349 & n4395 ) ;
  assign n4397 = n4349 | n4396 ;
  assign n4398 = ( x55 & ~n4342 ) | ( x55 & n4397 ) | ( ~n4342 & n4397 ) ;
  assign n4399 = ~x55 & n4398 ;
  assign n4400 = n2070 | n4330 ;
  assign n4401 = n4400 ^ x56 ^ 1'b0 ;
  assign n4402 = ( x55 & n2266 ) | ( x55 & n4301 ) | ( n2266 & n4301 ) ;
  assign n4403 = ( n4400 & ~n4401 ) | ( n4400 & n4402 ) | ( ~n4401 & n4402 ) ;
  assign n4404 = ( x56 & n4401 ) | ( x56 & n4403 ) | ( n4401 & n4403 ) ;
  assign n4405 = ( ~n4339 & n4399 ) | ( ~n4339 & n4404 ) | ( n4399 & n4404 ) ;
  assign n4406 = ~n4339 & n4405 ;
  assign n4407 = ( n2120 & ~n4333 ) | ( n2120 & n4406 ) | ( ~n4333 & n4406 ) ;
  assign n4408 = n4333 | n4407 ;
  assign n4409 = n4322 & n4408 ;
  assign n4410 = n2120 & ~n4207 ;
  assign n4411 = x245 | n4410 ;
  assign n4412 = ~n4409 & n4411 ;
  assign n4413 = ( n4319 & n4409 ) | ( n4319 & ~n4412 ) | ( n4409 & ~n4412 ) ;
  assign n4414 = x223 & x1135 ;
  assign n4415 = x1135 | n1208 ;
  assign n4416 = x222 & n4415 ;
  assign n4417 = x224 | x879 ;
  assign n4418 = n1224 | n4417 ;
  assign n4419 = x224 & ~x279 ;
  assign n4420 = ( x222 & n4418 ) | ( x222 & ~n4419 ) | ( n4418 & ~n4419 ) ;
  assign n4421 = ~x222 & n4420 ;
  assign n4422 = ~x938 & n1208 ;
  assign n4423 = ~n4421 & n4422 ;
  assign n4424 = ( n4416 & n4421 ) | ( n4416 & ~n4423 ) | ( n4421 & ~n4423 ) ;
  assign n4425 = ~x223 & n4424 ;
  assign n4426 = n4414 | n4425 ;
  assign n4427 = ~x299 & n4426 ;
  assign n4428 = x879 & ~n1224 ;
  assign n4429 = n1360 | n4428 ;
  assign n4430 = n4427 & n4429 ;
  assign n4431 = x215 & x1135 ;
  assign n4432 = ~x938 & n1315 ;
  assign n4433 = x1135 | n1315 ;
  assign n4434 = ( x221 & n4432 ) | ( x221 & n4433 ) | ( n4432 & n4433 ) ;
  assign n4435 = ~n4432 & n4434 ;
  assign n4436 = x279 ^ x216 ^ 1'b0 ;
  assign n4437 = x161 ^ x105 ^ 1'b0 ;
  assign n4438 = ( x161 & n4428 ) | ( x161 & n4437 ) | ( n4428 & n4437 ) ;
  assign n4439 = x228 & n4438 ;
  assign n4440 = x161 & ~x228 ;
  assign n4441 = n4439 | n4440 ;
  assign n4442 = ( x279 & ~n4436 ) | ( x279 & n4441 ) | ( ~n4436 & n4441 ) ;
  assign n4443 = x221 | n4442 ;
  assign n4444 = ( ~x221 & n4435 ) | ( ~x221 & n4443 ) | ( n4435 & n4443 ) ;
  assign n4445 = x215 | n4444 ;
  assign n4446 = ( ~x215 & n4431 ) | ( ~x215 & n4445 ) | ( n4431 & n4445 ) ;
  assign n4447 = x299 & n4446 ;
  assign n4448 = n4430 | n4447 ;
  assign n4449 = n1994 & ~n4448 ;
  assign n4450 = x100 & ~n4449 ;
  assign n4451 = x216 & x279 ;
  assign n4452 = x879 | n2197 ;
  assign n4453 = x161 & n4452 ;
  assign n4454 = x152 | x166 ;
  assign n4455 = n2195 & ~n4454 ;
  assign n4456 = n2197 & n4454 ;
  assign n4457 = ( x879 & n4455 ) | ( x879 & ~n4456 ) | ( n4455 & ~n4456 ) ;
  assign n4458 = ~n4455 & n4457 ;
  assign n4459 = ( ~x228 & n4453 ) | ( ~x228 & n4458 ) | ( n4453 & n4458 ) ;
  assign n4460 = ~x228 & n4459 ;
  assign n4461 = ( ~x216 & n4439 ) | ( ~x216 & n4460 ) | ( n4439 & n4460 ) ;
  assign n4462 = ( ~x221 & n4451 ) | ( ~x221 & n4461 ) | ( n4451 & n4461 ) ;
  assign n4463 = ~x221 & n4462 ;
  assign n4464 = ( ~x215 & n4435 ) | ( ~x215 & n4463 ) | ( n4435 & n4463 ) ;
  assign n4465 = ~x215 & n4464 ;
  assign n4466 = ( x299 & n4431 ) | ( x299 & n4465 ) | ( n4431 & n4465 ) ;
  assign n4467 = n4465 ^ n4431 ^ 1'b0 ;
  assign n4468 = ( x299 & n4466 ) | ( x299 & n4467 ) | ( n4466 & n4467 ) ;
  assign n4469 = ( n1994 & n4430 ) | ( n1994 & ~n4468 ) | ( n4430 & ~n4468 ) ;
  assign n4470 = n4468 | n4469 ;
  assign n4471 = n4450 & n4470 ;
  assign n4472 = n4233 & ~n4438 ;
  assign n4473 = x161 & n2319 ;
  assign n4474 = x161 | n2311 ;
  assign n4475 = ( x879 & n4473 ) | ( x879 & n4474 ) | ( n4473 & n4474 ) ;
  assign n4476 = ~n4473 & n4475 ;
  assign n4477 = x161 & ~x879 ;
  assign n4478 = ( ~n2230 & n4476 ) | ( ~n2230 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4479 = n4476 ^ n2230 ^ 1'b0 ;
  assign n4480 = ( n4476 & n4478 ) | ( n4476 & ~n4479 ) | ( n4478 & ~n4479 ) ;
  assign n4481 = ( ~n2318 & n2320 ) | ( ~n2318 & n4480 ) | ( n2320 & n4480 ) ;
  assign n4482 = ( x216 & ~n4472 ) | ( x216 & n4481 ) | ( ~n4472 & n4481 ) ;
  assign n4483 = ~x216 & n4482 ;
  assign n4484 = ( ~x221 & n4451 ) | ( ~x221 & n4483 ) | ( n4451 & n4483 ) ;
  assign n4485 = ~x221 & n4484 ;
  assign n4486 = ( ~x215 & n4435 ) | ( ~x215 & n4485 ) | ( n4435 & n4485 ) ;
  assign n4487 = ~x215 & n4486 ;
  assign n4488 = ( x299 & n4431 ) | ( x299 & ~n4487 ) | ( n4431 & ~n4487 ) ;
  assign n4489 = ~n4431 & n4488 ;
  assign n4490 = x299 | n4414 ;
  assign n4491 = ( x222 & n4415 ) | ( x222 & n4422 ) | ( n4415 & n4422 ) ;
  assign n4492 = ~n4422 & n4491 ;
  assign n4493 = n4254 & ~n4492 ;
  assign n4494 = n4425 & ~n4493 ;
  assign n4495 = n4490 | n4494 ;
  assign n4496 = ( x39 & ~n4489 ) | ( x39 & n4495 ) | ( ~n4489 & n4495 ) ;
  assign n4497 = ~x39 & n4496 ;
  assign n4498 = n2142 & ~n4440 ;
  assign n4499 = x879 | n1292 ;
  assign n4500 = ~n4498 & n4499 ;
  assign n4501 = n4439 | n4500 ;
  assign n4502 = ( x279 & ~n4436 ) | ( x279 & n4501 ) | ( ~n4436 & n4501 ) ;
  assign n4503 = x221 | n4502 ;
  assign n4504 = ( ~x221 & n4435 ) | ( ~x221 & n4503 ) | ( n4435 & n4503 ) ;
  assign n4505 = x215 | n4504 ;
  assign n4506 = ( ~x215 & n4431 ) | ( ~x215 & n4505 ) | ( n4431 & n4505 ) ;
  assign n4507 = x299 & n4506 ;
  assign n4508 = n4430 | n4507 ;
  assign n4509 = x39 & n4508 ;
  assign n4510 = ( x38 & ~n4497 ) | ( x38 & n4509 ) | ( ~n4497 & n4509 ) ;
  assign n4511 = n4497 | n4510 ;
  assign n4512 = x38 & ~n4448 ;
  assign n4513 = ( x100 & n4511 ) | ( x100 & ~n4512 ) | ( n4511 & ~n4512 ) ;
  assign n4514 = ~x100 & n4513 ;
  assign n4515 = ( ~x87 & n4471 ) | ( ~x87 & n4514 ) | ( n4471 & n4514 ) ;
  assign n4516 = ~x87 & n4515 ;
  assign n4517 = n4508 ^ n2036 ^ 1'b0 ;
  assign n4518 = ( n4448 & n4508 ) | ( n4448 & n4517 ) | ( n4508 & n4517 ) ;
  assign n4519 = x87 & n4518 ;
  assign n4520 = ( x75 & ~n4516 ) | ( x75 & n4519 ) | ( ~n4516 & n4519 ) ;
  assign n4521 = n4516 | n4520 ;
  assign n4522 = x75 & ~n4448 ;
  assign n4523 = ( x92 & n4521 ) | ( x92 & ~n4522 ) | ( n4521 & ~n4522 ) ;
  assign n4524 = ~x92 & n4523 ;
  assign n4525 = n2044 & ~n4448 ;
  assign n4526 = n2044 | n4518 ;
  assign n4527 = ( x92 & n4525 ) | ( x92 & n4526 ) | ( n4525 & n4526 ) ;
  assign n4528 = ~n4525 & n4527 ;
  assign n4529 = ( n2067 & ~n4524 ) | ( n2067 & n4528 ) | ( ~n4524 & n4528 ) ;
  assign n4530 = n4524 | n4529 ;
  assign n4531 = n2070 | n4506 ;
  assign n4532 = n4531 ^ x56 ^ 1'b0 ;
  assign n4533 = n2070 & ~n4446 ;
  assign n4534 = x55 & ~n4533 ;
  assign n4535 = ( n4531 & ~n4532 ) | ( n4531 & n4534 ) | ( ~n4532 & n4534 ) ;
  assign n4536 = ( x56 & n4532 ) | ( x56 & n4535 ) | ( n4532 & n4535 ) ;
  assign n4537 = n2067 & ~n4448 ;
  assign n4538 = x55 | n4537 ;
  assign n4539 = ~n4536 & n4538 ;
  assign n4540 = ( n4530 & n4536 ) | ( n4530 & ~n4539 ) | ( n4536 & ~n4539 ) ;
  assign n4541 = n2099 & n4446 ;
  assign n4542 = ~n2099 & n4506 ;
  assign n4543 = ( x56 & n4541 ) | ( x56 & ~n4542 ) | ( n4541 & ~n4542 ) ;
  assign n4544 = ~n4541 & n4543 ;
  assign n4545 = ( x62 & n4540 ) | ( x62 & ~n4544 ) | ( n4540 & ~n4544 ) ;
  assign n4546 = ~x62 & n4545 ;
  assign n4547 = n2151 & ~n4446 ;
  assign n4548 = n2151 | n4506 ;
  assign n4549 = ( x62 & n4547 ) | ( x62 & n4548 ) | ( n4547 & n4548 ) ;
  assign n4550 = ~n4547 & n4549 ;
  assign n4551 = ( n2120 & ~n4546 ) | ( n2120 & n4550 ) | ( ~n4546 & n4550 ) ;
  assign n4552 = n4546 | n4551 ;
  assign n4553 = n2266 | n4446 ;
  assign n4554 = n2120 & ~n4553 ;
  assign n4555 = x244 & ~n4554 ;
  assign n4556 = n2151 & ~n4553 ;
  assign n4557 = n2265 | n4439 ;
  assign n4558 = n4500 | n4557 ;
  assign n4559 = ( x279 & ~n4436 ) | ( x279 & n4558 ) | ( ~n4436 & n4558 ) ;
  assign n4560 = x221 | n4559 ;
  assign n4561 = ( ~x221 & n4435 ) | ( ~x221 & n4560 ) | ( n4435 & n4560 ) ;
  assign n4562 = x215 | n4561 ;
  assign n4563 = ( ~x215 & n4431 ) | ( ~x215 & n4562 ) | ( n4431 & n4562 ) ;
  assign n4564 = n2151 | n4563 ;
  assign n4565 = ( x62 & n4556 ) | ( x62 & n4564 ) | ( n4556 & n4564 ) ;
  assign n4566 = ~n4556 & n4565 ;
  assign n4567 = n2099 & n4553 ;
  assign n4568 = x56 & ~n4567 ;
  assign n4569 = ~n2099 & n4563 ;
  assign n4570 = ( x62 & n4568 ) | ( x62 & ~n4569 ) | ( n4568 & ~n4569 ) ;
  assign n4571 = n4570 ^ n4568 ^ 1'b0 ;
  assign n4572 = ( x62 & n4570 ) | ( x62 & ~n4571 ) | ( n4570 & ~n4571 ) ;
  assign n4573 = x299 & n4553 ;
  assign n4574 = n4427 | n4573 ;
  assign n4575 = n2067 & ~n4574 ;
  assign n4576 = n2044 & ~n4574 ;
  assign n4577 = x299 & n4563 ;
  assign n4578 = n4427 | n4577 ;
  assign n4579 = n4578 ^ n2036 ^ 1'b0 ;
  assign n4580 = ( n4574 & n4578 ) | ( n4574 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4581 = n2044 | n4580 ;
  assign n4582 = ( x92 & n4576 ) | ( x92 & n4581 ) | ( n4576 & n4581 ) ;
  assign n4583 = ~n4576 & n4582 ;
  assign n4584 = x75 & ~n4574 ;
  assign n4585 = x87 & n4580 ;
  assign n4586 = x38 & ~n4574 ;
  assign n4587 = x39 & n4578 ;
  assign n4588 = n4254 | n4424 ;
  assign n4589 = x223 | n4588 ;
  assign n4590 = ( ~x223 & n4490 ) | ( ~x223 & n4589 ) | ( n4490 & n4589 ) ;
  assign n4591 = x161 & n2311 ;
  assign n4592 = x161 | n2319 ;
  assign n4593 = ( x879 & ~n4591 ) | ( x879 & n4592 ) | ( ~n4591 & n4592 ) ;
  assign n4594 = ~x879 & n4593 ;
  assign n4595 = x161 | n2230 ;
  assign n4596 = x879 & n4595 ;
  assign n4597 = ( x228 & ~n4594 ) | ( x228 & n4596 ) | ( ~n4594 & n4596 ) ;
  assign n4598 = n4594 | n4597 ;
  assign n4599 = ( x216 & ~n4472 ) | ( x216 & n4598 ) | ( ~n4472 & n4598 ) ;
  assign n4600 = ~x216 & n4599 ;
  assign n4601 = ( ~x221 & n4451 ) | ( ~x221 & n4600 ) | ( n4451 & n4600 ) ;
  assign n4602 = ~x221 & n4601 ;
  assign n4603 = ( ~x215 & n4435 ) | ( ~x215 & n4602 ) | ( n4435 & n4602 ) ;
  assign n4604 = ~x215 & n4603 ;
  assign n4605 = ( x299 & n4431 ) | ( x299 & ~n4604 ) | ( n4431 & ~n4604 ) ;
  assign n4606 = ~n4431 & n4605 ;
  assign n4607 = ( x39 & n4590 ) | ( x39 & ~n4606 ) | ( n4590 & ~n4606 ) ;
  assign n4608 = ~x39 & n4607 ;
  assign n4609 = ( x38 & ~n4587 ) | ( x38 & n4608 ) | ( ~n4587 & n4608 ) ;
  assign n4610 = n4587 | n4609 ;
  assign n4611 = ( x100 & ~n4586 ) | ( x100 & n4610 ) | ( ~n4586 & n4610 ) ;
  assign n4612 = ~x100 & n4611 ;
  assign n4613 = n1994 & ~n4574 ;
  assign n4614 = x100 & ~n4613 ;
  assign n4615 = n4460 | n4557 ;
  assign n4616 = ~x216 & n4615 ;
  assign n4617 = ( ~x221 & n4451 ) | ( ~x221 & n4616 ) | ( n4451 & n4616 ) ;
  assign n4618 = ~x221 & n4617 ;
  assign n4619 = ( ~x215 & n4435 ) | ( ~x215 & n4618 ) | ( n4435 & n4618 ) ;
  assign n4620 = ~x215 & n4619 ;
  assign n4621 = ( x299 & n4431 ) | ( x299 & n4620 ) | ( n4431 & n4620 ) ;
  assign n4622 = n4620 ^ n4431 ^ 1'b0 ;
  assign n4623 = ( x299 & n4621 ) | ( x299 & n4622 ) | ( n4621 & n4622 ) ;
  assign n4624 = ( n1994 & n4427 ) | ( n1994 & ~n4623 ) | ( n4427 & ~n4623 ) ;
  assign n4625 = n4623 | n4624 ;
  assign n4626 = n4614 & n4625 ;
  assign n4627 = ( ~x87 & n4612 ) | ( ~x87 & n4626 ) | ( n4612 & n4626 ) ;
  assign n4628 = ~x87 & n4627 ;
  assign n4629 = ( x75 & ~n4585 ) | ( x75 & n4628 ) | ( ~n4585 & n4628 ) ;
  assign n4630 = n4585 | n4629 ;
  assign n4631 = ( x92 & ~n4584 ) | ( x92 & n4630 ) | ( ~n4584 & n4630 ) ;
  assign n4632 = ~x92 & n4631 ;
  assign n4633 = ( n2067 & ~n4583 ) | ( n2067 & n4632 ) | ( ~n4583 & n4632 ) ;
  assign n4634 = n4583 | n4633 ;
  assign n4635 = ( x55 & ~n4575 ) | ( x55 & n4634 ) | ( ~n4575 & n4634 ) ;
  assign n4636 = ~x55 & n4635 ;
  assign n4637 = n2070 | n4563 ;
  assign n4638 = n4637 ^ x56 ^ 1'b0 ;
  assign n4639 = ( x55 & n2266 ) | ( x55 & n4534 ) | ( n2266 & n4534 ) ;
  assign n4640 = ( n4637 & ~n4638 ) | ( n4637 & n4639 ) | ( ~n4638 & n4639 ) ;
  assign n4641 = ( x56 & n4638 ) | ( x56 & n4640 ) | ( n4638 & n4640 ) ;
  assign n4642 = ( ~n4572 & n4636 ) | ( ~n4572 & n4641 ) | ( n4636 & n4641 ) ;
  assign n4643 = ~n4572 & n4642 ;
  assign n4644 = ( n2120 & ~n4566 ) | ( n2120 & n4643 ) | ( ~n4566 & n4643 ) ;
  assign n4645 = n4566 | n4644 ;
  assign n4646 = n4555 & n4645 ;
  assign n4647 = n2120 & ~n4446 ;
  assign n4648 = x244 | n4647 ;
  assign n4649 = ~n4646 & n4648 ;
  assign n4650 = ( n4552 & n4646 ) | ( n4552 & ~n4649 ) | ( n4646 & ~n4649 ) ;
  assign n4651 = x833 & ~x930 ;
  assign n4652 = ~x216 & x221 ;
  assign n4653 = n4651 & n4652 ;
  assign n4654 = x846 & ~n1224 ;
  assign n4655 = x152 ^ x105 ^ 1'b0 ;
  assign n4656 = ( x152 & n4654 ) | ( x152 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = x228 ^ x152 ^ 1'b0 ;
  assign n4658 = ( x152 & n4656 ) | ( x152 & n4657 ) | ( n4656 & n4657 ) ;
  assign n4659 = x216 | n4658 ;
  assign n4660 = ( x221 & x278 ) | ( x221 & n2263 ) | ( x278 & n2263 ) ;
  assign n4661 = ( ~x216 & n4659 ) | ( ~x216 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = ~n4653 & n4661 ;
  assign n4663 = x215 | n4662 ;
  assign n4664 = n2266 | n4663 ;
  assign n4665 = n2120 & ~n4664 ;
  assign n4666 = x242 & ~n4665 ;
  assign n4667 = x228 & n4656 ;
  assign n4668 = n2265 | n4667 ;
  assign n4669 = ~x152 & n1292 ;
  assign n4670 = x228 | n4669 ;
  assign n4671 = ( x846 & n1292 ) | ( x846 & ~n4670 ) | ( n1292 & ~n4670 ) ;
  assign n4672 = ~n4670 & n4671 ;
  assign n4673 = n4668 | n4672 ;
  assign n4674 = x216 | n4673 ;
  assign n4675 = ( ~x216 & n4660 ) | ( ~x216 & n4674 ) | ( n4660 & n4674 ) ;
  assign n4676 = ~n4653 & n4675 ;
  assign n4677 = x215 | n4676 ;
  assign n4678 = n2151 | n4677 ;
  assign n4679 = n2151 & ~n4663 ;
  assign n4680 = x62 & ~n4679 ;
  assign n4681 = ( x62 & n2266 ) | ( x62 & n4680 ) | ( n2266 & n4680 ) ;
  assign n4682 = n4678 & n4681 ;
  assign n4683 = ~n2099 & n4677 ;
  assign n4684 = n2099 & n4664 ;
  assign n4685 = x56 & ~n4684 ;
  assign n4686 = n4685 ^ n4683 ^ 1'b0 ;
  assign n4687 = ( n4683 & n4685 ) | ( n4683 & n4686 ) | ( n4685 & n4686 ) ;
  assign n4688 = ( x62 & ~n4683 ) | ( x62 & n4687 ) | ( ~n4683 & n4687 ) ;
  assign n4689 = ~x224 & n4654 ;
  assign n4690 = ( x222 & x278 ) | ( x222 & n1359 ) | ( x278 & n1359 ) ;
  assign n4691 = n4689 | n4690 ;
  assign n4692 = x222 & ~x224 ;
  assign n4693 = n4651 & n4692 ;
  assign n4694 = n1220 | n4693 ;
  assign n4695 = n4691 & ~n4694 ;
  assign n4696 = x299 | n4695 ;
  assign n4697 = n2699 | n4696 ;
  assign n4698 = n1220 | n4697 ;
  assign n4699 = ~x299 & n4698 ;
  assign n4700 = ( n4664 & n4698 ) | ( n4664 & n4699 ) | ( n4698 & n4699 ) ;
  assign n4701 = n2067 & ~n4700 ;
  assign n4702 = n2044 & ~n4700 ;
  assign n4703 = x299 & n4677 ;
  assign n4704 = n4699 | n4703 ;
  assign n4705 = n4704 ^ n2036 ^ 1'b0 ;
  assign n4706 = ( n4700 & n4704 ) | ( n4700 & n4705 ) | ( n4704 & n4705 ) ;
  assign n4707 = n2044 | n4706 ;
  assign n4708 = ( x92 & n4702 ) | ( x92 & n4707 ) | ( n4702 & n4707 ) ;
  assign n4709 = ~n4702 & n4708 ;
  assign n4710 = x75 & ~n4700 ;
  assign n4711 = x87 & n4706 ;
  assign n4712 = x38 & ~n4700 ;
  assign n4713 = x39 & n4704 ;
  assign n4714 = x846 | n2314 ;
  assign n4715 = ~x224 & n4714 ;
  assign n4716 = n4690 | n4715 ;
  assign n4717 = ~n4693 & n4716 ;
  assign n4718 = n2290 | n4717 ;
  assign n4719 = ~x39 & n4718 ;
  assign n4720 = x105 & n4714 ;
  assign n4721 = ( x228 & n1323 ) | ( x228 & n4657 ) | ( n1323 & n4657 ) ;
  assign n4722 = ~n4720 & n4721 ;
  assign n4723 = ~x152 & x846 ;
  assign n4724 = ~n2230 & n4723 ;
  assign n4725 = ~x152 & n2319 ;
  assign n4726 = x152 & ~n2311 ;
  assign n4727 = ( x846 & ~n4725 ) | ( x846 & n4726 ) | ( ~n4725 & n4726 ) ;
  assign n4728 = n4725 | n4727 ;
  assign n4729 = n4728 ^ n4724 ^ 1'b0 ;
  assign n4730 = ( n4724 & n4728 ) | ( n4724 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = ( x228 & ~n4724 ) | ( x228 & n4730 ) | ( ~n4724 & n4730 ) ;
  assign n4732 = ( x216 & ~n4722 ) | ( x216 & n4731 ) | ( ~n4722 & n4731 ) ;
  assign n4733 = ~x216 & n4732 ;
  assign n4734 = ( ~n4653 & n4660 ) | ( ~n4653 & n4733 ) | ( n4660 & n4733 ) ;
  assign n4735 = ~n4653 & n4734 ;
  assign n4736 = ~x215 & x299 ;
  assign n4737 = ~n4735 & n4736 ;
  assign n4738 = n4719 & ~n4737 ;
  assign n4739 = ( x38 & ~n4713 ) | ( x38 & n4738 ) | ( ~n4713 & n4738 ) ;
  assign n4740 = n4713 | n4739 ;
  assign n4741 = ( x100 & ~n4712 ) | ( x100 & n4740 ) | ( ~n4712 & n4740 ) ;
  assign n4742 = ~x100 & n4741 ;
  assign n4743 = n1994 & ~n4700 ;
  assign n4744 = x100 & ~n4743 ;
  assign n4745 = x846 & ~n2203 ;
  assign n4746 = ( ~x228 & n2198 ) | ( ~x228 & n4745 ) | ( n2198 & n4745 ) ;
  assign n4747 = ~x228 & n4746 ;
  assign n4748 = n4668 | n4747 ;
  assign n4749 = x216 | n4748 ;
  assign n4750 = ( ~x216 & n4660 ) | ( ~x216 & n4749 ) | ( n4660 & n4749 ) ;
  assign n4751 = ~n4653 & n4750 ;
  assign n4752 = ( x215 & x299 ) | ( x215 & n4751 ) | ( x299 & n4751 ) ;
  assign n4753 = x299 & n4752 ;
  assign n4754 = ( n1994 & n4699 ) | ( n1994 & ~n4753 ) | ( n4699 & ~n4753 ) ;
  assign n4755 = n4753 | n4754 ;
  assign n4756 = n4744 & n4755 ;
  assign n4757 = ( ~x87 & n4742 ) | ( ~x87 & n4756 ) | ( n4742 & n4756 ) ;
  assign n4758 = ~x87 & n4757 ;
  assign n4759 = ( x75 & ~n4711 ) | ( x75 & n4758 ) | ( ~n4711 & n4758 ) ;
  assign n4760 = n4711 | n4759 ;
  assign n4761 = ( x92 & ~n4710 ) | ( x92 & n4760 ) | ( ~n4710 & n4760 ) ;
  assign n4762 = ~x92 & n4761 ;
  assign n4763 = ( n2067 & ~n4709 ) | ( n2067 & n4762 ) | ( ~n4709 & n4762 ) ;
  assign n4764 = n4709 | n4763 ;
  assign n4765 = ( x55 & ~n4701 ) | ( x55 & n4764 ) | ( ~n4701 & n4764 ) ;
  assign n4766 = ~x55 & n4765 ;
  assign n4767 = n2070 & ~n4663 ;
  assign n4768 = x55 & ~n4767 ;
  assign n4769 = ( x55 & n2266 ) | ( x55 & n4768 ) | ( n2266 & n4768 ) ;
  assign n4770 = n4769 ^ x56 ^ 1'b0 ;
  assign n4771 = n2070 | n4677 ;
  assign n4772 = ( n4769 & ~n4770 ) | ( n4769 & n4771 ) | ( ~n4770 & n4771 ) ;
  assign n4773 = ( x56 & n4770 ) | ( x56 & n4772 ) | ( n4770 & n4772 ) ;
  assign n4774 = ( ~n4688 & n4766 ) | ( ~n4688 & n4773 ) | ( n4766 & n4773 ) ;
  assign n4775 = ~n4688 & n4774 ;
  assign n4776 = ( n2120 & ~n4682 ) | ( n2120 & n4775 ) | ( ~n4682 & n4775 ) ;
  assign n4777 = n4682 | n4776 ;
  assign n4778 = n4666 & n4777 ;
  assign n4779 = x223 | n4691 ;
  assign n4780 = n4699 & n4779 ;
  assign n4781 = x299 & n4663 ;
  assign n4782 = n4780 | n4781 ;
  assign n4783 = x38 & ~n4782 ;
  assign n4784 = ( n4661 & n4672 ) | ( n4661 & n4675 ) | ( n4672 & n4675 ) ;
  assign n4785 = ( n4663 & n4677 ) | ( n4663 & n4784 ) | ( n4677 & n4784 ) ;
  assign n4786 = x299 & n4785 ;
  assign n4787 = n4780 | n4786 ;
  assign n4788 = x39 & n4787 ;
  assign n4789 = x216 | n4722 ;
  assign n4790 = n2314 & n4721 ;
  assign n4791 = x152 & ~x846 ;
  assign n4792 = ~n2230 & n4791 ;
  assign n4793 = x152 & n2319 ;
  assign n4794 = x846 & ~n4793 ;
  assign n4795 = ( n2311 & n4726 ) | ( n2311 & n4794 ) | ( n4726 & n4794 ) ;
  assign n4796 = ( x228 & ~n4792 ) | ( x228 & n4795 ) | ( ~n4792 & n4795 ) ;
  assign n4797 = n4792 | n4796 ;
  assign n4798 = ( n4789 & ~n4790 ) | ( n4789 & n4797 ) | ( ~n4790 & n4797 ) ;
  assign n4799 = ~n4789 & n4798 ;
  assign n4800 = ( ~n4653 & n4660 ) | ( ~n4653 & n4799 ) | ( n4660 & n4799 ) ;
  assign n4801 = ~n4653 & n4800 ;
  assign n4802 = n4736 & ~n4801 ;
  assign n4803 = ~n2313 & n4689 ;
  assign n4804 = n4690 | n4803 ;
  assign n4805 = n2290 | n4804 ;
  assign n4806 = ( n4719 & n4802 ) | ( n4719 & n4805 ) | ( n4802 & n4805 ) ;
  assign n4807 = ~n4802 & n4806 ;
  assign n4808 = ( x38 & ~n4788 ) | ( x38 & n4807 ) | ( ~n4788 & n4807 ) ;
  assign n4809 = n4788 | n4808 ;
  assign n4810 = ( x100 & ~n4783 ) | ( x100 & n4809 ) | ( ~n4783 & n4809 ) ;
  assign n4811 = ~x100 & n4810 ;
  assign n4812 = n1994 & ~n4782 ;
  assign n4813 = n4667 | n4747 ;
  assign n4814 = x216 | n4813 ;
  assign n4815 = ( ~x216 & n4660 ) | ( ~x216 & n4814 ) | ( n4660 & n4814 ) ;
  assign n4816 = ~n4653 & n4815 ;
  assign n4817 = ( x215 & x299 ) | ( x215 & n4816 ) | ( x299 & n4816 ) ;
  assign n4818 = x299 & n4817 ;
  assign n4819 = ( n1994 & n4780 ) | ( n1994 & ~n4818 ) | ( n4780 & ~n4818 ) ;
  assign n4820 = n4818 | n4819 ;
  assign n4821 = ( x100 & n4812 ) | ( x100 & n4820 ) | ( n4812 & n4820 ) ;
  assign n4822 = ~n4812 & n4821 ;
  assign n4823 = ( ~x87 & n4811 ) | ( ~x87 & n4822 ) | ( n4811 & n4822 ) ;
  assign n4824 = ~x87 & n4823 ;
  assign n4825 = n4787 ^ n2036 ^ 1'b0 ;
  assign n4826 = ( n4782 & n4787 ) | ( n4782 & n4825 ) | ( n4787 & n4825 ) ;
  assign n4827 = x87 & n4826 ;
  assign n4828 = ( x75 & ~n4824 ) | ( x75 & n4827 ) | ( ~n4824 & n4827 ) ;
  assign n4829 = n4824 | n4828 ;
  assign n4830 = ( x92 & n2046 ) | ( x92 & n4782 ) | ( n2046 & n4782 ) ;
  assign n4831 = n4830 ^ n2067 ^ 1'b0 ;
  assign n4832 = n2044 | n4826 ;
  assign n4833 = ( n4830 & ~n4831 ) | ( n4830 & n4832 ) | ( ~n4831 & n4832 ) ;
  assign n4834 = ( n2067 & n4831 ) | ( n2067 & n4833 ) | ( n4831 & n4833 ) ;
  assign n4835 = x75 & ~n4782 ;
  assign n4836 = x92 | n4835 ;
  assign n4837 = ~n4834 & n4836 ;
  assign n4838 = ( n4829 & n4834 ) | ( n4829 & ~n4837 ) | ( n4834 & ~n4837 ) ;
  assign n4839 = n4768 ^ x56 ^ 1'b0 ;
  assign n4840 = n2070 | n4785 ;
  assign n4841 = ( n4768 & ~n4839 ) | ( n4768 & n4840 ) | ( ~n4839 & n4840 ) ;
  assign n4842 = ( x56 & n4839 ) | ( x56 & n4841 ) | ( n4839 & n4841 ) ;
  assign n4843 = n2067 & ~n4782 ;
  assign n4844 = x55 | n4843 ;
  assign n4845 = ~n4842 & n4844 ;
  assign n4846 = ( n4838 & n4842 ) | ( n4838 & ~n4845 ) | ( n4842 & ~n4845 ) ;
  assign n4847 = n4680 ^ n2120 ^ 1'b0 ;
  assign n4848 = n2151 | n4785 ;
  assign n4849 = ( n4680 & ~n4847 ) | ( n4680 & n4848 ) | ( ~n4847 & n4848 ) ;
  assign n4850 = ( n2120 & n4847 ) | ( n2120 & n4849 ) | ( n4847 & n4849 ) ;
  assign n4851 = ~n2099 & n4785 ;
  assign n4852 = n2099 & n4663 ;
  assign n4853 = x56 & ~n4852 ;
  assign n4854 = n4853 ^ n4851 ^ 1'b0 ;
  assign n4855 = ( n4851 & n4853 ) | ( n4851 & n4854 ) | ( n4853 & n4854 ) ;
  assign n4856 = ( x62 & ~n4851 ) | ( x62 & n4855 ) | ( ~n4851 & n4855 ) ;
  assign n4857 = ~n4850 & n4856 ;
  assign n4858 = ( n4846 & n4850 ) | ( n4846 & ~n4857 ) | ( n4850 & ~n4857 ) ;
  assign n4859 = n2120 & ~n4663 ;
  assign n4860 = ( x242 & n4858 ) | ( x242 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  assign n4861 = ~x242 & n4860 ;
  assign n4862 = ( x1134 & n4778 ) | ( x1134 & ~n4861 ) | ( n4778 & ~n4861 ) ;
  assign n4863 = ~n4778 & n4862 ;
  assign n4864 = x221 & ~n1315 ;
  assign n4865 = x215 | n4864 ;
  assign n4866 = n4653 | n4865 ;
  assign n4867 = n4661 & ~n4866 ;
  assign n4868 = n2266 | n4867 ;
  assign n4869 = n2120 & n4868 ;
  assign n4870 = n1219 | n2290 ;
  assign n4871 = n4717 & ~n4870 ;
  assign n4872 = n4736 & ~n4864 ;
  assign n4873 = n4735 & n4872 ;
  assign n4874 = ( x39 & ~n4871 ) | ( x39 & n4873 ) | ( ~n4871 & n4873 ) ;
  assign n4875 = n4871 | n4874 ;
  assign n4876 = n4675 & ~n4866 ;
  assign n4877 = x299 & ~n4876 ;
  assign n4878 = n4697 & ~n4877 ;
  assign n4879 = x39 & ~n4878 ;
  assign n4880 = ( x38 & n4875 ) | ( x38 & ~n4879 ) | ( n4875 & ~n4879 ) ;
  assign n4881 = ~x38 & n4880 ;
  assign n4882 = x299 & ~n4868 ;
  assign n4883 = n4697 & ~n4882 ;
  assign n4884 = x38 & n4883 ;
  assign n4885 = ( x100 & ~n4881 ) | ( x100 & n4884 ) | ( ~n4881 & n4884 ) ;
  assign n4886 = n4881 | n4885 ;
  assign n4887 = n1994 & n4883 ;
  assign n4888 = n4750 & ~n4866 ;
  assign n4889 = x299 & ~n4888 ;
  assign n4890 = ( n1994 & n4697 ) | ( n1994 & ~n4889 ) | ( n4697 & ~n4889 ) ;
  assign n4891 = ~n1994 & n4890 ;
  assign n4892 = ( x100 & n4887 ) | ( x100 & ~n4891 ) | ( n4887 & ~n4891 ) ;
  assign n4893 = ~n4887 & n4892 ;
  assign n4894 = ( x87 & n4886 ) | ( x87 & ~n4893 ) | ( n4886 & ~n4893 ) ;
  assign n4895 = n4894 ^ n4886 ^ 1'b0 ;
  assign n4896 = ( x87 & n4894 ) | ( x87 & ~n4895 ) | ( n4894 & ~n4895 ) ;
  assign n4897 = n4878 ^ n2036 ^ 1'b0 ;
  assign n4898 = ( n4878 & n4883 ) | ( n4878 & n4897 ) | ( n4883 & n4897 ) ;
  assign n4899 = x87 & ~n4898 ;
  assign n4900 = ( x75 & n4896 ) | ( x75 & ~n4899 ) | ( n4896 & ~n4899 ) ;
  assign n4901 = ~x75 & n4900 ;
  assign n4902 = x75 & n4883 ;
  assign n4903 = ( x92 & ~n4901 ) | ( x92 & n4902 ) | ( ~n4901 & n4902 ) ;
  assign n4904 = n4901 | n4903 ;
  assign n4905 = ~n2044 & n4898 ;
  assign n4906 = n2044 & n4883 ;
  assign n4907 = ( x92 & n4905 ) | ( x92 & ~n4906 ) | ( n4905 & ~n4906 ) ;
  assign n4908 = ~n4905 & n4907 ;
  assign n4909 = ( n2067 & n4904 ) | ( n2067 & ~n4908 ) | ( n4904 & ~n4908 ) ;
  assign n4910 = ~n2067 & n4909 ;
  assign n4911 = n2067 & n4883 ;
  assign n4912 = ( x55 & ~n4910 ) | ( x55 & n4911 ) | ( ~n4910 & n4911 ) ;
  assign n4913 = n4910 | n4912 ;
  assign n4914 = n2099 | n4876 ;
  assign n4915 = n4914 ^ x62 ^ 1'b0 ;
  assign n4916 = n2099 & ~n4867 ;
  assign n4917 = x56 & ~n4916 ;
  assign n4918 = ( x56 & n2266 ) | ( x56 & n4917 ) | ( n2266 & n4917 ) ;
  assign n4919 = ( n4914 & ~n4915 ) | ( n4914 & n4918 ) | ( ~n4915 & n4918 ) ;
  assign n4920 = ( x62 & n4915 ) | ( x62 & n4919 ) | ( n4915 & n4919 ) ;
  assign n4921 = n2070 & n4868 ;
  assign n4922 = x55 & ~n4921 ;
  assign n4923 = ~n2070 & n4876 ;
  assign n4924 = ( x56 & n4922 ) | ( x56 & ~n4923 ) | ( n4922 & ~n4923 ) ;
  assign n4925 = n4924 ^ n4922 ^ 1'b0 ;
  assign n4926 = ( x56 & n4924 ) | ( x56 & ~n4925 ) | ( n4924 & ~n4925 ) ;
  assign n4927 = ~n4920 & n4926 ;
  assign n4928 = ( n4913 & n4920 ) | ( n4913 & ~n4927 ) | ( n4920 & ~n4927 ) ;
  assign n4929 = n2151 & n4868 ;
  assign n4930 = ~n2151 & n4876 ;
  assign n4931 = ( x62 & n4929 ) | ( x62 & ~n4930 ) | ( n4929 & ~n4930 ) ;
  assign n4932 = ~n4929 & n4931 ;
  assign n4933 = ( n2120 & n4928 ) | ( n2120 & ~n4932 ) | ( n4928 & ~n4932 ) ;
  assign n4934 = ~n2120 & n4933 ;
  assign n4935 = ( x242 & n4869 ) | ( x242 & ~n4934 ) | ( n4869 & ~n4934 ) ;
  assign n4936 = ~n4869 & n4935 ;
  assign n4937 = n2120 & n4867 ;
  assign n4938 = x242 | n4937 ;
  assign n4939 = n4801 & n4872 ;
  assign n4940 = n4693 | n4870 ;
  assign n4941 = n4804 & ~n4940 ;
  assign n4942 = ( x39 & ~n4939 ) | ( x39 & n4941 ) | ( ~n4939 & n4941 ) ;
  assign n4943 = n4939 | n4942 ;
  assign n4944 = n4784 & ~n4866 ;
  assign n4945 = ~x299 & n4695 ;
  assign n4946 = ( n4696 & n4944 ) | ( n4696 & n4945 ) | ( n4944 & n4945 ) ;
  assign n4947 = x39 & ~n4946 ;
  assign n4948 = ( x38 & n4943 ) | ( x38 & ~n4947 ) | ( n4943 & ~n4947 ) ;
  assign n4949 = ~x38 & n4948 ;
  assign n4950 = ( n4696 & n4867 ) | ( n4696 & n4945 ) | ( n4867 & n4945 ) ;
  assign n4951 = x38 & n4950 ;
  assign n4952 = ( x100 & ~n4949 ) | ( x100 & n4951 ) | ( ~n4949 & n4951 ) ;
  assign n4953 = n4949 | n4952 ;
  assign n4954 = n1994 & n4950 ;
  assign n4955 = n4815 & ~n4866 ;
  assign n4956 = x299 & ~n4955 ;
  assign n4957 = ( n1994 & n4696 ) | ( n1994 & ~n4956 ) | ( n4696 & ~n4956 ) ;
  assign n4958 = ~n1994 & n4957 ;
  assign n4959 = ( x100 & n4954 ) | ( x100 & ~n4958 ) | ( n4954 & ~n4958 ) ;
  assign n4960 = ~n4954 & n4959 ;
  assign n4961 = ( x87 & n4953 ) | ( x87 & ~n4960 ) | ( n4953 & ~n4960 ) ;
  assign n4962 = n4961 ^ n4953 ^ 1'b0 ;
  assign n4963 = ( x87 & n4961 ) | ( x87 & ~n4962 ) | ( n4961 & ~n4962 ) ;
  assign n4964 = n4946 ^ n2036 ^ 1'b0 ;
  assign n4965 = ( n4946 & n4950 ) | ( n4946 & n4964 ) | ( n4950 & n4964 ) ;
  assign n4966 = x87 & ~n4965 ;
  assign n4967 = ( x75 & n4963 ) | ( x75 & ~n4966 ) | ( n4963 & ~n4966 ) ;
  assign n4968 = ~x75 & n4967 ;
  assign n4969 = x75 & n4950 ;
  assign n4970 = ( x92 & ~n4968 ) | ( x92 & n4969 ) | ( ~n4968 & n4969 ) ;
  assign n4971 = n4968 | n4970 ;
  assign n4972 = ~n2044 & n4965 ;
  assign n4973 = n2044 & n4950 ;
  assign n4974 = ( x92 & n4972 ) | ( x92 & ~n4973 ) | ( n4972 & ~n4973 ) ;
  assign n4975 = ~n4972 & n4974 ;
  assign n4976 = ( n2067 & n4971 ) | ( n2067 & ~n4975 ) | ( n4971 & ~n4975 ) ;
  assign n4977 = ~n2067 & n4976 ;
  assign n4978 = n2067 & n4950 ;
  assign n4979 = ( x55 & ~n4977 ) | ( x55 & n4978 ) | ( ~n4977 & n4978 ) ;
  assign n4980 = n4977 | n4979 ;
  assign n4981 = n2099 | n4944 ;
  assign n4982 = n4981 ^ x62 ^ 1'b0 ;
  assign n4983 = ( n4917 & n4981 ) | ( n4917 & ~n4982 ) | ( n4981 & ~n4982 ) ;
  assign n4984 = ( x62 & n4982 ) | ( x62 & n4983 ) | ( n4982 & n4983 ) ;
  assign n4985 = n2070 & n4867 ;
  assign n4986 = x55 & ~n4985 ;
  assign n4987 = ~n2070 & n4944 ;
  assign n4988 = ( x56 & n4986 ) | ( x56 & ~n4987 ) | ( n4986 & ~n4987 ) ;
  assign n4989 = n4988 ^ n4986 ^ 1'b0 ;
  assign n4990 = ( x56 & n4988 ) | ( x56 & ~n4989 ) | ( n4988 & ~n4989 ) ;
  assign n4991 = ~n4984 & n4990 ;
  assign n4992 = ( n4980 & n4984 ) | ( n4980 & ~n4991 ) | ( n4984 & ~n4991 ) ;
  assign n4993 = n2151 & n4867 ;
  assign n4994 = ~n2151 & n4944 ;
  assign n4995 = ( x62 & n4993 ) | ( x62 & ~n4994 ) | ( n4993 & ~n4994 ) ;
  assign n4996 = ~n4993 & n4995 ;
  assign n4997 = ( n2120 & n4992 ) | ( n2120 & ~n4996 ) | ( n4992 & ~n4996 ) ;
  assign n4998 = ~n2120 & n4997 ;
  assign n4999 = ( ~n4936 & n4938 ) | ( ~n4936 & n4998 ) | ( n4938 & n4998 ) ;
  assign n5000 = ~n4936 & n4999 ;
  assign n5001 = ( x1134 & ~n4863 ) | ( x1134 & n5000 ) | ( ~n4863 & n5000 ) ;
  assign n5002 = ~n4863 & n5001 ;
  assign n5003 = n1276 | n2036 ;
  assign n5004 = n2150 | n5003 ;
  assign n5005 = x62 & n5004 ;
  assign n5006 = x59 | n5005 ;
  assign n5007 = n2098 | n5003 ;
  assign n5008 = x56 & n5007 ;
  assign n5009 = x54 | n2096 ;
  assign n5010 = n5003 | n5009 ;
  assign n5011 = x74 & n5010 ;
  assign n5012 = x55 | n5011 ;
  assign n5013 = x87 & n5003 ;
  assign n5014 = x75 | n5013 ;
  assign n5015 = x54 | x92 ;
  assign n5016 = n5014 | n5015 ;
  assign n5017 = x39 | n1292 ;
  assign n5018 = ~x38 & x100 ;
  assign n5019 = ~n5017 & n5018 ;
  assign n5020 = x950 & x1092 ;
  assign n5021 = x824 | x829 ;
  assign n5022 = n5020 & n5021 ;
  assign n5023 = ~x1093 & n5022 ;
  assign n5024 = x250 ^ x129 ^ 1'b0 ;
  assign n5025 = ( ~x129 & n5023 ) | ( ~x129 & n5024 ) | ( n5023 & n5024 ) ;
  assign n5026 = x41 | x99 ;
  assign n5027 = x101 | n5026 ;
  assign n5028 = x42 | x43 ;
  assign n5029 = x52 | n5028 ;
  assign n5030 = x113 | x116 ;
  assign n5031 = x114 | x115 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n5029 | n5032 ;
  assign n5034 = n5027 | n5033 ;
  assign n5035 = x44 | n5034 ;
  assign n5036 = ~x683 & n5035 ;
  assign n5037 = n5025 | n5036 ;
  assign n5038 = ~x299 & n1283 ;
  assign n5039 = x299 & n1329 ;
  assign n5040 = n5038 | n5039 ;
  assign n5041 = x146 & n5039 ;
  assign n5042 = x142 & n5038 ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = n5040 & ~n5043 ;
  assign n5045 = n5035 & n5044 ;
  assign n5046 = ~n5037 & n5045 ;
  assign n5047 = n2195 & ~n5044 ;
  assign n5048 = n5046 | n5047 ;
  assign n5049 = ( x87 & n5019 ) | ( x87 & ~n5048 ) | ( n5019 & ~n5048 ) ;
  assign n5050 = n5049 ^ n5019 ^ 1'b0 ;
  assign n5051 = ( x87 & n5049 ) | ( x87 & ~n5050 ) | ( n5049 & ~n5050 ) ;
  assign n5052 = x39 | n1276 ;
  assign n5053 = x38 & n5052 ;
  assign n5054 = x100 | n5053 ;
  assign n5055 = x907 | x947 ;
  assign n5056 = x975 | x978 ;
  assign n5057 = x960 | x963 ;
  assign n5058 = x970 | x972 ;
  assign n5059 = ( ~n5056 & n5057 ) | ( ~n5056 & n5058 ) | ( n5057 & n5058 ) ;
  assign n5060 = n5056 | n5059 ;
  assign n5061 = n5055 | n5060 ;
  assign n5062 = x824 & ~x1091 ;
  assign n5063 = x1093 & ~n1615 ;
  assign n5064 = ~n5062 & n5063 ;
  assign n5065 = n5021 & ~n5064 ;
  assign n5066 = x835 & x984 ;
  assign n5067 = x252 | x1001 ;
  assign n5068 = ~x979 & n5067 ;
  assign n5069 = ~n5066 & n5068 ;
  assign n5070 = ~x287 & n5069 ;
  assign n5071 = x835 & x950 ;
  assign n5072 = n5070 & n5071 ;
  assign n5073 = x1092 & n5072 ;
  assign n5074 = n5065 & n5073 ;
  assign n5075 = x332 | x468 ;
  assign n5076 = ~x662 & x680 ;
  assign n5077 = ~x661 & n5076 ;
  assign n5078 = ~x681 & n5077 ;
  assign n5079 = x603 & ~x642 ;
  assign n5080 = x614 | x616 ;
  assign n5081 = n5079 & ~n5080 ;
  assign n5082 = n5078 | n5081 ;
  assign n5083 = n5075 & ~n5082 ;
  assign n5084 = n5074 & ~n5083 ;
  assign n5085 = n1292 | n5084 ;
  assign n5086 = n5061 & ~n5085 ;
  assign n5087 = x215 & ~n5086 ;
  assign n5088 = n1276 | n5075 ;
  assign n5089 = n5082 & ~n5088 ;
  assign n5090 = ~n5074 & n5075 ;
  assign n5091 = n5082 & ~n5090 ;
  assign n5092 = ( n1292 & ~n5089 ) | ( n1292 & n5091 ) | ( ~n5089 & n5091 ) ;
  assign n5093 = ~n5089 & n5092 ;
  assign n5094 = n5061 | n5093 ;
  assign n5095 = n5087 & n5094 ;
  assign n5096 = n1670 & n5072 ;
  assign n5097 = x216 & x221 ;
  assign n5098 = n5096 & n5097 ;
  assign n5099 = n5075 & n5082 ;
  assign n5100 = ( n5061 & ~n5083 ) | ( n5061 & n5099 ) | ( ~n5083 & n5099 ) ;
  assign n5101 = n5098 & n5100 ;
  assign n5102 = ( ~x215 & n1292 ) | ( ~x215 & n5101 ) | ( n1292 & n5101 ) ;
  assign n5103 = ~x215 & n5102 ;
  assign n5104 = ( x299 & n5095 ) | ( x299 & ~n5103 ) | ( n5095 & ~n5103 ) ;
  assign n5105 = ~n5095 & n5104 ;
  assign n5106 = x222 & x224 ;
  assign n5107 = n5096 & n5106 ;
  assign n5108 = x961 | x967 ;
  assign n5109 = x969 | x971 ;
  assign n5110 = x974 | x977 ;
  assign n5111 = n5109 | n5110 ;
  assign n5112 = x587 | x602 ;
  assign n5113 = ( ~n5108 & n5111 ) | ( ~n5108 & n5112 ) | ( n5111 & n5112 ) ;
  assign n5114 = n5108 | n5113 ;
  assign n5115 = ( ~n5083 & n5099 ) | ( ~n5083 & n5114 ) | ( n5099 & n5114 ) ;
  assign n5116 = n5107 & n5115 ;
  assign n5117 = ( ~x223 & n1292 ) | ( ~x223 & n5116 ) | ( n1292 & n5116 ) ;
  assign n5118 = ~x223 & n5117 ;
  assign n5119 = ~n5085 & n5114 ;
  assign n5120 = n5093 | n5114 ;
  assign n5121 = ( x223 & n5119 ) | ( x223 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5122 = ~n5119 & n5121 ;
  assign n5123 = ( x299 & ~n5118 ) | ( x299 & n5122 ) | ( ~n5118 & n5122 ) ;
  assign n5124 = n5118 | n5123 ;
  assign n5125 = ( x39 & n5105 ) | ( x39 & n5124 ) | ( n5105 & n5124 ) ;
  assign n5126 = ~n5105 & n5125 ;
  assign n5127 = n1387 | n1456 ;
  assign n5128 = n1558 & ~n5127 ;
  assign n5129 = ( ~n1462 & n1467 ) | ( ~n1462 & n5128 ) | ( n1467 & n5128 ) ;
  assign n5130 = ~n1462 & n5129 ;
  assign n5131 = x108 | n5130 ;
  assign n5132 = ~n1704 & n5131 ;
  assign n5133 = ( x110 & n1841 ) | ( x110 & ~n5132 ) | ( n1841 & ~n5132 ) ;
  assign n5134 = n5132 | n5133 ;
  assign n5135 = n1446 | n1703 ;
  assign n5136 = ( x47 & n5134 ) | ( x47 & ~n5135 ) | ( n5134 & ~n5135 ) ;
  assign n5137 = n5136 ^ n5134 ^ 1'b0 ;
  assign n5138 = ( x47 & n5136 ) | ( x47 & ~n5137 ) | ( n5136 & ~n5137 ) ;
  assign n5139 = ( n1370 & ~n1449 ) | ( n1370 & n5138 ) | ( ~n1449 & n5138 ) ;
  assign n5140 = ~n1370 & n5139 ;
  assign n5141 = x58 & ~n1266 ;
  assign n5142 = ( x90 & ~n5140 ) | ( x90 & n5141 ) | ( ~n5140 & n5141 ) ;
  assign n5143 = n5140 | n5142 ;
  assign n5144 = n5143 ^ n1440 ^ 1'b0 ;
  assign n5145 = ( n1440 & n5143 ) | ( n1440 & n5144 ) | ( n5143 & n5144 ) ;
  assign n5146 = ( x93 & ~n1440 ) | ( x93 & n5145 ) | ( ~n1440 & n5145 ) ;
  assign n5147 = x93 & ~n1594 ;
  assign n5148 = n5147 ^ n1701 ^ x93 ;
  assign n5149 = ( x35 & n5146 ) | ( x35 & ~n5148 ) | ( n5146 & ~n5148 ) ;
  assign n5150 = n5149 ^ n5146 ^ 1'b0 ;
  assign n5151 = ( x35 & n5149 ) | ( x35 & ~n5150 ) | ( n5149 & ~n5150 ) ;
  assign n5152 = ( x70 & ~n1400 ) | ( x70 & n5151 ) | ( ~n1400 & n5151 ) ;
  assign n5153 = ~x70 & n5152 ;
  assign n5154 = x51 | n5153 ;
  assign n5155 = ~n1435 & n5154 ;
  assign n5156 = ( ~n1433 & n1773 ) | ( ~n1433 & n5155 ) | ( n1773 & n5155 ) ;
  assign n5157 = ~n1433 & n5156 ;
  assign n5158 = ( x32 & n1586 ) | ( x32 & ~n5157 ) | ( n1586 & ~n5157 ) ;
  assign n5159 = n5157 | n5158 ;
  assign n5160 = x35 | n1272 ;
  assign n5161 = x40 | n5160 ;
  assign n5162 = n1595 & ~n5161 ;
  assign n5163 = x32 & ~n5162 ;
  assign n5164 = x299 ^ x210 ^ 1'b0 ;
  assign n5165 = ( x198 & x210 ) | ( x198 & ~n5164 ) | ( x210 & ~n5164 ) ;
  assign n5166 = n5165 ^ n5163 ^ 1'b0 ;
  assign n5167 = ( n1381 & n5163 ) | ( n1381 & n5166 ) | ( n5163 & n5166 ) ;
  assign n5168 = ( x95 & n5159 ) | ( x95 & ~n5167 ) | ( n5159 & ~n5167 ) ;
  assign n5169 = ~x95 & n5168 ;
  assign n5170 = ( x39 & n1785 ) | ( x39 & ~n5169 ) | ( n1785 & ~n5169 ) ;
  assign n5171 = n5169 | n5170 ;
  assign n5172 = n5171 ^ n5126 ^ 1'b0 ;
  assign n5173 = ( n5126 & n5171 ) | ( n5126 & n5172 ) | ( n5171 & n5172 ) ;
  assign n5174 = ( x38 & ~n5126 ) | ( x38 & n5173 ) | ( ~n5126 & n5173 ) ;
  assign n5175 = n5174 ^ n5054 ^ 1'b0 ;
  assign n5176 = ( n5054 & n5174 ) | ( n5054 & n5175 ) | ( n5174 & n5175 ) ;
  assign n5177 = ( n5051 & ~n5054 ) | ( n5051 & n5176 ) | ( ~n5054 & n5176 ) ;
  assign n5178 = n5177 ^ n5016 ^ 1'b0 ;
  assign n5179 = ( n5016 & n5177 ) | ( n5016 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5180 = ( x74 & ~n5016 ) | ( x74 & n5179 ) | ( ~n5016 & n5179 ) ;
  assign n5181 = n5180 ^ n5012 ^ 1'b0 ;
  assign n5182 = ( n5012 & n5180 ) | ( n5012 & n5181 ) | ( n5180 & n5181 ) ;
  assign n5183 = ( x56 & ~n5012 ) | ( x56 & n5182 ) | ( ~n5012 & n5182 ) ;
  assign n5184 = n5183 ^ n5008 ^ 1'b0 ;
  assign n5185 = ( n5008 & n5183 ) | ( n5008 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5186 = ( x62 & ~n5008 ) | ( x62 & n5185 ) | ( ~n5008 & n5185 ) ;
  assign n5187 = ( x57 & ~n5006 ) | ( x57 & n5186 ) | ( ~n5006 & n5186 ) ;
  assign n5188 = ~x57 & n5187 ;
  assign n5189 = n1292 | n2110 ;
  assign n5190 = ( x57 & x59 ) | ( x57 & n5189 ) | ( x59 & n5189 ) ;
  assign n5191 = ( x57 & n5188 ) | ( x57 & ~n5190 ) | ( n5188 & ~n5190 ) ;
  assign n5192 = x55 | n2109 ;
  assign n5193 = x59 | n5192 ;
  assign n5194 = ~x228 & n5193 ;
  assign n5195 = x57 & ~n5194 ;
  assign n5196 = n5075 & n5078 ;
  assign n5197 = n5075 & ~n5078 ;
  assign n5198 = x468 & n5078 ;
  assign n5199 = ~x468 & x602 ;
  assign n5200 = n5198 | n5199 ;
  assign n5201 = ( n5196 & ~n5197 ) | ( n5196 & n5200 ) | ( ~n5197 & n5200 ) ;
  assign n5202 = x30 & x228 ;
  assign n5203 = x95 | n1274 ;
  assign n5204 = x35 | n5147 ;
  assign n5205 = x91 | x314 ;
  assign n5206 = n1452 | n1703 ;
  assign n5207 = x46 | n1258 ;
  assign n5208 = x102 | n1474 ;
  assign n5209 = n1227 | n5208 ;
  assign n5210 = x85 & n1511 ;
  assign n5211 = n1234 | n5210 ;
  assign n5212 = ~n1492 & n5211 ;
  assign n5213 = n1243 | n5212 ;
  assign n5214 = ( n1489 & ~n1491 ) | ( n1489 & n5213 ) | ( ~n1491 & n5213 ) ;
  assign n5215 = ~n1489 & n5214 ;
  assign n5216 = ~n1244 & n5215 ;
  assign n5217 = n1524 | n5216 ;
  assign n5218 = ~n1522 & n5217 ;
  assign n5219 = x67 & ~n1248 ;
  assign n5220 = ( n1485 & ~n5218 ) | ( n1485 & n5219 ) | ( ~n5218 & n5219 ) ;
  assign n5221 = n5218 | n5220 ;
  assign n5222 = n5221 ^ n1484 ^ 1'b0 ;
  assign n5223 = ( n1484 & n5221 ) | ( n1484 & n5222 ) | ( n5221 & n5222 ) ;
  assign n5224 = ( x71 & ~n1484 ) | ( x71 & n5223 ) | ( ~n1484 & n5223 ) ;
  assign n5225 = x64 | n1230 ;
  assign n5226 = n1537 | n5225 ;
  assign n5227 = ( x81 & n5224 ) | ( x81 & ~n5226 ) | ( n5224 & ~n5226 ) ;
  assign n5228 = n5227 ^ n5224 ^ 1'b0 ;
  assign n5229 = ( x81 & n5227 ) | ( x81 & ~n5228 ) | ( n5227 & ~n5228 ) ;
  assign n5230 = n1534 & ~n5226 ;
  assign n5231 = n5229 | n5230 ;
  assign n5232 = ~n5209 & n5231 ;
  assign n5233 = ( x50 & n1470 ) | ( x50 & ~n5232 ) | ( n1470 & ~n5232 ) ;
  assign n5234 = n5232 | n5233 ;
  assign n5235 = ( x60 & ~n1468 ) | ( x60 & n5234 ) | ( ~n1468 & n5234 ) ;
  assign n5236 = ~x60 & n5235 ;
  assign n5237 = ( x53 & n1385 ) | ( x53 & ~n5236 ) | ( n1385 & ~n5236 ) ;
  assign n5238 = n5236 | n5237 ;
  assign n5239 = n5238 ^ n1389 ^ 1'b0 ;
  assign n5240 = ( n1389 & n5238 ) | ( n1389 & n5239 ) | ( n5238 & n5239 ) ;
  assign n5241 = ( x86 & ~n1389 ) | ( x86 & n5240 ) | ( ~n1389 & n5240 ) ;
  assign n5242 = ( n1564 & ~n5207 ) | ( n1564 & n5241 ) | ( ~n5207 & n5241 ) ;
  assign n5243 = ~n1564 & n5242 ;
  assign n5244 = n1841 | n5243 ;
  assign n5245 = ~n5206 & n5244 ;
  assign n5246 = n5205 | n5245 ;
  assign n5247 = ~x91 & x314 ;
  assign n5248 = ~n5209 & n5229 ;
  assign n5249 = n1471 | n5248 ;
  assign n5250 = n5249 ^ n1469 ^ 1'b0 ;
  assign n5251 = ( n1469 & n5249 ) | ( n1469 & n5250 ) | ( n5249 & n5250 ) ;
  assign n5252 = ( n1386 & ~n1469 ) | ( n1386 & n5251 ) | ( ~n1469 & n5251 ) ;
  assign n5253 = n5252 ^ n1389 ^ 1'b0 ;
  assign n5254 = ( n1389 & n5252 ) | ( n1389 & n5253 ) | ( n5252 & n5253 ) ;
  assign n5255 = ( x86 & ~n1389 ) | ( x86 & n5254 ) | ( ~n1389 & n5254 ) ;
  assign n5256 = ( n1564 & ~n5207 ) | ( n1564 & n5255 ) | ( ~n5207 & n5255 ) ;
  assign n5257 = ~n1564 & n5256 ;
  assign n5258 = n1841 | n5257 ;
  assign n5259 = ~n5206 & n5258 ;
  assign n5260 = n5247 & ~n5259 ;
  assign n5261 = x91 & n1409 ;
  assign n5262 = ( x58 & ~n5260 ) | ( x58 & n5261 ) | ( ~n5260 & n5261 ) ;
  assign n5263 = n5260 | n5262 ;
  assign n5264 = ( x90 & n5246 ) | ( x90 & ~n5263 ) | ( n5246 & ~n5263 ) ;
  assign n5265 = n5264 ^ n5246 ^ 1'b0 ;
  assign n5266 = ( x90 & n5264 ) | ( x90 & ~n5265 ) | ( n5264 & ~n5265 ) ;
  assign n5267 = n5266 ^ n1440 ^ 1'b0 ;
  assign n5268 = ( n1440 & n5266 ) | ( n1440 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = ( x93 & ~n1440 ) | ( x93 & n5268 ) | ( ~n1440 & n5268 ) ;
  assign n5270 = n5269 ^ n5204 ^ 1'b0 ;
  assign n5271 = ( n5204 & n5269 ) | ( n5204 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5272 = ( x70 & ~n5204 ) | ( x70 & n5271 ) | ( ~n5204 & n5271 ) ;
  assign n5273 = n5272 ^ n1694 ^ 1'b0 ;
  assign n5274 = ( n1694 & n5272 ) | ( n1694 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5275 = ( x72 & ~n1694 ) | ( x72 & n5274 ) | ( ~n1694 & n5274 ) ;
  assign n5276 = ( n1432 & ~n5203 ) | ( n1432 & n5275 ) | ( ~n5203 & n5275 ) ;
  assign n5277 = ~n1432 & n5276 ;
  assign n5278 = ( n1224 & ~n1275 ) | ( n1224 & n5277 ) | ( ~n1275 & n5277 ) ;
  assign n5279 = n5277 ^ n1275 ^ 1'b0 ;
  assign n5280 = ( n5277 & n5278 ) | ( n5277 & ~n5279 ) | ( n5278 & ~n5279 ) ;
  assign n5281 = x841 | n1399 ;
  assign n5282 = n1411 | n5281 ;
  assign n5283 = n1652 | n5282 ;
  assign n5284 = x32 & ~n5283 ;
  assign n5285 = ~x95 & n5284 ;
  assign n5286 = ~x198 & n5285 ;
  assign n5287 = n5280 | n5286 ;
  assign n5288 = ~x30 & x228 ;
  assign n5289 = ( n5202 & n5287 ) | ( n5202 & ~n5288 ) | ( n5287 & ~n5288 ) ;
  assign n5290 = n5201 & n5289 ;
  assign n5291 = x299 | n5290 ;
  assign n5292 = ( x907 & n5196 ) | ( x907 & ~n5197 ) | ( n5196 & ~n5197 ) ;
  assign n5293 = n5202 & n5292 ;
  assign n5294 = x299 & ~n5293 ;
  assign n5295 = ~x210 & n5285 ;
  assign n5296 = n5280 | n5295 ;
  assign n5297 = n5292 & n5296 ;
  assign n5298 = ~x228 & n5297 ;
  assign n5299 = n5294 & ~n5298 ;
  assign n5300 = ( x232 & n5291 ) | ( x232 & ~n5299 ) | ( n5291 & ~n5299 ) ;
  assign n5301 = ~x232 & n5300 ;
  assign n5302 = x160 & x197 ;
  assign n5303 = x158 & x159 ;
  assign n5304 = n5302 & n5303 ;
  assign n5305 = n5297 | n5304 ;
  assign n5306 = x47 | n1257 ;
  assign n5307 = n1840 | n5243 ;
  assign n5308 = ~n5306 & n5307 ;
  assign n5309 = n5205 | n5308 ;
  assign n5310 = n1840 | n5257 ;
  assign n5311 = ~n5306 & n5310 ;
  assign n5312 = n5247 & ~n5311 ;
  assign n5313 = ( x58 & n5261 ) | ( x58 & ~n5312 ) | ( n5261 & ~n5312 ) ;
  assign n5314 = n5312 | n5313 ;
  assign n5315 = ( x90 & n5309 ) | ( x90 & ~n5314 ) | ( n5309 & ~n5314 ) ;
  assign n5316 = n5315 ^ n5309 ^ 1'b0 ;
  assign n5317 = ( x90 & n5315 ) | ( x90 & ~n5316 ) | ( n5315 & ~n5316 ) ;
  assign n5318 = n5317 ^ n1440 ^ 1'b0 ;
  assign n5319 = ( n1440 & n5317 ) | ( n1440 & n5318 ) | ( n5317 & n5318 ) ;
  assign n5320 = ( x93 & ~n1440 ) | ( x93 & n5319 ) | ( ~n1440 & n5319 ) ;
  assign n5321 = n5320 ^ n5204 ^ 1'b0 ;
  assign n5322 = ( n5204 & n5320 ) | ( n5204 & n5321 ) | ( n5320 & n5321 ) ;
  assign n5323 = ( x70 & ~n5204 ) | ( x70 & n5322 ) | ( ~n5204 & n5322 ) ;
  assign n5324 = n5323 ^ n1694 ^ 1'b0 ;
  assign n5325 = ( n1694 & n5323 ) | ( n1694 & n5324 ) | ( n5323 & n5324 ) ;
  assign n5326 = ( x72 & ~n1694 ) | ( x72 & n5325 ) | ( ~n1694 & n5325 ) ;
  assign n5327 = ( n1432 & ~n5203 ) | ( n1432 & n5326 ) | ( ~n5203 & n5326 ) ;
  assign n5328 = ~n1432 & n5327 ;
  assign n5329 = ( n1224 & ~n1275 ) | ( n1224 & n5328 ) | ( ~n1275 & n5328 ) ;
  assign n5330 = n5328 ^ n1275 ^ 1'b0 ;
  assign n5331 = ( n5328 & n5329 ) | ( n5328 & ~n5330 ) | ( n5329 & ~n5330 ) ;
  assign n5332 = n5295 | n5331 ;
  assign n5333 = ~n5075 & n5332 ;
  assign n5334 = n5075 & n5296 ;
  assign n5335 = n5333 | n5334 ;
  assign n5336 = n5292 & n5335 ;
  assign n5337 = n5304 & ~n5336 ;
  assign n5338 = ( x228 & n5305 ) | ( x228 & ~n5337 ) | ( n5305 & ~n5337 ) ;
  assign n5339 = ~x228 & n5338 ;
  assign n5340 = ( x299 & n5293 ) | ( x299 & ~n5339 ) | ( n5293 & ~n5339 ) ;
  assign n5341 = ~n5293 & n5340 ;
  assign n5342 = x145 & x180 ;
  assign n5343 = x181 & x182 ;
  assign n5344 = n5342 & n5343 ;
  assign n5345 = n5286 | n5331 ;
  assign n5346 = ~n5075 & n5345 ;
  assign n5347 = n5075 & n5287 ;
  assign n5348 = n5346 | n5347 ;
  assign n5349 = ~x228 & n5201 ;
  assign n5350 = n5348 & n5349 ;
  assign n5351 = n5201 & n5202 ;
  assign n5352 = ( n5344 & n5350 ) | ( n5344 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5353 = n5351 ^ n5350 ^ 1'b0 ;
  assign n5354 = ( n5344 & n5352 ) | ( n5344 & n5353 ) | ( n5352 & n5353 ) ;
  assign n5355 = ~x299 & n5344 ;
  assign n5356 = ~n5354 & n5355 ;
  assign n5357 = ( n5291 & n5354 ) | ( n5291 & ~n5356 ) | ( n5354 & ~n5356 ) ;
  assign n5358 = ( x232 & n5341 ) | ( x232 & n5357 ) | ( n5341 & n5357 ) ;
  assign n5359 = ~n5341 & n5358 ;
  assign n5360 = ( ~x39 & n5301 ) | ( ~x39 & n5359 ) | ( n5301 & n5359 ) ;
  assign n5361 = ~x39 & n5360 ;
  assign n5362 = x287 | n1292 ;
  assign n5363 = x835 & n5069 ;
  assign n5364 = ~n5362 & n5363 ;
  assign n5365 = x824 & x1093 ;
  assign n5366 = n5020 & n5365 ;
  assign n5367 = x1091 & n1614 ;
  assign n5368 = n5366 & ~n5367 ;
  assign n5369 = n1670 | n5368 ;
  assign n5370 = x1091 & n5369 ;
  assign n5371 = n5364 & n5370 ;
  assign n5372 = n5364 & n5366 ;
  assign n5373 = ~x1091 & n5372 ;
  assign n5374 = n5371 | n5373 ;
  assign n5375 = x224 & ~n5374 ;
  assign n5376 = x222 & ~x223 ;
  assign n5377 = x829 | n1614 ;
  assign n5378 = x1091 & n5377 ;
  assign n5379 = n5372 & ~n5378 ;
  assign n5380 = x224 | n5379 ;
  assign n5381 = ( n5375 & n5376 ) | ( n5375 & n5380 ) | ( n5376 & n5380 ) ;
  assign n5382 = ~n5375 & n5381 ;
  assign n5383 = ~x228 & n5382 ;
  assign n5384 = n5202 | n5383 ;
  assign n5385 = n5201 & n5384 ;
  assign n5386 = x299 | n5385 ;
  assign n5387 = n5374 ^ x216 ^ 1'b0 ;
  assign n5388 = ( n5374 & n5379 ) | ( n5374 & ~n5387 ) | ( n5379 & ~n5387 ) ;
  assign n5389 = x228 | n5388 ;
  assign n5390 = ~x215 & x221 ;
  assign n5391 = ~n5288 & n5390 ;
  assign n5392 = n5389 & n5391 ;
  assign n5393 = n5202 | n5392 ;
  assign n5394 = x299 & ~n5393 ;
  assign n5395 = ( x299 & ~n5292 ) | ( x299 & n5394 ) | ( ~n5292 & n5394 ) ;
  assign n5396 = x39 & ~n5395 ;
  assign n5397 = n5386 & n5396 ;
  assign n5398 = ( x38 & ~n5361 ) | ( x38 & n5397 ) | ( ~n5361 & n5397 ) ;
  assign n5399 = n5361 | n5398 ;
  assign n5400 = n5292 ^ x299 ^ 1'b0 ;
  assign n5401 = ( n5201 & n5292 ) | ( n5201 & ~n5400 ) | ( n5292 & ~n5400 ) ;
  assign n5402 = n2613 | n5288 ;
  assign n5403 = x39 | n5402 ;
  assign n5404 = n5401 & ~n5403 ;
  assign n5405 = n5202 & n5401 ;
  assign n5406 = x38 & ~n5405 ;
  assign n5407 = ~n5404 & n5406 ;
  assign n5408 = ( x100 & n5399 ) | ( x100 & ~n5407 ) | ( n5399 & ~n5407 ) ;
  assign n5409 = n5408 ^ n5399 ^ 1'b0 ;
  assign n5410 = ( x100 & n5408 ) | ( x100 & ~n5409 ) | ( n5408 & ~n5409 ) ;
  assign n5411 = n1994 & n5405 ;
  assign n5412 = ~x142 & n1283 ;
  assign n5413 = x252 & ~n5412 ;
  assign n5414 = x252 & ~n5088 ;
  assign n5415 = x252 & ~n1292 ;
  assign n5416 = n5414 ^ n5078 ^ 1'b0 ;
  assign n5417 = ( n5414 & n5415 ) | ( n5414 & n5416 ) | ( n5415 & n5416 ) ;
  assign n5418 = n5413 & n5417 ;
  assign n5419 = n1292 | n5025 ;
  assign n5420 = x683 & n5035 ;
  assign n5421 = ~n5419 & n5420 ;
  assign n5422 = ~n5197 & n5421 ;
  assign n5423 = n5412 & n5422 ;
  assign n5424 = n5418 | n5423 ;
  assign n5425 = x602 | n5075 ;
  assign n5426 = ( x228 & n5424 ) | ( x228 & n5425 ) | ( n5424 & n5425 ) ;
  assign n5427 = ~x228 & n5426 ;
  assign n5428 = ( x299 & n5351 ) | ( x299 & ~n5427 ) | ( n5351 & ~n5427 ) ;
  assign n5429 = n5427 | n5428 ;
  assign n5430 = n1330 & ~n5422 ;
  assign n5431 = x907 | n5075 ;
  assign n5432 = ( x228 & ~n5430 ) | ( x228 & n5431 ) | ( ~n5430 & n5431 ) ;
  assign n5433 = ~x228 & n5432 ;
  assign n5434 = n1330 | n5417 ;
  assign n5435 = n5294 & ~n5434 ;
  assign n5436 = ( n5294 & ~n5433 ) | ( n5294 & n5435 ) | ( ~n5433 & n5435 ) ;
  assign n5437 = ( n1994 & n5429 ) | ( n1994 & ~n5436 ) | ( n5429 & ~n5436 ) ;
  assign n5438 = ~n1994 & n5437 ;
  assign n5439 = ( x100 & n5411 ) | ( x100 & ~n5438 ) | ( n5411 & ~n5438 ) ;
  assign n5440 = ~n5411 & n5439 ;
  assign n5441 = ( x87 & n5410 ) | ( x87 & ~n5440 ) | ( n5410 & ~n5440 ) ;
  assign n5442 = ~x87 & n5441 ;
  assign n5443 = x87 & n5405 ;
  assign n5444 = ( x75 & ~n5442 ) | ( x75 & n5443 ) | ( ~n5442 & n5443 ) ;
  assign n5445 = n5442 | n5444 ;
  assign n5446 = x75 & ~n5405 ;
  assign n5447 = x92 & ~n5446 ;
  assign n5448 = n5447 ^ x54 ^ 1'b0 ;
  assign n5449 = n1207 & n5405 ;
  assign n5450 = ~n2052 & n5404 ;
  assign n5451 = n5449 | n5450 ;
  assign n5452 = x75 | n5451 ;
  assign n5453 = ( n5447 & ~n5448 ) | ( n5447 & n5452 ) | ( ~n5448 & n5452 ) ;
  assign n5454 = ( x54 & n5448 ) | ( x54 & n5453 ) | ( n5448 & n5453 ) ;
  assign n5455 = x75 & ~n5451 ;
  assign n5456 = x92 | n5455 ;
  assign n5457 = ~n5454 & n5456 ;
  assign n5458 = ( n5445 & n5454 ) | ( n5445 & ~n5457 ) | ( n5454 & ~n5457 ) ;
  assign n5459 = x54 | n2053 ;
  assign n5460 = ~n5405 & n5459 ;
  assign n5461 = x74 & ~n5460 ;
  assign n5462 = n5461 ^ x55 ^ 1'b0 ;
  assign n5463 = n2053 | n5451 ;
  assign n5464 = x54 | n5463 ;
  assign n5465 = ( n5461 & ~n5462 ) | ( n5461 & n5464 ) | ( ~n5462 & n5464 ) ;
  assign n5466 = ( x55 & n5462 ) | ( x55 & n5465 ) | ( n5462 & n5465 ) ;
  assign n5467 = n2053 & ~n5405 ;
  assign n5468 = x54 & ~n5463 ;
  assign n5469 = ( x54 & n5467 ) | ( x54 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5470 = x74 | n5469 ;
  assign n5471 = ~n5466 & n5470 ;
  assign n5472 = ( n5458 & n5466 ) | ( n5458 & ~n5471 ) | ( n5466 & ~n5471 ) ;
  assign n5473 = ~x228 & n2070 ;
  assign n5474 = n5402 | n5473 ;
  assign n5475 = n5292 & ~n5474 ;
  assign n5476 = x55 & ~n5475 ;
  assign n5477 = ( n2109 & n5472 ) | ( n2109 & ~n5476 ) | ( n5472 & ~n5476 ) ;
  assign n5478 = ~n2109 & n5477 ;
  assign n5479 = n2109 & n5293 ;
  assign n5480 = ( x59 & ~n5478 ) | ( x59 & n5479 ) | ( ~n5478 & n5479 ) ;
  assign n5481 = n5478 | n5480 ;
  assign n5482 = ~x228 & n5192 ;
  assign n5483 = n5475 & ~n5482 ;
  assign n5484 = x59 & ~n5483 ;
  assign n5485 = ( x57 & n5481 ) | ( x57 & ~n5484 ) | ( n5481 & ~n5484 ) ;
  assign n5486 = ~x57 & n5485 ;
  assign n5487 = n5486 ^ n5195 ^ 1'b0 ;
  assign n5488 = ( ~n5195 & n5475 ) | ( ~n5195 & n5487 ) | ( n5475 & n5487 ) ;
  assign n5489 = ( n5195 & n5486 ) | ( n5195 & n5488 ) | ( n5486 & n5488 ) ;
  assign n5490 = n5075 & ~n5081 ;
  assign n5491 = n5075 & n5081 ;
  assign n5492 = x587 | n5491 ;
  assign n5493 = ( ~n5490 & n5491 ) | ( ~n5490 & n5492 ) | ( n5491 & n5492 ) ;
  assign n5494 = n5289 & n5493 ;
  assign n5495 = x299 | n5494 ;
  assign n5496 = x947 | n5491 ;
  assign n5497 = ( ~n5490 & n5491 ) | ( ~n5490 & n5496 ) | ( n5491 & n5496 ) ;
  assign n5498 = n5202 & n5497 ;
  assign n5499 = x299 & ~n5498 ;
  assign n5500 = n5296 & n5497 ;
  assign n5501 = ~x228 & n5500 ;
  assign n5502 = n5499 & ~n5501 ;
  assign n5503 = ( x232 & n5495 ) | ( x232 & ~n5502 ) | ( n5495 & ~n5502 ) ;
  assign n5504 = ~x232 & n5503 ;
  assign n5505 = n5304 | n5500 ;
  assign n5506 = n5335 & n5497 ;
  assign n5507 = n5304 & ~n5506 ;
  assign n5508 = ( x228 & n5505 ) | ( x228 & ~n5507 ) | ( n5505 & ~n5507 ) ;
  assign n5509 = ~x228 & n5508 ;
  assign n5510 = ( x299 & n5498 ) | ( x299 & ~n5509 ) | ( n5498 & ~n5509 ) ;
  assign n5511 = ~n5498 & n5510 ;
  assign n5512 = ~x228 & n5493 ;
  assign n5513 = n5348 & n5512 ;
  assign n5514 = n5202 & n5493 ;
  assign n5515 = ( n5344 & n5513 ) | ( n5344 & n5514 ) | ( n5513 & n5514 ) ;
  assign n5516 = n5514 ^ n5513 ^ 1'b0 ;
  assign n5517 = ( n5344 & n5515 ) | ( n5344 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5518 = ~n5344 & n5494 ;
  assign n5519 = ( x299 & ~n5517 ) | ( x299 & n5518 ) | ( ~n5517 & n5518 ) ;
  assign n5520 = n5517 | n5519 ;
  assign n5521 = ( x232 & n5511 ) | ( x232 & n5520 ) | ( n5511 & n5520 ) ;
  assign n5522 = ~n5511 & n5521 ;
  assign n5523 = ( ~x39 & n5504 ) | ( ~x39 & n5522 ) | ( n5504 & n5522 ) ;
  assign n5524 = ~x39 & n5523 ;
  assign n5525 = x299 & n5390 ;
  assign n5526 = n5499 | n5525 ;
  assign n5527 = n5392 & n5497 ;
  assign n5528 = n5526 & ~n5527 ;
  assign n5529 = x39 & ~n5528 ;
  assign n5530 = x299 | n5493 ;
  assign n5531 = ( x299 & n5384 ) | ( x299 & n5530 ) | ( n5384 & n5530 ) ;
  assign n5532 = n5529 & n5531 ;
  assign n5533 = ( x38 & ~n5524 ) | ( x38 & n5532 ) | ( ~n5524 & n5532 ) ;
  assign n5534 = n5524 | n5533 ;
  assign n5535 = x587 ^ x299 ^ 1'b0 ;
  assign n5536 = ( x587 & x947 ) | ( x587 & n5535 ) | ( x947 & n5535 ) ;
  assign n5537 = n5081 ^ x468 ^ 1'b0 ;
  assign n5538 = ( n5081 & n5536 ) | ( n5081 & ~n5537 ) | ( n5536 & ~n5537 ) ;
  assign n5539 = ( n5493 & n5497 ) | ( n5493 & n5538 ) | ( n5497 & n5538 ) ;
  assign n5540 = ~n5403 & n5539 ;
  assign n5541 = n5202 & n5539 ;
  assign n5542 = x38 & ~n5541 ;
  assign n5543 = ~n5540 & n5542 ;
  assign n5544 = ( x100 & n5534 ) | ( x100 & ~n5543 ) | ( n5534 & ~n5543 ) ;
  assign n5545 = n5544 ^ n5534 ^ 1'b0 ;
  assign n5546 = ( x100 & n5544 ) | ( x100 & ~n5545 ) | ( n5544 & ~n5545 ) ;
  assign n5547 = n5414 ^ n5081 ^ 1'b0 ;
  assign n5548 = ( n5414 & n5415 ) | ( n5414 & n5547 ) | ( n5415 & n5547 ) ;
  assign n5549 = ( n1330 & n5496 ) | ( n1330 & n5548 ) | ( n5496 & n5548 ) ;
  assign n5550 = ~n1330 & n5549 ;
  assign n5551 = n5421 & ~n5490 ;
  assign n5552 = x947 | n5075 ;
  assign n5553 = ( ~n1330 & n5551 ) | ( ~n1330 & n5552 ) | ( n5551 & n5552 ) ;
  assign n5554 = n1330 & n5553 ;
  assign n5555 = ( ~x228 & n5550 ) | ( ~x228 & n5554 ) | ( n5550 & n5554 ) ;
  assign n5556 = ~x228 & n5555 ;
  assign n5557 = ( n1994 & n5499 ) | ( n1994 & ~n5556 ) | ( n5499 & ~n5556 ) ;
  assign n5558 = n5557 ^ n5499 ^ 1'b0 ;
  assign n5559 = ( n1994 & n5557 ) | ( n1994 & ~n5558 ) | ( n5557 & ~n5558 ) ;
  assign n5560 = x228 | n1283 ;
  assign n5561 = x142 | n5551 ;
  assign n5562 = ( x228 & n5492 ) | ( x228 & n5561 ) | ( n5492 & n5561 ) ;
  assign n5563 = ~x228 & n5562 ;
  assign n5564 = n5563 ^ n5548 ^ 1'b0 ;
  assign n5565 = ( ~x142 & n5548 ) | ( ~x142 & n5564 ) | ( n5548 & n5564 ) ;
  assign n5566 = ( n5563 & ~n5564 ) | ( n5563 & n5565 ) | ( ~n5564 & n5565 ) ;
  assign n5567 = ( n5514 & n5560 ) | ( n5514 & ~n5566 ) | ( n5560 & ~n5566 ) ;
  assign n5568 = ~n5514 & n5567 ;
  assign n5569 = x587 | n5075 ;
  assign n5570 = n5548 & n5569 ;
  assign n5571 = ( n5560 & ~n5568 ) | ( n5560 & n5570 ) | ( ~n5568 & n5570 ) ;
  assign n5572 = ~n5568 & n5571 ;
  assign n5573 = ( x299 & ~n5559 ) | ( x299 & n5572 ) | ( ~n5559 & n5572 ) ;
  assign n5574 = ~n5559 & n5573 ;
  assign n5575 = n1994 & n5541 ;
  assign n5576 = ( x100 & n5574 ) | ( x100 & ~n5575 ) | ( n5574 & ~n5575 ) ;
  assign n5577 = ~n5574 & n5576 ;
  assign n5578 = ( x87 & n5546 ) | ( x87 & ~n5577 ) | ( n5546 & ~n5577 ) ;
  assign n5579 = ~x87 & n5578 ;
  assign n5580 = x87 & n5541 ;
  assign n5581 = ( x75 & ~n5579 ) | ( x75 & n5580 ) | ( ~n5579 & n5580 ) ;
  assign n5582 = n5579 | n5581 ;
  assign n5583 = x75 & ~n5541 ;
  assign n5584 = x92 & ~n5583 ;
  assign n5585 = n5584 ^ x54 ^ 1'b0 ;
  assign n5586 = n1207 & n5541 ;
  assign n5587 = ~n2052 & n5540 ;
  assign n5588 = n5586 | n5587 ;
  assign n5589 = x75 | n5588 ;
  assign n5590 = ( n5584 & ~n5585 ) | ( n5584 & n5589 ) | ( ~n5585 & n5589 ) ;
  assign n5591 = ( x54 & n5585 ) | ( x54 & n5590 ) | ( n5585 & n5590 ) ;
  assign n5592 = x75 & ~n5588 ;
  assign n5593 = x92 | n5592 ;
  assign n5594 = ~n5591 & n5593 ;
  assign n5595 = ( n5582 & n5591 ) | ( n5582 & ~n5594 ) | ( n5591 & ~n5594 ) ;
  assign n5596 = n5459 & ~n5541 ;
  assign n5597 = x74 & ~n5596 ;
  assign n5598 = n5597 ^ x55 ^ 1'b0 ;
  assign n5599 = n2053 | n5588 ;
  assign n5600 = x54 | n5599 ;
  assign n5601 = ( n5597 & ~n5598 ) | ( n5597 & n5600 ) | ( ~n5598 & n5600 ) ;
  assign n5602 = ( x55 & n5598 ) | ( x55 & n5601 ) | ( n5598 & n5601 ) ;
  assign n5603 = n2053 & ~n5541 ;
  assign n5604 = x54 & ~n5599 ;
  assign n5605 = ( x54 & n5603 ) | ( x54 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5606 = x74 | n5605 ;
  assign n5607 = ~n5602 & n5606 ;
  assign n5608 = ( n5595 & n5602 ) | ( n5595 & ~n5607 ) | ( n5602 & ~n5607 ) ;
  assign n5609 = ~n5474 & n5497 ;
  assign n5610 = x55 & ~n5609 ;
  assign n5611 = ( n2109 & n5608 ) | ( n2109 & ~n5610 ) | ( n5608 & ~n5610 ) ;
  assign n5612 = ~n2109 & n5611 ;
  assign n5613 = n2109 & n5498 ;
  assign n5614 = ( x59 & ~n5612 ) | ( x59 & n5613 ) | ( ~n5612 & n5613 ) ;
  assign n5615 = n5612 | n5614 ;
  assign n5616 = ~n5482 & n5609 ;
  assign n5617 = x59 & ~n5616 ;
  assign n5618 = ( x57 & n5615 ) | ( x57 & ~n5617 ) | ( n5615 & ~n5617 ) ;
  assign n5619 = ~x57 & n5618 ;
  assign n5620 = n5619 ^ n5195 ^ 1'b0 ;
  assign n5621 = ( ~n5195 & n5609 ) | ( ~n5195 & n5620 ) | ( n5609 & n5620 ) ;
  assign n5622 = ( n5195 & n5619 ) | ( n5195 & n5621 ) | ( n5619 & n5621 ) ;
  assign n5623 = x30 & ~n5075 ;
  assign n5624 = x228 & n5623 ;
  assign n5625 = x970 & n5624 ;
  assign n5626 = x299 & ~n5625 ;
  assign n5627 = ~x228 & x970 ;
  assign n5628 = ~n5075 & n5296 ;
  assign n5629 = n5627 & n5628 ;
  assign n5630 = n5626 & ~n5629 ;
  assign n5631 = ~n5075 & n5289 ;
  assign n5632 = x967 & n5631 ;
  assign n5633 = x299 | n5632 ;
  assign n5634 = ( x232 & ~n5630 ) | ( x232 & n5633 ) | ( ~n5630 & n5633 ) ;
  assign n5635 = ~x232 & n5634 ;
  assign n5636 = n5344 | n5631 ;
  assign n5637 = ~x228 & n5346 ;
  assign n5638 = n5287 & ~n5344 ;
  assign n5639 = n5624 | n5638 ;
  assign n5640 = ( n5636 & n5637 ) | ( n5636 & n5639 ) | ( n5637 & n5639 ) ;
  assign n5641 = n5639 ^ n5637 ^ 1'b0 ;
  assign n5642 = ( n5636 & n5640 ) | ( n5636 & n5641 ) | ( n5640 & n5641 ) ;
  assign n5643 = x967 & n5642 ;
  assign n5644 = x299 | n5643 ;
  assign n5645 = n5333 ^ n5302 ^ 1'b0 ;
  assign n5646 = ( n5296 & n5333 ) | ( n5296 & ~n5645 ) | ( n5333 & ~n5645 ) ;
  assign n5647 = ~n5075 & n5646 ;
  assign n5648 = n5627 & n5647 ;
  assign n5649 = n5625 | n5648 ;
  assign n5650 = n5303 & n5649 ;
  assign n5651 = x299 & n5303 ;
  assign n5652 = ( n5630 & ~n5650 ) | ( n5630 & n5651 ) | ( ~n5650 & n5651 ) ;
  assign n5653 = ~n5650 & n5652 ;
  assign n5654 = x232 & ~n5653 ;
  assign n5655 = n5644 & n5654 ;
  assign n5656 = ( ~x39 & n5635 ) | ( ~x39 & n5655 ) | ( n5635 & n5655 ) ;
  assign n5657 = ~x39 & n5656 ;
  assign n5658 = x228 & ~n5623 ;
  assign n5659 = ~x299 & x967 ;
  assign n5660 = ~n5075 & n5382 ;
  assign n5661 = x228 | n5660 ;
  assign n5662 = n5659 & n5661 ;
  assign n5663 = x299 & x970 ;
  assign n5664 = n5388 & n5390 ;
  assign n5665 = ~n5075 & n5664 ;
  assign n5666 = x228 | n5665 ;
  assign n5667 = n5663 & n5666 ;
  assign n5668 = n5662 | n5667 ;
  assign n5669 = ( x39 & n5658 ) | ( x39 & n5668 ) | ( n5658 & n5668 ) ;
  assign n5670 = ~n5658 & n5669 ;
  assign n5671 = ( x38 & ~n5657 ) | ( x38 & n5670 ) | ( ~n5657 & n5670 ) ;
  assign n5672 = n5657 | n5671 ;
  assign n5673 = ( n5088 & ~n5624 ) | ( n5088 & n5658 ) | ( ~n5624 & n5658 ) ;
  assign n5674 = x967 & ~n5673 ;
  assign n5675 = x299 | n5674 ;
  assign n5676 = ~n5088 & n5627 ;
  assign n5677 = n5626 & ~n5676 ;
  assign n5678 = ( x39 & n5675 ) | ( x39 & ~n5677 ) | ( n5675 & ~n5677 ) ;
  assign n5679 = ~x39 & n5678 ;
  assign n5680 = ( n5624 & n5659 ) | ( n5624 & n5663 ) | ( n5659 & n5663 ) ;
  assign n5681 = x39 & n5680 ;
  assign n5682 = x38 & ~n5681 ;
  assign n5683 = ~n5679 & n5682 ;
  assign n5684 = ( x100 & n5672 ) | ( x100 & ~n5683 ) | ( n5672 & ~n5683 ) ;
  assign n5685 = n5684 ^ n5672 ^ 1'b0 ;
  assign n5686 = ( x100 & n5684 ) | ( x100 & ~n5685 ) | ( n5684 & ~n5685 ) ;
  assign n5687 = n1994 & n5680 ;
  assign n5688 = ~n5075 & n5421 ;
  assign n5689 = n5412 & n5688 ;
  assign n5690 = ~n5412 & n5414 ;
  assign n5691 = x228 | n5690 ;
  assign n5692 = ( ~n5658 & n5689 ) | ( ~n5658 & n5691 ) | ( n5689 & n5691 ) ;
  assign n5693 = ~n5658 & n5692 ;
  assign n5694 = x967 & n5693 ;
  assign n5695 = x299 | n5694 ;
  assign n5696 = n1330 | n5414 ;
  assign n5697 = n1330 & ~n5688 ;
  assign n5698 = ( x228 & n5696 ) | ( x228 & ~n5697 ) | ( n5696 & ~n5697 ) ;
  assign n5699 = ~x228 & n5698 ;
  assign n5700 = x970 & n5699 ;
  assign n5701 = n5626 & ~n5700 ;
  assign n5702 = ( n1994 & n5695 ) | ( n1994 & ~n5701 ) | ( n5695 & ~n5701 ) ;
  assign n5703 = ~n1994 & n5702 ;
  assign n5704 = ( x100 & n5687 ) | ( x100 & ~n5703 ) | ( n5687 & ~n5703 ) ;
  assign n5705 = ~n5687 & n5704 ;
  assign n5706 = ( x87 & n5686 ) | ( x87 & ~n5705 ) | ( n5686 & ~n5705 ) ;
  assign n5707 = ~x87 & n5706 ;
  assign n5708 = x87 & n5680 ;
  assign n5709 = ( x75 & ~n5707 ) | ( x75 & n5708 ) | ( ~n5707 & n5708 ) ;
  assign n5710 = n5707 | n5709 ;
  assign n5711 = x75 & ~n5680 ;
  assign n5712 = x92 & ~n5711 ;
  assign n5713 = n5712 ^ x54 ^ 1'b0 ;
  assign n5714 = n1207 & n5680 ;
  assign n5715 = ~n2052 & n5679 ;
  assign n5716 = n5714 | n5715 ;
  assign n5717 = x75 | n5716 ;
  assign n5718 = ( n5712 & ~n5713 ) | ( n5712 & n5717 ) | ( ~n5713 & n5717 ) ;
  assign n5719 = ( x54 & n5713 ) | ( x54 & n5718 ) | ( n5713 & n5718 ) ;
  assign n5720 = x75 & ~n5716 ;
  assign n5721 = x92 | n5720 ;
  assign n5722 = ~n5719 & n5721 ;
  assign n5723 = ( n5710 & n5719 ) | ( n5710 & ~n5722 ) | ( n5719 & ~n5722 ) ;
  assign n5724 = n5459 & ~n5680 ;
  assign n5725 = x74 & ~n5724 ;
  assign n5726 = n5725 ^ x55 ^ 1'b0 ;
  assign n5727 = n2053 | n5716 ;
  assign n5728 = x54 | n5727 ;
  assign n5729 = ( n5725 & ~n5726 ) | ( n5725 & n5728 ) | ( ~n5726 & n5728 ) ;
  assign n5730 = ( x55 & n5726 ) | ( x55 & n5729 ) | ( n5726 & n5729 ) ;
  assign n5731 = n2053 & ~n5680 ;
  assign n5732 = x54 & ~n5727 ;
  assign n5733 = ( x54 & n5731 ) | ( x54 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5734 = x74 | n5733 ;
  assign n5735 = ~n5730 & n5734 ;
  assign n5736 = ( n5723 & n5730 ) | ( n5723 & ~n5735 ) | ( n5730 & ~n5735 ) ;
  assign n5737 = ~n2070 & n5676 ;
  assign n5738 = x55 & ~n5625 ;
  assign n5739 = ~n5737 & n5738 ;
  assign n5740 = ( n2109 & n5736 ) | ( n2109 & ~n5739 ) | ( n5736 & ~n5739 ) ;
  assign n5741 = ~n2109 & n5740 ;
  assign n5742 = n2109 & n5625 ;
  assign n5743 = ( x59 & ~n5741 ) | ( x59 & n5742 ) | ( ~n5741 & n5742 ) ;
  assign n5744 = n5741 | n5743 ;
  assign n5745 = x59 & ~n5625 ;
  assign n5746 = ~n5192 & n5737 ;
  assign n5747 = n5745 & ~n5746 ;
  assign n5748 = ( x57 & n5744 ) | ( x57 & ~n5747 ) | ( n5744 & ~n5747 ) ;
  assign n5749 = ~x57 & n5748 ;
  assign n5750 = ~n5193 & n5737 ;
  assign n5751 = n5625 | n5750 ;
  assign n5752 = n5749 ^ x57 ^ 1'b0 ;
  assign n5753 = ( ~x57 & n5751 ) | ( ~x57 & n5752 ) | ( n5751 & n5752 ) ;
  assign n5754 = ( x57 & n5749 ) | ( x57 & n5753 ) | ( n5749 & n5753 ) ;
  assign n5755 = x972 & n5624 ;
  assign n5756 = x299 & ~n5755 ;
  assign n5757 = ~x228 & x972 ;
  assign n5758 = n5628 & n5757 ;
  assign n5759 = n5756 & ~n5758 ;
  assign n5760 = x961 & n5631 ;
  assign n5761 = x299 | n5760 ;
  assign n5762 = ( x232 & ~n5759 ) | ( x232 & n5761 ) | ( ~n5759 & n5761 ) ;
  assign n5763 = ~x232 & n5762 ;
  assign n5764 = x961 & n5642 ;
  assign n5765 = x299 | n5764 ;
  assign n5766 = n5647 & n5757 ;
  assign n5767 = n5755 | n5766 ;
  assign n5768 = n5303 & n5767 ;
  assign n5769 = ( n5651 & n5759 ) | ( n5651 & ~n5768 ) | ( n5759 & ~n5768 ) ;
  assign n5770 = ~n5768 & n5769 ;
  assign n5771 = x232 & ~n5770 ;
  assign n5772 = n5765 & n5771 ;
  assign n5773 = ( ~x39 & n5763 ) | ( ~x39 & n5772 ) | ( n5763 & n5772 ) ;
  assign n5774 = ~x39 & n5773 ;
  assign n5775 = x39 & ~n5658 ;
  assign n5776 = x299 & x972 ;
  assign n5777 = n5666 & n5776 ;
  assign n5778 = ~x299 & x961 ;
  assign n5779 = n5661 & n5778 ;
  assign n5780 = n5777 | n5779 ;
  assign n5781 = n5775 & n5780 ;
  assign n5782 = ( x38 & ~n5774 ) | ( x38 & n5781 ) | ( ~n5774 & n5781 ) ;
  assign n5783 = n5774 | n5782 ;
  assign n5784 = x961 & ~n5673 ;
  assign n5785 = x299 | n5784 ;
  assign n5786 = ~n5088 & n5757 ;
  assign n5787 = n5756 & ~n5786 ;
  assign n5788 = ( x39 & n5785 ) | ( x39 & ~n5787 ) | ( n5785 & ~n5787 ) ;
  assign n5789 = ~x39 & n5788 ;
  assign n5790 = ( n5624 & n5776 ) | ( n5624 & n5778 ) | ( n5776 & n5778 ) ;
  assign n5791 = x39 & n5790 ;
  assign n5792 = x38 & ~n5791 ;
  assign n5793 = ~n5789 & n5792 ;
  assign n5794 = ( x100 & n5783 ) | ( x100 & ~n5793 ) | ( n5783 & ~n5793 ) ;
  assign n5795 = n5794 ^ n5783 ^ 1'b0 ;
  assign n5796 = ( x100 & n5794 ) | ( x100 & ~n5795 ) | ( n5794 & ~n5795 ) ;
  assign n5797 = n1994 & n5790 ;
  assign n5798 = x961 & n5693 ;
  assign n5799 = x299 | n5798 ;
  assign n5800 = x972 & n5699 ;
  assign n5801 = n5756 & ~n5800 ;
  assign n5802 = ( n1994 & n5799 ) | ( n1994 & ~n5801 ) | ( n5799 & ~n5801 ) ;
  assign n5803 = ~n1994 & n5802 ;
  assign n5804 = ( x100 & n5797 ) | ( x100 & ~n5803 ) | ( n5797 & ~n5803 ) ;
  assign n5805 = ~n5797 & n5804 ;
  assign n5806 = ( x87 & n5796 ) | ( x87 & ~n5805 ) | ( n5796 & ~n5805 ) ;
  assign n5807 = ~x87 & n5806 ;
  assign n5808 = x87 & n5790 ;
  assign n5809 = ( x75 & ~n5807 ) | ( x75 & n5808 ) | ( ~n5807 & n5808 ) ;
  assign n5810 = n5807 | n5809 ;
  assign n5811 = x75 & ~n5790 ;
  assign n5812 = x92 & ~n5811 ;
  assign n5813 = n5812 ^ x54 ^ 1'b0 ;
  assign n5814 = n1207 & n5790 ;
  assign n5815 = ~n2052 & n5789 ;
  assign n5816 = n5814 | n5815 ;
  assign n5817 = x75 | n5816 ;
  assign n5818 = ( n5812 & ~n5813 ) | ( n5812 & n5817 ) | ( ~n5813 & n5817 ) ;
  assign n5819 = ( x54 & n5813 ) | ( x54 & n5818 ) | ( n5813 & n5818 ) ;
  assign n5820 = x75 & ~n5816 ;
  assign n5821 = x92 | n5820 ;
  assign n5822 = ~n5819 & n5821 ;
  assign n5823 = ( n5810 & n5819 ) | ( n5810 & ~n5822 ) | ( n5819 & ~n5822 ) ;
  assign n5824 = n5459 & ~n5790 ;
  assign n5825 = x74 & ~n5824 ;
  assign n5826 = n5825 ^ x55 ^ 1'b0 ;
  assign n5827 = n2053 | n5816 ;
  assign n5828 = x54 | n5827 ;
  assign n5829 = ( n5825 & ~n5826 ) | ( n5825 & n5828 ) | ( ~n5826 & n5828 ) ;
  assign n5830 = ( x55 & n5826 ) | ( x55 & n5829 ) | ( n5826 & n5829 ) ;
  assign n5831 = n2053 & ~n5790 ;
  assign n5832 = x54 & ~n5827 ;
  assign n5833 = ( x54 & n5831 ) | ( x54 & n5832 ) | ( n5831 & n5832 ) ;
  assign n5834 = x74 | n5833 ;
  assign n5835 = ~n5830 & n5834 ;
  assign n5836 = ( n5823 & n5830 ) | ( n5823 & ~n5835 ) | ( n5830 & ~n5835 ) ;
  assign n5837 = ~n2070 & n5786 ;
  assign n5838 = x55 & ~n5755 ;
  assign n5839 = ~n5837 & n5838 ;
  assign n5840 = ( n2109 & n5836 ) | ( n2109 & ~n5839 ) | ( n5836 & ~n5839 ) ;
  assign n5841 = ~n2109 & n5840 ;
  assign n5842 = n2109 & n5755 ;
  assign n5843 = ( x59 & ~n5841 ) | ( x59 & n5842 ) | ( ~n5841 & n5842 ) ;
  assign n5844 = n5841 | n5843 ;
  assign n5845 = x59 & ~n5755 ;
  assign n5846 = ~n5192 & n5837 ;
  assign n5847 = n5845 & ~n5846 ;
  assign n5848 = ( x57 & n5844 ) | ( x57 & ~n5847 ) | ( n5844 & ~n5847 ) ;
  assign n5849 = ~x57 & n5848 ;
  assign n5850 = ~n5193 & n5837 ;
  assign n5851 = n5755 | n5850 ;
  assign n5852 = n5849 ^ x57 ^ 1'b0 ;
  assign n5853 = ( ~x57 & n5851 ) | ( ~x57 & n5852 ) | ( n5851 & n5852 ) ;
  assign n5854 = ( x57 & n5849 ) | ( x57 & n5853 ) | ( n5849 & n5853 ) ;
  assign n5855 = x960 & n5624 ;
  assign n5856 = x299 & ~n5855 ;
  assign n5857 = ~x228 & x960 ;
  assign n5858 = n5628 & n5857 ;
  assign n5859 = n5856 & ~n5858 ;
  assign n5860 = x977 & n5631 ;
  assign n5861 = x299 | n5860 ;
  assign n5862 = ( x232 & ~n5859 ) | ( x232 & n5861 ) | ( ~n5859 & n5861 ) ;
  assign n5863 = ~x232 & n5862 ;
  assign n5864 = x977 & n5642 ;
  assign n5865 = x299 | n5864 ;
  assign n5866 = n5647 & n5857 ;
  assign n5867 = n5855 | n5866 ;
  assign n5868 = n5303 & n5867 ;
  assign n5869 = ( n5651 & n5859 ) | ( n5651 & ~n5868 ) | ( n5859 & ~n5868 ) ;
  assign n5870 = ~n5868 & n5869 ;
  assign n5871 = x232 & ~n5870 ;
  assign n5872 = n5865 & n5871 ;
  assign n5873 = ( ~x39 & n5863 ) | ( ~x39 & n5872 ) | ( n5863 & n5872 ) ;
  assign n5874 = ~x39 & n5873 ;
  assign n5875 = x299 & x960 ;
  assign n5876 = n5666 & n5875 ;
  assign n5877 = ~x299 & x977 ;
  assign n5878 = n5661 & n5877 ;
  assign n5879 = n5876 | n5878 ;
  assign n5880 = n5775 & n5879 ;
  assign n5881 = ( x38 & ~n5874 ) | ( x38 & n5880 ) | ( ~n5874 & n5880 ) ;
  assign n5882 = n5874 | n5881 ;
  assign n5883 = x977 & ~n5673 ;
  assign n5884 = x299 | n5883 ;
  assign n5885 = ~n5088 & n5857 ;
  assign n5886 = n5856 & ~n5885 ;
  assign n5887 = ( x39 & n5884 ) | ( x39 & ~n5886 ) | ( n5884 & ~n5886 ) ;
  assign n5888 = ~x39 & n5887 ;
  assign n5889 = ( n5624 & n5875 ) | ( n5624 & n5877 ) | ( n5875 & n5877 ) ;
  assign n5890 = x39 & n5889 ;
  assign n5891 = x38 & ~n5890 ;
  assign n5892 = ~n5888 & n5891 ;
  assign n5893 = ( x100 & n5882 ) | ( x100 & ~n5892 ) | ( n5882 & ~n5892 ) ;
  assign n5894 = n5893 ^ n5882 ^ 1'b0 ;
  assign n5895 = ( x100 & n5893 ) | ( x100 & ~n5894 ) | ( n5893 & ~n5894 ) ;
  assign n5896 = n1994 & n5889 ;
  assign n5897 = x977 & n5693 ;
  assign n5898 = x299 | n5897 ;
  assign n5899 = x960 & n5699 ;
  assign n5900 = n5856 & ~n5899 ;
  assign n5901 = ( n1994 & n5898 ) | ( n1994 & ~n5900 ) | ( n5898 & ~n5900 ) ;
  assign n5902 = ~n1994 & n5901 ;
  assign n5903 = ( x100 & n5896 ) | ( x100 & ~n5902 ) | ( n5896 & ~n5902 ) ;
  assign n5904 = ~n5896 & n5903 ;
  assign n5905 = ( x87 & n5895 ) | ( x87 & ~n5904 ) | ( n5895 & ~n5904 ) ;
  assign n5906 = ~x87 & n5905 ;
  assign n5907 = x87 & n5889 ;
  assign n5908 = ( x75 & ~n5906 ) | ( x75 & n5907 ) | ( ~n5906 & n5907 ) ;
  assign n5909 = n5906 | n5908 ;
  assign n5910 = x75 & ~n5889 ;
  assign n5911 = x92 & ~n5910 ;
  assign n5912 = n5911 ^ x54 ^ 1'b0 ;
  assign n5913 = n1207 & n5889 ;
  assign n5914 = ~n2052 & n5888 ;
  assign n5915 = n5913 | n5914 ;
  assign n5916 = x75 | n5915 ;
  assign n5917 = ( n5911 & ~n5912 ) | ( n5911 & n5916 ) | ( ~n5912 & n5916 ) ;
  assign n5918 = ( x54 & n5912 ) | ( x54 & n5917 ) | ( n5912 & n5917 ) ;
  assign n5919 = x75 & ~n5915 ;
  assign n5920 = x92 | n5919 ;
  assign n5921 = ~n5918 & n5920 ;
  assign n5922 = ( n5909 & n5918 ) | ( n5909 & ~n5921 ) | ( n5918 & ~n5921 ) ;
  assign n5923 = n5459 & ~n5889 ;
  assign n5924 = x74 & ~n5923 ;
  assign n5925 = n5924 ^ x55 ^ 1'b0 ;
  assign n5926 = n2053 | n5915 ;
  assign n5927 = x54 | n5926 ;
  assign n5928 = ( n5924 & ~n5925 ) | ( n5924 & n5927 ) | ( ~n5925 & n5927 ) ;
  assign n5929 = ( x55 & n5925 ) | ( x55 & n5928 ) | ( n5925 & n5928 ) ;
  assign n5930 = n2053 & ~n5889 ;
  assign n5931 = x54 & ~n5926 ;
  assign n5932 = ( x54 & n5930 ) | ( x54 & n5931 ) | ( n5930 & n5931 ) ;
  assign n5933 = x74 | n5932 ;
  assign n5934 = ~n5929 & n5933 ;
  assign n5935 = ( n5922 & n5929 ) | ( n5922 & ~n5934 ) | ( n5929 & ~n5934 ) ;
  assign n5936 = ~n2070 & n5885 ;
  assign n5937 = x55 & ~n5855 ;
  assign n5938 = ~n5936 & n5937 ;
  assign n5939 = ( n2109 & n5935 ) | ( n2109 & ~n5938 ) | ( n5935 & ~n5938 ) ;
  assign n5940 = ~n2109 & n5939 ;
  assign n5941 = n2109 & n5855 ;
  assign n5942 = ( x59 & ~n5940 ) | ( x59 & n5941 ) | ( ~n5940 & n5941 ) ;
  assign n5943 = n5940 | n5942 ;
  assign n5944 = x59 & ~n5855 ;
  assign n5945 = ~n5192 & n5936 ;
  assign n5946 = n5944 & ~n5945 ;
  assign n5947 = ( x57 & n5943 ) | ( x57 & ~n5946 ) | ( n5943 & ~n5946 ) ;
  assign n5948 = ~x57 & n5947 ;
  assign n5949 = ~n5193 & n5936 ;
  assign n5950 = n5855 | n5949 ;
  assign n5951 = n5948 ^ x57 ^ 1'b0 ;
  assign n5952 = ( ~x57 & n5950 ) | ( ~x57 & n5951 ) | ( n5950 & n5951 ) ;
  assign n5953 = ( x57 & n5948 ) | ( x57 & n5952 ) | ( n5948 & n5952 ) ;
  assign n5954 = x963 & n5624 ;
  assign n5955 = x299 & ~n5954 ;
  assign n5956 = ~x228 & x963 ;
  assign n5957 = n5628 & n5956 ;
  assign n5958 = n5955 & ~n5957 ;
  assign n5959 = x969 & n5631 ;
  assign n5960 = x299 | n5959 ;
  assign n5961 = ( x232 & ~n5958 ) | ( x232 & n5960 ) | ( ~n5958 & n5960 ) ;
  assign n5962 = ~x232 & n5961 ;
  assign n5963 = x969 & n5642 ;
  assign n5964 = x299 | n5963 ;
  assign n5965 = n5647 & n5956 ;
  assign n5966 = n5954 | n5965 ;
  assign n5967 = n5303 & n5966 ;
  assign n5968 = ( n5651 & n5958 ) | ( n5651 & ~n5967 ) | ( n5958 & ~n5967 ) ;
  assign n5969 = ~n5967 & n5968 ;
  assign n5970 = x232 & ~n5969 ;
  assign n5971 = n5964 & n5970 ;
  assign n5972 = ( ~x39 & n5962 ) | ( ~x39 & n5971 ) | ( n5962 & n5971 ) ;
  assign n5973 = ~x39 & n5972 ;
  assign n5974 = x299 & x963 ;
  assign n5975 = n5666 & n5974 ;
  assign n5976 = ~x299 & x969 ;
  assign n5977 = n5661 & n5976 ;
  assign n5978 = n5975 | n5977 ;
  assign n5979 = n5775 & n5978 ;
  assign n5980 = ( x38 & ~n5973 ) | ( x38 & n5979 ) | ( ~n5973 & n5979 ) ;
  assign n5981 = n5973 | n5980 ;
  assign n5982 = x969 & ~n5673 ;
  assign n5983 = x299 | n5982 ;
  assign n5984 = ~n5088 & n5956 ;
  assign n5985 = n5955 & ~n5984 ;
  assign n5986 = ( x39 & n5983 ) | ( x39 & ~n5985 ) | ( n5983 & ~n5985 ) ;
  assign n5987 = ~x39 & n5986 ;
  assign n5988 = ( n5624 & n5974 ) | ( n5624 & n5976 ) | ( n5974 & n5976 ) ;
  assign n5989 = x39 & n5988 ;
  assign n5990 = x38 & ~n5989 ;
  assign n5991 = ~n5987 & n5990 ;
  assign n5992 = ( x100 & n5981 ) | ( x100 & ~n5991 ) | ( n5981 & ~n5991 ) ;
  assign n5993 = n5992 ^ n5981 ^ 1'b0 ;
  assign n5994 = ( x100 & n5992 ) | ( x100 & ~n5993 ) | ( n5992 & ~n5993 ) ;
  assign n5995 = n1994 & n5988 ;
  assign n5996 = x969 & n5693 ;
  assign n5997 = x299 | n5996 ;
  assign n5998 = x963 & n5699 ;
  assign n5999 = n5955 & ~n5998 ;
  assign n6000 = ( n1994 & n5997 ) | ( n1994 & ~n5999 ) | ( n5997 & ~n5999 ) ;
  assign n6001 = ~n1994 & n6000 ;
  assign n6002 = ( x100 & n5995 ) | ( x100 & ~n6001 ) | ( n5995 & ~n6001 ) ;
  assign n6003 = ~n5995 & n6002 ;
  assign n6004 = ( x87 & n5994 ) | ( x87 & ~n6003 ) | ( n5994 & ~n6003 ) ;
  assign n6005 = ~x87 & n6004 ;
  assign n6006 = x87 & n5988 ;
  assign n6007 = ( x75 & ~n6005 ) | ( x75 & n6006 ) | ( ~n6005 & n6006 ) ;
  assign n6008 = n6005 | n6007 ;
  assign n6009 = x75 & ~n5988 ;
  assign n6010 = x92 & ~n6009 ;
  assign n6011 = n6010 ^ x54 ^ 1'b0 ;
  assign n6012 = n1207 & n5988 ;
  assign n6013 = ~n2052 & n5987 ;
  assign n6014 = n6012 | n6013 ;
  assign n6015 = x75 | n6014 ;
  assign n6016 = ( n6010 & ~n6011 ) | ( n6010 & n6015 ) | ( ~n6011 & n6015 ) ;
  assign n6017 = ( x54 & n6011 ) | ( x54 & n6016 ) | ( n6011 & n6016 ) ;
  assign n6018 = x75 & ~n6014 ;
  assign n6019 = x92 | n6018 ;
  assign n6020 = ~n6017 & n6019 ;
  assign n6021 = ( n6008 & n6017 ) | ( n6008 & ~n6020 ) | ( n6017 & ~n6020 ) ;
  assign n6022 = n5459 & ~n5988 ;
  assign n6023 = x74 & ~n6022 ;
  assign n6024 = n6023 ^ x55 ^ 1'b0 ;
  assign n6025 = n2053 | n6014 ;
  assign n6026 = x54 | n6025 ;
  assign n6027 = ( n6023 & ~n6024 ) | ( n6023 & n6026 ) | ( ~n6024 & n6026 ) ;
  assign n6028 = ( x55 & n6024 ) | ( x55 & n6027 ) | ( n6024 & n6027 ) ;
  assign n6029 = n2053 & ~n5988 ;
  assign n6030 = x54 & ~n6025 ;
  assign n6031 = ( x54 & n6029 ) | ( x54 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6032 = x74 | n6031 ;
  assign n6033 = ~n6028 & n6032 ;
  assign n6034 = ( n6021 & n6028 ) | ( n6021 & ~n6033 ) | ( n6028 & ~n6033 ) ;
  assign n6035 = ~n2070 & n5984 ;
  assign n6036 = x55 & ~n5954 ;
  assign n6037 = ~n6035 & n6036 ;
  assign n6038 = ( n2109 & n6034 ) | ( n2109 & ~n6037 ) | ( n6034 & ~n6037 ) ;
  assign n6039 = ~n2109 & n6038 ;
  assign n6040 = n2109 & n5954 ;
  assign n6041 = ( x59 & ~n6039 ) | ( x59 & n6040 ) | ( ~n6039 & n6040 ) ;
  assign n6042 = n6039 | n6041 ;
  assign n6043 = x59 & ~n5954 ;
  assign n6044 = ~n5192 & n6035 ;
  assign n6045 = n6043 & ~n6044 ;
  assign n6046 = ( x57 & n6042 ) | ( x57 & ~n6045 ) | ( n6042 & ~n6045 ) ;
  assign n6047 = ~x57 & n6046 ;
  assign n6048 = ~n5193 & n6035 ;
  assign n6049 = n5954 | n6048 ;
  assign n6050 = n6047 ^ x57 ^ 1'b0 ;
  assign n6051 = ( ~x57 & n6049 ) | ( ~x57 & n6050 ) | ( n6049 & n6050 ) ;
  assign n6052 = ( x57 & n6047 ) | ( x57 & n6051 ) | ( n6047 & n6051 ) ;
  assign n6053 = x975 & n5624 ;
  assign n6054 = x299 & ~n6053 ;
  assign n6055 = ~x228 & x975 ;
  assign n6056 = n5628 & n6055 ;
  assign n6057 = n6054 & ~n6056 ;
  assign n6058 = x971 & n5631 ;
  assign n6059 = x299 | n6058 ;
  assign n6060 = ( x232 & ~n6057 ) | ( x232 & n6059 ) | ( ~n6057 & n6059 ) ;
  assign n6061 = ~x232 & n6060 ;
  assign n6062 = x971 & n5642 ;
  assign n6063 = x299 | n6062 ;
  assign n6064 = n5647 & n6055 ;
  assign n6065 = n6053 | n6064 ;
  assign n6066 = n5303 & n6065 ;
  assign n6067 = ( n5651 & n6057 ) | ( n5651 & ~n6066 ) | ( n6057 & ~n6066 ) ;
  assign n6068 = ~n6066 & n6067 ;
  assign n6069 = x232 & ~n6068 ;
  assign n6070 = n6063 & n6069 ;
  assign n6071 = ( ~x39 & n6061 ) | ( ~x39 & n6070 ) | ( n6061 & n6070 ) ;
  assign n6072 = ~x39 & n6071 ;
  assign n6073 = x299 & x975 ;
  assign n6074 = n5666 & n6073 ;
  assign n6075 = ~x299 & x971 ;
  assign n6076 = n5661 & n6075 ;
  assign n6077 = n6074 | n6076 ;
  assign n6078 = n5775 & n6077 ;
  assign n6079 = ( x38 & ~n6072 ) | ( x38 & n6078 ) | ( ~n6072 & n6078 ) ;
  assign n6080 = n6072 | n6079 ;
  assign n6081 = x971 & ~n5673 ;
  assign n6082 = x299 | n6081 ;
  assign n6083 = ~n5088 & n6055 ;
  assign n6084 = n6054 & ~n6083 ;
  assign n6085 = ( x39 & n6082 ) | ( x39 & ~n6084 ) | ( n6082 & ~n6084 ) ;
  assign n6086 = ~x39 & n6085 ;
  assign n6087 = ( n5624 & n6073 ) | ( n5624 & n6075 ) | ( n6073 & n6075 ) ;
  assign n6088 = x39 & n6087 ;
  assign n6089 = x38 & ~n6088 ;
  assign n6090 = ~n6086 & n6089 ;
  assign n6091 = ( x100 & n6080 ) | ( x100 & ~n6090 ) | ( n6080 & ~n6090 ) ;
  assign n6092 = n6091 ^ n6080 ^ 1'b0 ;
  assign n6093 = ( x100 & n6091 ) | ( x100 & ~n6092 ) | ( n6091 & ~n6092 ) ;
  assign n6094 = n1994 & n6087 ;
  assign n6095 = x971 & n5693 ;
  assign n6096 = x299 | n6095 ;
  assign n6097 = x975 & n5699 ;
  assign n6098 = n6054 & ~n6097 ;
  assign n6099 = ( n1994 & n6096 ) | ( n1994 & ~n6098 ) | ( n6096 & ~n6098 ) ;
  assign n6100 = ~n1994 & n6099 ;
  assign n6101 = ( x100 & n6094 ) | ( x100 & ~n6100 ) | ( n6094 & ~n6100 ) ;
  assign n6102 = ~n6094 & n6101 ;
  assign n6103 = ( x87 & n6093 ) | ( x87 & ~n6102 ) | ( n6093 & ~n6102 ) ;
  assign n6104 = ~x87 & n6103 ;
  assign n6105 = x87 & n6087 ;
  assign n6106 = ( x75 & ~n6104 ) | ( x75 & n6105 ) | ( ~n6104 & n6105 ) ;
  assign n6107 = n6104 | n6106 ;
  assign n6108 = x75 & ~n6087 ;
  assign n6109 = x92 & ~n6108 ;
  assign n6110 = n6109 ^ x54 ^ 1'b0 ;
  assign n6111 = n1207 & n6087 ;
  assign n6112 = ~n2052 & n6086 ;
  assign n6113 = n6111 | n6112 ;
  assign n6114 = x75 | n6113 ;
  assign n6115 = ( n6109 & ~n6110 ) | ( n6109 & n6114 ) | ( ~n6110 & n6114 ) ;
  assign n6116 = ( x54 & n6110 ) | ( x54 & n6115 ) | ( n6110 & n6115 ) ;
  assign n6117 = x75 & ~n6113 ;
  assign n6118 = x92 | n6117 ;
  assign n6119 = ~n6116 & n6118 ;
  assign n6120 = ( n6107 & n6116 ) | ( n6107 & ~n6119 ) | ( n6116 & ~n6119 ) ;
  assign n6121 = n5459 & ~n6087 ;
  assign n6122 = x74 & ~n6121 ;
  assign n6123 = n6122 ^ x55 ^ 1'b0 ;
  assign n6124 = n2053 | n6113 ;
  assign n6125 = x54 | n6124 ;
  assign n6126 = ( n6122 & ~n6123 ) | ( n6122 & n6125 ) | ( ~n6123 & n6125 ) ;
  assign n6127 = ( x55 & n6123 ) | ( x55 & n6126 ) | ( n6123 & n6126 ) ;
  assign n6128 = n2053 & ~n6087 ;
  assign n6129 = x54 & ~n6124 ;
  assign n6130 = ( x54 & n6128 ) | ( x54 & n6129 ) | ( n6128 & n6129 ) ;
  assign n6131 = x74 | n6130 ;
  assign n6132 = ~n6127 & n6131 ;
  assign n6133 = ( n6120 & n6127 ) | ( n6120 & ~n6132 ) | ( n6127 & ~n6132 ) ;
  assign n6134 = ~n2070 & n6083 ;
  assign n6135 = x55 & ~n6053 ;
  assign n6136 = ~n6134 & n6135 ;
  assign n6137 = ( n2109 & n6133 ) | ( n2109 & ~n6136 ) | ( n6133 & ~n6136 ) ;
  assign n6138 = ~n2109 & n6137 ;
  assign n6139 = n2109 & n6053 ;
  assign n6140 = ( x59 & ~n6138 ) | ( x59 & n6139 ) | ( ~n6138 & n6139 ) ;
  assign n6141 = n6138 | n6140 ;
  assign n6142 = x59 & ~n6053 ;
  assign n6143 = ~n5192 & n6134 ;
  assign n6144 = n6142 & ~n6143 ;
  assign n6145 = ( x57 & n6141 ) | ( x57 & ~n6144 ) | ( n6141 & ~n6144 ) ;
  assign n6146 = ~x57 & n6145 ;
  assign n6147 = ~n5193 & n6134 ;
  assign n6148 = n6053 | n6147 ;
  assign n6149 = n6146 ^ x57 ^ 1'b0 ;
  assign n6150 = ( ~x57 & n6148 ) | ( ~x57 & n6149 ) | ( n6148 & n6149 ) ;
  assign n6151 = ( x57 & n6146 ) | ( x57 & n6150 ) | ( n6146 & n6150 ) ;
  assign n6152 = ~x299 & x974 ;
  assign n6153 = x299 & x978 ;
  assign n6154 = n6152 | n6153 ;
  assign n6155 = n5624 & n6154 ;
  assign n6156 = x39 & n6155 ;
  assign n6157 = ~n5673 & n6154 ;
  assign n6158 = ~x39 & n6157 ;
  assign n6159 = ( x38 & n6156 ) | ( x38 & ~n6158 ) | ( n6156 & ~n6158 ) ;
  assign n6160 = ~n6156 & n6159 ;
  assign n6161 = x978 & n5624 ;
  assign n6162 = x299 & ~n6161 ;
  assign n6163 = ~x228 & x978 ;
  assign n6164 = n5628 & n6163 ;
  assign n6165 = n6162 & ~n6164 ;
  assign n6166 = x974 & n5631 ;
  assign n6167 = x299 | n6166 ;
  assign n6168 = ( x232 & ~n6165 ) | ( x232 & n6167 ) | ( ~n6165 & n6167 ) ;
  assign n6169 = ~x232 & n6168 ;
  assign n6170 = x974 & n5642 ;
  assign n6171 = x299 | n6170 ;
  assign n6172 = n5647 & n6163 ;
  assign n6173 = n6161 | n6172 ;
  assign n6174 = n5303 & n6173 ;
  assign n6175 = ( n5651 & n6165 ) | ( n5651 & ~n6174 ) | ( n6165 & ~n6174 ) ;
  assign n6176 = ~n6174 & n6175 ;
  assign n6177 = x232 & ~n6176 ;
  assign n6178 = n6171 & n6177 ;
  assign n6179 = ( ~x39 & n6169 ) | ( ~x39 & n6178 ) | ( n6169 & n6178 ) ;
  assign n6180 = ~x39 & n6179 ;
  assign n6181 = n5666 & n6153 ;
  assign n6182 = n5661 & n6152 ;
  assign n6183 = n6181 | n6182 ;
  assign n6184 = n5775 & n6183 ;
  assign n6185 = ( x38 & ~n6180 ) | ( x38 & n6184 ) | ( ~n6180 & n6184 ) ;
  assign n6186 = n6180 | n6185 ;
  assign n6187 = n6186 ^ n6160 ^ 1'b0 ;
  assign n6188 = ( n6160 & n6186 ) | ( n6160 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6189 = ( x100 & ~n6160 ) | ( x100 & n6188 ) | ( ~n6160 & n6188 ) ;
  assign n6190 = n1994 & n6155 ;
  assign n6191 = x974 & n5693 ;
  assign n6192 = x299 | n6191 ;
  assign n6193 = x978 & n5699 ;
  assign n6194 = n6162 & ~n6193 ;
  assign n6195 = ( n1994 & n6192 ) | ( n1994 & ~n6194 ) | ( n6192 & ~n6194 ) ;
  assign n6196 = ~n1994 & n6195 ;
  assign n6197 = ( x100 & n6190 ) | ( x100 & ~n6196 ) | ( n6190 & ~n6196 ) ;
  assign n6198 = ~n6190 & n6197 ;
  assign n6199 = ( x87 & n6189 ) | ( x87 & ~n6198 ) | ( n6189 & ~n6198 ) ;
  assign n6200 = ~x87 & n6199 ;
  assign n6201 = x87 & n6155 ;
  assign n6202 = ( x75 & ~n6200 ) | ( x75 & n6201 ) | ( ~n6200 & n6201 ) ;
  assign n6203 = n6200 | n6202 ;
  assign n6204 = ~x228 & n1207 ;
  assign n6205 = n6157 & ~n6204 ;
  assign n6206 = x75 | n6205 ;
  assign n6207 = n6206 ^ x54 ^ 1'b0 ;
  assign n6208 = x75 & ~n6155 ;
  assign n6209 = x92 & ~n6208 ;
  assign n6210 = ( n6206 & ~n6207 ) | ( n6206 & n6209 ) | ( ~n6207 & n6209 ) ;
  assign n6211 = ( x54 & n6207 ) | ( x54 & n6210 ) | ( n6207 & n6210 ) ;
  assign n6212 = x75 & ~n6205 ;
  assign n6213 = x92 | n6212 ;
  assign n6214 = ~n6211 & n6213 ;
  assign n6215 = ( n6203 & n6211 ) | ( n6203 & ~n6214 ) | ( n6211 & ~n6214 ) ;
  assign n6216 = n5459 & ~n6155 ;
  assign n6217 = x74 & ~n6216 ;
  assign n6218 = n6217 ^ x55 ^ 1'b0 ;
  assign n6219 = n2053 | n6205 ;
  assign n6220 = x54 | n6219 ;
  assign n6221 = ( n6217 & ~n6218 ) | ( n6217 & n6220 ) | ( ~n6218 & n6220 ) ;
  assign n6222 = ( x55 & n6218 ) | ( x55 & n6221 ) | ( n6218 & n6221 ) ;
  assign n6223 = n2053 & ~n6155 ;
  assign n6224 = x54 & ~n6219 ;
  assign n6225 = ( x54 & n6223 ) | ( x54 & n6224 ) | ( n6223 & n6224 ) ;
  assign n6226 = x74 | n6225 ;
  assign n6227 = ~n6222 & n6226 ;
  assign n6228 = ( n6215 & n6222 ) | ( n6215 & ~n6227 ) | ( n6222 & ~n6227 ) ;
  assign n6229 = ~n2070 & n6163 ;
  assign n6230 = ~n5088 & n6229 ;
  assign n6231 = x55 & ~n6161 ;
  assign n6232 = ~n6230 & n6231 ;
  assign n6233 = ( n2109 & n6228 ) | ( n2109 & ~n6232 ) | ( n6228 & ~n6232 ) ;
  assign n6234 = ~n2109 & n6233 ;
  assign n6235 = n2109 & n6161 ;
  assign n6236 = ( x59 & ~n6234 ) | ( x59 & n6235 ) | ( ~n6234 & n6235 ) ;
  assign n6237 = n6234 | n6236 ;
  assign n6238 = x59 & ~n6161 ;
  assign n6239 = ~n5192 & n6230 ;
  assign n6240 = n6238 & ~n6239 ;
  assign n6241 = ( x57 & n6237 ) | ( x57 & ~n6240 ) | ( n6237 & ~n6240 ) ;
  assign n6242 = ~x57 & n6241 ;
  assign n6243 = ~n5193 & n6230 ;
  assign n6244 = n6161 | n6243 ;
  assign n6245 = n6242 ^ x57 ^ 1'b0 ;
  assign n6246 = ( ~x57 & n6244 ) | ( ~x57 & n6245 ) | ( n6244 & n6245 ) ;
  assign n6247 = ( x57 & n6242 ) | ( x57 & n6246 ) | ( n6242 & n6246 ) ;
  assign n6248 = n2097 | n5003 ;
  assign n6249 = x55 & n6248 ;
  assign n6250 = x56 | n6249 ;
  assign n6251 = n1205 | n2044 ;
  assign n6252 = n5017 | n6251 ;
  assign n6253 = x92 | n6252 ;
  assign n6254 = x54 & n6253 ;
  assign n6255 = n2052 | n5017 ;
  assign n6256 = x75 & n6255 ;
  assign n6257 = x92 & n6252 ;
  assign n6258 = n6256 | n6257 ;
  assign n6259 = x38 | n5017 ;
  assign n6260 = x100 & n6259 ;
  assign n6261 = ~x299 & n5115 ;
  assign n6262 = n5382 & n6261 ;
  assign n6263 = x299 & n5100 ;
  assign n6264 = n5664 & n6263 ;
  assign n6265 = ( x39 & n6262 ) | ( x39 & ~n6264 ) | ( n6262 & ~n6264 ) ;
  assign n6266 = ~n6262 & n6265 ;
  assign n6267 = x299 | n5287 ;
  assign n6268 = x299 & ~n5296 ;
  assign n6269 = x232 | n6268 ;
  assign n6270 = n6267 & ~n6269 ;
  assign n6271 = ~n5334 & n5651 ;
  assign n6272 = ~n5646 & n6271 ;
  assign n6273 = ~n5303 & n6268 ;
  assign n6274 = x232 & ~n6273 ;
  assign n6275 = x299 | n5347 ;
  assign n6276 = n5344 & n5346 ;
  assign n6277 = ( n5638 & ~n6275 ) | ( n5638 & n6276 ) | ( ~n6275 & n6276 ) ;
  assign n6278 = n6275 | n6277 ;
  assign n6279 = ( n6272 & n6274 ) | ( n6272 & n6278 ) | ( n6274 & n6278 ) ;
  assign n6280 = ~n6272 & n6279 ;
  assign n6281 = ( x39 & ~n6270 ) | ( x39 & n6280 ) | ( ~n6270 & n6280 ) ;
  assign n6282 = n6270 | n6281 ;
  assign n6283 = n6282 ^ n6266 ^ 1'b0 ;
  assign n6284 = ( n6266 & n6282 ) | ( n6266 & n6283 ) | ( n6282 & n6283 ) ;
  assign n6285 = ( x38 & ~n6266 ) | ( x38 & n6284 ) | ( ~n6266 & n6284 ) ;
  assign n6286 = n6285 ^ n5053 ^ 1'b0 ;
  assign n6287 = ( n5053 & n6285 ) | ( n5053 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = ( x100 & ~n5053 ) | ( x100 & n6287 ) | ( ~n5053 & n6287 ) ;
  assign n6289 = ( n5051 & ~n6260 ) | ( n5051 & n6288 ) | ( ~n6260 & n6288 ) ;
  assign n6290 = ~n5051 & n6289 ;
  assign n6291 = ( x75 & x92 ) | ( x75 & ~n6290 ) | ( x92 & ~n6290 ) ;
  assign n6292 = n6290 | n6291 ;
  assign n6293 = n6292 ^ n6258 ^ 1'b0 ;
  assign n6294 = ( n6258 & n6292 ) | ( n6258 & n6293 ) | ( n6292 & n6293 ) ;
  assign n6295 = ( x54 & ~n6258 ) | ( x54 & n6294 ) | ( ~n6258 & n6294 ) ;
  assign n6296 = n6295 ^ n6254 ^ 1'b0 ;
  assign n6297 = ( n6254 & n6295 ) | ( n6254 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6298 = ( x74 & ~n6254 ) | ( x74 & n6297 ) | ( ~n6254 & n6297 ) ;
  assign n6299 = n6298 ^ n5011 ^ 1'b0 ;
  assign n6300 = ( n5011 & n6298 ) | ( n5011 & n6299 ) | ( n6298 & n6299 ) ;
  assign n6301 = ( x55 & ~n5011 ) | ( x55 & n6300 ) | ( ~n5011 & n6300 ) ;
  assign n6302 = ( x62 & ~n6250 ) | ( x62 & n6301 ) | ( ~n6250 & n6301 ) ;
  assign n6303 = ~x62 & n6302 ;
  assign n6304 = n2120 | n6303 ;
  assign n6305 = ~n5190 & n6304 ;
  assign n6306 = x954 ^ x24 ^ 1'b0 ;
  assign n6307 = ( ~x24 & n6305 ) | ( ~x24 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6308 = ~x228 & n2230 ;
  assign n6309 = ~x100 & n6308 ;
  assign n6310 = n1292 | n5413 ;
  assign n6311 = n2404 ^ x299 ^ 1'b0 ;
  assign n6312 = ( n2404 & n6310 ) | ( n2404 & ~n6311 ) | ( n6310 & ~n6311 ) ;
  assign n6313 = x100 & ~n2142 ;
  assign n6314 = ~n6312 & n6313 ;
  assign n6315 = ( x39 & ~n6309 ) | ( x39 & n6314 ) | ( ~n6309 & n6314 ) ;
  assign n6316 = n6309 | n6315 ;
  assign n6317 = x100 | n2142 ;
  assign n6318 = x39 & n6317 ;
  assign n6319 = ( x38 & n6316 ) | ( x38 & ~n6318 ) | ( n6316 & ~n6318 ) ;
  assign n6320 = ~x38 & n6319 ;
  assign n6321 = ( ~x87 & n1323 ) | ( ~x87 & n6320 ) | ( n1323 & n6320 ) ;
  assign n6322 = ~x87 & n6321 ;
  assign n6323 = n2095 | n2142 ;
  assign n6324 = ~n1323 & n6323 ;
  assign n6325 = x87 & ~n6324 ;
  assign n6326 = ( x75 & ~n6322 ) | ( x75 & n6325 ) | ( ~n6322 & n6325 ) ;
  assign n6327 = n6322 | n6326 ;
  assign n6328 = x75 & ~n1323 ;
  assign n6329 = ( x92 & n6327 ) | ( x92 & ~n6328 ) | ( n6327 & ~n6328 ) ;
  assign n6330 = ~x92 & n6329 ;
  assign n6331 = n2142 | n2177 ;
  assign n6332 = ~n1323 & n6331 ;
  assign n6333 = x92 & ~n6332 ;
  assign n6334 = ( n2067 & ~n6330 ) | ( n2067 & n6333 ) | ( ~n6330 & n6333 ) ;
  assign n6335 = n6330 | n6334 ;
  assign n6336 = n2095 | n5009 ;
  assign n6337 = n2142 | n6336 ;
  assign n6338 = x74 | n6337 ;
  assign n6339 = ~n1323 & n6338 ;
  assign n6340 = ( x55 & x56 ) | ( x55 & ~n6339 ) | ( x56 & ~n6339 ) ;
  assign n6341 = n6339 ^ x56 ^ 1'b0 ;
  assign n6342 = ( x56 & n6340 ) | ( x56 & ~n6341 ) | ( n6340 & ~n6341 ) ;
  assign n6343 = ~n1323 & n2067 ;
  assign n6344 = x55 | n6343 ;
  assign n6345 = ~n6342 & n6344 ;
  assign n6346 = ( n6335 & n6342 ) | ( n6335 & ~n6345 ) | ( n6342 & ~n6345 ) ;
  assign n6347 = n2099 | n2142 ;
  assign n6348 = x56 & ~n1323 ;
  assign n6349 = n6347 & n6348 ;
  assign n6350 = ( x62 & n6346 ) | ( x62 & ~n6349 ) | ( n6346 & ~n6349 ) ;
  assign n6351 = ~x62 & n6350 ;
  assign n6352 = n2150 | n6323 ;
  assign n6353 = ~n1323 & n6352 ;
  assign n6354 = ~n6351 & n6353 ;
  assign n6355 = ( x62 & n6351 ) | ( x62 & ~n6354 ) | ( n6351 & ~n6354 ) ;
  assign n6356 = n2120 ^ n1323 ^ 1'b0 ;
  assign n6357 = ( n1323 & n6355 ) | ( n1323 & ~n6356 ) | ( n6355 & ~n6356 ) ;
  assign n6358 = x119 & x1056 ;
  assign n6359 = ~x228 & x252 ;
  assign n6360 = x119 | n6359 ;
  assign n6361 = ~x468 & n6360 ;
  assign n6362 = ~n6358 & n6361 ;
  assign n6363 = x119 & x1077 ;
  assign n6364 = n6361 & ~n6363 ;
  assign n6365 = x119 & x1073 ;
  assign n6366 = n6361 & ~n6365 ;
  assign n6367 = x119 & x1041 ;
  assign n6368 = n6361 & ~n6367 ;
  assign n6369 = x75 | n2095 ;
  assign n6370 = ~n1292 & n5023 ;
  assign n6371 = x87 & ~n6370 ;
  assign n6372 = n6369 | n6371 ;
  assign n6373 = n1410 | n5148 ;
  assign n6374 = x841 | n1373 ;
  assign n6375 = x90 & ~n6374 ;
  assign n6376 = x93 | n6375 ;
  assign n6377 = ~n6373 & n6376 ;
  assign n6378 = x51 | n6377 ;
  assign n6379 = x50 | x77 ;
  assign n6380 = x94 | n6379 ;
  assign n6381 = n1454 | n6380 ;
  assign n6382 = ~x88 & x98 ;
  assign n6383 = ~n1261 & n6382 ;
  assign n6384 = ~n6381 & n6383 ;
  assign n6385 = x97 | n6384 ;
  assign n6386 = ~n1395 & n6385 ;
  assign n6387 = x35 | n1374 ;
  assign n6388 = x70 | n6387 ;
  assign n6389 = n6386 & ~n6388 ;
  assign n6390 = ( ~n1434 & n6378 ) | ( ~n1434 & n6389 ) | ( n6378 & n6389 ) ;
  assign n6391 = ~n1434 & n6390 ;
  assign n6392 = x96 | n6391 ;
  assign n6393 = x96 & n5282 ;
  assign n6394 = n1290 | n6393 ;
  assign n6395 = ~x122 & x829 ;
  assign n6396 = n5020 & n6395 ;
  assign n6397 = ~n6394 & n6396 ;
  assign n6398 = n6392 & n6397 ;
  assign n6399 = x96 | n1290 ;
  assign n6400 = n6391 & ~n6399 ;
  assign n6401 = n5022 & n6400 ;
  assign n6402 = ~n6395 & n6401 ;
  assign n6403 = n6398 | n6402 ;
  assign n6404 = ~x1093 & n6403 ;
  assign n6405 = x87 | n6404 ;
  assign n6406 = n6405 ^ n6372 ^ 1'b0 ;
  assign n6407 = ( n6372 & n6405 ) | ( n6372 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6408 = ( x567 & ~n6372 ) | ( x567 & n6407 ) | ( ~n6372 & n6407 ) ;
  assign n6409 = ( x74 & ~n5015 ) | ( x74 & n6408 ) | ( ~n5015 & n6408 ) ;
  assign n6410 = ~x74 & n6409 ;
  assign n6411 = x232 & ~n5075 ;
  assign n6412 = ~n5040 & n6411 ;
  assign n6413 = n1207 | n6412 ;
  assign n6414 = ~x24 & n5415 ;
  assign n6415 = ~n1614 & n5035 ;
  assign n6416 = x1091 & n6415 ;
  assign n6417 = n6396 & n6416 ;
  assign n6418 = n6414 & n6417 ;
  assign n6419 = x1093 & n6418 ;
  assign n6420 = ~n6413 & n6419 ;
  assign n6421 = x75 & ~n6420 ;
  assign n6422 = x1093 & ~n1614 ;
  assign n6423 = n1434 | n6399 ;
  assign n6424 = n6378 & ~n6423 ;
  assign n6425 = x824 & n5020 ;
  assign n6426 = n6424 & n6425 ;
  assign n6427 = ~x829 & n6426 ;
  assign n6428 = ~x24 & n1443 ;
  assign n6429 = ~x46 & x97 ;
  assign n6430 = ~x108 & n6429 ;
  assign n6431 = ( ~n1459 & n5306 ) | ( ~n1459 & n6430 ) | ( n5306 & n6430 ) ;
  assign n6432 = ~n5306 & n6431 ;
  assign n6433 = ~x91 & n6432 ;
  assign n6434 = n6428 | n6433 ;
  assign n6435 = ( n1225 & ~n6373 ) | ( n1225 & n6434 ) | ( ~n6373 & n6434 ) ;
  assign n6436 = ~n1225 & n6435 ;
  assign n6437 = ( x51 & n6377 ) | ( x51 & ~n6436 ) | ( n6377 & ~n6436 ) ;
  assign n6438 = n6436 | n6437 ;
  assign n6439 = n6438 ^ n1434 ^ 1'b0 ;
  assign n6440 = ( n1434 & n6438 ) | ( n1434 & n6439 ) | ( n6438 & n6439 ) ;
  assign n6441 = ( x96 & ~n1434 ) | ( x96 & n6440 ) | ( ~n1434 & n6440 ) ;
  assign n6442 = x829 & n5020 ;
  assign n6443 = ~n6394 & n6442 ;
  assign n6444 = n6441 & n6443 ;
  assign n6445 = ( ~x122 & n6427 ) | ( ~x122 & n6444 ) | ( n6427 & n6444 ) ;
  assign n6446 = ~x122 & n6445 ;
  assign n6447 = x122 & n5022 ;
  assign n6448 = n6446 ^ n6424 ^ 1'b0 ;
  assign n6449 = ( ~n6424 & n6447 ) | ( ~n6424 & n6448 ) | ( n6447 & n6448 ) ;
  assign n6450 = ( n6424 & n6446 ) | ( n6424 & n6449 ) | ( n6446 & n6449 ) ;
  assign n6451 = x1091 & ~n6450 ;
  assign n6452 = ( x1091 & ~n6422 ) | ( x1091 & n6451 ) | ( ~n6422 & n6451 ) ;
  assign n6453 = ~n6404 & n6452 ;
  assign n6454 = x1091 | n6404 ;
  assign n6455 = ~n6453 & n6454 ;
  assign n6456 = x39 | n6455 ;
  assign n6457 = n1610 & ~n1614 ;
  assign n6458 = n5364 & n6457 ;
  assign n6459 = n1611 & n6458 ;
  assign n6460 = x1091 & n6459 ;
  assign n6461 = n5115 & n6460 ;
  assign n6462 = ~x299 & n5376 ;
  assign n6463 = ~x224 & n6462 ;
  assign n6464 = n6461 & n6463 ;
  assign n6465 = n5100 & n6460 ;
  assign n6466 = ~x216 & n5525 ;
  assign n6467 = n6465 & n6466 ;
  assign n6468 = x39 & ~n6467 ;
  assign n6469 = n6468 ^ n6464 ^ 1'b0 ;
  assign n6470 = ( n6464 & n6468 ) | ( n6464 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = ( x38 & ~n6464 ) | ( x38 & n6470 ) | ( ~n6464 & n6470 ) ;
  assign n6472 = ( x100 & n6456 ) | ( x100 & ~n6471 ) | ( n6456 & ~n6471 ) ;
  assign n6473 = n6472 ^ n6456 ^ 1'b0 ;
  assign n6474 = ( x100 & n6472 ) | ( x100 & ~n6473 ) | ( n6472 & ~n6473 ) ;
  assign n6475 = n5366 & n6424 ;
  assign n6476 = ( n6452 & ~n6471 ) | ( n6452 & n6475 ) | ( ~n6471 & n6475 ) ;
  assign n6477 = ~n6452 & n6476 ;
  assign n6478 = n6474 | n6477 ;
  assign n6479 = n1994 | n6412 ;
  assign n6480 = x1093 & n6396 ;
  assign n6481 = n6415 & n6480 ;
  assign n6482 = ~n1292 & n6481 ;
  assign n6483 = x1091 & n6482 ;
  assign n6484 = x228 & n6483 ;
  assign n6485 = x100 & ~n6484 ;
  assign n6486 = ( x100 & n6479 ) | ( x100 & n6485 ) | ( n6479 & n6485 ) ;
  assign n6487 = n6478 & ~n6486 ;
  assign n6488 = n6487 ^ x87 ^ 1'b0 ;
  assign n6489 = ~x1091 & x1093 ;
  assign n6490 = x1093 & n1614 ;
  assign n6491 = n5022 & ~n6490 ;
  assign n6492 = ~n1292 & n6491 ;
  assign n6493 = n6489 | n6492 ;
  assign n6494 = ~n2036 & n6493 ;
  assign n6495 = ~n1292 & n6425 ;
  assign n6496 = n6492 ^ n6489 ^ 1'b0 ;
  assign n6497 = ( n6492 & n6495 ) | ( n6492 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6498 = n6497 ^ n2036 ^ 1'b0 ;
  assign n6499 = ( n6494 & n6497 ) | ( n6494 & n6498 ) | ( n6497 & n6498 ) ;
  assign n6500 = ( n6487 & n6488 ) | ( n6487 & n6499 ) | ( n6488 & n6499 ) ;
  assign n6501 = x75 | n6500 ;
  assign n6502 = ~n6421 & n6501 ;
  assign n6503 = x567 & ~n6502 ;
  assign n6504 = n6410 & ~n6503 ;
  assign n6505 = x591 & n6504 ;
  assign n6506 = x353 ^ x352 ^ 1'b0 ;
  assign n6507 = n6506 ^ x462 ^ x360 ;
  assign n6508 = n6507 ^ x354 ^ 1'b0 ;
  assign n6509 = n6410 ^ x567 ^ 1'b0 ;
  assign n6510 = x1091 | n6370 ;
  assign n6511 = x1091 & ~n6492 ;
  assign n6512 = x87 & ~x100 ;
  assign n6513 = ~n1994 & n6512 ;
  assign n6514 = ~n6511 & n6513 ;
  assign n6515 = n6510 & n6514 ;
  assign n6516 = x75 | n6515 ;
  assign n6517 = x87 | n6486 ;
  assign n6518 = n6474 & ~n6517 ;
  assign n6519 = ( ~n6421 & n6516 ) | ( ~n6421 & n6518 ) | ( n6516 & n6518 ) ;
  assign n6520 = ~n6421 & n6519 ;
  assign n6521 = ( ~x567 & n6410 ) | ( ~x567 & n6520 ) | ( n6410 & n6520 ) ;
  assign n6522 = ( n6410 & n6509 ) | ( n6410 & n6521 ) | ( n6509 & n6521 ) ;
  assign n6523 = x592 & n6522 ;
  assign n6524 = ~x592 & n6504 ;
  assign n6525 = n6523 | n6524 ;
  assign n6526 = n6525 ^ n6522 ^ n6504 ;
  assign n6527 = x1199 & ~n6526 ;
  assign n6528 = x351 & n6527 ;
  assign n6529 = x351 & x1199 ;
  assign n6533 = x455 ^ x452 ^ 1'b0 ;
  assign n6534 = n6533 ^ x355 ^ 1'b0 ;
  assign n6530 = x460 ^ x342 ^ x320 ;
  assign n6531 = n6530 ^ x441 ^ x361 ;
  assign n6532 = n6531 ^ x458 ^ 1'b0 ;
  assign n6535 = n6534 ^ n6532 ^ 1'b0 ;
  assign n6536 = x1196 & n6535 ;
  assign n6537 = ~n6526 & n6536 ;
  assign n6538 = x1198 & ~n6537 ;
  assign n6539 = x1196 | n6504 ;
  assign n6540 = n6504 ^ x455 ^ 1'b0 ;
  assign n6541 = ( n6504 & n6526 ) | ( n6504 & ~n6540 ) | ( n6526 & ~n6540 ) ;
  assign n6542 = ( n6504 & n6526 ) | ( n6504 & n6540 ) | ( n6526 & n6540 ) ;
  assign n6543 = n6541 ^ x452 ^ 1'b0 ;
  assign n6544 = ( n6541 & n6542 ) | ( n6541 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6545 = ( n6541 & n6542 ) | ( n6541 & ~n6543 ) | ( n6542 & ~n6543 ) ;
  assign n6546 = n6544 ^ x355 ^ 1'b0 ;
  assign n6547 = ( n6544 & n6545 ) | ( n6544 & ~n6546 ) | ( n6545 & ~n6546 ) ;
  assign n6548 = x458 & ~n6547 ;
  assign n6549 = n6531 & ~n6548 ;
  assign n6550 = ( n6544 & n6545 ) | ( n6544 & n6546 ) | ( n6545 & n6546 ) ;
  assign n6551 = x458 | n6550 ;
  assign n6552 = n6549 & n6551 ;
  assign n6553 = x458 | n6547 ;
  assign n6554 = x458 & ~n6550 ;
  assign n6555 = ( n6531 & n6553 ) | ( n6531 & ~n6554 ) | ( n6553 & ~n6554 ) ;
  assign n6556 = ~n6531 & n6555 ;
  assign n6557 = ( x1196 & n6552 ) | ( x1196 & ~n6556 ) | ( n6552 & ~n6556 ) ;
  assign n6558 = ~n6552 & n6557 ;
  assign n6559 = ( x1198 & n6539 ) | ( x1198 & ~n6558 ) | ( n6539 & ~n6558 ) ;
  assign n6560 = ~x1198 & n6559 ;
  assign n6561 = x350 | x592 ;
  assign n6562 = ~n6504 & n6561 ;
  assign n6564 = x349 ^ x316 ^ 1'b0 ;
  assign n6563 = x359 ^ x322 ^ x315 ;
  assign n6565 = n6564 ^ n6563 ^ x348 ;
  assign n6566 = n6565 ^ x347 ^ x321 ;
  assign n6567 = n6522 | n6561 ;
  assign n6568 = n6566 & n6567 ;
  assign n6569 = ~n6562 & n6568 ;
  assign n6570 = x350 & ~x592 ;
  assign n6571 = ~n6522 & n6570 ;
  assign n6572 = n6566 | n6571 ;
  assign n6573 = n6504 | n6570 ;
  assign n6574 = ~n6572 & n6573 ;
  assign n6575 = ( n6536 & ~n6569 ) | ( n6536 & n6574 ) | ( ~n6569 & n6574 ) ;
  assign n6576 = n6569 | n6575 ;
  assign n6577 = n6560 ^ n6538 ^ 1'b0 ;
  assign n6578 = ( ~n6538 & n6576 ) | ( ~n6538 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6579 = ( n6538 & n6560 ) | ( n6538 & n6578 ) | ( n6560 & n6578 ) ;
  assign n6582 = x346 ^ x345 ^ x323 ;
  assign n6583 = n6582 ^ x450 ^ x358 ;
  assign n6580 = x344 ^ x343 ^ 1'b0 ;
  assign n6581 = n6580 ^ x362 ^ x327 ;
  assign n6584 = n6583 ^ n6581 ^ 1'b0 ;
  assign n6585 = x1197 & n6584 ;
  assign n6586 = n6585 ^ n6526 ^ 1'b0 ;
  assign n6587 = ( n6526 & n6579 ) | ( n6526 & ~n6586 ) | ( n6579 & ~n6586 ) ;
  assign n6588 = n6529 | n6587 ;
  assign n6589 = ~n6528 & n6588 ;
  assign n6590 = ~x351 & x1199 ;
  assign n6591 = n6587 | n6590 ;
  assign n6592 = ~x351 & n6527 ;
  assign n6593 = n6591 & ~n6592 ;
  assign n6594 = n6589 ^ x461 ^ 1'b0 ;
  assign n6595 = ( n6589 & n6593 ) | ( n6589 & n6594 ) | ( n6593 & n6594 ) ;
  assign n6596 = ( n6589 & n6593 ) | ( n6589 & ~n6594 ) | ( n6593 & ~n6594 ) ;
  assign n6597 = n6595 ^ x357 ^ 1'b0 ;
  assign n6598 = ( n6595 & n6596 ) | ( n6595 & n6597 ) | ( n6596 & n6597 ) ;
  assign n6599 = ( n6595 & n6596 ) | ( n6595 & ~n6597 ) | ( n6596 & ~n6597 ) ;
  assign n6600 = n6598 ^ x356 ^ 1'b0 ;
  assign n6601 = ( n6598 & n6599 ) | ( n6598 & ~n6600 ) | ( n6599 & ~n6600 ) ;
  assign n6602 = ( x591 & n6508 ) | ( x591 & ~n6601 ) | ( n6508 & ~n6601 ) ;
  assign n6603 = n6602 ^ n6508 ^ 1'b0 ;
  assign n6604 = ( x591 & n6602 ) | ( x591 & ~n6603 ) | ( n6602 & ~n6603 ) ;
  assign n6605 = ( n6598 & n6599 ) | ( n6598 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6606 = ( n6508 & ~n6604 ) | ( n6508 & n6605 ) | ( ~n6604 & n6605 ) ;
  assign n6607 = ~n6604 & n6606 ;
  assign n6608 = ( x590 & n6505 ) | ( x590 & ~n6607 ) | ( n6505 & ~n6607 ) ;
  assign n6609 = ~n6505 & n6608 ;
  assign n6610 = x285 | x286 ;
  assign n6611 = x289 | n6610 ;
  assign n6612 = x288 | n6611 ;
  assign n6616 = x372 ^ x363 ^ 1'b0 ;
  assign n6613 = x339 ^ x337 ^ 1'b0 ;
  assign n6614 = n6613 ^ x387 ^ x380 ;
  assign n6615 = n6614 ^ x388 ^ x338 ;
  assign n6617 = n6616 ^ n6615 ^ x386 ;
  assign n6622 = x389 ^ x368 ^ 1'b0 ;
  assign n6620 = x447 ^ x365 ^ 1'b0 ;
  assign n6618 = x366 ^ x364 ^ 1'b0 ;
  assign n6619 = n6618 ^ x383 ^ x336 ;
  assign n6621 = n6620 ^ n6619 ^ 1'b0 ;
  assign n6623 = n6622 ^ n6621 ^ x367 ;
  assign n6624 = x1197 & n6623 ;
  assign n6625 = n6624 ^ n6504 ^ 1'b0 ;
  assign n6626 = ( n6504 & n6525 ) | ( n6504 & n6625 ) | ( n6525 & n6625 ) ;
  assign n6627 = ~n6617 & n6626 ;
  assign n6628 = x1196 | n6624 ;
  assign n6629 = n6525 & n6628 ;
  assign n6630 = n6504 & ~n6624 ;
  assign n6631 = ~x1196 & n6630 ;
  assign n6632 = ( n6617 & n6629 ) | ( n6617 & n6631 ) | ( n6629 & n6631 ) ;
  assign n6633 = n6631 ^ n6629 ^ 1'b0 ;
  assign n6634 = ( n6617 & n6632 ) | ( n6617 & n6633 ) | ( n6632 & n6633 ) ;
  assign n6635 = ( x1199 & ~n6627 ) | ( x1199 & n6634 ) | ( ~n6627 & n6634 ) ;
  assign n6636 = n6627 | n6635 ;
  assign n6637 = x377 & x592 ;
  assign n6638 = n6504 | n6637 ;
  assign n6639 = ~x377 & x592 ;
  assign n6640 = n6504 | n6639 ;
  assign n6642 = x439 ^ x376 ^ 1'b0 ;
  assign n6641 = x385 ^ x378 ^ x317 ;
  assign n6643 = n6642 ^ n6641 ^ x381 ;
  assign n6644 = n6643 ^ x382 ^ x379 ;
  assign n6645 = ~n6522 & n6639 ;
  assign n6646 = n6644 & ~n6645 ;
  assign n6647 = n6640 & n6646 ;
  assign n6648 = ~n6522 & n6637 ;
  assign n6649 = n6644 | n6648 ;
  assign n6650 = ~n6647 & n6649 ;
  assign n6651 = ( n6638 & n6647 ) | ( n6638 & ~n6650 ) | ( n6647 & ~n6650 ) ;
  assign n6652 = x1196 & n6617 ;
  assign n6653 = n6624 | n6652 ;
  assign n6654 = n6653 ^ n6651 ^ 1'b0 ;
  assign n6655 = ( n6525 & n6651 ) | ( n6525 & n6654 ) | ( n6651 & n6654 ) ;
  assign n6656 = x1199 & ~n6655 ;
  assign n6657 = n6636 & ~n6656 ;
  assign n6658 = ~x1198 & x1199 ;
  assign n6659 = ~n6655 & n6658 ;
  assign n6660 = x1198 | n6636 ;
  assign n6661 = x1198 & ~n6525 ;
  assign n6662 = ( n6659 & n6660 ) | ( n6659 & ~n6661 ) | ( n6660 & ~n6661 ) ;
  assign n6663 = ~n6659 & n6662 ;
  assign n6664 = n6657 ^ x374 ^ 1'b0 ;
  assign n6665 = ( n6657 & n6663 ) | ( n6657 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = ( n6657 & n6663 ) | ( n6657 & ~n6664 ) | ( n6663 & ~n6664 ) ;
  assign n6667 = n6665 ^ x369 ^ 1'b0 ;
  assign n6668 = ( n6665 & n6666 ) | ( n6665 & n6667 ) | ( n6666 & n6667 ) ;
  assign n6669 = ( n6665 & n6666 ) | ( n6665 & ~n6667 ) | ( n6666 & ~n6667 ) ;
  assign n6670 = n6668 ^ x370 ^ 1'b0 ;
  assign n6671 = ( n6668 & n6669 ) | ( n6668 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6672 = ( n6668 & n6669 ) | ( n6668 & ~n6670 ) | ( n6669 & ~n6670 ) ;
  assign n6673 = n6671 ^ x371 ^ 1'b0 ;
  assign n6674 = ( n6671 & n6672 ) | ( n6671 & n6673 ) | ( n6672 & n6673 ) ;
  assign n6675 = ( n6671 & n6672 ) | ( n6671 & ~n6673 ) | ( n6672 & ~n6673 ) ;
  assign n6676 = n6674 ^ x373 ^ 1'b0 ;
  assign n6677 = ( n6674 & n6675 ) | ( n6674 & n6676 ) | ( n6675 & n6676 ) ;
  assign n6678 = ~x375 & n6677 ;
  assign n6679 = x442 ^ x440 ^ x384 ;
  assign n6680 = ( n6674 & n6675 ) | ( n6674 & ~n6676 ) | ( n6675 & ~n6676 ) ;
  assign n6681 = x375 & n6680 ;
  assign n6682 = ( ~n6678 & n6679 ) | ( ~n6678 & n6681 ) | ( n6679 & n6681 ) ;
  assign n6683 = n6678 | n6682 ;
  assign n6687 = x408 ^ x328 ^ 1'b0 ;
  assign n6686 = x396 ^ x394 ^ 1'b0 ;
  assign n6684 = x399 ^ x398 ^ x395 ;
  assign n6685 = n6684 ^ x400 ^ x329 ;
  assign n6688 = n6687 ^ n6686 ^ n6685 ;
  assign n6689 = x1198 & n6688 ;
  assign n6691 = x412 ^ x404 ^ x397 ;
  assign n6690 = x456 ^ x324 ^ x319 ;
  assign n6692 = n6691 ^ n6690 ^ 1'b0 ;
  assign n6693 = n6692 ^ x410 ^ x390 ;
  assign n6694 = n6693 ^ x411 ^ 1'b0 ;
  assign n6695 = n6495 & ~n6694 ;
  assign n6696 = n6489 & ~n6695 ;
  assign n6697 = n6493 & n6513 ;
  assign n6700 = x402 ^ x401 ^ 1'b0 ;
  assign n6698 = x326 ^ x325 ^ 1'b0 ;
  assign n6699 = n6698 ^ x405 ^ x403 ;
  assign n6701 = n6700 ^ n6699 ^ x406 ;
  assign n6702 = n6701 ^ x409 ^ x318 ;
  assign n6703 = n6495 & ~n6702 ;
  assign n6704 = n6489 & ~n6703 ;
  assign n6705 = n6697 & ~n6704 ;
  assign n6706 = ~n6696 & n6705 ;
  assign n6707 = x75 | x592 ;
  assign n6708 = x1199 & ~n6707 ;
  assign n6709 = ~x1196 & n6705 ;
  assign n6710 = ( n6706 & n6708 ) | ( n6706 & ~n6709 ) | ( n6708 & ~n6709 ) ;
  assign n6711 = ~n6706 & n6710 ;
  assign n6712 = n6711 ^ n6517 ^ 1'b0 ;
  assign n6713 = x1196 & n6694 ;
  assign n6714 = ~x75 & n6713 ;
  assign n6715 = ( n6477 & n6702 ) | ( n6477 & ~n6714 ) | ( n6702 & ~n6714 ) ;
  assign n6716 = ~n6702 & n6715 ;
  assign n6717 = n6474 | n6716 ;
  assign n6718 = ( n6517 & n6712 ) | ( n6517 & ~n6717 ) | ( n6712 & ~n6717 ) ;
  assign n6719 = ( n6711 & ~n6712 ) | ( n6711 & n6718 ) | ( ~n6712 & n6718 ) ;
  assign n6720 = ( ~n6502 & n6707 ) | ( ~n6502 & n6719 ) | ( n6707 & n6719 ) ;
  assign n6721 = n6719 ^ n6502 ^ 1'b0 ;
  assign n6722 = ( n6719 & n6720 ) | ( n6719 & ~n6721 ) | ( n6720 & ~n6721 ) ;
  assign n6723 = ~n6696 & n6697 ;
  assign n6724 = x1196 & ~n6707 ;
  assign n6725 = n6477 & ~n6694 ;
  assign n6726 = n6474 | n6725 ;
  assign n6727 = ~n6517 & n6726 ;
  assign n6728 = ( n6723 & n6724 ) | ( n6723 & ~n6727 ) | ( n6724 & ~n6727 ) ;
  assign n6729 = ~n6723 & n6728 ;
  assign n6730 = x1196 | n6501 ;
  assign n6731 = n6730 ^ n6729 ^ 1'b0 ;
  assign n6732 = ( n6729 & n6730 ) | ( n6729 & n6731 ) | ( n6730 & n6731 ) ;
  assign n6733 = ( x1199 & ~n6729 ) | ( x1199 & n6732 ) | ( ~n6729 & n6732 ) ;
  assign n6734 = x567 & ~n6733 ;
  assign n6735 = ( x567 & n6722 ) | ( x567 & n6734 ) | ( n6722 & n6734 ) ;
  assign n6736 = ( n6410 & n6689 ) | ( n6410 & ~n6735 ) | ( n6689 & ~n6735 ) ;
  assign n6737 = ~n6689 & n6736 ;
  assign n6738 = n6737 ^ n6526 ^ 1'b0 ;
  assign n6739 = ( ~n6526 & n6689 ) | ( ~n6526 & n6738 ) | ( n6689 & n6738 ) ;
  assign n6740 = ( n6526 & n6737 ) | ( n6526 & n6739 ) | ( n6737 & n6739 ) ;
  assign n6741 = n6526 ^ x1197 ^ 1'b0 ;
  assign n6742 = ( n6526 & n6740 ) | ( n6526 & ~n6741 ) | ( n6740 & ~n6741 ) ;
  assign n6743 = n6740 ^ x333 ^ 1'b0 ;
  assign n6744 = ( n6740 & n6742 ) | ( n6740 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6745 = ( n6740 & n6742 ) | ( n6740 & ~n6743 ) | ( n6742 & ~n6743 ) ;
  assign n6746 = n6744 ^ x391 ^ 1'b0 ;
  assign n6747 = ( n6744 & n6745 ) | ( n6744 & ~n6746 ) | ( n6745 & ~n6746 ) ;
  assign n6748 = ( n6744 & n6745 ) | ( n6744 & n6746 ) | ( n6745 & n6746 ) ;
  assign n6749 = n6747 ^ x392 ^ 1'b0 ;
  assign n6750 = ( n6747 & n6748 ) | ( n6747 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = ( n6747 & n6748 ) | ( n6747 & ~n6749 ) | ( n6748 & ~n6749 ) ;
  assign n6752 = n6750 ^ x393 ^ 1'b0 ;
  assign n6753 = ( n6750 & n6751 ) | ( n6750 & n6752 ) | ( n6751 & n6752 ) ;
  assign n6754 = x334 & n6753 ;
  assign n6755 = x413 ^ x335 ^ 1'b0 ;
  assign n6756 = n6755 ^ x463 ^ x407 ;
  assign n6757 = ( n6750 & n6751 ) | ( n6750 & ~n6752 ) | ( n6751 & ~n6752 ) ;
  assign n6758 = ~x334 & n6757 ;
  assign n6759 = ( ~n6754 & n6756 ) | ( ~n6754 & n6758 ) | ( n6756 & n6758 ) ;
  assign n6760 = n6754 | n6759 ;
  assign n6761 = n6760 ^ x590 ^ 1'b0 ;
  assign n6764 = x334 & n6757 ;
  assign n6762 = ~x334 & n6753 ;
  assign n6763 = n6756 & ~n6762 ;
  assign n6765 = n6764 ^ n6763 ^ 1'b0 ;
  assign n6766 = ( x591 & ~n6763 ) | ( x591 & n6764 ) | ( ~n6763 & n6764 ) ;
  assign n6767 = ( x591 & ~n6765 ) | ( x591 & n6766 ) | ( ~n6765 & n6766 ) ;
  assign n6768 = ( n6760 & ~n6761 ) | ( n6760 & n6767 ) | ( ~n6761 & n6767 ) ;
  assign n6769 = ( x590 & n6761 ) | ( x590 & n6768 ) | ( n6761 & n6768 ) ;
  assign n6770 = x375 & n6677 ;
  assign n6771 = ~x375 & n6680 ;
  assign n6772 = n6679 & ~n6771 ;
  assign n6773 = n6772 ^ n6770 ^ 1'b0 ;
  assign n6774 = ( n6770 & n6772 ) | ( n6770 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6775 = ( x591 & ~n6770 ) | ( x591 & n6774 ) | ( ~n6770 & n6774 ) ;
  assign n6776 = ~n6769 & n6775 ;
  assign n6777 = ( n6683 & n6769 ) | ( n6683 & ~n6776 ) | ( n6769 & ~n6776 ) ;
  assign n6778 = ( n6609 & ~n6612 ) | ( n6609 & n6777 ) | ( ~n6612 & n6777 ) ;
  assign n6779 = ~n6609 & n6778 ;
  assign n6780 = n6756 ^ x334 ^ 1'b0 ;
  assign n6781 = n6780 ^ x393 ^ 1'b0 ;
  assign n6782 = x74 | n5015 ;
  assign n6783 = ~x122 & x1093 ;
  assign n6784 = ~x98 & n6425 ;
  assign n6785 = n6783 & n6784 ;
  assign n6786 = ~x1091 & n6785 ;
  assign n6787 = x567 & n6786 ;
  assign n6788 = n6782 & n6787 ;
  assign n6844 = n6413 & n6786 ;
  assign n6845 = n6414 & n6481 ;
  assign n6846 = x1091 & ~n6845 ;
  assign n6847 = n6413 | n6846 ;
  assign n6848 = ( x1091 & n6786 ) | ( x1091 & ~n6847 ) | ( n6786 & ~n6847 ) ;
  assign n6849 = ( x75 & n6844 ) | ( x75 & ~n6848 ) | ( n6844 & ~n6848 ) ;
  assign n6850 = ~n6844 & n6849 ;
  assign n6789 = n6454 ^ x1093 ^ 1'b0 ;
  assign n6790 = x122 & n6426 ;
  assign n6791 = ~x122 & n6784 ;
  assign n6792 = n6790 | n6791 ;
  assign n6793 = ( x1093 & ~n6789 ) | ( x1093 & n6792 ) | ( ~n6789 & n6792 ) ;
  assign n6794 = ( n6454 & n6789 ) | ( n6454 & n6793 ) | ( n6789 & n6793 ) ;
  assign n6795 = ( x39 & ~n6453 ) | ( x39 & n6794 ) | ( ~n6453 & n6794 ) ;
  assign n6796 = ~x39 & n6795 ;
  assign n6797 = n6460 | n6786 ;
  assign n6798 = ~n5083 & n6460 ;
  assign n6799 = ( n6786 & n6797 ) | ( n6786 & n6798 ) | ( n6797 & n6798 ) ;
  assign n6800 = n5114 & ~n6799 ;
  assign n6801 = ~x223 & n4692 ;
  assign n6802 = ( n5099 & n6786 ) | ( n5099 & n6797 ) | ( n6786 & n6797 ) ;
  assign n6803 = n5114 | n6802 ;
  assign n6804 = ( n6800 & n6801 ) | ( n6800 & n6803 ) | ( n6801 & n6803 ) ;
  assign n6805 = ~n6800 & n6804 ;
  assign n6806 = n6786 & ~n6801 ;
  assign n6807 = ( x299 & ~n6805 ) | ( x299 & n6806 ) | ( ~n6805 & n6806 ) ;
  assign n6808 = n6805 | n6807 ;
  assign n6809 = n5061 & ~n6799 ;
  assign n6810 = ~x216 & n5390 ;
  assign n6811 = n5061 | n6802 ;
  assign n6812 = ( n6809 & n6810 ) | ( n6809 & n6811 ) | ( n6810 & n6811 ) ;
  assign n6813 = ~n6809 & n6812 ;
  assign n6814 = n6786 & ~n6810 ;
  assign n6815 = ( x299 & n6813 ) | ( x299 & ~n6814 ) | ( n6813 & ~n6814 ) ;
  assign n6816 = ~n6813 & n6815 ;
  assign n6817 = x39 & ~n6816 ;
  assign n6818 = n6808 & n6817 ;
  assign n6819 = ( ~x38 & n6796 ) | ( ~x38 & n6818 ) | ( n6796 & n6818 ) ;
  assign n6820 = ~x38 & n6819 ;
  assign n6821 = x38 & n6786 ;
  assign n6822 = ( x100 & ~n6820 ) | ( x100 & n6821 ) | ( ~n6820 & n6821 ) ;
  assign n6823 = n6820 | n6822 ;
  assign n6824 = x228 & ~n6412 ;
  assign n6825 = n6786 | n6824 ;
  assign n6826 = n6483 | n6786 ;
  assign n6827 = n6824 & ~n6826 ;
  assign n6828 = ( n1994 & n6825 ) | ( n1994 & ~n6827 ) | ( n6825 & ~n6827 ) ;
  assign n6829 = ~n1994 & n6828 ;
  assign n6830 = n1994 & n6786 ;
  assign n6831 = ( x100 & n6829 ) | ( x100 & ~n6830 ) | ( n6829 & ~n6830 ) ;
  assign n6832 = ~n6829 & n6831 ;
  assign n6833 = ( x87 & n6823 ) | ( x87 & ~n6832 ) | ( n6823 & ~n6832 ) ;
  assign n6834 = ~x87 & n6833 ;
  assign n6835 = x122 & n6495 ;
  assign n6836 = ( x1093 & n6785 ) | ( x1093 & n6835 ) | ( n6785 & n6835 ) ;
  assign n6837 = n6510 | n6836 ;
  assign n6838 = ( n2036 & ~n6511 ) | ( n2036 & n6837 ) | ( ~n6511 & n6837 ) ;
  assign n6839 = ~n2036 & n6838 ;
  assign n6840 = n6786 | n6839 ;
  assign n6841 = x87 & n6840 ;
  assign n6842 = ( x75 & ~n6834 ) | ( x75 & n6841 ) | ( ~n6834 & n6841 ) ;
  assign n6843 = n6834 | n6842 ;
  assign n6851 = n6850 ^ n6843 ^ 1'b0 ;
  assign n6852 = ( x567 & ~n6843 ) | ( x567 & n6850 ) | ( ~n6843 & n6850 ) ;
  assign n6853 = ( x567 & ~n6851 ) | ( x567 & n6852 ) | ( ~n6851 & n6852 ) ;
  assign n6854 = ~n6788 & n6853 ;
  assign n6855 = ( n6410 & n6788 ) | ( n6410 & ~n6854 ) | ( n6788 & ~n6854 ) ;
  assign n6856 = x592 & ~n6855 ;
  assign n6857 = x1196 | n6855 ;
  assign n6858 = ~n6694 & n6785 ;
  assign n6859 = ~x1091 & n6858 ;
  assign n6860 = x567 & n6859 ;
  assign n6861 = n6782 & n6860 ;
  assign n6862 = ~x592 & x1196 ;
  assign n6863 = x38 & n6859 ;
  assign n6864 = x100 | n6863 ;
  assign n6865 = n6798 | n6859 ;
  assign n6866 = n5061 & ~n6865 ;
  assign n6867 = n5099 & n6460 ;
  assign n6868 = n6859 | n6867 ;
  assign n6869 = n5061 | n6868 ;
  assign n6870 = ( n6810 & n6866 ) | ( n6810 & n6869 ) | ( n6866 & n6869 ) ;
  assign n6871 = ~n6866 & n6870 ;
  assign n6872 = ~n6810 & n6859 ;
  assign n6873 = x299 & ~n6872 ;
  assign n6874 = x39 & ~n6873 ;
  assign n6875 = ( x39 & n6871 ) | ( x39 & n6874 ) | ( n6871 & n6874 ) ;
  assign n6880 = ~n6801 & n6859 ;
  assign n6881 = x299 | n6880 ;
  assign n6876 = n5114 & ~n6865 ;
  assign n6877 = n5114 | n6868 ;
  assign n6878 = ( n6801 & n6876 ) | ( n6801 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6879 = ~n6876 & n6878 ;
  assign n6882 = n6881 ^ n6879 ^ 1'b0 ;
  assign n6883 = ( n6879 & n6881 ) | ( n6879 & ~n6882 ) | ( n6881 & ~n6882 ) ;
  assign n6884 = ( n6875 & n6882 ) | ( n6875 & n6883 ) | ( n6882 & n6883 ) ;
  assign n6885 = ~n6454 & n6694 ;
  assign n6886 = ~n6884 & n6885 ;
  assign n6887 = ( n6796 & n6884 ) | ( n6796 & ~n6886 ) | ( n6884 & ~n6886 ) ;
  assign n6888 = x38 | n6887 ;
  assign n6889 = ( ~x38 & n6864 ) | ( ~x38 & n6888 ) | ( n6864 & n6888 ) ;
  assign n6890 = n6486 & ~n6859 ;
  assign n6891 = ( x87 & n6889 ) | ( x87 & ~n6890 ) | ( n6889 & ~n6890 ) ;
  assign n6892 = n6891 ^ n6889 ^ 1'b0 ;
  assign n6893 = ( x87 & n6891 ) | ( x87 & ~n6892 ) | ( n6891 & ~n6892 ) ;
  assign n6894 = n2036 & n6859 ;
  assign n6895 = x87 & ~n6894 ;
  assign n6896 = ~n6510 & n6694 ;
  assign n6897 = n6839 & ~n6896 ;
  assign n6898 = n6895 & ~n6897 ;
  assign n6899 = ( x75 & n6893 ) | ( x75 & ~n6898 ) | ( n6893 & ~n6898 ) ;
  assign n6900 = n6899 ^ n6893 ^ 1'b0 ;
  assign n6901 = ( x75 & n6899 ) | ( x75 & ~n6900 ) | ( n6899 & ~n6900 ) ;
  assign n6902 = n6413 & n6859 ;
  assign n6903 = x75 & ~n6902 ;
  assign n6904 = ( x1091 & ~n6847 ) | ( x1091 & n6859 ) | ( ~n6847 & n6859 ) ;
  assign n6905 = ( n6901 & ~n6903 ) | ( n6901 & n6904 ) | ( ~n6903 & n6904 ) ;
  assign n6906 = n6903 ^ n6901 ^ 1'b0 ;
  assign n6907 = ( n6901 & n6905 ) | ( n6901 & n6906 ) | ( n6905 & n6906 ) ;
  assign n6908 = ( ~x567 & n6410 ) | ( ~x567 & n6907 ) | ( n6410 & n6907 ) ;
  assign n6909 = ( n6410 & n6509 ) | ( n6410 & n6908 ) | ( n6509 & n6908 ) ;
  assign n6910 = ( n6861 & n6862 ) | ( n6861 & ~n6909 ) | ( n6862 & ~n6909 ) ;
  assign n6911 = ~n6861 & n6910 ;
  assign n6912 = ( x1199 & n6857 ) | ( x1199 & ~n6911 ) | ( n6857 & ~n6911 ) ;
  assign n6913 = ~x1199 & n6912 ;
  assign n6914 = ~n6702 & n6784 ;
  assign n6915 = n6861 & n6914 ;
  assign n6916 = n6862 & ~n6915 ;
  assign n6917 = x592 | x1196 ;
  assign n6918 = ~n6702 & n6785 ;
  assign n6919 = ~x1091 & n6918 ;
  assign n6920 = x567 & n6919 ;
  assign n6921 = n6782 & n6920 ;
  assign n6922 = n6917 | n6921 ;
  assign n6923 = ~n6916 & n6922 ;
  assign n6924 = n6410 | n6923 ;
  assign n6978 = ~n6702 & n6859 ;
  assign n6979 = n6867 | n6978 ;
  assign n6980 = n5061 | n6979 ;
  assign n6981 = n6798 | n6978 ;
  assign n6982 = n5061 & ~n6981 ;
  assign n6983 = n6810 & ~n6982 ;
  assign n6984 = n6980 & n6983 ;
  assign n6933 = ~n6810 & n6919 ;
  assign n6934 = x299 & ~n6933 ;
  assign n6985 = ( n6873 & n6934 ) | ( n6873 & ~n6984 ) | ( n6934 & ~n6984 ) ;
  assign n6986 = ~n6984 & n6985 ;
  assign n6987 = n5114 | n6979 ;
  assign n6988 = n5114 & ~n6981 ;
  assign n6989 = n6801 & ~n6988 ;
  assign n6990 = n6987 & n6989 ;
  assign n6946 = ~n6801 & n6919 ;
  assign n6991 = x299 | n6946 ;
  assign n6992 = n6990 ^ n6881 ^ 1'b0 ;
  assign n6993 = ( ~n6881 & n6991 ) | ( ~n6881 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6994 = ( n6881 & n6990 ) | ( n6881 & n6993 ) | ( n6990 & n6993 ) ;
  assign n6995 = ( x39 & n6986 ) | ( x39 & n6994 ) | ( n6986 & n6994 ) ;
  assign n6996 = ~n6986 & n6995 ;
  assign n6951 = x122 | n6914 ;
  assign n6952 = n6426 & ~n6702 ;
  assign n6953 = x122 & ~n6952 ;
  assign n6954 = x1093 & ~n6953 ;
  assign n6955 = n6951 & n6954 ;
  assign n6956 = ( x1091 & n6404 ) | ( x1091 & ~n6955 ) | ( n6404 & ~n6955 ) ;
  assign n6957 = n6955 | n6956 ;
  assign n6997 = n6796 & ~n6885 ;
  assign n6998 = n6957 & n6997 ;
  assign n6999 = ( ~x38 & n6996 ) | ( ~x38 & n6998 ) | ( n6996 & n6998 ) ;
  assign n7000 = ~x38 & n6999 ;
  assign n6931 = x38 & n6919 ;
  assign n6932 = x100 | n6931 ;
  assign n7001 = n7000 ^ n6864 ^ 1'b0 ;
  assign n7002 = ( ~n6864 & n6932 ) | ( ~n6864 & n7001 ) | ( n6932 & n7001 ) ;
  assign n7003 = ( n6864 & n7000 ) | ( n6864 & n7002 ) | ( n7000 & n7002 ) ;
  assign n7004 = n5038 & n6483 ;
  assign n7005 = x1091 & ~n6482 ;
  assign n7006 = x1091 | n6978 ;
  assign n7007 = ( ~n5038 & n5039 ) | ( ~n5038 & n5075 ) | ( n5039 & n5075 ) ;
  assign n7008 = n7006 & n7007 ;
  assign n7009 = ~n7005 & n7008 ;
  assign n7010 = ( x228 & n7004 ) | ( x228 & n7009 ) | ( n7004 & n7009 ) ;
  assign n7011 = n7009 ^ n7004 ^ 1'b0 ;
  assign n7012 = ( x228 & n7010 ) | ( x228 & n7011 ) | ( n7010 & n7011 ) ;
  assign n7013 = x228 & n7007 ;
  assign n7014 = n6978 & ~n7013 ;
  assign n7015 = ( x232 & n7012 ) | ( x232 & ~n7014 ) | ( n7012 & ~n7014 ) ;
  assign n7016 = ~n7012 & n7015 ;
  assign n7017 = x232 | n6978 ;
  assign n7018 = n6484 | n7017 ;
  assign n7019 = ( n1994 & ~n7016 ) | ( n1994 & n7018 ) | ( ~n7016 & n7018 ) ;
  assign n7020 = ~n1994 & n7019 ;
  assign n7021 = n1994 & n6978 ;
  assign n7022 = ( x100 & n7020 ) | ( x100 & ~n7021 ) | ( n7020 & ~n7021 ) ;
  assign n7023 = ~n7020 & n7022 ;
  assign n7024 = ( x87 & n7003 ) | ( x87 & ~n7023 ) | ( n7003 & ~n7023 ) ;
  assign n7025 = n7024 ^ n7003 ^ 1'b0 ;
  assign n7026 = ( x87 & n7024 ) | ( x87 & ~n7025 ) | ( n7024 & ~n7025 ) ;
  assign n6925 = ~n6510 & n6702 ;
  assign n6926 = n6839 & ~n6925 ;
  assign n7027 = ~n6896 & n6926 ;
  assign n6927 = n2036 & n6919 ;
  assign n6928 = x87 & ~n6927 ;
  assign n7028 = n6895 | n6928 ;
  assign n7029 = ~n7027 & n7028 ;
  assign n7030 = ( x75 & n7026 ) | ( x75 & ~n7029 ) | ( n7026 & ~n7029 ) ;
  assign n7031 = n7030 ^ n7026 ^ 1'b0 ;
  assign n7032 = ( x75 & n7030 ) | ( x75 & ~n7031 ) | ( n7030 & ~n7031 ) ;
  assign n7033 = ~n6847 & n7006 ;
  assign n6970 = n6413 & n6919 ;
  assign n6971 = x75 & ~n6970 ;
  assign n7034 = n6903 | n6971 ;
  assign n7035 = n7032 & ~n7034 ;
  assign n7036 = ( n7032 & n7033 ) | ( n7032 & n7035 ) | ( n7033 & n7035 ) ;
  assign n7037 = ( n6862 & n6915 ) | ( n6862 & ~n7036 ) | ( n6915 & ~n7036 ) ;
  assign n7038 = ~n6915 & n7037 ;
  assign n6929 = ~n6926 & n6928 ;
  assign n6930 = n6486 & ~n6919 ;
  assign n6935 = n6867 | n6919 ;
  assign n6936 = n5061 | n6935 ;
  assign n6937 = n6798 | n6919 ;
  assign n6938 = n5061 & ~n6937 ;
  assign n6939 = n6810 & ~n6938 ;
  assign n6940 = n6934 & ~n6939 ;
  assign n6941 = ( n6934 & ~n6936 ) | ( n6934 & n6940 ) | ( ~n6936 & n6940 ) ;
  assign n6942 = n5114 & ~n6937 ;
  assign n6943 = n5114 | n6935 ;
  assign n6944 = ( n6801 & n6942 ) | ( n6801 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6945 = ~n6942 & n6944 ;
  assign n6947 = ( x299 & ~n6945 ) | ( x299 & n6946 ) | ( ~n6945 & n6946 ) ;
  assign n6948 = n6945 | n6947 ;
  assign n6949 = ( x39 & n6941 ) | ( x39 & n6948 ) | ( n6941 & n6948 ) ;
  assign n6950 = ~n6941 & n6949 ;
  assign n6958 = x39 | n6453 ;
  assign n6959 = ( n6950 & n6957 ) | ( n6950 & ~n6958 ) | ( n6957 & ~n6958 ) ;
  assign n6960 = n6958 ^ n6950 ^ 1'b0 ;
  assign n6961 = ( n6950 & n6959 ) | ( n6950 & ~n6960 ) | ( n6959 & ~n6960 ) ;
  assign n6962 = x38 | n6961 ;
  assign n6963 = ( ~x38 & n6932 ) | ( ~x38 & n6962 ) | ( n6932 & n6962 ) ;
  assign n6964 = n6963 ^ n6930 ^ 1'b0 ;
  assign n6965 = ( n6930 & n6963 ) | ( n6930 & n6964 ) | ( n6963 & n6964 ) ;
  assign n6966 = ( x87 & ~n6930 ) | ( x87 & n6965 ) | ( ~n6930 & n6965 ) ;
  assign n6967 = n6966 ^ n6929 ^ 1'b0 ;
  assign n6968 = ( n6929 & n6966 ) | ( n6929 & n6967 ) | ( n6966 & n6967 ) ;
  assign n6969 = ( x75 & ~n6929 ) | ( x75 & n6968 ) | ( ~n6929 & n6968 ) ;
  assign n6972 = ( x1091 & ~n6847 ) | ( x1091 & n6919 ) | ( ~n6847 & n6919 ) ;
  assign n6973 = ( n6969 & ~n6971 ) | ( n6969 & n6972 ) | ( ~n6971 & n6972 ) ;
  assign n6974 = n6971 ^ n6969 ^ 1'b0 ;
  assign n6975 = ( n6969 & n6973 ) | ( n6969 & n6974 ) | ( n6973 & n6974 ) ;
  assign n6976 = ( n6917 & n6921 ) | ( n6917 & ~n6975 ) | ( n6921 & ~n6975 ) ;
  assign n6977 = n6975 | n6976 ;
  assign n7039 = n7038 ^ n6977 ^ 1'b0 ;
  assign n7040 = ( x567 & ~n6977 ) | ( x567 & n7038 ) | ( ~n6977 & n7038 ) ;
  assign n7041 = ( x567 & ~n7039 ) | ( x567 & n7040 ) | ( ~n7039 & n7040 ) ;
  assign n7042 = x1199 & ~n7041 ;
  assign n7043 = n6924 & n7042 ;
  assign n7044 = ( n6689 & ~n6913 ) | ( n6689 & n7043 ) | ( ~n6913 & n7043 ) ;
  assign n7045 = n6913 | n7044 ;
  assign n7046 = x592 | n6522 ;
  assign n7047 = n6689 & ~n7046 ;
  assign n7048 = ( n6856 & n7045 ) | ( n6856 & ~n7047 ) | ( n7045 & ~n7047 ) ;
  assign n7049 = ~n6856 & n7048 ;
  assign n7050 = ~x592 & n6855 ;
  assign n7051 = n6523 | n7050 ;
  assign n7052 = n7051 ^ n6855 ^ n6522 ;
  assign n7053 = n7052 ^ x1197 ^ 1'b0 ;
  assign n7054 = ( n7049 & n7052 ) | ( n7049 & ~n7053 ) | ( n7052 & ~n7053 ) ;
  assign n7055 = n7049 ^ x333 ^ 1'b0 ;
  assign n7056 = ( n7049 & n7054 ) | ( n7049 & n7055 ) | ( n7054 & n7055 ) ;
  assign n7057 = ( n7049 & n7054 ) | ( n7049 & ~n7055 ) | ( n7054 & ~n7055 ) ;
  assign n7058 = n7056 ^ x391 ^ 1'b0 ;
  assign n7059 = ( n7056 & n7057 ) | ( n7056 & n7058 ) | ( n7057 & n7058 ) ;
  assign n7060 = ( n7056 & n7057 ) | ( n7056 & ~n7058 ) | ( n7057 & ~n7058 ) ;
  assign n7061 = n7059 ^ x392 ^ 1'b0 ;
  assign n7062 = ( n7059 & n7060 ) | ( n7059 & ~n7061 ) | ( n7060 & ~n7061 ) ;
  assign n7063 = n6781 & ~n7062 ;
  assign n7064 = ( n7059 & n7060 ) | ( n7059 & n7061 ) | ( n7060 & n7061 ) ;
  assign n7065 = n6781 | n7064 ;
  assign n7066 = ( x591 & n7063 ) | ( x591 & n7065 ) | ( n7063 & n7065 ) ;
  assign n7067 = ~n7063 & n7066 ;
  assign n7068 = n6679 ^ x375 ^ x373 ;
  assign n7069 = n6653 & n7051 ;
  assign n7070 = n6639 | n6855 ;
  assign n7071 = n6646 & n7070 ;
  assign n7072 = n6637 | n6855 ;
  assign n7073 = ~n6649 & n7072 ;
  assign n7074 = ( ~n6653 & n7071 ) | ( ~n6653 & n7073 ) | ( n7071 & n7073 ) ;
  assign n7075 = ~n6653 & n7074 ;
  assign n7076 = ( x1199 & n7069 ) | ( x1199 & ~n7075 ) | ( n7069 & ~n7075 ) ;
  assign n7077 = ~n7069 & n7076 ;
  assign n7078 = ~n6653 & n6855 ;
  assign n7079 = x1199 | n7078 ;
  assign n7080 = ( n7069 & ~n7077 ) | ( n7069 & n7079 ) | ( ~n7077 & n7079 ) ;
  assign n7081 = ~n7077 & n7080 ;
  assign n7082 = n7051 ^ x1198 ^ 1'b0 ;
  assign n7083 = ( n7051 & n7081 ) | ( n7051 & ~n7082 ) | ( n7081 & ~n7082 ) ;
  assign n7084 = n7081 ^ x374 ^ 1'b0 ;
  assign n7085 = ( n7081 & n7083 ) | ( n7081 & n7084 ) | ( n7083 & n7084 ) ;
  assign n7086 = ( n7081 & n7083 ) | ( n7081 & ~n7084 ) | ( n7083 & ~n7084 ) ;
  assign n7087 = n7085 ^ x369 ^ 1'b0 ;
  assign n7088 = ( n7085 & n7086 ) | ( n7085 & n7087 ) | ( n7086 & n7087 ) ;
  assign n7089 = ( n7085 & n7086 ) | ( n7085 & ~n7087 ) | ( n7086 & ~n7087 ) ;
  assign n7090 = n7088 ^ x370 ^ 1'b0 ;
  assign n7091 = ( n7088 & n7089 ) | ( n7088 & n7090 ) | ( n7089 & n7090 ) ;
  assign n7092 = ( n7088 & n7089 ) | ( n7088 & ~n7090 ) | ( n7089 & ~n7090 ) ;
  assign n7093 = n7091 ^ x371 ^ 1'b0 ;
  assign n7094 = ( n7091 & n7092 ) | ( n7091 & ~n7093 ) | ( n7092 & ~n7093 ) ;
  assign n7095 = ( x591 & n7068 ) | ( x591 & ~n7094 ) | ( n7068 & ~n7094 ) ;
  assign n7096 = n7095 ^ n7068 ^ 1'b0 ;
  assign n7097 = ( x591 & n7095 ) | ( x591 & ~n7096 ) | ( n7095 & ~n7096 ) ;
  assign n7098 = ( n7091 & n7092 ) | ( n7091 & n7093 ) | ( n7092 & n7093 ) ;
  assign n7099 = ( n7068 & ~n7097 ) | ( n7068 & n7098 ) | ( ~n7097 & n7098 ) ;
  assign n7100 = ~n7097 & n7099 ;
  assign n7101 = ( x590 & ~n7067 ) | ( x590 & n7100 ) | ( ~n7067 & n7100 ) ;
  assign n7102 = n7067 | n7101 ;
  assign n7103 = x591 & n6855 ;
  assign n7104 = x1199 & ~n7052 ;
  assign n7105 = x351 & n7104 ;
  assign n7106 = n6536 & ~n7052 ;
  assign n7107 = x1198 & ~n7106 ;
  assign n7108 = n6570 | n6855 ;
  assign n7109 = n6572 | n7108 ;
  assign n7110 = ( n6536 & ~n6572 ) | ( n6536 & n7109 ) | ( ~n6572 & n7109 ) ;
  assign n7111 = n6561 & ~n6855 ;
  assign n7112 = ~n7110 & n7111 ;
  assign n7113 = ( n6568 & n7110 ) | ( n6568 & ~n7112 ) | ( n7110 & ~n7112 ) ;
  assign n7114 = n7107 & n7113 ;
  assign n7115 = n6855 ^ x455 ^ 1'b0 ;
  assign n7116 = ( n6855 & n7052 ) | ( n6855 & n7115 ) | ( n7052 & n7115 ) ;
  assign n7117 = x452 & ~n7116 ;
  assign n7118 = n6532 ^ x355 ^ 1'b0 ;
  assign n7119 = ( n6855 & n7052 ) | ( n6855 & ~n7115 ) | ( n7052 & ~n7115 ) ;
  assign n7120 = x452 | n7119 ;
  assign n7121 = ( n7117 & n7118 ) | ( n7117 & n7120 ) | ( n7118 & n7120 ) ;
  assign n7122 = ~n7117 & n7121 ;
  assign n7123 = x452 & ~n7119 ;
  assign n7124 = x452 | n7116 ;
  assign n7125 = ( n7118 & ~n7123 ) | ( n7118 & n7124 ) | ( ~n7123 & n7124 ) ;
  assign n7126 = ~n7118 & n7125 ;
  assign n7127 = ( x1196 & n7122 ) | ( x1196 & ~n7126 ) | ( n7122 & ~n7126 ) ;
  assign n7128 = ~n7122 & n7127 ;
  assign n7129 = ( x1198 & n6857 ) | ( x1198 & ~n7128 ) | ( n6857 & ~n7128 ) ;
  assign n7130 = ~x1198 & n7129 ;
  assign n7131 = ( n6585 & ~n7114 ) | ( n6585 & n7130 ) | ( ~n7114 & n7130 ) ;
  assign n7132 = n7114 | n7131 ;
  assign n7133 = n7132 ^ n7052 ^ 1'b0 ;
  assign n7134 = ( ~n6585 & n7052 ) | ( ~n6585 & n7133 ) | ( n7052 & n7133 ) ;
  assign n7135 = ( n7132 & ~n7133 ) | ( n7132 & n7134 ) | ( ~n7133 & n7134 ) ;
  assign n7136 = n6529 | n7135 ;
  assign n7137 = ~n7105 & n7136 ;
  assign n7138 = ~x351 & n7104 ;
  assign n7139 = n6590 | n7135 ;
  assign n7140 = ~n7138 & n7139 ;
  assign n7141 = n7137 ^ x461 ^ 1'b0 ;
  assign n7142 = ( n7137 & n7140 ) | ( n7137 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7143 = ( n7137 & n7140 ) | ( n7137 & ~n7141 ) | ( n7140 & ~n7141 ) ;
  assign n7144 = n7142 ^ x357 ^ 1'b0 ;
  assign n7145 = ( n7142 & n7143 ) | ( n7142 & n7144 ) | ( n7143 & n7144 ) ;
  assign n7146 = ( n7142 & n7143 ) | ( n7142 & ~n7144 ) | ( n7143 & ~n7144 ) ;
  assign n7147 = n7145 ^ x356 ^ 1'b0 ;
  assign n7148 = ( n7145 & n7146 ) | ( n7145 & ~n7147 ) | ( n7146 & ~n7147 ) ;
  assign n7149 = ( x591 & n6508 ) | ( x591 & ~n7148 ) | ( n6508 & ~n7148 ) ;
  assign n7150 = n7149 ^ n6508 ^ 1'b0 ;
  assign n7151 = ( x591 & n7149 ) | ( x591 & ~n7150 ) | ( n7149 & ~n7150 ) ;
  assign n7152 = ( n7145 & n7146 ) | ( n7145 & n7147 ) | ( n7146 & n7147 ) ;
  assign n7153 = ( n6508 & ~n7151 ) | ( n6508 & n7152 ) | ( ~n7151 & n7152 ) ;
  assign n7154 = ~n7151 & n7153 ;
  assign n7155 = ( x590 & n7103 ) | ( x590 & ~n7154 ) | ( n7103 & ~n7154 ) ;
  assign n7156 = ~n7103 & n7155 ;
  assign n7157 = n6612 & ~n7156 ;
  assign n7158 = n7102 & n7157 ;
  assign n7159 = ( x588 & ~n6779 ) | ( x588 & n7158 ) | ( ~n6779 & n7158 ) ;
  assign n7160 = n6779 | n7159 ;
  assign n7161 = x592 & n6787 ;
  assign n7162 = x1199 & ~n7161 ;
  assign n7163 = ~x351 & n7162 ;
  assign n7164 = ~x592 & n6535 ;
  assign n7165 = ~n6530 & n6787 ;
  assign n7166 = ~n7164 & n7165 ;
  assign n7167 = n6534 ^ x458 ^ x361 ;
  assign n7168 = ~x441 & n7167 ;
  assign n7169 = x592 | n7168 ;
  assign n7170 = n7167 & ~n7169 ;
  assign n7171 = ( x441 & n7169 ) | ( x441 & ~n7170 ) | ( n7169 & ~n7170 ) ;
  assign n7172 = n6530 & n6787 ;
  assign n7173 = x1196 & ~n7172 ;
  assign n7174 = ( x1196 & ~n7171 ) | ( x1196 & n7173 ) | ( ~n7171 & n7173 ) ;
  assign n7175 = n7174 ^ n7166 ^ 1'b0 ;
  assign n7176 = ( n7166 & n7174 ) | ( n7166 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7177 = ( x1198 & ~n7166 ) | ( x1198 & n7176 ) | ( ~n7166 & n7176 ) ;
  assign n7178 = n6566 ^ x350 ^ 1'b0 ;
  assign n7179 = n6536 | n7178 ;
  assign n7180 = ~x592 & n6787 ;
  assign n7181 = x1198 & n7180 ;
  assign n7182 = ~n7179 & n7181 ;
  assign n7183 = ( n6585 & n7177 ) | ( n6585 & ~n7182 ) | ( n7177 & ~n7182 ) ;
  assign n7184 = n7183 ^ n7177 ^ 1'b0 ;
  assign n7185 = ( n6585 & n7183 ) | ( n6585 & ~n7184 ) | ( n7183 & ~n7184 ) ;
  assign n7186 = ~x592 & n7185 ;
  assign n7187 = n6787 & ~n7186 ;
  assign n7188 = n6590 | n7187 ;
  assign n7189 = ~n7163 & n7188 ;
  assign n7190 = x351 & n7162 ;
  assign n7191 = n6529 | n7187 ;
  assign n7192 = ~n7190 & n7191 ;
  assign n7193 = n7189 ^ x461 ^ 1'b0 ;
  assign n7194 = ( n7189 & n7192 ) | ( n7189 & n7193 ) | ( n7192 & n7193 ) ;
  assign n7195 = ( n7189 & n7192 ) | ( n7189 & ~n7193 ) | ( n7192 & ~n7193 ) ;
  assign n7196 = n7194 ^ x357 ^ 1'b0 ;
  assign n7197 = ( n7194 & n7195 ) | ( n7194 & n7196 ) | ( n7195 & n7196 ) ;
  assign n7198 = x356 | n7197 ;
  assign n7199 = ( n7194 & n7195 ) | ( n7194 & ~n7196 ) | ( n7195 & ~n7196 ) ;
  assign n7200 = x356 & ~n7199 ;
  assign n7201 = n6508 & ~n7200 ;
  assign n7202 = n7198 & n7201 ;
  assign n7203 = x356 & ~n7197 ;
  assign n7204 = x356 | n7199 ;
  assign n7205 = ( n6508 & ~n7203 ) | ( n6508 & n7204 ) | ( ~n7203 & n7204 ) ;
  assign n7206 = ~n6508 & n7205 ;
  assign n7207 = ( x590 & n7202 ) | ( x590 & n7206 ) | ( n7202 & n7206 ) ;
  assign n7208 = n7206 ^ n7202 ^ 1'b0 ;
  assign n7209 = ( x590 & n7207 ) | ( x590 & n7208 ) | ( n7207 & n7208 ) ;
  assign n7222 = n7161 ^ x1198 ^ 1'b0 ;
  assign n7210 = n6644 ^ x377 ^ 1'b0 ;
  assign n7211 = n6653 | n7210 ;
  assign n7212 = x592 & n7211 ;
  assign n7213 = x1199 & ~n6787 ;
  assign n7214 = ( x1199 & n7212 ) | ( x1199 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7215 = n7214 ^ x592 ^ 1'b0 ;
  assign n7216 = ( ~x592 & n6653 ) | ( ~x592 & n7215 ) | ( n6653 & n7215 ) ;
  assign n7217 = ( x592 & n7214 ) | ( x592 & n7216 ) | ( n7214 & n7216 ) ;
  assign n7223 = n6787 & n7217 ;
  assign n7224 = ( n7161 & ~n7222 ) | ( n7161 & n7223 ) | ( ~n7222 & n7223 ) ;
  assign n7225 = n7224 ^ n7180 ^ 1'b0 ;
  assign n7226 = n7225 ^ n7180 ^ n7161 ;
  assign n7218 = x374 ^ x370 ^ x369 ;
  assign n7219 = n7218 ^ n7068 ^ x371 ;
  assign n7220 = ( n7161 & n7217 ) | ( n7161 & ~n7219 ) | ( n7217 & ~n7219 ) ;
  assign n7221 = ~n7217 & n7220 ;
  assign n7227 = ( n7180 & n7221 ) | ( n7180 & ~n7226 ) | ( n7221 & ~n7226 ) ;
  assign n7228 = n7226 | n7227 ;
  assign n7229 = ~x590 & n7228 ;
  assign n7230 = ( x591 & ~n7209 ) | ( x591 & n7229 ) | ( ~n7209 & n7229 ) ;
  assign n7231 = n7209 | n7230 ;
  assign n7232 = x590 & n6787 ;
  assign n7233 = n6860 & n6862 ;
  assign n7234 = n6787 & ~n6862 ;
  assign n7235 = ( x1199 & ~n7233 ) | ( x1199 & n7234 ) | ( ~n7233 & n7234 ) ;
  assign n7236 = n7233 | n7235 ;
  assign n7237 = ~x592 & n6920 ;
  assign n7238 = ~n6713 & n7237 ;
  assign n7239 = n7238 ^ n7236 ^ 1'b0 ;
  assign n7240 = ( ~n7162 & n7238 ) | ( ~n7162 & n7239 ) | ( n7238 & n7239 ) ;
  assign n7241 = ( n7236 & ~n7239 ) | ( n7236 & n7240 ) | ( ~n7239 & n7240 ) ;
  assign n7242 = x1198 & ~n7161 ;
  assign n7243 = n6688 & ~n7241 ;
  assign n7244 = ( n6688 & n7242 ) | ( n6688 & n7243 ) | ( n7242 & n7243 ) ;
  assign n7245 = n7241 & ~n7244 ;
  assign n7246 = n7161 ^ x1197 ^ 1'b0 ;
  assign n7247 = ( n7161 & n7241 ) | ( n7161 & ~n7246 ) | ( n7241 & ~n7246 ) ;
  assign n7248 = x333 | n7247 ;
  assign n7249 = n7245 & n7248 ;
  assign n7250 = x333 & ~n7247 ;
  assign n7251 = x333 | n7241 ;
  assign n7252 = ( n7244 & ~n7250 ) | ( n7244 & n7251 ) | ( ~n7250 & n7251 ) ;
  assign n7253 = ~n7244 & n7252 ;
  assign n7254 = n7249 ^ x391 ^ 1'b0 ;
  assign n7255 = ( n7249 & n7253 ) | ( n7249 & n7254 ) | ( n7253 & n7254 ) ;
  assign n7256 = ( n7249 & n7253 ) | ( n7249 & ~n7254 ) | ( n7253 & ~n7254 ) ;
  assign n7257 = n7255 ^ x392 ^ 1'b0 ;
  assign n7258 = ( n7255 & n7256 ) | ( n7255 & n7257 ) | ( n7256 & n7257 ) ;
  assign n7259 = x393 | n7258 ;
  assign n7260 = ( n7255 & n7256 ) | ( n7255 & ~n7257 ) | ( n7256 & ~n7257 ) ;
  assign n7261 = x393 & ~n7260 ;
  assign n7262 = n6780 & ~n7261 ;
  assign n7263 = n7259 & n7262 ;
  assign n7264 = x393 & ~n7258 ;
  assign n7265 = x393 | n7260 ;
  assign n7266 = ( n6780 & ~n7264 ) | ( n6780 & n7265 ) | ( ~n7264 & n7265 ) ;
  assign n7267 = ~n6780 & n7266 ;
  assign n7268 = ( ~x590 & n7263 ) | ( ~x590 & n7267 ) | ( n7263 & n7267 ) ;
  assign n7269 = ~x590 & n7268 ;
  assign n7270 = ( x591 & n7232 ) | ( x591 & ~n7269 ) | ( n7232 & ~n7269 ) ;
  assign n7271 = ~n7232 & n7270 ;
  assign n7272 = ( x588 & n7231 ) | ( x588 & ~n7271 ) | ( n7231 & ~n7271 ) ;
  assign n7273 = n7272 ^ n7231 ^ 1'b0 ;
  assign n7274 = ( x588 & n7272 ) | ( x588 & ~n7273 ) | ( n7272 & ~n7273 ) ;
  assign n7275 = n7274 ^ x217 ^ 1'b0 ;
  assign n7276 = x590 | x591 ;
  assign n7280 = x444 ^ x436 ^ 1'b0 ;
  assign n7277 = x422 ^ x414 ^ 1'b0 ;
  assign n7278 = n7277 ^ x446 ^ x434 ;
  assign n7279 = n7278 ^ x435 ^ x429 ;
  assign n7281 = n7280 ^ n7279 ^ x443 ;
  assign n7282 = n6862 & n7281 ;
  assign n7285 = x437 ^ x418 ^ x417 ;
  assign n7286 = n7285 ^ x464 ^ x453 ;
  assign n7283 = x438 ^ x416 ^ 1'b0 ;
  assign n7284 = n7283 ^ x431 ^ x415 ;
  assign n7287 = n7286 ^ n7284 ^ 1'b0 ;
  assign n7288 = x1197 & n7287 ;
  assign n7292 = x454 ^ x421 ^ 1'b0 ;
  assign n7291 = x459 ^ x432 ^ 1'b0 ;
  assign n7289 = x424 ^ x423 ^ 1'b0 ;
  assign n7290 = n7289 ^ x420 ^ x419 ;
  assign n7293 = n7292 ^ n7291 ^ n7290 ;
  assign n7294 = x1198 ^ x425 ^ 1'b0 ;
  assign n7295 = ( x425 & ~n7293 ) | ( x425 & n7294 ) | ( ~n7293 & n7294 ) ;
  assign n7296 = n7295 ^ n7294 ^ 1'b0 ;
  assign n7297 = ( ~n7282 & n7288 ) | ( ~n7282 & n7296 ) | ( n7288 & n7296 ) ;
  assign n7298 = n7282 | n7297 ;
  assign n7299 = n7180 & ~n7298 ;
  assign n7300 = x1199 | n7161 ;
  assign n7301 = n7299 | n7300 ;
  assign n7302 = x451 ^ x449 ^ x433 ;
  assign n7303 = x428 ^ x427 ^ 1'b0 ;
  assign n7304 = n7303 ^ x430 ^ x426 ;
  assign n7305 = n7304 ^ x448 ^ x445 ;
  assign n7306 = n7299 & ~n7305 ;
  assign n7307 = n7306 ^ n7299 ^ n7161 ;
  assign n7308 = n7302 & n7307 ;
  assign n7309 = ( n7161 & ~n7302 ) | ( n7161 & n7306 ) | ( ~n7302 & n7306 ) ;
  assign n7310 = ~n7302 & n7309 ;
  assign n7311 = ( x1199 & n7308 ) | ( x1199 & ~n7310 ) | ( n7308 & ~n7310 ) ;
  assign n7312 = ~n7308 & n7311 ;
  assign n7313 = ( n7276 & n7301 ) | ( n7276 & ~n7312 ) | ( n7301 & ~n7312 ) ;
  assign n7314 = ~n7276 & n7313 ;
  assign n7315 = n6787 & n7276 ;
  assign n7316 = ( x588 & n7314 ) | ( x588 & ~n7315 ) | ( n7314 & ~n7315 ) ;
  assign n7317 = ~n7314 & n7316 ;
  assign n7318 = x57 | n5193 ;
  assign n7319 = ( n6612 & n7317 ) | ( n6612 & n7318 ) | ( n7317 & n7318 ) ;
  assign n7320 = ~n7317 & n7319 ;
  assign n7321 = ( n7274 & ~n7275 ) | ( n7274 & n7320 ) | ( ~n7275 & n7320 ) ;
  assign n7322 = ( x217 & n7275 ) | ( x217 & n7321 ) | ( n7275 & n7321 ) ;
  assign n7378 = n6855 & n7276 ;
  assign n7379 = n7280 ^ n7279 ^ 1'b0 ;
  assign n7331 = x443 & ~x592 ;
  assign n7380 = ~n6522 & n7331 ;
  assign n7381 = n7379 | n7380 ;
  assign n7382 = ( n6855 & n7331 ) | ( n6855 & ~n7381 ) | ( n7331 & ~n7381 ) ;
  assign n7383 = ~n7381 & n7382 ;
  assign n7328 = x443 | x592 ;
  assign n7384 = ~n6855 & n7328 ;
  assign n7385 = n6522 | n7328 ;
  assign n7386 = ( n7379 & n7384 ) | ( n7379 & n7385 ) | ( n7384 & n7385 ) ;
  assign n7387 = ~n7384 & n7386 ;
  assign n7388 = ( x1196 & n7383 ) | ( x1196 & ~n7387 ) | ( n7383 & ~n7387 ) ;
  assign n7389 = ~n7383 & n7388 ;
  assign n7390 = ( x1196 & n6855 ) | ( x1196 & ~n7389 ) | ( n6855 & ~n7389 ) ;
  assign n7391 = ~n7389 & n7390 ;
  assign n7324 = n7284 & n7286 ;
  assign n7325 = ~n7296 & n7324 ;
  assign n7326 = ( x1197 & n7284 ) | ( x1197 & n7288 ) | ( n7284 & n7288 ) ;
  assign n7327 = ( n7296 & ~n7325 ) | ( n7296 & n7326 ) | ( ~n7325 & n7326 ) ;
  assign n7392 = n7391 ^ n7327 ^ 1'b0 ;
  assign n7393 = ( n7052 & n7391 ) | ( n7052 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7394 = n7393 ^ n7303 ^ 1'b0 ;
  assign n7395 = ( n7052 & n7393 ) | ( n7052 & ~n7394 ) | ( n7393 & ~n7394 ) ;
  assign n7396 = n7395 ^ n7393 ^ n7052 ;
  assign n7397 = n7396 ^ x430 ^ 1'b0 ;
  assign n7398 = ( n7395 & n7396 ) | ( n7395 & ~n7397 ) | ( n7396 & ~n7397 ) ;
  assign n7399 = ( n7395 & n7396 ) | ( n7395 & n7397 ) | ( n7396 & n7397 ) ;
  assign n7400 = n7398 ^ x426 ^ 1'b0 ;
  assign n7401 = ( n7398 & n7399 ) | ( n7398 & n7400 ) | ( n7399 & n7400 ) ;
  assign n7402 = ( n7398 & n7399 ) | ( n7398 & ~n7400 ) | ( n7399 & ~n7400 ) ;
  assign n7403 = n7401 ^ x445 ^ 1'b0 ;
  assign n7406 = ( n7401 & n7402 ) | ( n7401 & ~n7403 ) | ( n7402 & ~n7403 ) ;
  assign n7410 = x448 & n7406 ;
  assign n7404 = ( n7401 & n7402 ) | ( n7401 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7411 = ~x448 & n7404 ;
  assign n7412 = ( n7302 & n7410 ) | ( n7302 & ~n7411 ) | ( n7410 & ~n7411 ) ;
  assign n7413 = ~n7410 & n7412 ;
  assign n7405 = x448 & n7404 ;
  assign n7407 = ~x448 & n7406 ;
  assign n7408 = ( n7302 & ~n7405 ) | ( n7302 & n7407 ) | ( ~n7405 & n7407 ) ;
  assign n7409 = n7405 | n7408 ;
  assign n7414 = n7413 ^ n7409 ^ 1'b0 ;
  assign n7415 = ( x1199 & ~n7409 ) | ( x1199 & n7413 ) | ( ~n7409 & n7413 ) ;
  assign n7416 = ( x1199 & ~n7414 ) | ( x1199 & n7415 ) | ( ~n7414 & n7415 ) ;
  assign n7417 = x1199 | n7393 ;
  assign n7418 = ( n7276 & ~n7416 ) | ( n7276 & n7417 ) | ( ~n7416 & n7417 ) ;
  assign n7419 = ~n7276 & n7418 ;
  assign n7420 = ( n6612 & n7378 ) | ( n6612 & ~n7419 ) | ( n7378 & ~n7419 ) ;
  assign n7421 = ~n7378 & n7420 ;
  assign n7323 = n6504 & n7276 ;
  assign n7329 = n7328 ^ n6504 ^ 1'b0 ;
  assign n7330 = ( n6504 & n6522 ) | ( n6504 & ~n7329 ) | ( n6522 & ~n7329 ) ;
  assign n7332 = n7331 ^ n6522 ^ 1'b0 ;
  assign n7333 = ( n6504 & n6522 ) | ( n6504 & ~n7332 ) | ( n6522 & ~n7332 ) ;
  assign n7334 = n7330 ^ x444 ^ 1'b0 ;
  assign n7335 = ( n7330 & n7333 ) | ( n7330 & n7334 ) | ( n7333 & n7334 ) ;
  assign n7336 = x436 & ~n7335 ;
  assign n7337 = ( n7330 & n7333 ) | ( n7330 & ~n7334 ) | ( n7333 & ~n7334 ) ;
  assign n7338 = x436 | n7337 ;
  assign n7339 = ( ~n7279 & n7336 ) | ( ~n7279 & n7338 ) | ( n7336 & n7338 ) ;
  assign n7340 = ~n7336 & n7339 ;
  assign n7341 = x436 | n7335 ;
  assign n7342 = x436 & ~n7337 ;
  assign n7343 = n7279 & ~n7342 ;
  assign n7344 = n7341 & n7343 ;
  assign n7345 = ( x1196 & n7340 ) | ( x1196 & ~n7344 ) | ( n7340 & ~n7344 ) ;
  assign n7346 = ~n7340 & n7345 ;
  assign n7347 = ( n6539 & n7327 ) | ( n6539 & ~n7346 ) | ( n7327 & ~n7346 ) ;
  assign n7348 = ~n7327 & n7347 ;
  assign n7349 = n7348 ^ n6526 ^ 1'b0 ;
  assign n7350 = ( ~n6526 & n7327 ) | ( ~n6526 & n7349 ) | ( n7327 & n7349 ) ;
  assign n7351 = ( n6526 & n7348 ) | ( n6526 & n7350 ) | ( n7348 & n7350 ) ;
  assign n7352 = x1199 | n7351 ;
  assign n7353 = n7302 ^ x448 ^ 1'b0 ;
  assign n7354 = n6526 ^ x428 ^ 1'b0 ;
  assign n7355 = ( n6526 & n7351 ) | ( n6526 & ~n7354 ) | ( n7351 & ~n7354 ) ;
  assign n7356 = ( n6526 & n7351 ) | ( n6526 & n7354 ) | ( n7351 & n7354 ) ;
  assign n7357 = n7355 ^ x427 ^ 1'b0 ;
  assign n7358 = ( n7355 & n7356 ) | ( n7355 & n7357 ) | ( n7356 & n7357 ) ;
  assign n7359 = ( n7355 & n7356 ) | ( n7355 & ~n7357 ) | ( n7356 & ~n7357 ) ;
  assign n7360 = n7358 ^ x430 ^ 1'b0 ;
  assign n7361 = ( n7358 & n7359 ) | ( n7358 & ~n7360 ) | ( n7359 & ~n7360 ) ;
  assign n7362 = ( n7358 & n7359 ) | ( n7358 & n7360 ) | ( n7359 & n7360 ) ;
  assign n7363 = n7361 ^ x426 ^ 1'b0 ;
  assign n7364 = ( n7361 & n7362 ) | ( n7361 & ~n7363 ) | ( n7362 & ~n7363 ) ;
  assign n7365 = ( n7361 & n7362 ) | ( n7361 & n7363 ) | ( n7362 & n7363 ) ;
  assign n7366 = n7364 ^ x445 ^ 1'b0 ;
  assign n7367 = ( n7364 & n7365 ) | ( n7364 & ~n7366 ) | ( n7365 & ~n7366 ) ;
  assign n7368 = n7353 & n7367 ;
  assign n7369 = ( n7364 & n7365 ) | ( n7364 & n7366 ) | ( n7365 & n7366 ) ;
  assign n7370 = n7369 ^ n7353 ^ 1'b0 ;
  assign n7371 = ( ~n7353 & n7369 ) | ( ~n7353 & n7370 ) | ( n7369 & n7370 ) ;
  assign n7372 = ( x1199 & n7368 ) | ( x1199 & ~n7371 ) | ( n7368 & ~n7371 ) ;
  assign n7373 = ~n7368 & n7372 ;
  assign n7374 = ( n7276 & n7352 ) | ( n7276 & ~n7373 ) | ( n7352 & ~n7373 ) ;
  assign n7375 = ~n7276 & n7374 ;
  assign n7376 = ( n6612 & ~n7323 ) | ( n6612 & n7375 ) | ( ~n7323 & n7375 ) ;
  assign n7377 = n7323 | n7376 ;
  assign n7422 = n7421 ^ n7377 ^ 1'b0 ;
  assign n7423 = ( x588 & ~n7377 ) | ( x588 & n7421 ) | ( ~n7377 & n7421 ) ;
  assign n7424 = ( x588 & ~n7422 ) | ( x588 & n7423 ) | ( ~n7422 & n7423 ) ;
  assign n7425 = ( x57 & n5193 ) | ( x57 & ~n7424 ) | ( n5193 & ~n7424 ) ;
  assign n7426 = n7424 | n7425 ;
  assign n7427 = ~n7322 & n7426 ;
  assign n7428 = ( n7160 & n7322 ) | ( n7160 & ~n7427 ) | ( n7322 & ~n7427 ) ;
  assign n7429 = x1161 & ~x1163 ;
  assign n7430 = n1611 & n7429 ;
  assign n7431 = ~x31 & x1162 ;
  assign n7432 = n7430 & n7431 ;
  assign n7433 = n6612 & ~n6855 ;
  assign n7434 = n7318 | n7433 ;
  assign n7435 = ( n6504 & n6612 ) | ( n6504 & ~n7434 ) | ( n6612 & ~n7434 ) ;
  assign n7436 = ~n7434 & n7435 ;
  assign n7437 = n6612 & n7318 ;
  assign n7438 = n6787 & n7437 ;
  assign n7439 = ( x217 & n7436 ) | ( x217 & ~n7438 ) | ( n7436 & ~n7438 ) ;
  assign n7440 = ~n7436 & n7439 ;
  assign n7441 = x1161 | x1162 ;
  assign n7442 = ( x1163 & ~n7440 ) | ( x1163 & n7441 ) | ( ~n7440 & n7441 ) ;
  assign n7443 = n7440 | n7442 ;
  assign n7444 = ~n7432 & n7443 ;
  assign n7445 = ( n7428 & n7432 ) | ( n7428 & ~n7444 ) | ( n7432 & ~n7444 ) ;
  assign n7446 = n2109 | n2120 ;
  assign n7447 = x55 | x74 ;
  assign n7448 = n7446 | n7447 ;
  assign n7449 = x829 & ~x1093 ;
  assign n7450 = n5020 & n7449 ;
  assign n7451 = n1670 | n7450 ;
  assign n7452 = x24 | n1269 ;
  assign n7453 = n1290 | n1375 ;
  assign n7454 = x51 | n7453 ;
  assign n7455 = n7452 | n7454 ;
  assign n7456 = n7451 | n7455 ;
  assign n7457 = n5035 & ~n6412 ;
  assign n7458 = x252 & ~n7457 ;
  assign n7459 = x87 | n1994 ;
  assign n7460 = x75 & ~x100 ;
  assign n7461 = ~n7459 & n7460 ;
  assign n7462 = ~x137 & n7461 ;
  assign n7463 = ~n5045 & n7462 ;
  assign n7464 = ( n7456 & ~n7458 ) | ( n7456 & n7463 ) | ( ~n7458 & n7463 ) ;
  assign n7465 = ~n7456 & n7464 ;
  assign n7466 = x100 & ~n1994 ;
  assign n7467 = x24 | x90 ;
  assign n7468 = n5161 | n7467 ;
  assign n7469 = x50 & ~n1463 ;
  assign n7470 = ~n1261 & n7469 ;
  assign n7471 = n1259 | n1392 ;
  assign n7472 = n1371 | n7471 ;
  assign n7473 = x93 | n7472 ;
  assign n7474 = n7470 & ~n7473 ;
  assign n7475 = ~n7468 & n7474 ;
  assign n7476 = x32 | n7475 ;
  assign n7477 = x24 | x841 ;
  assign n7478 = x32 & n7477 ;
  assign n7479 = ~n1380 & n7478 ;
  assign n7480 = x137 | n6387 ;
  assign n7481 = n6612 & ~n7451 ;
  assign n7482 = n1271 | n1652 ;
  assign n7483 = ( ~n7480 & n7481 ) | ( ~n7480 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7484 = n7480 | n7483 ;
  assign n7485 = n1226 | n1522 ;
  assign n7486 = x103 | n1236 ;
  assign n7487 = n7485 | n7486 ;
  assign n7488 = x89 | x102 ;
  assign n7489 = n6379 | n7488 ;
  assign n7490 = x68 | x73 ;
  assign n7491 = x76 & ~x84 ;
  assign n7492 = ~n1244 & n7491 ;
  assign n7493 = x49 | x66 ;
  assign n7494 = ( n7490 & n7492 ) | ( n7490 & ~n7493 ) | ( n7492 & ~n7493 ) ;
  assign n7495 = ~n7490 & n7494 ;
  assign n7496 = x64 | x81 ;
  assign n7497 = n1230 | n7496 ;
  assign n7498 = ( n7489 & n7495 ) | ( n7489 & ~n7497 ) | ( n7495 & ~n7497 ) ;
  assign n7499 = ~n7489 & n7498 ;
  assign n7500 = n1231 | n1485 ;
  assign n7501 = x45 | x48 ;
  assign n7502 = x61 | x104 ;
  assign n7503 = n7501 | n7502 ;
  assign n7504 = n7500 | n7503 ;
  assign n7505 = ( n7487 & n7499 ) | ( n7487 & ~n7504 ) | ( n7499 & ~n7504 ) ;
  assign n7506 = ~n7487 & n7505 ;
  assign n7507 = ~n1261 & n7506 ;
  assign n7508 = ~n7472 & n7507 ;
  assign n7509 = ~n7484 & n7508 ;
  assign n7510 = ( x24 & n7484 ) | ( x24 & ~n7509 ) | ( n7484 & ~n7509 ) ;
  assign n7511 = n1263 | n1372 ;
  assign n7512 = n7469 | n7506 ;
  assign n7513 = ~n7511 & n7512 ;
  assign n7514 = ( x24 & ~n7510 ) | ( x24 & n7513 ) | ( ~n7510 & n7513 ) ;
  assign n7515 = ~n7510 & n7514 ;
  assign n7516 = x137 | n7481 ;
  assign n7517 = n7475 & n7516 ;
  assign n7518 = ( ~x32 & n7515 ) | ( ~x32 & n7517 ) | ( n7515 & n7517 ) ;
  assign n7519 = ~x32 & n7518 ;
  assign n7520 = ( ~n5165 & n7479 ) | ( ~n5165 & n7519 ) | ( n7479 & n7519 ) ;
  assign n7521 = ~n5165 & n7520 ;
  assign n7522 = ~n5163 & n5165 ;
  assign n7523 = n7521 ^ n7476 ^ 1'b0 ;
  assign n7524 = ( ~n7476 & n7522 ) | ( ~n7476 & n7523 ) | ( n7522 & n7523 ) ;
  assign n7525 = ( n7476 & n7521 ) | ( n7476 & n7524 ) | ( n7521 & n7524 ) ;
  assign n7526 = ( x95 & ~n2095 ) | ( x95 & n7525 ) | ( ~n2095 & n7525 ) ;
  assign n7527 = ~x95 & n7526 ;
  assign n7528 = x129 & ~n1292 ;
  assign n7529 = ~x137 & x252 ;
  assign n7530 = n5044 | n7457 ;
  assign n7531 = n7529 & ~n7530 ;
  assign n7532 = n7528 & n7531 ;
  assign n7533 = ~n5035 & n5044 ;
  assign n7534 = ~n5419 & n7533 ;
  assign n7535 = ( ~x137 & n7532 ) | ( ~x137 & n7534 ) | ( n7532 & n7534 ) ;
  assign n7536 = n7532 ^ x137 ^ 1'b0 ;
  assign n7537 = ( n7532 & n7535 ) | ( n7532 & ~n7536 ) | ( n7535 & ~n7536 ) ;
  assign n7538 = n7527 ^ n7466 ^ 1'b0 ;
  assign n7539 = ( ~n7466 & n7537 ) | ( ~n7466 & n7538 ) | ( n7537 & n7538 ) ;
  assign n7540 = ( n7466 & n7527 ) | ( n7466 & n7539 ) | ( n7527 & n7539 ) ;
  assign n7541 = ( ~n2044 & n7465 ) | ( ~n2044 & n7540 ) | ( n7465 & n7540 ) ;
  assign n7542 = n7465 ^ n2044 ^ 1'b0 ;
  assign n7543 = ( n7465 & n7541 ) | ( n7465 & ~n7542 ) | ( n7541 & ~n7542 ) ;
  assign n7544 = ( n5015 & ~n7448 ) | ( n5015 & n7543 ) | ( ~n7448 & n7543 ) ;
  assign n7545 = ~n5015 & n7544 ;
  assign n7546 = n2120 ^ n2109 ^ 1'b0 ;
  assign n7547 = x149 | x157 ;
  assign n7548 = ~n5075 & n7547 ;
  assign n7549 = x149 & x157 ;
  assign n7550 = n7548 & ~n7549 ;
  assign n7551 = x232 & n7550 ;
  assign n7552 = x75 & ~n7551 ;
  assign n7553 = x100 & ~n7551 ;
  assign n7554 = n7552 | n7553 ;
  assign n7555 = x75 | x100 ;
  assign n7556 = n6411 & ~n7555 ;
  assign n7557 = x169 & n7556 ;
  assign n7558 = n7554 | n7557 ;
  assign n7559 = x74 & n7558 ;
  assign n7560 = x164 & n7556 ;
  assign n7561 = n7554 | n7560 ;
  assign n7562 = x54 & n7561 ;
  assign n7563 = ( x38 & n7554 ) | ( x38 & n7561 ) | ( n7554 & n7561 ) ;
  assign n7564 = n7562 | n7563 ;
  assign n7565 = x74 | n7564 ;
  assign n7566 = ( ~x74 & n7559 ) | ( ~x74 & n7565 ) | ( n7559 & n7565 ) ;
  assign n7567 = ( n2109 & ~n7546 ) | ( n2109 & n7566 ) | ( ~n7546 & n7566 ) ;
  assign n7568 = ( n2120 & n7546 ) | ( n2120 & n7567 ) | ( n7546 & n7567 ) ;
  assign n7569 = x40 | n1230 ;
  assign n7570 = x38 | n7569 ;
  assign n7571 = n7555 | n7570 ;
  assign n7572 = n2067 | n7571 ;
  assign n7573 = n2109 & ~n7572 ;
  assign n7574 = ~x38 & n7569 ;
  assign n7575 = x164 & n6411 ;
  assign n7576 = x38 & ~n7575 ;
  assign n7577 = ( x100 & ~n7574 ) | ( x100 & n7576 ) | ( ~n7574 & n7576 ) ;
  assign n7578 = n7574 | n7577 ;
  assign n7579 = x75 | n7578 ;
  assign n7580 = n7579 ^ x54 ^ 1'b0 ;
  assign n7581 = x92 & ~n7554 ;
  assign n7582 = ( n7579 & ~n7580 ) | ( n7579 & n7581 ) | ( ~n7580 & n7581 ) ;
  assign n7583 = ( x54 & n7580 ) | ( x54 & n7582 ) | ( n7580 & n7582 ) ;
  assign n7584 = x92 | n7552 ;
  assign n7585 = n2051 | n7576 ;
  assign n7586 = x102 | n7496 ;
  assign n7587 = n1231 | n7586 ;
  assign n7588 = n1228 | n7587 ;
  assign n7589 = n1250 | n7588 ;
  assign n7590 = x60 | n7589 ;
  assign n7591 = n1387 | n1394 ;
  assign n7592 = x53 | n7591 ;
  assign n7593 = n7590 | n7592 ;
  assign n7594 = x58 | n7593 ;
  assign n7595 = n6387 | n7594 ;
  assign n7596 = x32 | n1272 ;
  assign n7597 = n7595 | n7596 ;
  assign n7598 = x95 | n7597 ;
  assign n7599 = x149 & n6411 ;
  assign n7600 = x39 | n7599 ;
  assign n7601 = ( ~n7569 & n7598 ) | ( ~n7569 & n7600 ) | ( n7598 & n7600 ) ;
  assign n7602 = ~n7569 & n7601 ;
  assign n7603 = x38 | n7602 ;
  assign n7604 = ~n7585 & n7603 ;
  assign n7605 = x87 & ~n7578 ;
  assign n7606 = n7553 | n7605 ;
  assign n7607 = ( ~x75 & n7604 ) | ( ~x75 & n7606 ) | ( n7604 & n7606 ) ;
  assign n7608 = ~x75 & n7607 ;
  assign n7609 = ( ~n7583 & n7584 ) | ( ~n7583 & n7608 ) | ( n7584 & n7608 ) ;
  assign n7610 = ~n7583 & n7609 ;
  assign n7611 = ( ~x74 & n7562 ) | ( ~x74 & n7610 ) | ( n7562 & n7610 ) ;
  assign n7612 = ~x74 & n7611 ;
  assign n7613 = ( x55 & n7559 ) | ( x55 & ~n7612 ) | ( n7559 & ~n7612 ) ;
  assign n7614 = ~n7559 & n7613 ;
  assign n7615 = x74 ^ x55 ^ 1'b0 ;
  assign n7616 = x299 & ~n7550 ;
  assign n7617 = x178 & x183 ;
  assign n7618 = x178 | x183 ;
  assign n7619 = ~n5075 & n7618 ;
  assign n7620 = ~n7617 & n7619 ;
  assign n7621 = x299 | n7620 ;
  assign n7622 = ( x232 & n7616 ) | ( x232 & n7621 ) | ( n7616 & n7621 ) ;
  assign n7623 = ~n7616 & n7622 ;
  assign n7624 = x100 & ~n7623 ;
  assign n7625 = x75 & ~n7623 ;
  assign n7626 = n7624 | n7625 ;
  assign n7627 = x191 & ~x299 ;
  assign n7628 = x169 & x299 ;
  assign n7629 = n7627 | n7628 ;
  assign n7630 = n7556 & n7629 ;
  assign n7631 = n7626 | n7630 ;
  assign n7632 = ( x74 & ~n7615 ) | ( x74 & n7631 ) | ( ~n7615 & n7631 ) ;
  assign n7633 = ( x55 & n7615 ) | ( x55 & n7632 ) | ( n7615 & n7632 ) ;
  assign n7634 = x299 ^ x164 ^ 1'b0 ;
  assign n7635 = ( x164 & x186 ) | ( x164 & ~n7634 ) | ( x186 & ~n7634 ) ;
  assign n7636 = n6411 & n7635 ;
  assign n7637 = ~n7555 & n7636 ;
  assign n7638 = n7626 | n7637 ;
  assign n7639 = ~x75 & x92 ;
  assign n7640 = x38 & n7636 ;
  assign n7641 = n7640 ^ x100 ^ 1'b0 ;
  assign n7642 = ( ~n7623 & n7640 ) | ( ~n7623 & n7641 ) | ( n7640 & n7641 ) ;
  assign n7643 = n1205 | n7569 ;
  assign n7644 = x232 & ~n2206 ;
  assign n7645 = x176 | x299 ;
  assign n7646 = ~n5075 & n7645 ;
  assign n7647 = n7644 & n7646 ;
  assign n7648 = n1206 | n7598 ;
  assign n7649 = n7647 | n7648 ;
  assign n7650 = ~n7643 & n7649 ;
  assign n7651 = ( n7639 & n7642 ) | ( n7639 & n7650 ) | ( n7642 & n7650 ) ;
  assign n7652 = n7639 & n7651 ;
  assign n7653 = x87 & n7643 ;
  assign n7654 = ~n7642 & n7653 ;
  assign n7655 = ~x299 & n6411 ;
  assign n7656 = n5052 & n7655 ;
  assign n7657 = ~x164 & x186 ;
  assign n7658 = n7656 & n7657 ;
  assign n7659 = n5017 & n6411 ;
  assign n7660 = x186 & ~n7659 ;
  assign n7661 = x299 & n6411 ;
  assign n7662 = n5052 & n7661 ;
  assign n7663 = x186 | n7662 ;
  assign n7664 = ( x164 & n7660 ) | ( x164 & n7663 ) | ( n7660 & n7663 ) ;
  assign n7665 = ~n7660 & n7664 ;
  assign n7666 = ( x38 & n7658 ) | ( x38 & n7665 ) | ( n7658 & n7665 ) ;
  assign n7667 = n7665 ^ n7658 ^ 1'b0 ;
  assign n7668 = ( x38 & n7666 ) | ( x38 & n7667 ) | ( n7666 & n7667 ) ;
  assign n7669 = x216 & n5390 ;
  assign n7670 = n7569 | n7669 ;
  assign n7671 = x299 & n7670 ;
  assign n7672 = n5365 & ~n5378 ;
  assign n7673 = n5073 & n7672 ;
  assign n7674 = n5096 | n7673 ;
  assign n7675 = ~n7598 & n7674 ;
  assign n7676 = n5099 & n7675 ;
  assign n7677 = n7569 | n7676 ;
  assign n7678 = x224 & n5376 ;
  assign n7679 = n7569 | n7678 ;
  assign n7680 = n7677 & n7679 ;
  assign n7681 = ~n7598 & n7673 ;
  assign n7682 = ~n5075 & n7681 ;
  assign n7683 = n7569 | n7682 ;
  assign n7684 = n5114 & n7683 ;
  assign n7685 = n7679 & n7684 ;
  assign n7686 = x174 & n7685 ;
  assign n7687 = ( ~x299 & n7680 ) | ( ~x299 & n7686 ) | ( n7680 & n7686 ) ;
  assign n7688 = ~x299 & n7687 ;
  assign n7689 = n5061 & ~n5075 ;
  assign n7690 = n7569 | n7681 ;
  assign n7691 = n7689 & n7690 ;
  assign n7692 = x152 & n7691 ;
  assign n7693 = n7677 | n7692 ;
  assign n7694 = ( x154 & ~n7669 ) | ( x154 & n7693 ) | ( ~n7669 & n7693 ) ;
  assign n7695 = n7669 ^ x154 ^ 1'b0 ;
  assign n7696 = ( n7669 & ~n7694 ) | ( n7669 & n7695 ) | ( ~n7694 & n7695 ) ;
  assign n7697 = n5096 & ~n7598 ;
  assign n7698 = ~n5083 & n7697 ;
  assign n7699 = n7569 | n7698 ;
  assign n7700 = n5075 | n7699 ;
  assign n7701 = x152 | n7700 ;
  assign n7702 = ~n5075 & n7675 ;
  assign n7703 = n7569 | n7702 ;
  assign n7704 = n5061 & n7703 ;
  assign n7705 = n7677 | n7704 ;
  assign n7706 = ~x154 & n7705 ;
  assign n7707 = ( ~n7696 & n7701 ) | ( ~n7696 & n7706 ) | ( n7701 & n7706 ) ;
  assign n7708 = n7707 ^ n7696 ^ 1'b0 ;
  assign n7709 = ( n7696 & ~n7707 ) | ( n7696 & n7708 ) | ( ~n7707 & n7708 ) ;
  assign n7710 = ~n7688 & n7709 ;
  assign n7711 = ( n7671 & n7688 ) | ( n7671 & ~n7710 ) | ( n7688 & ~n7710 ) ;
  assign n7712 = x176 & x232 ;
  assign n7713 = n7711 & n7712 ;
  assign n7714 = n7671 & n7705 ;
  assign n7715 = n5114 & n7703 ;
  assign n7716 = ( n7679 & n7680 ) | ( n7679 & n7715 ) | ( n7680 & n7715 ) ;
  assign n7717 = ~x299 & n7716 ;
  assign n7718 = ( ~x232 & n7714 ) | ( ~x232 & n7717 ) | ( n7714 & n7717 ) ;
  assign n7719 = ~x232 & n7718 ;
  assign n7720 = x39 & ~n7719 ;
  assign n7721 = ~x176 & x232 ;
  assign n7722 = ~n7569 & n7678 ;
  assign n7723 = ~n5075 & n5114 ;
  assign n7724 = n7697 & n7723 ;
  assign n7725 = n7722 & ~n7724 ;
  assign n7726 = n7679 & ~n7725 ;
  assign n7727 = ~x299 & n7726 ;
  assign n7728 = n7711 | n7727 ;
  assign n7729 = n7721 & n7728 ;
  assign n7730 = ( n7713 & n7720 ) | ( n7713 & ~n7729 ) | ( n7720 & ~n7729 ) ;
  assign n7731 = ~n7713 & n7730 ;
  assign n7732 = x40 | x479 ;
  assign n7733 = ~n1230 & n7597 ;
  assign n7734 = ~n7732 & n7733 ;
  assign n7735 = x95 & n7569 ;
  assign n7736 = n1224 | n7735 ;
  assign n7737 = ~n7734 & n7736 ;
  assign n7738 = x32 & n7569 ;
  assign n7739 = ~n1230 & n1270 ;
  assign n7740 = ~n1230 & n7595 ;
  assign n7741 = x70 & ~n7740 ;
  assign n7742 = ~n1230 & n1268 ;
  assign n7743 = x70 | n7742 ;
  assign n7744 = x841 | n7594 ;
  assign n7745 = ~n1230 & n7744 ;
  assign n7746 = x90 & ~n7745 ;
  assign n7747 = n1268 | n7746 ;
  assign n7748 = ~n1230 & n7593 ;
  assign n7749 = x58 & ~n7748 ;
  assign n7750 = ~x60 & n7469 ;
  assign n7751 = n1386 | n7750 ;
  assign n7752 = x53 & n7590 ;
  assign n7753 = n7751 & ~n7752 ;
  assign n7754 = x111 | n1232 ;
  assign n7755 = x68 | n1233 ;
  assign n7756 = x36 | n7755 ;
  assign n7757 = n7754 | n7756 ;
  assign n7758 = x66 | x84 ;
  assign n7759 = x73 & ~x82 ;
  assign n7760 = ~n7758 & n7759 ;
  assign n7761 = ~n7757 & n7760 ;
  assign n7762 = ( n1242 & ~n7588 ) | ( n1242 & n7761 ) | ( ~n7588 & n7761 ) ;
  assign n7763 = ~n1242 & n7762 ;
  assign n7764 = ~n1260 & n7763 ;
  assign n7765 = n1230 | n7764 ;
  assign n7766 = ( ~n1387 & n7753 ) | ( ~n1387 & n7765 ) | ( n7753 & n7765 ) ;
  assign n7767 = ~n1387 & n7766 ;
  assign n7768 = ( n1230 & n1394 ) | ( n1230 & n7591 ) | ( n1394 & n7591 ) ;
  assign n7769 = n7767 | n7768 ;
  assign n7770 = ~n1230 & n1394 ;
  assign n7771 = ( x58 & n7769 ) | ( x58 & ~n7770 ) | ( n7769 & ~n7770 ) ;
  assign n7772 = ~x58 & n7771 ;
  assign n7773 = ( ~x90 & n7749 ) | ( ~x90 & n7772 ) | ( n7749 & n7772 ) ;
  assign n7774 = ( ~n7743 & n7747 ) | ( ~n7743 & n7773 ) | ( n7747 & n7773 ) ;
  assign n7775 = ~n7743 & n7774 ;
  assign n7776 = ( ~x51 & n7741 ) | ( ~x51 & n7775 ) | ( n7741 & n7775 ) ;
  assign n7777 = ~x51 & n7776 ;
  assign n7778 = x51 & n1230 ;
  assign n7779 = n1270 | n7778 ;
  assign n7780 = ( ~n7739 & n7777 ) | ( ~n7739 & n7779 ) | ( n7777 & n7779 ) ;
  assign n7781 = ~n7739 & n7780 ;
  assign n7782 = ( ~x32 & x40 ) | ( ~x32 & n7781 ) | ( x40 & n7781 ) ;
  assign n7783 = ~x32 & n7782 ;
  assign n7784 = ( ~x95 & n7738 ) | ( ~x95 & n7783 ) | ( n7738 & n7783 ) ;
  assign n7785 = n7737 | n7784 ;
  assign n7786 = n1374 | n5160 ;
  assign n7787 = n7744 | n7786 ;
  assign n7788 = ~n7569 & n7787 ;
  assign n7789 = x32 & ~n7788 ;
  assign n7790 = ( ~x95 & n7783 ) | ( ~x95 & n7789 ) | ( n7783 & n7789 ) ;
  assign n7791 = ~n5165 & n7790 ;
  assign n7792 = ( ~x232 & n7785 ) | ( ~x232 & n7791 ) | ( n7785 & n7791 ) ;
  assign n7793 = ~x232 & n7792 ;
  assign n7794 = ~x198 & n7790 ;
  assign n7795 = n7785 | n7794 ;
  assign n7796 = n5075 & ~n7795 ;
  assign n7797 = ~n7591 & n7753 ;
  assign n7798 = ( ~x58 & n1230 ) | ( ~x58 & n7797 ) | ( n1230 & n7797 ) ;
  assign n7799 = ~x58 & n7798 ;
  assign n7800 = ( ~x90 & n7749 ) | ( ~x90 & n7799 ) | ( n7749 & n7799 ) ;
  assign n7801 = n7747 | n7800 ;
  assign n7802 = ~n7743 & n7801 ;
  assign n7803 = ( ~x51 & n7741 ) | ( ~x51 & n7802 ) | ( n7741 & n7802 ) ;
  assign n7804 = ~x51 & n7803 ;
  assign n7805 = ( ~n7739 & n7779 ) | ( ~n7739 & n7804 ) | ( n7779 & n7804 ) ;
  assign n7806 = ~n7739 & n7805 ;
  assign n7807 = ~x40 & n7806 ;
  assign n7808 = ( ~x32 & x40 ) | ( ~x32 & n7807 ) | ( x40 & n7807 ) ;
  assign n7809 = ( ~x95 & n7789 ) | ( ~x95 & n7808 ) | ( n7789 & n7808 ) ;
  assign n7810 = ~x198 & n7809 ;
  assign n7811 = n5075 | n7735 ;
  assign n7819 = ~x95 & n7569 ;
  assign n7812 = ~x40 & n1230 ;
  assign n7813 = x95 & ~n7812 ;
  assign n7814 = x32 & ~n7812 ;
  assign n7815 = x32 | n7807 ;
  assign n7816 = ~n7814 & n7815 ;
  assign n7817 = x95 | n7816 ;
  assign n7818 = ~n7813 & n7817 ;
  assign n7820 = n7819 ^ n7818 ^ n7812 ;
  assign n7821 = n7811 | n7820 ;
  assign n7822 = n7810 | n7821 ;
  assign n7823 = ~n7796 & n7822 ;
  assign n7824 = ~n1230 & n5160 ;
  assign n7825 = x32 | n7824 ;
  assign n7826 = x93 & n1230 ;
  assign n7827 = n5160 | n7826 ;
  assign n7828 = n1230 | n7749 ;
  assign n7829 = n7828 ^ x90 ^ 1'b0 ;
  assign n7830 = ( ~n7745 & n7828 ) | ( ~n7745 & n7829 ) | ( n7828 & n7829 ) ;
  assign n7831 = ~x93 & n7830 ;
  assign n7832 = n7827 | n7831 ;
  assign n7833 = ~n7825 & n7832 ;
  assign n7834 = ( x40 & n7738 ) | ( x40 & ~n7833 ) | ( n7738 & ~n7833 ) ;
  assign n7835 = n7833 | n7834 ;
  assign n7836 = ~x95 & n7835 ;
  assign n7837 = n7811 | n7836 ;
  assign n7838 = ~n7796 & n7837 ;
  assign n7839 = n7823 ^ x183 ^ 1'b0 ;
  assign n7840 = ( n7823 & n7838 ) | ( n7823 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7841 = x174 | n7840 ;
  assign n7842 = ~n7511 & n7763 ;
  assign n7843 = ~x90 & n7842 ;
  assign n7844 = ( ~x93 & n7830 ) | ( ~x93 & n7843 ) | ( n7830 & n7843 ) ;
  assign n7845 = ~x93 & n7844 ;
  assign n7846 = ( ~n7825 & n7827 ) | ( ~n7825 & n7845 ) | ( n7827 & n7845 ) ;
  assign n7847 = ~n7825 & n7846 ;
  assign n7848 = ( x40 & n7738 ) | ( x40 & ~n7847 ) | ( n7738 & ~n7847 ) ;
  assign n7849 = n7847 | n7848 ;
  assign n7850 = ~x95 & n7849 ;
  assign n7851 = n7811 | n7850 ;
  assign n7852 = ~n7796 & n7851 ;
  assign n7853 = x40 | n5075 ;
  assign n7854 = n7735 | n7784 ;
  assign n7855 = n7794 | n7854 ;
  assign n7856 = n7853 | n7855 ;
  assign n7857 = ~n7796 & n7856 ;
  assign n7858 = n7852 ^ x183 ^ 1'b0 ;
  assign n7859 = ( n7852 & n7857 ) | ( n7852 & ~n7858 ) | ( n7857 & ~n7858 ) ;
  assign n7860 = x174 & ~n7859 ;
  assign n7861 = x180 & ~n7860 ;
  assign n7862 = n7841 & n7861 ;
  assign n7863 = x183 & ~n5075 ;
  assign n7864 = n7795 & ~n7863 ;
  assign n7865 = n7737 | n7850 ;
  assign n7866 = ~n5075 & n7865 ;
  assign n7867 = x183 & n7866 ;
  assign n7868 = x174 & ~n7867 ;
  assign n7869 = n7868 ^ n7864 ^ 1'b0 ;
  assign n7870 = ( n7864 & n7868 ) | ( n7864 & n7869 ) | ( n7868 & n7869 ) ;
  assign n7871 = ( x180 & ~n7864 ) | ( x180 & n7870 ) | ( ~n7864 & n7870 ) ;
  assign n7872 = x174 | n7737 ;
  assign n7873 = ~x95 & n7840 ;
  assign n7874 = ( ~n7871 & n7872 ) | ( ~n7871 & n7873 ) | ( n7872 & n7873 ) ;
  assign n7875 = ~n7871 & n7874 ;
  assign n7876 = ( ~x193 & n7862 ) | ( ~x193 & n7875 ) | ( n7862 & n7875 ) ;
  assign n7877 = ~x193 & n7876 ;
  assign n7878 = n1225 | n1268 ;
  assign n7879 = n1230 & n7878 ;
  assign n7880 = ~n6387 & n7799 ;
  assign n7881 = ( ~x70 & n7879 ) | ( ~x70 & n7880 ) | ( n7879 & n7880 ) ;
  assign n7882 = ~x70 & n7881 ;
  assign n7883 = ( ~x51 & n7741 ) | ( ~x51 & n7882 ) | ( n7741 & n7882 ) ;
  assign n7884 = ~x51 & n7883 ;
  assign n7885 = ( ~n7739 & n7779 ) | ( ~n7739 & n7884 ) | ( n7779 & n7884 ) ;
  assign n7886 = ~n7739 & n7885 ;
  assign n7887 = ~x40 & n7886 ;
  assign n7888 = ( ~x32 & x40 ) | ( ~x32 & n7887 ) | ( x40 & n7887 ) ;
  assign n7889 = ( ~x95 & n7738 ) | ( ~x95 & n7888 ) | ( n7738 & n7888 ) ;
  assign n7890 = n7735 | n7889 ;
  assign n7891 = n7890 ^ n7813 ^ x40 ;
  assign n7892 = ~n7813 & n7891 ;
  assign n7893 = x32 | n7887 ;
  assign n7894 = n7814 ^ n7789 ^ n7738 ;
  assign n7895 = n7893 & ~n7894 ;
  assign n7896 = x95 | n7895 ;
  assign n7897 = ~n7813 & n7896 ;
  assign n7898 = n7892 ^ x198 ^ 1'b0 ;
  assign n7899 = ( n7892 & n7897 ) | ( n7892 & ~n7898 ) | ( n7897 & ~n7898 ) ;
  assign n7900 = n7853 | n7899 ;
  assign n7901 = ~n7796 & n7900 ;
  assign n7902 = x183 | n7901 ;
  assign n7903 = n5075 | n7569 ;
  assign n7904 = ~n7796 & n7903 ;
  assign n7905 = x183 & ~n7904 ;
  assign n7906 = ( x174 & n7902 ) | ( x174 & ~n7905 ) | ( n7902 & ~n7905 ) ;
  assign n7907 = ~x174 & n7906 ;
  assign n7908 = n7511 | n7786 ;
  assign n7909 = x32 | n7908 ;
  assign n7910 = n7763 & ~n7909 ;
  assign n7911 = n7569 | n7910 ;
  assign n7912 = ~x95 & n7911 ;
  assign n7913 = n7811 | n7912 ;
  assign n7914 = ~n7796 & n7913 ;
  assign n7915 = x183 & ~n7914 ;
  assign n7916 = ~n6387 & n7772 ;
  assign n7917 = n7879 | n7916 ;
  assign n7918 = x70 | n7917 ;
  assign n7919 = ( ~x70 & n7741 ) | ( ~x70 & n7918 ) | ( n7741 & n7918 ) ;
  assign n7920 = x51 | n7919 ;
  assign n7921 = ( ~x51 & n7779 ) | ( ~x51 & n7920 ) | ( n7779 & n7920 ) ;
  assign n7922 = x40 | n7739 ;
  assign n7923 = ( x32 & n7921 ) | ( x32 & ~n7922 ) | ( n7921 & ~n7922 ) ;
  assign n7924 = n7923 ^ n7921 ^ 1'b0 ;
  assign n7925 = ( x32 & n7923 ) | ( x32 & ~n7924 ) | ( n7923 & ~n7924 ) ;
  assign n7926 = ~n7814 & n7925 ;
  assign n7927 = n1652 & n7569 ;
  assign n7928 = ( ~x95 & n7926 ) | ( ~x95 & n7927 ) | ( n7926 & n7927 ) ;
  assign n7929 = ~x95 & n7928 ;
  assign n7930 = n7735 | n7929 ;
  assign n7931 = ~n7894 & n7925 ;
  assign n7932 = x95 | n7931 ;
  assign n7933 = ~n7813 & n7932 ;
  assign n7934 = n7930 | n7933 ;
  assign n7935 = ~x198 & n7934 ;
  assign n7936 = n5075 | n7935 ;
  assign n7937 = n7930 | n7936 ;
  assign n7938 = ~n7796 & n7937 ;
  assign n7939 = x183 | n7938 ;
  assign n7940 = ( x174 & n7915 ) | ( x174 & n7939 ) | ( n7915 & n7939 ) ;
  assign n7941 = ~n7915 & n7940 ;
  assign n7942 = ( x180 & n7907 ) | ( x180 & ~n7941 ) | ( n7907 & ~n7941 ) ;
  assign n7943 = ~n7907 & n7942 ;
  assign n7944 = n7737 | n7819 ;
  assign n7945 = n5075 | n7944 ;
  assign n7946 = ~n7796 & n7945 ;
  assign n7947 = x183 & ~n7946 ;
  assign n7948 = n7737 | n7889 ;
  assign n7949 = ( ~x95 & n7789 ) | ( ~x95 & n7888 ) | ( n7789 & n7888 ) ;
  assign n7950 = ~x198 & n7949 ;
  assign n7951 = n7948 | n7950 ;
  assign n7952 = n7795 ^ n5075 ^ 1'b0 ;
  assign n7953 = ( n7795 & n7951 ) | ( n7795 & ~n7952 ) | ( n7951 & ~n7952 ) ;
  assign n7954 = x183 | n7953 ;
  assign n7955 = ( x174 & ~n7947 ) | ( x174 & n7954 ) | ( ~n7947 & n7954 ) ;
  assign n7956 = ~x174 & n7955 ;
  assign n7957 = n5075 | n7912 ;
  assign n7958 = n7737 | n7957 ;
  assign n7959 = ~n7796 & n7958 ;
  assign n7960 = x183 & ~n7959 ;
  assign n7961 = x174 & ~n7960 ;
  assign n7962 = n7737 | n7929 ;
  assign n7963 = ~n5075 & n7569 ;
  assign n7964 = n7936 & ~n7963 ;
  assign n7965 = n7962 | n7964 ;
  assign n7966 = ~n7796 & n7965 ;
  assign n7967 = x183 | n7966 ;
  assign n7968 = n7961 & n7967 ;
  assign n7969 = ( x180 & ~n7956 ) | ( x180 & n7968 ) | ( ~n7956 & n7968 ) ;
  assign n7970 = n7956 | n7969 ;
  assign n7971 = ( x193 & n7943 ) | ( x193 & n7970 ) | ( n7943 & n7970 ) ;
  assign n7972 = ~n7943 & n7971 ;
  assign n7973 = ( ~x299 & n7877 ) | ( ~x299 & n7972 ) | ( n7877 & n7972 ) ;
  assign n7974 = ~x299 & n7973 ;
  assign n7975 = ~x210 & n7790 ;
  assign n7976 = n7785 | n7975 ;
  assign n7977 = n5075 & ~n7976 ;
  assign n7978 = n7945 & ~n7977 ;
  assign n7979 = x152 | n7978 ;
  assign n7980 = ~n5075 & n7976 ;
  assign n7981 = n7980 ^ n7976 ^ n7866 ;
  assign n7982 = x152 & ~n7981 ;
  assign n7983 = n7737 | n7836 ;
  assign n7984 = n5075 | n7983 ;
  assign n7985 = ~n7977 & n7984 ;
  assign n7986 = x152 | n7985 ;
  assign n7987 = ( x172 & ~n7982 ) | ( x172 & n7986 ) | ( ~n7982 & n7986 ) ;
  assign n7988 = ~x172 & n7987 ;
  assign n7989 = n7958 & ~n7977 ;
  assign n7990 = x152 & ~n7989 ;
  assign n7991 = x172 & ~n7990 ;
  assign n7992 = n7988 ^ n7979 ^ 1'b0 ;
  assign n7993 = ( ~n7979 & n7991 ) | ( ~n7979 & n7992 ) | ( n7991 & n7992 ) ;
  assign n7994 = ( n7979 & n7988 ) | ( n7979 & n7993 ) | ( n7988 & n7993 ) ;
  assign n7995 = ( x158 & x299 ) | ( x158 & n7994 ) | ( x299 & n7994 ) ;
  assign n7996 = ~x158 & n7995 ;
  assign n7997 = n7837 & ~n7977 ;
  assign n7998 = x152 | n7997 ;
  assign n7999 = n7913 & ~n7977 ;
  assign n8000 = x152 & ~n7999 ;
  assign n8001 = n7903 & ~n7977 ;
  assign n8002 = x152 | n8001 ;
  assign n8003 = ( x172 & n8000 ) | ( x172 & n8002 ) | ( n8000 & n8002 ) ;
  assign n8004 = ~n8000 & n8003 ;
  assign n8005 = n7851 & ~n7977 ;
  assign n8006 = x152 & ~n8005 ;
  assign n8007 = x172 | n8006 ;
  assign n8008 = ~n8004 & n8007 ;
  assign n8009 = ( n7998 & n8004 ) | ( n7998 & ~n8008 ) | ( n8004 & ~n8008 ) ;
  assign n8010 = ( ~x158 & x299 ) | ( ~x158 & n8009 ) | ( x299 & n8009 ) ;
  assign n8011 = x158 & n8010 ;
  assign n8012 = ( x149 & n7996 ) | ( x149 & ~n8011 ) | ( n7996 & ~n8011 ) ;
  assign n8013 = ~n7996 & n8012 ;
  assign n8014 = ~x210 & n7809 ;
  assign n8015 = n7821 | n8014 ;
  assign n8016 = ~n7977 & n8015 ;
  assign n8017 = x152 | n8016 ;
  assign n8018 = ~x172 & n8017 ;
  assign n8019 = ~x210 & n7934 ;
  assign n8020 = n5075 | n8019 ;
  assign n8021 = n7930 | n8020 ;
  assign n8022 = ~n7977 & n8021 ;
  assign n8023 = x152 & ~n8022 ;
  assign n8024 = n7735 | n7949 ;
  assign n8025 = x210 | n8024 ;
  assign n8026 = ( ~x210 & n5075 ) | ( ~x210 & n8025 ) | ( n5075 & n8025 ) ;
  assign n8027 = ( n7890 & ~n7977 ) | ( n7890 & n8026 ) | ( ~n7977 & n8026 ) ;
  assign n8028 = ~n7977 & n8027 ;
  assign n8029 = x152 | n8028 ;
  assign n8030 = ( x172 & n8023 ) | ( x172 & n8029 ) | ( n8023 & n8029 ) ;
  assign n8031 = ~n8023 & n8030 ;
  assign n8032 = n7854 | n7975 ;
  assign n8033 = n5075 | n8032 ;
  assign n8034 = ~n7977 & n8033 ;
  assign n8035 = x152 & ~n8034 ;
  assign n8036 = ~n8031 & n8035 ;
  assign n8037 = ( n8018 & n8031 ) | ( n8018 & ~n8036 ) | ( n8031 & ~n8036 ) ;
  assign n8038 = ( ~x158 & x299 ) | ( ~x158 & n8037 ) | ( x299 & n8037 ) ;
  assign n8039 = x158 & n8038 ;
  assign n8040 = ~n7963 & n8026 ;
  assign n8041 = n7948 | n8040 ;
  assign n8042 = ~x152 & n8041 ;
  assign n8043 = ~n7963 & n8020 ;
  assign n8044 = n7962 | n8043 ;
  assign n8045 = x152 & n8044 ;
  assign n8046 = ( x172 & n8042 ) | ( x172 & ~n8045 ) | ( n8042 & ~n8045 ) ;
  assign n8047 = ~n8042 & n8046 ;
  assign n8048 = ~x158 & x299 ;
  assign n8049 = n7737 | n7820 ;
  assign n8050 = n8014 | n8049 ;
  assign n8051 = n5075 | n8050 ;
  assign n8052 = ~x152 & n8051 ;
  assign n8053 = x152 & n7976 ;
  assign n8054 = ( x172 & ~n8052 ) | ( x172 & n8053 ) | ( ~n8052 & n8053 ) ;
  assign n8055 = n8052 | n8054 ;
  assign n8056 = ( n7977 & n8048 ) | ( n7977 & n8055 ) | ( n8048 & n8055 ) ;
  assign n8057 = ~n7977 & n8056 ;
  assign n8058 = n8057 ^ n8047 ^ 1'b0 ;
  assign n8059 = ( n8047 & n8057 ) | ( n8047 & n8058 ) | ( n8057 & n8058 ) ;
  assign n8060 = ( x149 & ~n8047 ) | ( x149 & n8059 ) | ( ~n8047 & n8059 ) ;
  assign n8061 = ( ~n8013 & n8039 ) | ( ~n8013 & n8060 ) | ( n8039 & n8060 ) ;
  assign n8062 = ~n8013 & n8061 ;
  assign n8063 = ( x232 & n7974 ) | ( x232 & n8062 ) | ( n7974 & n8062 ) ;
  assign n8064 = n8062 ^ n7974 ^ 1'b0 ;
  assign n8065 = ( x232 & n8063 ) | ( x232 & n8064 ) | ( n8063 & n8064 ) ;
  assign n8066 = ( x39 & ~n7793 ) | ( x39 & n8065 ) | ( ~n7793 & n8065 ) ;
  assign n8067 = n7793 | n8066 ;
  assign n8068 = n8067 ^ n7731 ^ 1'b0 ;
  assign n8069 = ( n7731 & n8067 ) | ( n7731 & n8068 ) | ( n8067 & n8068 ) ;
  assign n8070 = ( x38 & ~n7731 ) | ( x38 & n8069 ) | ( ~n7731 & n8069 ) ;
  assign n8071 = n8070 ^ n7668 ^ 1'b0 ;
  assign n8072 = ( n7668 & n8070 ) | ( n7668 & n8071 ) | ( n8070 & n8071 ) ;
  assign n8073 = ( x100 & ~n7668 ) | ( x100 & n8072 ) | ( ~n7668 & n8072 ) ;
  assign n8074 = ( x87 & ~n7624 ) | ( x87 & n8073 ) | ( ~n7624 & n8073 ) ;
  assign n8075 = ~x87 & n8074 ;
  assign n8076 = ( n2053 & ~n7654 ) | ( n2053 & n8075 ) | ( ~n7654 & n8075 ) ;
  assign n8077 = n7654 | n8076 ;
  assign n8078 = ( n7625 & ~n7652 ) | ( n7625 & n8077 ) | ( ~n7652 & n8077 ) ;
  assign n8079 = ~n7625 & n8078 ;
  assign n8080 = n8079 ^ x54 ^ 1'b0 ;
  assign n8081 = ( ~n7638 & n8079 ) | ( ~n7638 & n8080 ) | ( n8079 & n8080 ) ;
  assign n8082 = x74 | n8081 ;
  assign n8083 = ~n7633 & n8082 ;
  assign n8084 = ( n2109 & ~n7614 ) | ( n2109 & n8083 ) | ( ~n7614 & n8083 ) ;
  assign n8085 = n7614 | n8084 ;
  assign n8086 = ( n7568 & ~n7573 ) | ( n7568 & n8085 ) | ( ~n7573 & n8085 ) ;
  assign n8087 = ~n7568 & n8086 ;
  assign n8088 = ~x74 & n7561 ;
  assign n8089 = n2120 & ~n8088 ;
  assign n8090 = ( ~n7559 & n8087 ) | ( ~n7559 & n8089 ) | ( n8087 & n8089 ) ;
  assign n8091 = n8087 ^ n7559 ^ 1'b0 ;
  assign n8092 = ( n8087 & n8090 ) | ( n8087 & ~n8091 ) | ( n8090 & ~n8091 ) ;
  assign n8093 = ~x33 & n8092 ;
  assign n8094 = ~n7559 & n8089 ;
  assign n8095 = x54 & n7638 ;
  assign n8096 = n1788 & ~n5075 ;
  assign n8097 = x180 & n8096 ;
  assign n8098 = n1289 | n5075 ;
  assign n8099 = x40 | n8098 ;
  assign n8100 = x90 | n5141 ;
  assign n8101 = x72 | x93 ;
  assign n8102 = n1377 | n8101 ;
  assign n8103 = x90 & n6374 ;
  assign n8104 = n8102 | n8103 ;
  assign n8105 = n8100 & ~n8104 ;
  assign n8106 = ~n8099 & n8105 ;
  assign n8107 = ~x183 & n8106 ;
  assign n8108 = n1290 | n1694 ;
  assign n8109 = ~n1268 & n8100 ;
  assign n8110 = ~n8103 & n8109 ;
  assign n8111 = x90 | n1395 ;
  assign n8112 = n1268 | n8111 ;
  assign n8113 = n1390 | n8112 ;
  assign n8114 = n7751 & ~n8113 ;
  assign n8115 = x70 | n8114 ;
  assign n8116 = ~n8108 & n8115 ;
  assign n8117 = ( ~n8108 & n8110 ) | ( ~n8108 & n8116 ) | ( n8110 & n8116 ) ;
  assign n8118 = n5286 | n8117 ;
  assign n8119 = ~n5075 & n8118 ;
  assign n8120 = x183 & n8119 ;
  assign n8121 = ( x174 & n8107 ) | ( x174 & ~n8120 ) | ( n8107 & ~n8120 ) ;
  assign n8122 = ~n8107 & n8121 ;
  assign n8123 = n1230 | n8113 ;
  assign n8124 = n7767 & ~n8123 ;
  assign n8125 = x70 | n8124 ;
  assign n8126 = ~n8108 & n8125 ;
  assign n8127 = n5285 | n8126 ;
  assign n8128 = ~x198 & n8127 ;
  assign n8129 = ( ~n8108 & n8110 ) | ( ~n8108 & n8126 ) | ( n8110 & n8126 ) ;
  assign n8130 = n8128 | n8129 ;
  assign n8131 = n7863 & n8130 ;
  assign n8132 = ~n1230 & n7842 ;
  assign n8133 = ( ~n8104 & n8105 ) | ( ~n8104 & n8132 ) | ( n8105 & n8132 ) ;
  assign n8134 = ~n8099 & n8133 ;
  assign n8135 = ~x183 & n8134 ;
  assign n8136 = ( x174 & ~n8131 ) | ( x174 & n8135 ) | ( ~n8131 & n8135 ) ;
  assign n8137 = n8131 | n8136 ;
  assign n8138 = x193 & ~n8137 ;
  assign n8139 = ( x193 & n8122 ) | ( x193 & n8138 ) | ( n8122 & n8138 ) ;
  assign n8140 = n5286 | n8116 ;
  assign n8141 = x174 & ~n8140 ;
  assign n8142 = n7863 & ~n8141 ;
  assign n8143 = n5286 | n8126 ;
  assign n8144 = x174 | n8143 ;
  assign n8145 = n8142 & n8144 ;
  assign n8146 = ~n7786 & n8132 ;
  assign n8147 = ~n1289 & n8146 ;
  assign n8148 = ~n7853 & n8147 ;
  assign n8149 = x174 | x183 ;
  assign n8150 = n8148 & ~n8149 ;
  assign n8151 = x193 | n8150 ;
  assign n8152 = ( ~n8139 & n8145 ) | ( ~n8139 & n8151 ) | ( n8145 & n8151 ) ;
  assign n8153 = ~n8139 & n8152 ;
  assign n8154 = ( x299 & ~n8097 ) | ( x299 & n8153 ) | ( ~n8097 & n8153 ) ;
  assign n8155 = n8097 | n8154 ;
  assign n8156 = ~x39 & x232 ;
  assign n8157 = n5295 | n8116 ;
  assign n8158 = x172 & n8117 ;
  assign n8159 = x152 & ~n8158 ;
  assign n8160 = ~n8157 & n8159 ;
  assign n8161 = ( x149 & n5075 ) | ( x149 & ~n8160 ) | ( n5075 & ~n8160 ) ;
  assign n8162 = ~n5075 & n8161 ;
  assign n8165 = x172 & n8129 ;
  assign n8163 = n5295 | n8126 ;
  assign n8164 = x152 | n8163 ;
  assign n8166 = n8165 ^ n8164 ^ 1'b0 ;
  assign n8167 = ( n8164 & n8165 ) | ( n8164 & ~n8166 ) | ( n8165 & ~n8166 ) ;
  assign n8168 = ( n8162 & n8166 ) | ( n8162 & n8167 ) | ( n8166 & n8167 ) ;
  assign n8169 = x158 & n8096 ;
  assign n8170 = x299 & ~n8169 ;
  assign n8171 = x152 | x172 ;
  assign n8172 = n8148 & ~n8171 ;
  assign n8173 = ~x152 & n8134 ;
  assign n8174 = n8106 | n8173 ;
  assign n8175 = x172 & n8174 ;
  assign n8176 = ( ~x149 & n8172 ) | ( ~x149 & n8175 ) | ( n8172 & n8175 ) ;
  assign n8177 = ~x149 & n8176 ;
  assign n8178 = ( n8168 & n8170 ) | ( n8168 & ~n8177 ) | ( n8170 & ~n8177 ) ;
  assign n8179 = ~n8168 & n8178 ;
  assign n8180 = n8156 & ~n8179 ;
  assign n8181 = n8155 & n8180 ;
  assign n8182 = n5379 & n7689 ;
  assign n8183 = x154 | n8182 ;
  assign n8184 = n5374 & n7689 ;
  assign n8185 = x154 & ~n8184 ;
  assign n8186 = ( x152 & n8183 ) | ( x152 & ~n8185 ) | ( n8183 & ~n8185 ) ;
  assign n8187 = ~x152 & n8186 ;
  assign n8188 = ~n5075 & n6460 ;
  assign n8189 = n5061 & n8188 ;
  assign n8190 = n8189 ^ n8187 ^ 1'b0 ;
  assign n8191 = x152 & x154 ;
  assign n8192 = ( n8189 & ~n8190 ) | ( n8189 & n8191 ) | ( ~n8190 & n8191 ) ;
  assign n8193 = ( n8187 & n8190 ) | ( n8187 & n8192 ) | ( n8190 & n8192 ) ;
  assign n8194 = x299 & ~n8193 ;
  assign n8195 = ( x299 & ~n7669 ) | ( x299 & n8194 ) | ( ~n7669 & n8194 ) ;
  assign n8196 = n5379 & n7723 ;
  assign n8197 = n7678 & n8196 ;
  assign n8198 = ~x174 & n8197 ;
  assign n8199 = ( x299 & n7721 ) | ( x299 & n8198 ) | ( n7721 & n8198 ) ;
  assign n8200 = n7721 & n8199 ;
  assign n8201 = n5374 & n7678 ;
  assign n8202 = n7723 & n8201 ;
  assign n8203 = ~x174 & n8202 ;
  assign n8204 = n7678 & n7723 ;
  assign n8205 = n6460 & n8204 ;
  assign n8206 = x174 & n8205 ;
  assign n8207 = ( x299 & ~n8203 ) | ( x299 & n8206 ) | ( ~n8203 & n8206 ) ;
  assign n8208 = n8203 | n8207 ;
  assign n8209 = n8200 ^ n7712 ^ 1'b0 ;
  assign n8210 = ( ~n7712 & n8208 ) | ( ~n7712 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = ( n7712 & n8200 ) | ( n7712 & n8210 ) | ( n8200 & n8210 ) ;
  assign n8212 = ( x39 & n8195 ) | ( x39 & n8211 ) | ( n8195 & n8211 ) ;
  assign n8213 = ~n8195 & n8212 ;
  assign n8214 = ( ~x38 & n8181 ) | ( ~x38 & n8213 ) | ( n8181 & n8213 ) ;
  assign n8215 = ~x38 & n8214 ;
  assign n8216 = ( x87 & n7668 ) | ( x87 & ~n8215 ) | ( n7668 & ~n8215 ) ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = x87 & ~n7640 ;
  assign n8219 = ( x100 & n8217 ) | ( x100 & ~n8218 ) | ( n8217 & ~n8218 ) ;
  assign n8220 = ~x100 & n8219 ;
  assign n8221 = ( ~n2053 & n7624 ) | ( ~n2053 & n8220 ) | ( n7624 & n8220 ) ;
  assign n8222 = ~n2053 & n8221 ;
  assign n8223 = x38 | x87 ;
  assign n8224 = x100 | n8223 ;
  assign n8225 = ( n5052 & n7647 ) | ( n5052 & ~n8224 ) | ( n7647 & ~n8224 ) ;
  assign n8226 = ~n5052 & n8225 ;
  assign n8227 = ( n7639 & n7642 ) | ( n7639 & n8226 ) | ( n7642 & n8226 ) ;
  assign n8228 = n7639 & n8227 ;
  assign n8229 = ( n7625 & ~n8222 ) | ( n7625 & n8228 ) | ( ~n8222 & n8228 ) ;
  assign n8230 = n8222 | n8229 ;
  assign n8231 = x54 | n8230 ;
  assign n8232 = ( ~x54 & n8095 ) | ( ~x54 & n8231 ) | ( n8095 & n8231 ) ;
  assign n8233 = x74 | n8232 ;
  assign n8234 = ( ~x74 & n7633 ) | ( ~x74 & n8233 ) | ( n7633 & n8233 ) ;
  assign n8235 = ~n5052 & n7599 ;
  assign n8236 = x38 | n8235 ;
  assign n8237 = ~n7585 & n8236 ;
  assign n8238 = x38 & n7575 ;
  assign n8239 = n6512 & n8238 ;
  assign n8240 = ( n7553 & ~n8237 ) | ( n7553 & n8239 ) | ( ~n8237 & n8239 ) ;
  assign n8241 = n8237 | n8240 ;
  assign n8242 = x75 | n8241 ;
  assign n8243 = ( ~x75 & n7584 ) | ( ~x75 & n8242 ) | ( n7584 & n8242 ) ;
  assign n8244 = x92 & ~n7563 ;
  assign n8245 = ( x54 & n8243 ) | ( x54 & ~n8244 ) | ( n8243 & ~n8244 ) ;
  assign n8246 = ~x54 & n8245 ;
  assign n8247 = ( ~x74 & n7562 ) | ( ~x74 & n8246 ) | ( n7562 & n8246 ) ;
  assign n8248 = ~x74 & n8247 ;
  assign n8249 = ( x55 & n7559 ) | ( x55 & ~n8248 ) | ( n7559 & ~n8248 ) ;
  assign n8250 = ~n7559 & n8249 ;
  assign n8251 = ( n2109 & n8234 ) | ( n2109 & ~n8250 ) | ( n8234 & ~n8250 ) ;
  assign n8252 = ~n2109 & n8251 ;
  assign n8253 = ( n7568 & ~n8094 ) | ( n7568 & n8252 ) | ( ~n8094 & n8252 ) ;
  assign n8254 = ~n8094 & n8253 ;
  assign n8255 = x33 & ~n8254 ;
  assign n8256 = ( x954 & n8093 ) | ( x954 & ~n8255 ) | ( n8093 & ~n8255 ) ;
  assign n8257 = ~n8093 & n8256 ;
  assign n8258 = x195 | x196 ;
  assign n8259 = x138 | n8258 ;
  assign n8260 = x139 | n8259 ;
  assign n8261 = x118 | n8260 ;
  assign n8262 = x79 | n8261 ;
  assign n8263 = x34 | n8262 ;
  assign n8264 = ~x33 & n8263 ;
  assign n8265 = n8092 & ~n8264 ;
  assign n8266 = ~n8254 & n8264 ;
  assign n8267 = x954 | n8266 ;
  assign n8268 = ( ~n8257 & n8265 ) | ( ~n8257 & n8267 ) | ( n8265 & n8267 ) ;
  assign n8269 = ~n8257 & n8268 ;
  assign n8270 = x162 & ~n5075 ;
  assign n8271 = x197 & ~n7547 ;
  assign n8272 = n8270 & n8271 ;
  assign n8273 = x162 | x197 ;
  assign n8274 = n7548 & n8273 ;
  assign n8275 = n5075 | n8274 ;
  assign n8276 = n8272 | n8275 ;
  assign n8277 = n8270 ^ n7547 ^ x197 ;
  assign n8278 = ( n8270 & ~n8276 ) | ( n8270 & n8277 ) | ( ~n8276 & n8277 ) ;
  assign n8279 = x232 & n8278 ;
  assign n8280 = n7555 & n8279 ;
  assign n8281 = x148 & n7556 ;
  assign n8282 = ( x74 & n8280 ) | ( x74 & ~n8281 ) | ( n8280 & ~n8281 ) ;
  assign n8283 = ~n8280 & n8282 ;
  assign n8284 = x167 & n6411 ;
  assign n8285 = ~n7555 & n8284 ;
  assign n8286 = n8280 | n8285 ;
  assign n8287 = x74 | n8286 ;
  assign n8288 = ~n8283 & n8287 ;
  assign n8289 = n2120 & n8288 ;
  assign n8290 = x54 | n8280 ;
  assign n8291 = x38 & n8285 ;
  assign n8292 = n8290 | n8291 ;
  assign n8293 = x74 | n8292 ;
  assign n8294 = n2109 & ~n8293 ;
  assign n8295 = ( n2109 & ~n8288 ) | ( n2109 & n8294 ) | ( ~n8288 & n8294 ) ;
  assign n8296 = ( x57 & x59 ) | ( x57 & ~n8295 ) | ( x59 & ~n8295 ) ;
  assign n8297 = n8295 | n8296 ;
  assign n8298 = ( n2120 & n7446 ) | ( n2120 & n7572 ) | ( n7446 & n7572 ) ;
  assign n8299 = n8297 & n8298 ;
  assign n8300 = x140 & x145 ;
  assign n8301 = x140 | x145 ;
  assign n8302 = ~n8300 & n8301 ;
  assign n8303 = n7619 & ~n8302 ;
  assign n8304 = n7618 | n8300 ;
  assign n8305 = ~n5075 & n8301 ;
  assign n8306 = ~n8304 & n8305 ;
  assign n8307 = x299 | n8306 ;
  assign n8308 = ( x232 & n8303 ) | ( x232 & n8307 ) | ( n8303 & n8307 ) ;
  assign n8309 = n8307 ^ n8303 ^ 1'b0 ;
  assign n8310 = ( x232 & n8308 ) | ( x232 & n8309 ) | ( n8308 & n8309 ) ;
  assign n8311 = n8310 ^ n8278 ^ 1'b0 ;
  assign n8312 = ( ~x299 & n8278 ) | ( ~x299 & n8311 ) | ( n8278 & n8311 ) ;
  assign n8313 = ( n8310 & ~n8311 ) | ( n8310 & n8312 ) | ( ~n8311 & n8312 ) ;
  assign n8314 = x100 & ~n8313 ;
  assign n8315 = x75 & ~n8313 ;
  assign n8316 = n8314 | n8315 ;
  assign n8317 = x141 & ~x299 ;
  assign n8318 = x148 & x299 ;
  assign n8319 = n8317 | n8318 ;
  assign n8320 = n6411 & n8319 ;
  assign n8321 = n7555 | n8320 ;
  assign n8322 = ~n8316 & n8321 ;
  assign n8323 = ( x55 & x74 ) | ( x55 & ~n8322 ) | ( x74 & ~n8322 ) ;
  assign n8324 = n8323 ^ x74 ^ 1'b0 ;
  assign n8325 = ( x55 & n8323 ) | ( x55 & ~n8324 ) | ( n8323 & ~n8324 ) ;
  assign n8326 = x299 ^ x167 ^ 1'b0 ;
  assign n8327 = ( x167 & x188 ) | ( x167 & ~n8326 ) | ( x188 & ~n8326 ) ;
  assign n8328 = n6411 & n8327 ;
  assign n8329 = x38 & n8328 ;
  assign n8330 = n7570 & ~n8329 ;
  assign n8331 = x87 & ~n8330 ;
  assign n8332 = x188 & n7656 ;
  assign n8333 = x167 | n8332 ;
  assign n8334 = x167 & x188 ;
  assign n8335 = ~n7659 & n8334 ;
  assign n8336 = ( x188 & n7662 ) | ( x188 & ~n8335 ) | ( n7662 & ~n8335 ) ;
  assign n8337 = ~n8335 & n8336 ;
  assign n8338 = x38 & ~n8337 ;
  assign n8339 = ( x38 & ~n8333 ) | ( x38 & n8338 ) | ( ~n8333 & n8338 ) ;
  assign n8340 = x87 | n8339 ;
  assign n8341 = x142 & ~n7852 ;
  assign n8342 = x142 | n7914 ;
  assign n8343 = ( x140 & n8341 ) | ( x140 & n8342 ) | ( n8341 & n8342 ) ;
  assign n8344 = ~n8341 & n8343 ;
  assign n8345 = x142 | n7938 ;
  assign n8346 = x142 & ~n7857 ;
  assign n8347 = ( x140 & n8345 ) | ( x140 & ~n8346 ) | ( n8345 & ~n8346 ) ;
  assign n8348 = ~x140 & n8347 ;
  assign n8349 = ( x181 & n8344 ) | ( x181 & n8348 ) | ( n8344 & n8348 ) ;
  assign n8350 = n8348 ^ n8344 ^ 1'b0 ;
  assign n8351 = ( x181 & n8349 ) | ( x181 & n8350 ) | ( n8349 & n8350 ) ;
  assign n8352 = x142 & ~n7795 ;
  assign n8353 = x140 | n8352 ;
  assign n8354 = ( x142 & n7966 ) | ( x142 & ~n8353 ) | ( n7966 & ~n8353 ) ;
  assign n8355 = ~n8353 & n8354 ;
  assign n8356 = n5075 & n7795 ;
  assign n8357 = x142 & ~n7866 ;
  assign n8358 = ~n8356 & n8357 ;
  assign n8359 = x140 & ~n8358 ;
  assign n8360 = x142 | n7959 ;
  assign n8361 = n8359 & n8360 ;
  assign n8362 = ( ~x181 & n8355 ) | ( ~x181 & n8361 ) | ( n8355 & n8361 ) ;
  assign n8363 = ~x181 & n8362 ;
  assign n8364 = ( x144 & n8351 ) | ( x144 & ~n8363 ) | ( n8351 & ~n8363 ) ;
  assign n8365 = ~n8351 & n8364 ;
  assign n8366 = x142 | n7953 ;
  assign n8367 = n7810 | n8049 ;
  assign n8368 = ~n5075 & n8367 ;
  assign n8369 = ( x142 & n8356 ) | ( x142 & ~n8368 ) | ( n8356 & ~n8368 ) ;
  assign n8370 = ~n8356 & n8369 ;
  assign n8371 = ( x140 & n8366 ) | ( x140 & ~n8370 ) | ( n8366 & ~n8370 ) ;
  assign n8372 = ~x140 & n8371 ;
  assign n8373 = ( x142 & n7796 ) | ( x142 & ~n7984 ) | ( n7796 & ~n7984 ) ;
  assign n8374 = x140 & ~n8373 ;
  assign n8375 = x142 | n7946 ;
  assign n8376 = n8374 & n8375 ;
  assign n8377 = ( ~x181 & n8372 ) | ( ~x181 & n8376 ) | ( n8372 & n8376 ) ;
  assign n8378 = ~x181 & n8377 ;
  assign n8379 = x142 & ~n7823 ;
  assign n8380 = x140 | n8379 ;
  assign n8381 = ( x142 & n7901 ) | ( x142 & ~n8380 ) | ( n7901 & ~n8380 ) ;
  assign n8382 = ~n8380 & n8381 ;
  assign n8383 = x142 & ~n7838 ;
  assign n8384 = x142 | n7904 ;
  assign n8385 = ( x140 & n8383 ) | ( x140 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8386 = ~n8383 & n8385 ;
  assign n8387 = ( x181 & n8382 ) | ( x181 & n8386 ) | ( n8382 & n8386 ) ;
  assign n8388 = n8386 ^ n8382 ^ 1'b0 ;
  assign n8389 = ( x181 & n8387 ) | ( x181 & n8388 ) | ( n8387 & n8388 ) ;
  assign n8390 = ( x144 & ~n8378 ) | ( x144 & n8389 ) | ( ~n8378 & n8389 ) ;
  assign n8391 = n8378 | n8390 ;
  assign n8392 = ( x299 & ~n8365 ) | ( x299 & n8391 ) | ( ~n8365 & n8391 ) ;
  assign n8393 = ~x299 & n8392 ;
  assign n8394 = x146 | n7978 ;
  assign n8395 = x146 & ~n7985 ;
  assign n8396 = ( x161 & n8394 ) | ( x161 & ~n8395 ) | ( n8394 & ~n8395 ) ;
  assign n8397 = ~x161 & n8396 ;
  assign n8398 = x146 & ~n7981 ;
  assign n8399 = x146 | n7989 ;
  assign n8400 = ( x161 & n8398 ) | ( x161 & n8399 ) | ( n8398 & n8399 ) ;
  assign n8401 = ~n8398 & n8400 ;
  assign n8402 = ( x162 & n8397 ) | ( x162 & n8401 ) | ( n8397 & n8401 ) ;
  assign n8403 = n8401 ^ n8397 ^ 1'b0 ;
  assign n8404 = ( x162 & n8402 ) | ( x162 & n8403 ) | ( n8402 & n8403 ) ;
  assign n8405 = x161 & n8044 ;
  assign n8406 = ~x161 & n8041 ;
  assign n8407 = ( x146 & ~n8405 ) | ( x146 & n8406 ) | ( ~n8405 & n8406 ) ;
  assign n8408 = n8405 | n8407 ;
  assign n8409 = x161 & n7976 ;
  assign n8410 = ~x161 & n8051 ;
  assign n8411 = ( x146 & n8409 ) | ( x146 & ~n8410 ) | ( n8409 & ~n8410 ) ;
  assign n8412 = ~n8409 & n8411 ;
  assign n8413 = ( x162 & n7977 ) | ( x162 & ~n8412 ) | ( n7977 & ~n8412 ) ;
  assign n8414 = n8412 | n8413 ;
  assign n8415 = ( n8404 & n8408 ) | ( n8404 & ~n8414 ) | ( n8408 & ~n8414 ) ;
  assign n8416 = n8415 ^ n8408 ^ 1'b0 ;
  assign n8417 = ( n8404 & n8415 ) | ( n8404 & ~n8416 ) | ( n8415 & ~n8416 ) ;
  assign n8418 = ( x159 & x299 ) | ( x159 & n8417 ) | ( x299 & n8417 ) ;
  assign n8419 = ~x159 & n8418 ;
  assign n8420 = x146 & ~n7997 ;
  assign n8421 = x146 | n8001 ;
  assign n8422 = ( x161 & ~n8420 ) | ( x161 & n8421 ) | ( ~n8420 & n8421 ) ;
  assign n8423 = ~x161 & n8422 ;
  assign n8424 = x146 & ~n8005 ;
  assign n8425 = x146 | n7999 ;
  assign n8426 = ( x161 & n8424 ) | ( x161 & n8425 ) | ( n8424 & n8425 ) ;
  assign n8427 = ~n8424 & n8426 ;
  assign n8428 = ( x162 & n8423 ) | ( x162 & ~n8427 ) | ( n8423 & ~n8427 ) ;
  assign n8429 = ~n8423 & n8428 ;
  assign n8430 = x146 | n8022 ;
  assign n8431 = ~x146 & x161 ;
  assign n8432 = ( x161 & n8034 ) | ( x161 & n8431 ) | ( n8034 & n8431 ) ;
  assign n8433 = n8430 & n8432 ;
  assign n8434 = x146 | n8028 ;
  assign n8435 = x146 & ~n8016 ;
  assign n8436 = ( x161 & n8434 ) | ( x161 & ~n8435 ) | ( n8434 & ~n8435 ) ;
  assign n8437 = ~x161 & n8436 ;
  assign n8438 = ( x162 & ~n8433 ) | ( x162 & n8437 ) | ( ~n8433 & n8437 ) ;
  assign n8439 = n8433 | n8438 ;
  assign n8440 = ( ~x159 & x299 ) | ( ~x159 & n8439 ) | ( x299 & n8439 ) ;
  assign n8441 = x159 & n8440 ;
  assign n8442 = n8441 ^ n8429 ^ 1'b0 ;
  assign n8443 = ( n8429 & n8441 ) | ( n8429 & n8442 ) | ( n8441 & n8442 ) ;
  assign n8444 = ( n8419 & ~n8429 ) | ( n8419 & n8443 ) | ( ~n8429 & n8443 ) ;
  assign n8445 = ( x232 & n8393 ) | ( x232 & n8444 ) | ( n8393 & n8444 ) ;
  assign n8446 = n8444 ^ n8393 ^ 1'b0 ;
  assign n8447 = ( x232 & n8445 ) | ( x232 & n8446 ) | ( n8445 & n8446 ) ;
  assign n8448 = ( ~n1994 & n7793 ) | ( ~n1994 & n8447 ) | ( n7793 & n8447 ) ;
  assign n8449 = ~n1994 & n8448 ;
  assign n8450 = x177 | x299 ;
  assign n8451 = x144 | n7680 ;
  assign n8452 = n7726 | n8451 ;
  assign n8453 = x144 & ~n7716 ;
  assign n8454 = ( n8450 & n8452 ) | ( n8450 & ~n8453 ) | ( n8452 & ~n8453 ) ;
  assign n8455 = ~n8450 & n8454 ;
  assign n8456 = x177 & ~x299 ;
  assign n8457 = n8451 & n8456 ;
  assign n8458 = n7680 | n7685 ;
  assign n8459 = n8457 & n8458 ;
  assign n8460 = ( x232 & n8455 ) | ( x232 & n8459 ) | ( n8455 & n8459 ) ;
  assign n8461 = n8459 ^ n8455 ^ 1'b0 ;
  assign n8462 = ( x232 & n8460 ) | ( x232 & n8461 ) | ( n8460 & n8461 ) ;
  assign n8463 = ( ~x38 & n7719 ) | ( ~x38 & n8462 ) | ( n7719 & n8462 ) ;
  assign n8464 = ~x38 & n8463 ;
  assign n8465 = ~x38 & x155 ;
  assign n8466 = n7669 & ~n7677 ;
  assign n8467 = x161 & n7691 ;
  assign n8468 = n8466 & ~n8467 ;
  assign n8469 = n7671 & ~n8468 ;
  assign n8470 = n8465 & n8469 ;
  assign n8471 = x161 | n7700 ;
  assign n8472 = n7669 & ~n8471 ;
  assign n8473 = ( n7669 & ~n7705 ) | ( n7669 & n8472 ) | ( ~n7705 & n8472 ) ;
  assign n8474 = x38 | x155 ;
  assign n8475 = ( n7671 & n8473 ) | ( n7671 & ~n8474 ) | ( n8473 & ~n8474 ) ;
  assign n8476 = ~n8473 & n8475 ;
  assign n8477 = ( x232 & n8470 ) | ( x232 & n8476 ) | ( n8470 & n8476 ) ;
  assign n8478 = n8476 ^ n8470 ^ 1'b0 ;
  assign n8479 = ( x232 & n8477 ) | ( x232 & n8478 ) | ( n8477 & n8478 ) ;
  assign n8480 = ( x39 & n8464 ) | ( x39 & n8479 ) | ( n8464 & n8479 ) ;
  assign n8481 = n8479 ^ n8464 ^ 1'b0 ;
  assign n8482 = ( x39 & n8480 ) | ( x39 & n8481 ) | ( n8480 & n8481 ) ;
  assign n8483 = ( ~n8340 & n8449 ) | ( ~n8340 & n8482 ) | ( n8449 & n8482 ) ;
  assign n8484 = n8340 | n8483 ;
  assign n8485 = ( x100 & ~n8331 ) | ( x100 & n8484 ) | ( ~n8331 & n8484 ) ;
  assign n8486 = ~x100 & n8485 ;
  assign n8487 = ( ~n2053 & n8314 ) | ( ~n2053 & n8486 ) | ( n8314 & n8486 ) ;
  assign n8488 = ~n2053 & n8487 ;
  assign n8489 = n8313 ^ x100 ^ 1'b0 ;
  assign n8490 = ( x155 & n8450 ) | ( x155 & n8456 ) | ( n8450 & n8456 ) ;
  assign n8491 = x38 | n8490 ;
  assign n8492 = n6411 & n8491 ;
  assign n8493 = n7648 | n8492 ;
  assign n8494 = ~n8330 & n8493 ;
  assign n8495 = ( n8313 & ~n8489 ) | ( n8313 & n8494 ) | ( ~n8489 & n8494 ) ;
  assign n8496 = ( n7639 & n8315 ) | ( n7639 & ~n8495 ) | ( n8315 & ~n8495 ) ;
  assign n8497 = n8495 ^ n8315 ^ 1'b0 ;
  assign n8498 = ( n8315 & n8496 ) | ( n8315 & ~n8497 ) | ( n8496 & ~n8497 ) ;
  assign n8499 = ( ~x54 & n8488 ) | ( ~x54 & n8498 ) | ( n8488 & n8498 ) ;
  assign n8500 = ~x54 & n8499 ;
  assign n8501 = x100 | n8328 ;
  assign n8502 = x75 | n8501 ;
  assign n8503 = ~n8316 & n8502 ;
  assign n8504 = ~n8500 & n8503 ;
  assign n8505 = ( x54 & n8500 ) | ( x54 & ~n8504 ) | ( n8500 & ~n8504 ) ;
  assign n8506 = x74 | n8505 ;
  assign n8507 = ( ~x74 & n8325 ) | ( ~x74 & n8506 ) | ( n8325 & n8506 ) ;
  assign n8508 = x55 & ~n8283 ;
  assign n8509 = x54 & ~n8286 ;
  assign n8510 = x75 & ~n8279 ;
  assign n8511 = n7648 | n8270 ;
  assign n8512 = ~n7570 & n8511 ;
  assign n8513 = x100 | n8512 ;
  assign n8514 = n7648 ^ x232 ^ 1'b0 ;
  assign n8515 = ( x232 & n7648 ) | ( x232 & ~n8514 ) | ( n7648 & ~n8514 ) ;
  assign n8516 = ( n8513 & n8514 ) | ( n8513 & n8515 ) | ( n8514 & n8515 ) ;
  assign n8517 = n8516 ^ x38 ^ 1'b0 ;
  assign n8518 = ( ~x38 & n8284 ) | ( ~x38 & n8517 ) | ( n8284 & n8517 ) ;
  assign n8519 = ( x38 & n8516 ) | ( x38 & n8518 ) | ( n8516 & n8518 ) ;
  assign n8520 = x100 & ~n8279 ;
  assign n8521 = ( x75 & n8519 ) | ( x75 & ~n8520 ) | ( n8519 & ~n8520 ) ;
  assign n8522 = n8521 ^ n8519 ^ 1'b0 ;
  assign n8523 = ( x75 & n8521 ) | ( x75 & ~n8522 ) | ( n8521 & ~n8522 ) ;
  assign n8524 = ( x92 & ~n8510 ) | ( x92 & n8523 ) | ( ~n8510 & n8523 ) ;
  assign n8525 = ~x92 & n8524 ;
  assign n8526 = n7571 & ~n8292 ;
  assign n8527 = ~n8525 & n8526 ;
  assign n8528 = ( n5015 & n8525 ) | ( n5015 & ~n8527 ) | ( n8525 & ~n8527 ) ;
  assign n8529 = n8528 ^ n8509 ^ 1'b0 ;
  assign n8530 = ( n8509 & n8528 ) | ( n8509 & n8529 ) | ( n8528 & n8529 ) ;
  assign n8531 = ( x74 & ~n8509 ) | ( x74 & n8530 ) | ( ~n8509 & n8530 ) ;
  assign n8532 = n8508 & n8531 ;
  assign n8533 = ( n2109 & n8507 ) | ( n2109 & ~n8532 ) | ( n8507 & ~n8532 ) ;
  assign n8534 = ~n2109 & n8533 ;
  assign n8535 = ( ~n8289 & n8299 ) | ( ~n8289 & n8534 ) | ( n8299 & n8534 ) ;
  assign n8536 = ~n8289 & n8535 ;
  assign n8537 = ~x34 & n8536 ;
  assign n8538 = x54 & ~n8503 ;
  assign n8539 = n1205 & n8501 ;
  assign n8540 = ~n8314 & n8539 ;
  assign n8541 = n8540 ^ x87 ^ 1'b0 ;
  assign n8542 = ~n1994 & n8490 ;
  assign n8543 = ~n1276 & n8542 ;
  assign n8544 = x38 & n8327 ;
  assign n8545 = n8543 | n8544 ;
  assign n8546 = n6411 & n8545 ;
  assign n8547 = ( n8313 & ~n8489 ) | ( n8313 & n8546 ) | ( ~n8489 & n8546 ) ;
  assign n8548 = ( n8540 & ~n8541 ) | ( n8540 & n8547 ) | ( ~n8541 & n8547 ) ;
  assign n8549 = ( n7639 & n8315 ) | ( n7639 & ~n8548 ) | ( n8315 & ~n8548 ) ;
  assign n8550 = n8548 ^ n8315 ^ 1'b0 ;
  assign n8551 = ( n8315 & n8549 ) | ( n8315 & ~n8550 ) | ( n8549 & ~n8550 ) ;
  assign n8555 = x161 | n8184 ;
  assign n8552 = ~x161 & n7669 ;
  assign n8556 = ( n7669 & n8189 ) | ( n7669 & n8552 ) | ( n8189 & n8552 ) ;
  assign n8557 = n8555 & n8556 ;
  assign n8558 = ( x38 & x155 ) | ( x38 & ~n8557 ) | ( x155 & ~n8557 ) ;
  assign n8559 = ~x38 & n8558 ;
  assign n8553 = n8182 & n8552 ;
  assign n8554 = n8474 | n8553 ;
  assign n8560 = n8559 ^ n8554 ^ 1'b0 ;
  assign n8561 = ( x299 & ~n8554 ) | ( x299 & n8559 ) | ( ~n8554 & n8559 ) ;
  assign n8562 = ( x299 & ~n8560 ) | ( x299 & n8561 ) | ( ~n8560 & n8561 ) ;
  assign n8563 = ~x144 & n8197 ;
  assign n8564 = n8450 | n8563 ;
  assign n8565 = ~x144 & n8202 ;
  assign n8566 = x144 & n8205 ;
  assign n8567 = ( n8456 & n8565 ) | ( n8456 & ~n8566 ) | ( n8565 & ~n8566 ) ;
  assign n8568 = ~n8565 & n8567 ;
  assign n8569 = x232 & ~n8568 ;
  assign n8570 = n8564 & n8569 ;
  assign n8571 = x38 | n8570 ;
  assign n8572 = ~n8562 & n8571 ;
  assign n8573 = ( x39 & n8339 ) | ( x39 & ~n8572 ) | ( n8339 & ~n8572 ) ;
  assign n8574 = n8572 ^ n8339 ^ 1'b0 ;
  assign n8575 = ( n8339 & n8573 ) | ( n8339 & ~n8574 ) | ( n8573 & ~n8574 ) ;
  assign n8576 = n8106 & n8431 ;
  assign n8577 = x146 | n8134 ;
  assign n8578 = x146 & ~n8148 ;
  assign n8579 = ( x161 & n8577 ) | ( x161 & ~n8578 ) | ( n8577 & ~n8578 ) ;
  assign n8580 = ~x161 & n8579 ;
  assign n8581 = ( ~x162 & n8576 ) | ( ~x162 & n8580 ) | ( n8576 & n8580 ) ;
  assign n8582 = ~x162 & n8581 ;
  assign n8583 = ~x146 & n8129 ;
  assign n8584 = ( ~x161 & n8163 ) | ( ~x161 & n8583 ) | ( n8163 & n8583 ) ;
  assign n8585 = ~x161 & n8584 ;
  assign n8586 = x159 & n1788 ;
  assign n8587 = x299 & ~n8586 ;
  assign n8588 = ~x146 & n8117 ;
  assign n8589 = n8157 | n8588 ;
  assign n8590 = x161 & n8589 ;
  assign n8591 = ( n8585 & n8587 ) | ( n8585 & ~n8590 ) | ( n8587 & ~n8590 ) ;
  assign n8592 = ~n8585 & n8591 ;
  assign n8593 = ~x162 & n8096 ;
  assign n8594 = x159 & n8593 ;
  assign n8595 = ( x299 & n8270 ) | ( x299 & ~n8594 ) | ( n8270 & ~n8594 ) ;
  assign n8596 = ~n8270 & n8595 ;
  assign n8597 = ( ~n8582 & n8592 ) | ( ~n8582 & n8596 ) | ( n8592 & n8596 ) ;
  assign n8598 = ~n8582 & n8597 ;
  assign n8599 = ~x142 & n8117 ;
  assign n8600 = ( x140 & n8140 ) | ( x140 & ~n8599 ) | ( n8140 & ~n8599 ) ;
  assign n8601 = ~n8140 & n8600 ;
  assign n8602 = ~x142 & n8106 ;
  assign n8603 = x140 | n8602 ;
  assign n8604 = x144 & ~n8603 ;
  assign n8605 = ( x144 & n8601 ) | ( x144 & n8604 ) | ( n8601 & n8604 ) ;
  assign n8606 = ~x142 & n8134 ;
  assign n8607 = x142 & n8148 ;
  assign n8608 = ( x140 & ~n8606 ) | ( x140 & n8607 ) | ( ~n8606 & n8607 ) ;
  assign n8609 = n8606 | n8608 ;
  assign n8610 = x140 & ~n8143 ;
  assign n8611 = ~x142 & n8129 ;
  assign n8612 = n8610 & ~n8611 ;
  assign n8613 = ( x144 & n8609 ) | ( x144 & ~n8612 ) | ( n8609 & ~n8612 ) ;
  assign n8614 = n8613 ^ n8609 ^ 1'b0 ;
  assign n8615 = ( x144 & n8613 ) | ( x144 & ~n8614 ) | ( n8613 & ~n8614 ) ;
  assign n8616 = x140 & n5075 ;
  assign n8617 = ( n8605 & n8615 ) | ( n8605 & ~n8616 ) | ( n8615 & ~n8616 ) ;
  assign n8618 = ~n8605 & n8617 ;
  assign n8619 = x181 & n8096 ;
  assign n8620 = ( x299 & ~n8618 ) | ( x299 & n8619 ) | ( ~n8618 & n8619 ) ;
  assign n8621 = n8618 | n8620 ;
  assign n8622 = ( x232 & n8598 ) | ( x232 & n8621 ) | ( n8598 & n8621 ) ;
  assign n8623 = ~n8598 & n8622 ;
  assign n8624 = ( n1994 & ~n8575 ) | ( n1994 & n8623 ) | ( ~n8575 & n8623 ) ;
  assign n8625 = ~n8575 & n8624 ;
  assign n8626 = ( n8313 & ~n8489 ) | ( n8313 & n8625 ) | ( ~n8489 & n8625 ) ;
  assign n8627 = n8626 ^ x87 ^ 1'b0 ;
  assign n8628 = ( n8540 & n8626 ) | ( n8540 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8629 = ( n2053 & ~n8551 ) | ( n2053 & n8628 ) | ( ~n8551 & n8628 ) ;
  assign n8630 = ~n8551 & n8629 ;
  assign n8631 = x54 | n8630 ;
  assign n8632 = ~n8538 & n8631 ;
  assign n8633 = x74 | n8632 ;
  assign n8634 = ~n8325 & n8633 ;
  assign n8635 = x38 & n8284 ;
  assign n8636 = ~x92 & x162 ;
  assign n8637 = n8156 & ~n8223 ;
  assign n8638 = n8636 & n8637 ;
  assign n8639 = n5088 | n8638 ;
  assign n8640 = ( ~n5088 & n8635 ) | ( ~n5088 & n8639 ) | ( n8635 & n8639 ) ;
  assign n8641 = n7555 | n8640 ;
  assign n8642 = ( ~n7555 & n8290 ) | ( ~n7555 & n8641 ) | ( n8290 & n8641 ) ;
  assign n8643 = n8642 ^ n8509 ^ 1'b0 ;
  assign n8644 = ( n8509 & n8642 ) | ( n8509 & n8643 ) | ( n8642 & n8643 ) ;
  assign n8645 = ( x74 & ~n8509 ) | ( x74 & n8644 ) | ( ~n8509 & n8644 ) ;
  assign n8646 = n8508 & n8645 ;
  assign n8647 = ( n2109 & ~n8634 ) | ( n2109 & n8646 ) | ( ~n8634 & n8646 ) ;
  assign n8648 = n8634 | n8647 ;
  assign n8649 = n8648 ^ n8297 ^ 1'b0 ;
  assign n8650 = ( n8297 & n8648 ) | ( n8297 & n8649 ) | ( n8648 & n8649 ) ;
  assign n8651 = ( n8289 & ~n8297 ) | ( n8289 & n8650 ) | ( ~n8297 & n8650 ) ;
  assign n8652 = x34 & ~n8651 ;
  assign n8653 = x33 | x954 ;
  assign n8654 = ( n8537 & ~n8652 ) | ( n8537 & n8653 ) | ( ~n8652 & n8653 ) ;
  assign n8655 = ~n8537 & n8654 ;
  assign n8656 = ~x34 & n8262 ;
  assign n8657 = n8536 & ~n8656 ;
  assign n8658 = ~n8651 & n8656 ;
  assign n8659 = n8653 | n8658 ;
  assign n8660 = ( ~n8655 & n8657 ) | ( ~n8655 & n8659 ) | ( n8657 & n8659 ) ;
  assign n8661 = ~n8655 & n8660 ;
  assign n8662 = n2070 | n2109 ;
  assign n8663 = n7455 | n8662 ;
  assign n8664 = x55 | n8663 ;
  assign n8665 = x59 & n8664 ;
  assign n8666 = ( x24 & x54 ) | ( x24 & n6254 ) | ( x54 & n6254 ) ;
  assign n8667 = ( n2109 & n7447 ) | ( n2109 & ~n8666 ) | ( n7447 & ~n8666 ) ;
  assign n8668 = n8666 | n8667 ;
  assign n8669 = x137 & n7534 ;
  assign n8670 = x1091 & x1093 ;
  assign n8671 = n1614 & n8670 ;
  assign n8672 = n6425 & ~n8671 ;
  assign n8673 = x683 & n8672 ;
  assign n8674 = x252 & n5035 ;
  assign n8675 = ~n8673 & n8674 ;
  assign n8676 = ( n5044 & n7530 ) | ( n5044 & n8675 ) | ( n7530 & n8675 ) ;
  assign n8677 = n8676 ^ n7533 ^ n7457 ;
  assign n8678 = ( n7529 & n8676 ) | ( n7529 & ~n8677 ) | ( n8676 & ~n8677 ) ;
  assign n8679 = ~n8677 & n8678 ;
  assign n8680 = ~n8669 & n8679 ;
  assign n8681 = ( n7528 & n8669 ) | ( n7528 & ~n8680 ) | ( n8669 & ~n8680 ) ;
  assign n8682 = n7466 & n8681 ;
  assign n8683 = x39 | x100 ;
  assign n8684 = x38 & n7455 ;
  assign n8685 = n1615 & n6480 ;
  assign n8686 = x122 | n5023 ;
  assign n8687 = x137 | n5165 ;
  assign n8688 = ~n6612 & n8687 ;
  assign n8689 = ~n8686 & n8688 ;
  assign n8690 = n6612 & n8687 ;
  assign n8691 = n8689 ^ n8685 ^ 1'b0 ;
  assign n8692 = ( ~n8685 & n8690 ) | ( ~n8685 & n8691 ) | ( n8690 & n8691 ) ;
  assign n8693 = ( n8685 & n8689 ) | ( n8685 & n8692 ) | ( n8689 & n8692 ) ;
  assign n8694 = ( ~x90 & x93 ) | ( ~x90 & n8100 ) | ( x93 & n8100 ) ;
  assign n8695 = n8694 ^ n5148 ^ 1'b0 ;
  assign n8696 = ( n5148 & n8694 ) | ( n5148 & n8695 ) | ( n8694 & n8695 ) ;
  assign n8697 = ( x35 & ~n5148 ) | ( x35 & n8696 ) | ( ~n5148 & n8696 ) ;
  assign n8698 = n8693 ^ n5165 ^ 1'b0 ;
  assign n8699 = ( ~n5165 & n8697 ) | ( ~n5165 & n8698 ) | ( n8697 & n8698 ) ;
  assign n8700 = ( n5165 & n8693 ) | ( n5165 & n8699 ) | ( n8693 & n8699 ) ;
  assign n8701 = n8700 ^ x38 ^ 1'b0 ;
  assign n8702 = x35 & ~n1595 ;
  assign n8703 = n7482 | n8702 ;
  assign n8704 = ~n1374 & n7508 ;
  assign n8705 = n8697 | n8704 ;
  assign n8706 = ( n1289 & ~n8703 ) | ( n1289 & n8705 ) | ( ~n8703 & n8705 ) ;
  assign n8707 = ~n1289 & n8706 ;
  assign n8708 = ( n8700 & ~n8701 ) | ( n8700 & n8707 ) | ( ~n8701 & n8707 ) ;
  assign n8709 = ( x38 & n8701 ) | ( x38 & n8708 ) | ( n8701 & n8708 ) ;
  assign n8710 = x32 & ~x93 ;
  assign n8711 = ( n6374 & ~n7468 ) | ( n6374 & n8710 ) | ( ~n7468 & n8710 ) ;
  assign n8712 = ~n6374 & n8711 ;
  assign n8713 = n8697 & ~n8703 ;
  assign n8714 = ( ~x32 & n8712 ) | ( ~x32 & n8713 ) | ( n8712 & n8713 ) ;
  assign n8715 = n8712 ^ x32 ^ 1'b0 ;
  assign n8716 = ( n8712 & n8714 ) | ( n8712 & ~n8715 ) | ( n8714 & ~n8715 ) ;
  assign n8717 = ( x95 & ~n5165 ) | ( x95 & n8716 ) | ( ~n5165 & n8716 ) ;
  assign n8718 = ~x95 & n8717 ;
  assign n8719 = x1082 & ~n1289 ;
  assign n8720 = n1586 | n8713 ;
  assign n8721 = n8719 & n8720 ;
  assign n8722 = ( ~n8709 & n8718 ) | ( ~n8709 & n8721 ) | ( n8718 & n8721 ) ;
  assign n8723 = n8709 | n8722 ;
  assign n8724 = ( n8683 & ~n8684 ) | ( n8683 & n8723 ) | ( ~n8684 & n8723 ) ;
  assign n8725 = ~n8683 & n8724 ;
  assign n8726 = ( ~n2044 & n8682 ) | ( ~n2044 & n8725 ) | ( n8682 & n8725 ) ;
  assign n8727 = ~n2044 & n8726 ;
  assign n8728 = x137 & ~n7451 ;
  assign n8729 = ~n5045 & n8728 ;
  assign n8730 = ( n7458 & n7461 ) | ( n7458 & n8729 ) | ( n7461 & n8729 ) ;
  assign n8731 = n7461 & n8730 ;
  assign n8732 = n7455 | n8731 ;
  assign n8733 = ( ~n7455 & n8727 ) | ( ~n7455 & n8732 ) | ( n8727 & n8732 ) ;
  assign n8734 = n8733 ^ x92 ^ 1'b0 ;
  assign n8735 = ( x92 & n8733 ) | ( x92 & n8734 ) | ( n8733 & n8734 ) ;
  assign n8736 = ( x54 & ~x92 ) | ( x54 & n8735 ) | ( ~x92 & n8735 ) ;
  assign n8737 = n8736 ^ n8668 ^ 1'b0 ;
  assign n8738 = ( n8668 & n8736 ) | ( n8668 & n8737 ) | ( n8736 & n8737 ) ;
  assign n8739 = ( x59 & ~n8668 ) | ( x59 & n8738 ) | ( ~n8668 & n8738 ) ;
  assign n8740 = ( x57 & ~n8665 ) | ( x57 & n8739 ) | ( ~n8665 & n8739 ) ;
  assign n8741 = ~x57 & n8740 ;
  assign n8742 = n1395 | n1458 ;
  assign n8743 = x83 | n1527 ;
  assign n8744 = x65 | n1226 ;
  assign n8745 = ( n1230 & n7586 ) | ( n1230 & ~n8744 ) | ( n7586 & ~n8744 ) ;
  assign n8746 = n8744 | n8745 ;
  assign n8747 = x69 | n8746 ;
  assign n8748 = x67 | x71 ;
  assign n8749 = x36 & ~x103 ;
  assign n8750 = ~n8748 & n8749 ;
  assign n8751 = ( n8743 & ~n8747 ) | ( n8743 & n8750 ) | ( ~n8747 & n8750 ) ;
  assign n8752 = ~n8743 & n8751 ;
  assign n8753 = ~n8742 & n8752 ;
  assign n8754 = ~x58 & n6428 ;
  assign n8755 = n8753 | n8754 ;
  assign n8756 = n1374 | n5203 ;
  assign n8757 = n5160 | n8756 ;
  assign n8758 = n2067 | n7318 ;
  assign n8759 = n2177 | n8758 ;
  assign n8760 = x92 | n8759 ;
  assign n8761 = n8757 | n8760 ;
  assign n8762 = n5023 & ~n8761 ;
  assign n8763 = n8755 & n8762 ;
  assign n8764 = x39 | n1290 ;
  assign n8765 = x24 & ~n8764 ;
  assign n8766 = ~n1379 & n8765 ;
  assign n8767 = x38 & ~n8766 ;
  assign n8768 = x81 | n1477 ;
  assign n8769 = n5203 | n7878 ;
  assign n8770 = n1265 | n8769 ;
  assign n8771 = x71 | n1230 ;
  assign n8772 = x104 | n1237 ;
  assign n8773 = x45 | x73 ;
  assign n8774 = n7493 | n8773 ;
  assign n8775 = x48 | x65 ;
  assign n8776 = x82 | x84 ;
  assign n8777 = ( x89 & n8775 ) | ( x89 & ~n8776 ) | ( n8775 & ~n8776 ) ;
  assign n8778 = ~n8775 & n8777 ;
  assign n8779 = ( n7757 & ~n8774 ) | ( n7757 & n8778 ) | ( ~n8774 & n8778 ) ;
  assign n8780 = ~n7757 & n8779 ;
  assign n8781 = ( n8771 & ~n8772 ) | ( n8771 & n8780 ) | ( ~n8772 & n8780 ) ;
  assign n8782 = ~n8771 & n8781 ;
  assign n8783 = x332 & n8782 ;
  assign n8784 = x64 | n8783 ;
  assign n8785 = x39 | x841 ;
  assign n8786 = ( n1229 & n8784 ) | ( n1229 & ~n8785 ) | ( n8784 & ~n8785 ) ;
  assign n8787 = ~n1229 & n8786 ;
  assign n8788 = ( n1272 & ~n8770 ) | ( n1272 & n8787 ) | ( ~n8770 & n8787 ) ;
  assign n8789 = ~n1272 & n8788 ;
  assign n8790 = n8789 ^ n8768 ^ 1'b0 ;
  assign n8791 = ( n8768 & n8789 ) | ( n8768 & n8790 ) | ( n8789 & n8790 ) ;
  assign n8792 = ( x38 & ~n8768 ) | ( x38 & n8791 ) | ( ~n8768 & n8791 ) ;
  assign n8793 = n2069 | n7318 ;
  assign n8794 = ( n8767 & n8792 ) | ( n8767 & ~n8793 ) | ( n8792 & ~n8793 ) ;
  assign n8795 = ~n8767 & n8794 ;
  assign n8796 = n7485 | n7489 ;
  assign n8797 = n7496 | n7758 ;
  assign n8798 = x65 | x69 ;
  assign n8799 = x48 & ~x49 ;
  assign n8800 = x68 | x82 ;
  assign n8801 = ( n8773 & n8799 ) | ( n8773 & ~n8800 ) | ( n8799 & ~n8800 ) ;
  assign n8802 = ~n8773 & n8801 ;
  assign n8803 = ( n8797 & ~n8798 ) | ( n8797 & n8802 ) | ( ~n8798 & n8802 ) ;
  assign n8804 = ~n8797 & n8803 ;
  assign n8805 = ( n7754 & ~n8796 ) | ( n7754 & n8804 ) | ( ~n8796 & n8804 ) ;
  assign n8806 = ~n7754 & n8805 ;
  assign n8807 = ( n8771 & ~n8772 ) | ( n8771 & n8806 ) | ( ~n8772 & n8806 ) ;
  assign n8808 = ~n8771 & n8807 ;
  assign n8809 = x47 | x841 ;
  assign n8810 = n8808 & ~n8809 ;
  assign n8811 = n1447 | n8810 ;
  assign n8812 = n1370 | n1449 ;
  assign n8813 = n1392 | n1461 ;
  assign n8814 = x841 | n1260 ;
  assign n8815 = n1387 | n8814 ;
  assign n8816 = x97 | n8815 ;
  assign n8817 = n8808 & ~n8816 ;
  assign n8818 = ~n8813 & n8817 ;
  assign n8819 = x108 & ~n1392 ;
  assign n8820 = ~n1460 & n8819 ;
  assign n8821 = ( x47 & ~n8818 ) | ( x47 & n8820 ) | ( ~n8818 & n8820 ) ;
  assign n8822 = n8818 | n8821 ;
  assign n8823 = x986 | n5023 ;
  assign n8824 = x252 & n8823 ;
  assign n8825 = x314 & ~n8824 ;
  assign n8826 = ( n8812 & n8822 ) | ( n8812 & n8825 ) | ( n8822 & n8825 ) ;
  assign n8827 = ~n8812 & n8826 ;
  assign n8828 = n1264 | n1370 ;
  assign n8829 = n8825 | n8828 ;
  assign n8830 = ~n8827 & n8829 ;
  assign n8831 = ( n8811 & n8827 ) | ( n8811 & ~n8830 ) | ( n8827 & ~n8830 ) ;
  assign n8832 = n8831 ^ n1374 ^ 1'b0 ;
  assign n8833 = ( n1374 & n8831 ) | ( n1374 & n8832 ) | ( n8831 & n8832 ) ;
  assign n8834 = ( x35 & ~n1374 ) | ( x35 & n8833 ) | ( ~n1374 & n8833 ) ;
  assign n8835 = ( n1272 & n5160 ) | ( n1272 & n5281 ) | ( n5160 & n5281 ) ;
  assign n8836 = ( n1274 & n8834 ) | ( n1274 & ~n8835 ) | ( n8834 & ~n8835 ) ;
  assign n8837 = ~n1274 & n8836 ;
  assign n8838 = n8837 ^ n5284 ^ 1'b0 ;
  assign n8839 = ( n5165 & ~n5284 ) | ( n5165 & n8838 ) | ( ~n5284 & n8838 ) ;
  assign n8840 = ( n5284 & n8837 ) | ( n5284 & n8839 ) | ( n8837 & n8839 ) ;
  assign n8841 = ( x39 & ~x95 ) | ( x39 & n8840 ) | ( ~x95 & n8840 ) ;
  assign n8842 = ~x39 & n8841 ;
  assign n8843 = x786 & ~x1082 ;
  assign n8844 = n5023 & n8843 ;
  assign n8845 = n4736 & n5100 ;
  assign n8846 = ~n2290 & n5115 ;
  assign n8847 = n8845 | n8846 ;
  assign n8848 = ( ~n5364 & n8844 ) | ( ~n5364 & n8847 ) | ( n8844 & n8847 ) ;
  assign n8849 = n5364 & n8848 ;
  assign n8850 = n5069 & ~n5362 ;
  assign n8851 = ( x835 & n5020 ) | ( x835 & n5066 ) | ( n5020 & n5066 ) ;
  assign n8852 = n5068 & ~n8851 ;
  assign n8853 = n5065 & ~n8852 ;
  assign n8854 = n5099 & n8853 ;
  assign n8855 = n8850 & ~n8854 ;
  assign n8856 = ~n5061 & n8855 ;
  assign n8857 = ~n5083 & n8853 ;
  assign n8858 = n8850 & ~n8857 ;
  assign n8859 = n5061 & n8858 ;
  assign n8860 = ( x299 & n8856 ) | ( x299 & ~n8859 ) | ( n8856 & ~n8859 ) ;
  assign n8861 = ~n8856 & n8860 ;
  assign n8862 = x1093 & n8853 ;
  assign n8863 = n8850 & ~n8862 ;
  assign n8864 = ~x215 & n8863 ;
  assign n8865 = n8861 & ~n8864 ;
  assign n8866 = ~x223 & n8863 ;
  assign n8867 = n5114 & n8858 ;
  assign n8868 = ~n5114 & n8855 ;
  assign n8869 = ( x299 & ~n8867 ) | ( x299 & n8868 ) | ( ~n8867 & n8868 ) ;
  assign n8870 = n8867 | n8869 ;
  assign n8871 = n8866 | n8870 ;
  assign n8872 = ~n8843 & n8871 ;
  assign n8873 = ( n8849 & ~n8865 ) | ( n8849 & n8872 ) | ( ~n8865 & n8872 ) ;
  assign n8874 = n8865 ^ n8849 ^ 1'b0 ;
  assign n8875 = ( n8849 & n8873 ) | ( n8849 & ~n8874 ) | ( n8873 & ~n8874 ) ;
  assign n8876 = n8842 ^ x39 ^ 1'b0 ;
  assign n8877 = ( ~x39 & n8875 ) | ( ~x39 & n8876 ) | ( n8875 & n8876 ) ;
  assign n8878 = ( x39 & n8842 ) | ( x39 & n8877 ) | ( n8842 & n8877 ) ;
  assign n8879 = ( x38 & ~n8793 ) | ( x38 & n8878 ) | ( ~n8793 & n8878 ) ;
  assign n8880 = ~x38 & n8879 ;
  assign n8881 = ~x93 & x102 ;
  assign n8882 = ~n1225 & n8881 ;
  assign n8883 = ( n1228 & ~n5160 ) | ( n1228 & n8882 ) | ( ~n5160 & n8882 ) ;
  assign n8884 = ~n1228 & n8883 ;
  assign n8885 = ( n1254 & ~n1265 ) | ( n1254 & n8884 ) | ( ~n1265 & n8884 ) ;
  assign n8886 = ~n1254 & n8885 ;
  assign n8887 = ~n5203 & n8886 ;
  assign n8888 = x1082 & ~n8887 ;
  assign n8889 = n8760 | n8888 ;
  assign n8890 = n1289 | n2218 ;
  assign n8891 = x40 | n8886 ;
  assign n8892 = ~n8890 & n8891 ;
  assign n8893 = ( x1082 & ~n8889 ) | ( x1082 & n8892 ) | ( ~n8889 & n8892 ) ;
  assign n8894 = ~n8889 & n8893 ;
  assign n8895 = x41 | x72 ;
  assign n8896 = ~x39 & n8895 ;
  assign n8897 = x72 | n8896 ;
  assign n8898 = x166 | n5075 ;
  assign n8899 = x161 & ~n8898 ;
  assign n8900 = ~x152 & n8899 ;
  assign n8901 = x39 & x232 ;
  assign n8902 = n8900 & n8901 ;
  assign n8903 = ( n7318 & n8897 ) | ( n7318 & ~n8902 ) | ( n8897 & ~n8902 ) ;
  assign n8904 = ~n8897 & n8903 ;
  assign n8905 = x189 | n5075 ;
  assign n8906 = x144 & ~n8905 ;
  assign n8907 = ~x174 & n8906 ;
  assign n8908 = x299 | n8907 ;
  assign n8909 = n5038 | n8900 ;
  assign n8910 = ( ~x232 & n8908 ) | ( ~x232 & n8909 ) | ( n8908 & n8909 ) ;
  assign n8911 = x232 & n8910 ;
  assign n8912 = x72 | n8911 ;
  assign n8913 = x39 & ~n8912 ;
  assign n8914 = n8913 ^ n8896 ^ x39 ;
  assign n8915 = n2052 & ~n8914 ;
  assign n8916 = x75 & ~n8915 ;
  assign n8917 = x39 & n8912 ;
  assign n8918 = ~n6824 & n8895 ;
  assign n8919 = x44 | n1292 ;
  assign n8920 = x101 | n8919 ;
  assign n8921 = n6480 & ~n8920 ;
  assign n8922 = n6414 & n8921 ;
  assign n8923 = x41 & ~n8922 ;
  assign n8924 = ~x41 & x72 ;
  assign n8925 = n1615 & ~n8924 ;
  assign n8926 = x99 | n5033 ;
  assign n8927 = ~x72 & x101 ;
  assign n8928 = x41 | n8927 ;
  assign n8929 = x24 | n1379 ;
  assign n8930 = x252 & ~n5203 ;
  assign n8931 = n6480 & n8930 ;
  assign n8932 = ~n8929 & n8931 ;
  assign n8933 = ~x44 & n8932 ;
  assign n8934 = ~n8928 & n8933 ;
  assign n8935 = n8926 & n8934 ;
  assign n8936 = ( n8923 & n8925 ) | ( n8923 & ~n8935 ) | ( n8925 & ~n8935 ) ;
  assign n8937 = ~n8923 & n8936 ;
  assign n8938 = n1615 | n8895 ;
  assign n8939 = ( n6824 & n8937 ) | ( n6824 & n8938 ) | ( n8937 & n8938 ) ;
  assign n8940 = ~n8937 & n8939 ;
  assign n8941 = ( ~x39 & n8918 ) | ( ~x39 & n8940 ) | ( n8918 & n8940 ) ;
  assign n8942 = ~x39 & n8941 ;
  assign n8943 = ( n2052 & ~n8917 ) | ( n2052 & n8942 ) | ( ~n8917 & n8942 ) ;
  assign n8944 = n8917 | n8943 ;
  assign n8945 = n8916 & n8944 ;
  assign n8946 = x228 | n8895 ;
  assign n8947 = x41 & n8920 ;
  assign n8948 = n1379 | n5203 ;
  assign n8949 = x44 | n8948 ;
  assign n8950 = n8928 | n8949 ;
  assign n8951 = ~n8924 & n8950 ;
  assign n8952 = x228 & n8951 ;
  assign n8953 = ~n8947 & n8952 ;
  assign n8954 = ( n2036 & n8946 ) | ( n2036 & ~n8953 ) | ( n8946 & ~n8953 ) ;
  assign n8955 = ~n2036 & n8954 ;
  assign n8956 = n1205 & n8896 ;
  assign n8957 = ( x87 & n8917 ) | ( x87 & ~n8956 ) | ( n8917 & ~n8956 ) ;
  assign n8958 = ~n8917 & n8957 ;
  assign n8959 = n8958 ^ n8955 ^ 1'b0 ;
  assign n8960 = ( n8955 & n8958 ) | ( n8955 & n8959 ) | ( n8958 & n8959 ) ;
  assign n8961 = ( x75 & ~n8955 ) | ( x75 & n8960 ) | ( ~n8955 & n8960 ) ;
  assign n8962 = x287 & ~n1292 ;
  assign n8963 = n8911 & n8962 ;
  assign n8964 = ( x39 & n8913 ) | ( x39 & n8963 ) | ( n8913 & n8963 ) ;
  assign n8965 = n1371 | n1445 ;
  assign n8966 = x110 & ~n8965 ;
  assign n8967 = ~n8757 & n8966 ;
  assign n8968 = ~x480 & x949 ;
  assign n8969 = ~x250 & x252 ;
  assign n8970 = n8968 & ~n8969 ;
  assign n8971 = n8967 & n8970 ;
  assign n8972 = n1370 | n1446 ;
  assign n8973 = ~n1378 & n8968 ;
  assign n8974 = ~x47 & n8973 ;
  assign n8975 = x109 | n5207 ;
  assign n8976 = n1466 & ~n8975 ;
  assign n8977 = x110 | n8976 ;
  assign n8978 = ( n8972 & n8974 ) | ( n8972 & n8977 ) | ( n8974 & n8977 ) ;
  assign n8979 = ~n8972 & n8978 ;
  assign n8980 = x901 & ~x959 ;
  assign n8981 = ~n1395 & n1466 ;
  assign n8982 = ~n1378 & n8981 ;
  assign n8983 = ~n8968 & n8982 ;
  assign n8984 = ( n8979 & n8980 ) | ( n8979 & ~n8983 ) | ( n8980 & ~n8983 ) ;
  assign n8985 = ~n8979 & n8984 ;
  assign n8986 = ~n5203 & n8969 ;
  assign n8987 = n8966 & n8973 ;
  assign n8988 = n8980 | n8987 ;
  assign n8989 = ( n8985 & n8986 ) | ( n8985 & n8988 ) | ( n8986 & n8988 ) ;
  assign n8990 = ~n8985 & n8989 ;
  assign n8991 = ~x72 & n8990 ;
  assign n8992 = n8971 | n8991 ;
  assign n8993 = ~x44 & n8992 ;
  assign n8994 = ~x101 & n8993 ;
  assign n8995 = x41 & ~n8994 ;
  assign n8996 = x44 & ~x72 ;
  assign n8997 = n5203 | n8969 ;
  assign n8998 = n8987 & ~n8997 ;
  assign n8999 = ( x72 & n8990 ) | ( x72 & ~n8998 ) | ( n8990 & ~n8998 ) ;
  assign n9000 = n8998 | n8999 ;
  assign n9001 = x44 & x72 ;
  assign n9002 = ( ~n8996 & n9000 ) | ( ~n8996 & n9001 ) | ( n9000 & n9001 ) ;
  assign n9003 = x101 & ~n9002 ;
  assign n9004 = ( ~n8928 & n9002 ) | ( ~n8928 & n9003 ) | ( n9002 & n9003 ) ;
  assign n9005 = ( ~x228 & n8995 ) | ( ~x228 & n9004 ) | ( n8995 & n9004 ) ;
  assign n9006 = ~x228 & n9005 ;
  assign n9007 = ~n6396 & n6400 ;
  assign n9008 = x1093 | n6398 ;
  assign n9009 = ( ~x44 & n9007 ) | ( ~x44 & n9008 ) | ( n9007 & n9008 ) ;
  assign n9010 = ~x44 & n9009 ;
  assign n9011 = x96 & ~x1093 ;
  assign n9012 = ( n6400 & n9010 ) | ( n6400 & n9011 ) | ( n9010 & n9011 ) ;
  assign n9013 = ~x101 & n9012 ;
  assign n9014 = x41 & ~n9013 ;
  assign n9015 = n1615 | n9014 ;
  assign n9016 = x72 | n6400 ;
  assign n9017 = ~x72 & n6396 ;
  assign n9018 = n5203 | n6393 ;
  assign n9019 = n6392 & ~n9018 ;
  assign n9020 = n9017 & ~n9019 ;
  assign n9021 = n6396 | n9016 ;
  assign n9022 = ( x1093 & ~n9020 ) | ( x1093 & n9021 ) | ( ~n9020 & n9021 ) ;
  assign n9023 = ~x1093 & n9022 ;
  assign n9024 = n9016 | n9023 ;
  assign n9025 = ( ~n8996 & n9001 ) | ( ~n8996 & n9024 ) | ( n9001 & n9024 ) ;
  assign n9026 = x101 & ~n9025 ;
  assign n9027 = ( ~n8928 & n9025 ) | ( ~n8928 & n9026 ) | ( n9025 & n9026 ) ;
  assign n9028 = ( x228 & n9015 ) | ( x228 & n9027 ) | ( n9015 & n9027 ) ;
  assign n9029 = n9027 ^ n9015 ^ 1'b0 ;
  assign n9030 = ( x228 & n9028 ) | ( x228 & n9029 ) | ( n9028 & n9029 ) ;
  assign n9031 = ~n1625 & n6385 ;
  assign n9032 = n1623 | n9031 ;
  assign n9033 = ( ~n1623 & n6428 ) | ( ~n1623 & n9032 ) | ( n6428 & n9032 ) ;
  assign n9034 = n1225 | n9033 ;
  assign n9035 = ( ~n1225 & n6376 ) | ( ~n1225 & n9034 ) | ( n6376 & n9034 ) ;
  assign n9036 = n9035 ^ n6373 ^ 1'b0 ;
  assign n9037 = ( n6373 & n9035 ) | ( n6373 & n9036 ) | ( n9035 & n9036 ) ;
  assign n9038 = ( x51 & ~n6373 ) | ( x51 & n9037 ) | ( ~n6373 & n9037 ) ;
  assign n9039 = n9038 ^ n1434 ^ 1'b0 ;
  assign n9040 = ( n1434 & n9038 ) | ( n1434 & n9039 ) | ( n9038 & n9039 ) ;
  assign n9041 = ( x96 & ~n1434 ) | ( x96 & n9040 ) | ( ~n1434 & n9040 ) ;
  assign n9042 = n9017 & ~n9018 ;
  assign n9043 = n9041 & n9042 ;
  assign n9044 = n9007 | n9043 ;
  assign n9045 = x1093 & ~n9044 ;
  assign n9046 = n9010 & ~n9045 ;
  assign n9047 = ~x101 & n9046 ;
  assign n9048 = x41 & ~n9047 ;
  assign n9049 = n9048 ^ n9030 ^ 1'b0 ;
  assign n9050 = x72 | n9044 ;
  assign n9051 = x1093 & n9050 ;
  assign n9052 = n9023 | n9051 ;
  assign n9053 = x44 & ~n9052 ;
  assign n9054 = n9053 ^ n9052 ^ n8996 ;
  assign n9055 = x101 & ~n9054 ;
  assign n9056 = ( ~n8928 & n9054 ) | ( ~n8928 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9057 = n1615 & ~n9056 ;
  assign n9058 = ( n9048 & n9049 ) | ( n9048 & ~n9057 ) | ( n9049 & ~n9057 ) ;
  assign n9059 = ( n9030 & ~n9049 ) | ( n9030 & n9058 ) | ( ~n9049 & n9058 ) ;
  assign n9060 = ( x39 & ~n9006 ) | ( x39 & n9059 ) | ( ~n9006 & n9059 ) ;
  assign n9061 = n9006 | n9060 ;
  assign n9062 = ( n1205 & ~n8964 ) | ( n1205 & n9061 ) | ( ~n8964 & n9061 ) ;
  assign n9063 = ~n1205 & n9062 ;
  assign n9064 = n6824 & n8938 ;
  assign n9065 = x72 | n6480 ;
  assign n9066 = ~n8951 & n9065 ;
  assign n9067 = n8926 & n9066 ;
  assign n9068 = n1615 & n8926 ;
  assign n9069 = n8925 | n9068 ;
  assign n9070 = x41 & ~n8921 ;
  assign n9071 = ( n9067 & n9069 ) | ( n9067 & ~n9070 ) | ( n9069 & ~n9070 ) ;
  assign n9072 = ~n9067 & n9071 ;
  assign n9073 = ( n8918 & n9064 ) | ( n8918 & ~n9072 ) | ( n9064 & ~n9072 ) ;
  assign n9074 = n9073 ^ n9064 ^ 1'b0 ;
  assign n9075 = ( n8918 & n9073 ) | ( n8918 & ~n9074 ) | ( n9073 & ~n9074 ) ;
  assign n9076 = x39 | n9075 ;
  assign n9077 = ( ~x39 & n8917 ) | ( ~x39 & n9076 ) | ( n8917 & n9076 ) ;
  assign n9078 = ( x38 & x100 ) | ( x38 & n9077 ) | ( x100 & n9077 ) ;
  assign n9079 = ~x38 & n9078 ;
  assign n9080 = x38 & n8914 ;
  assign n9081 = ( x87 & ~n9079 ) | ( x87 & n9080 ) | ( ~n9079 & n9080 ) ;
  assign n9082 = n9079 | n9081 ;
  assign n9083 = ( ~n8961 & n9063 ) | ( ~n8961 & n9082 ) | ( n9063 & n9082 ) ;
  assign n9084 = ~n8961 & n9083 ;
  assign n9085 = ( ~n6782 & n8945 ) | ( ~n6782 & n9084 ) | ( n8945 & n9084 ) ;
  assign n9086 = ~n6782 & n9085 ;
  assign n9087 = n6782 & n8914 ;
  assign n9088 = n7318 | n9087 ;
  assign n9089 = ( ~n8904 & n9086 ) | ( ~n8904 & n9088 ) | ( n9086 & n9088 ) ;
  assign n9090 = ~n8904 & n9089 ;
  assign n9091 = x42 & ~x72 ;
  assign n9092 = n6824 | n9091 ;
  assign n9093 = ~x115 & n1615 ;
  assign n9094 = x114 & ~n9091 ;
  assign n9095 = n9093 & ~n9094 ;
  assign n9109 = n6824 & n9093 ;
  assign n9110 = ( ~n9091 & n9092 ) | ( ~n9091 & n9109 ) | ( n9092 & n9109 ) ;
  assign n9096 = n5026 | n8920 ;
  assign n9097 = n5030 | n9096 ;
  assign n9098 = n6480 & ~n9097 ;
  assign n9099 = ~x114 & n5029 ;
  assign n9100 = n9098 & n9099 ;
  assign n9101 = ~x42 & n9100 ;
  assign n9102 = n5027 | n8949 ;
  assign n9103 = n5030 | n9102 ;
  assign n9104 = ~x72 & n9103 ;
  assign n9105 = n9065 & ~n9104 ;
  assign n9106 = x42 & ~n9105 ;
  assign n9107 = ( x114 & ~n9101 ) | ( x114 & n9106 ) | ( ~n9101 & n9106 ) ;
  assign n9108 = n9101 | n9107 ;
  assign n9111 = ~n9108 & n9110 ;
  assign n9112 = ( ~n9095 & n9110 ) | ( ~n9095 & n9111 ) | ( n9110 & n9111 ) ;
  assign n9113 = ( x39 & n9092 ) | ( x39 & ~n9112 ) | ( n9092 & ~n9112 ) ;
  assign n9114 = n9113 ^ n9092 ^ 1'b0 ;
  assign n9115 = ( x39 & n9113 ) | ( x39 & ~n9114 ) | ( n9113 & ~n9114 ) ;
  assign n9116 = ~x72 & x199 ;
  assign n9117 = x232 | n9116 ;
  assign n9118 = ~x299 & n9117 ;
  assign n9119 = ~x72 & n8905 ;
  assign n9120 = x199 & n9119 ;
  assign n9121 = x232 & ~n9120 ;
  assign n9122 = n9118 & ~n9121 ;
  assign n9123 = x39 & ~n9122 ;
  assign n9124 = n9115 & ~n9123 ;
  assign n9125 = n5018 & ~n9124 ;
  assign n9126 = x115 & ~n9091 ;
  assign n9127 = x42 & ~x114 ;
  assign n9135 = ~x72 & x116 ;
  assign n9132 = ~x72 & x113 ;
  assign n9128 = x72 & n5026 ;
  assign n9129 = ~x99 & n9004 ;
  assign n9130 = n9128 | n9129 ;
  assign n9131 = x113 & ~n9130 ;
  assign n9133 = n9132 ^ n9131 ^ n9130 ;
  assign n9134 = x116 & ~n9133 ;
  assign n9136 = n9135 ^ n9134 ^ n9133 ;
  assign n9137 = n9127 & n9136 ;
  assign n9138 = ~n5026 & n8994 ;
  assign n9139 = ~x113 & n9138 ;
  assign n9140 = ~x116 & n9139 ;
  assign n9141 = x42 | n9140 ;
  assign n9142 = ~n9094 & n9141 ;
  assign n9143 = n9142 ^ n9137 ^ 1'b0 ;
  assign n9144 = ( n9137 & n9142 ) | ( n9137 & n9143 ) | ( n9142 & n9143 ) ;
  assign n9145 = ( x115 & ~n9137 ) | ( x115 & n9144 ) | ( ~n9137 & n9144 ) ;
  assign n9146 = ( x228 & ~n9126 ) | ( x228 & n9145 ) | ( ~n9126 & n9145 ) ;
  assign n9147 = ~x228 & n9146 ;
  assign n9148 = ~n5026 & n9047 ;
  assign n9149 = ~n5030 & n9148 ;
  assign n9150 = x42 | n9149 ;
  assign n9151 = ~x99 & n9056 ;
  assign n9152 = n9128 | n9151 ;
  assign n9153 = n9152 ^ x113 ^ 1'b0 ;
  assign n9154 = ( x72 & n9152 ) | ( x72 & n9153 ) | ( n9152 & n9153 ) ;
  assign n9155 = x116 | n9154 ;
  assign n9156 = ~n9135 & n9155 ;
  assign n9157 = n9127 & n9156 ;
  assign n9158 = ( n9094 & n9150 ) | ( n9094 & ~n9157 ) | ( n9150 & ~n9157 ) ;
  assign n9159 = ~n9094 & n9158 ;
  assign n9160 = ( x115 & n1615 ) | ( x115 & ~n9159 ) | ( n1615 & ~n9159 ) ;
  assign n9161 = ~x115 & n9160 ;
  assign n9162 = ~n5026 & n9013 ;
  assign n9163 = ~n5030 & n9162 ;
  assign n9164 = ~x42 & n9163 ;
  assign n9165 = x114 | n9164 ;
  assign n9166 = ~x99 & n9027 ;
  assign n9167 = n9128 | n9166 ;
  assign n9168 = n9167 ^ x113 ^ 1'b0 ;
  assign n9169 = ( x72 & n9167 ) | ( x72 & n9168 ) | ( n9167 & n9168 ) ;
  assign n9170 = x116 & ~n9169 ;
  assign n9171 = n9170 ^ n9169 ^ n9135 ;
  assign n9172 = x42 & ~n9171 ;
  assign n9173 = ( ~n9094 & n9165 ) | ( ~n9094 & n9172 ) | ( n9165 & n9172 ) ;
  assign n9174 = ~n9094 & n9173 ;
  assign n9175 = ( x115 & n1615 ) | ( x115 & ~n9174 ) | ( n1615 & ~n9174 ) ;
  assign n9176 = n9174 | n9175 ;
  assign n9177 = x228 & ~n9126 ;
  assign n9178 = ( n9161 & n9176 ) | ( n9161 & n9177 ) | ( n9176 & n9177 ) ;
  assign n9179 = ~n9161 & n9178 ;
  assign n9180 = ( x39 & ~n9147 ) | ( x39 & n9179 ) | ( ~n9147 & n9179 ) ;
  assign n9181 = n9147 | n9180 ;
  assign n9182 = ~n5075 & n8962 ;
  assign n9183 = ~x189 & n9182 ;
  assign n9184 = n9119 | n9183 ;
  assign n9185 = x199 & n9184 ;
  assign n9186 = x232 & ~n9185 ;
  assign n9187 = n9118 & ~n9186 ;
  assign n9188 = x39 & ~n9187 ;
  assign n9189 = ( n1205 & n9181 ) | ( n1205 & ~n9188 ) | ( n9181 & ~n9188 ) ;
  assign n9190 = n9189 ^ n9181 ^ 1'b0 ;
  assign n9191 = ( n1205 & n9189 ) | ( n1205 & ~n9190 ) | ( n9189 & ~n9190 ) ;
  assign n9192 = n9091 ^ x39 ^ 1'b0 ;
  assign n9193 = ( n9091 & n9122 ) | ( n9091 & n9192 ) | ( n9122 & n9192 ) ;
  assign n9194 = x38 & ~n9193 ;
  assign n9195 = x87 | n9194 ;
  assign n9196 = ( n9125 & n9191 ) | ( n9125 & ~n9195 ) | ( n9191 & ~n9195 ) ;
  assign n9197 = ~n9125 & n9196 ;
  assign n9198 = x228 & ~n9097 ;
  assign n9199 = ~x115 & n9198 ;
  assign n9200 = ~x114 & n9199 ;
  assign n9201 = ~x42 & n9200 ;
  assign n9202 = x228 & ~n9102 ;
  assign n9203 = ~n5032 & n9202 ;
  assign n9204 = n9091 & ~n9203 ;
  assign n9205 = ( n2036 & ~n9201 ) | ( n2036 & n9204 ) | ( ~n9201 & n9204 ) ;
  assign n9206 = n9201 | n9205 ;
  assign n9207 = x39 | n9091 ;
  assign n9208 = n1205 & ~n9207 ;
  assign n9209 = x87 & ~n9208 ;
  assign n9210 = n9206 & n9209 ;
  assign n9211 = ~n9123 & n9210 ;
  assign n9212 = ( x75 & ~n9197 ) | ( x75 & n9211 ) | ( ~n9197 & n9211 ) ;
  assign n9213 = n9197 | n9212 ;
  assign n9214 = ~n5027 & n8933 ;
  assign n9215 = ~x113 & n9214 ;
  assign n9216 = ~x116 & n9215 ;
  assign n9217 = n9091 & ~n9216 ;
  assign n9218 = n6414 & n9100 ;
  assign n9219 = ~x42 & n9218 ;
  assign n9220 = ( x114 & ~n9217 ) | ( x114 & n9219 ) | ( ~n9217 & n9219 ) ;
  assign n9221 = n9217 | n9220 ;
  assign n9222 = n9110 & ~n9221 ;
  assign n9223 = ( ~n9095 & n9110 ) | ( ~n9095 & n9222 ) | ( n9110 & n9222 ) ;
  assign n9224 = ( n2052 & n9092 ) | ( n2052 & ~n9223 ) | ( n9092 & ~n9223 ) ;
  assign n9225 = ~n2052 & n9224 ;
  assign n9226 = n2052 & n9091 ;
  assign n9227 = ( x39 & ~n9225 ) | ( x39 & n9226 ) | ( ~n9225 & n9226 ) ;
  assign n9228 = n9225 | n9227 ;
  assign n9229 = ~n9123 & n9228 ;
  assign n9230 = x75 & ~n9229 ;
  assign n9231 = ( n6782 & n9213 ) | ( n6782 & ~n9230 ) | ( n9213 & ~n9230 ) ;
  assign n9232 = ~n6782 & n9231 ;
  assign n9233 = x207 & x208 ;
  assign n9234 = n6782 & n9193 ;
  assign n9235 = ( ~n9232 & n9233 ) | ( ~n9232 & n9234 ) | ( n9233 & n9234 ) ;
  assign n9236 = n9232 | n9235 ;
  assign n9237 = ~x72 & x200 ;
  assign n9238 = x232 | n9237 ;
  assign n9239 = ~x299 & n9238 ;
  assign n9240 = x200 & n9119 ;
  assign n9241 = x232 & ~n9240 ;
  assign n9242 = n9239 & ~n9241 ;
  assign n9243 = x39 & ~n9242 ;
  assign n9244 = ~n9122 & n9243 ;
  assign n9245 = n9207 & ~n9244 ;
  assign n9246 = x38 & ~n9245 ;
  assign n9247 = x87 | n9246 ;
  assign n9248 = n9181 ^ x39 ^ 1'b0 ;
  assign n9249 = x200 & n9184 ;
  assign n9250 = n9186 & ~n9249 ;
  assign n9251 = n9118 | n9239 ;
  assign n9252 = ~n9250 & n9251 ;
  assign n9253 = ( n9181 & n9248 ) | ( n9181 & n9252 ) | ( n9248 & n9252 ) ;
  assign n9254 = ( x38 & x100 ) | ( x38 & ~n9253 ) | ( x100 & ~n9253 ) ;
  assign n9255 = n9253 | n9254 ;
  assign n9256 = n9115 & ~n9244 ;
  assign n9257 = n5018 & ~n9256 ;
  assign n9258 = ( n9247 & n9255 ) | ( n9247 & ~n9257 ) | ( n9255 & ~n9257 ) ;
  assign n9259 = ~n9247 & n9258 ;
  assign n9260 = n9210 & ~n9244 ;
  assign n9261 = ( x75 & ~n9259 ) | ( x75 & n9260 ) | ( ~n9259 & n9260 ) ;
  assign n9262 = n9259 | n9261 ;
  assign n9263 = n9228 & ~n9244 ;
  assign n9264 = x75 & ~n9263 ;
  assign n9265 = ( n6782 & n9262 ) | ( n6782 & ~n9264 ) | ( n9262 & ~n9264 ) ;
  assign n9266 = ~n6782 & n9265 ;
  assign n9267 = n6782 & n9245 ;
  assign n9268 = n9233 & ~n9267 ;
  assign n9269 = n9236 & ~n9268 ;
  assign n9270 = ( n9236 & n9266 ) | ( n9236 & n9269 ) | ( n9266 & n9269 ) ;
  assign n9271 = x211 & x214 ;
  assign n9272 = x212 & n9271 ;
  assign n9273 = ( x219 & ~n9270 ) | ( x219 & n9272 ) | ( ~n9270 & n9272 ) ;
  assign n9274 = n9270 | n9273 ;
  assign n9275 = x219 | n9272 ;
  assign n9276 = ~x166 & n6411 ;
  assign n9277 = x72 | n9276 ;
  assign n9278 = n9275 & ~n9277 ;
  assign n9279 = x39 & ~n9278 ;
  assign n9280 = ( n7318 & n9207 ) | ( n7318 & n9279 ) | ( n9207 & n9279 ) ;
  assign n9281 = ~n9279 & n9280 ;
  assign n9282 = x299 & ~n9277 ;
  assign n9283 = x39 & ~n9282 ;
  assign n9284 = ~n9122 & n9283 ;
  assign n9285 = n9243 & n9284 ;
  assign n9286 = n9228 & ~n9285 ;
  assign n9287 = x75 & ~n9286 ;
  assign n9288 = n9209 & ~n9285 ;
  assign n9289 = n9206 & n9288 ;
  assign n9290 = n9207 & ~n9284 ;
  assign n9291 = x38 & ~n9290 ;
  assign n9292 = x87 | n9291 ;
  assign n9293 = n9247 & n9292 ;
  assign n9294 = n9115 & ~n9285 ;
  assign n9295 = ~n9293 & n9294 ;
  assign n9296 = ( n5018 & n9293 ) | ( n5018 & ~n9295 ) | ( n9293 & ~n9295 ) ;
  assign n9297 = x232 & x299 ;
  assign n9298 = n9277 & n9297 ;
  assign n9299 = ~n8898 & n8962 ;
  assign n9300 = n9298 & ~n9299 ;
  assign n9301 = x72 & ~x232 ;
  assign n9302 = x299 & ~n9301 ;
  assign n9303 = n9117 | n9302 ;
  assign n9304 = n9237 | n9303 ;
  assign n9305 = ~x299 & n9250 ;
  assign n9306 = ( n9300 & n9304 ) | ( n9300 & ~n9305 ) | ( n9304 & ~n9305 ) ;
  assign n9307 = ~n9300 & n9306 ;
  assign n9308 = ( n9181 & n9248 ) | ( n9181 & n9307 ) | ( n9248 & n9307 ) ;
  assign n9309 = ( n1205 & ~n9296 ) | ( n1205 & n9308 ) | ( ~n9296 & n9308 ) ;
  assign n9310 = ~n9296 & n9309 ;
  assign n9311 = ( x75 & ~n9289 ) | ( x75 & n9310 ) | ( ~n9289 & n9310 ) ;
  assign n9312 = n9289 | n9311 ;
  assign n9313 = ( n6782 & ~n9287 ) | ( n6782 & n9312 ) | ( ~n9287 & n9312 ) ;
  assign n9314 = ~n6782 & n9313 ;
  assign n9315 = ( n9233 & n9267 ) | ( n9233 & ~n9314 ) | ( n9267 & ~n9314 ) ;
  assign n9316 = ~n9267 & n9315 ;
  assign n9317 = n9228 & ~n9284 ;
  assign n9318 = x75 & ~n9317 ;
  assign n9319 = n9210 & ~n9284 ;
  assign n9320 = n9115 & ~n9284 ;
  assign n9321 = n5018 & ~n9320 ;
  assign n9322 = n9292 | n9321 ;
  assign n9323 = x232 & ~x299 ;
  assign n9324 = ~n9185 & n9323 ;
  assign n9325 = ~n9300 & n9303 ;
  assign n9326 = ~n9324 & n9325 ;
  assign n9327 = ( n9181 & n9248 ) | ( n9181 & n9326 ) | ( n9248 & n9326 ) ;
  assign n9328 = ( n1205 & ~n9322 ) | ( n1205 & n9327 ) | ( ~n9322 & n9327 ) ;
  assign n9329 = ~n9322 & n9328 ;
  assign n9330 = ( x75 & ~n9319 ) | ( x75 & n9329 ) | ( ~n9319 & n9329 ) ;
  assign n9331 = n9319 | n9330 ;
  assign n9332 = ( n6782 & ~n9318 ) | ( n6782 & n9331 ) | ( ~n9318 & n9331 ) ;
  assign n9333 = ~n6782 & n9332 ;
  assign n9334 = ( n9233 & ~n9316 ) | ( n9233 & n9333 ) | ( ~n9316 & n9333 ) ;
  assign n9335 = ~n9316 & n9334 ;
  assign n9336 = n6782 & n9290 ;
  assign n9337 = ( n9275 & n9335 ) | ( n9275 & ~n9336 ) | ( n9335 & ~n9336 ) ;
  assign n9338 = ~n9335 & n9337 ;
  assign n9339 = ( x57 & n5193 ) | ( x57 & ~n9338 ) | ( n5193 & ~n9338 ) ;
  assign n9340 = n9338 | n9339 ;
  assign n9341 = ~n9281 & n9340 ;
  assign n9342 = ( n9274 & n9281 ) | ( n9274 & ~n9341 ) | ( n9281 & ~n9341 ) ;
  assign n9343 = x211 | x219 ;
  assign n9344 = x212 & x214 ;
  assign n9345 = n9344 ^ n9343 ^ 1'b0 ;
  assign n9346 = ( x211 & ~n9343 ) | ( x211 & n9345 ) | ( ~n9343 & n9345 ) ;
  assign n9347 = ~n9277 & n9346 ;
  assign n9348 = x39 & ~n9347 ;
  assign n9349 = x43 & ~x72 ;
  assign n9350 = x39 | n9349 ;
  assign n9351 = ( n7318 & n9348 ) | ( n7318 & n9350 ) | ( n9348 & n9350 ) ;
  assign n9352 = ~n9348 & n9351 ;
  assign n9353 = x199 | x200 ;
  assign n9354 = ~x299 & n9353 ;
  assign n9355 = ( ~x232 & n9301 ) | ( ~x232 & n9354 ) | ( n9301 & n9354 ) ;
  assign n9356 = x299 | n9355 ;
  assign n9357 = n9119 & ~n9353 ;
  assign n9358 = x232 & ~n9357 ;
  assign n9359 = n9356 | n9358 ;
  assign n9360 = x39 & n9359 ;
  assign n9361 = ~n9282 & n9360 ;
  assign n9362 = n9350 & ~n9361 ;
  assign n9363 = n6782 & n9362 ;
  assign n9364 = x38 & ~n9362 ;
  assign n9365 = n6824 | n9349 ;
  assign n9366 = x42 | n5031 ;
  assign n9367 = n1615 & ~n9366 ;
  assign n9368 = n9349 & ~n9367 ;
  assign n9369 = ~x43 & x52 ;
  assign n9370 = n9098 & n9369 ;
  assign n9371 = x43 & ~n9105 ;
  assign n9372 = n9370 | n9371 ;
  assign n9373 = n9367 & n9372 ;
  assign n9374 = ( n6824 & n9368 ) | ( n6824 & ~n9373 ) | ( n9368 & ~n9373 ) ;
  assign n9375 = ~n9368 & n9374 ;
  assign n9376 = ( x39 & n9365 ) | ( x39 & ~n9375 ) | ( n9365 & ~n9375 ) ;
  assign n9377 = n9376 ^ n9365 ^ 1'b0 ;
  assign n9378 = ( x39 & n9376 ) | ( x39 & ~n9377 ) | ( n9376 & ~n9377 ) ;
  assign n9379 = ~n9361 & n9378 ;
  assign n9380 = n5018 & ~n9379 ;
  assign n9381 = ( x87 & ~n9364 ) | ( x87 & n9380 ) | ( ~n9364 & n9380 ) ;
  assign n9382 = n9364 | n9381 ;
  assign n9383 = ~n9349 & n9366 ;
  assign n9384 = n1615 & ~n9148 ;
  assign n9385 = n1615 | n9162 ;
  assign n9386 = ~n9384 & n9385 ;
  assign n9387 = ~n5030 & n9386 ;
  assign n9388 = n9140 ^ x228 ^ 1'b0 ;
  assign n9389 = ( n9140 & n9387 ) | ( n9140 & n9388 ) | ( n9387 & n9388 ) ;
  assign n9390 = x43 | n9389 ;
  assign n9391 = ~n9383 & n9390 ;
  assign n9392 = n9156 ^ n1615 ^ 1'b0 ;
  assign n9393 = ( n9156 & n9171 ) | ( n9156 & ~n9392 ) | ( n9171 & ~n9392 ) ;
  assign n9394 = n9136 ^ x228 ^ 1'b0 ;
  assign n9395 = ( n9136 & n9393 ) | ( n9136 & n9394 ) | ( n9393 & n9394 ) ;
  assign n9396 = x43 & ~n9366 ;
  assign n9397 = n9395 & n9396 ;
  assign n9398 = ( x39 & n9391 ) | ( x39 & ~n9397 ) | ( n9391 & ~n9397 ) ;
  assign n9399 = n9398 ^ n9391 ^ 1'b0 ;
  assign n9400 = ( x39 & n9398 ) | ( x39 & ~n9399 ) | ( n9398 & ~n9399 ) ;
  assign n9401 = n9184 & ~n9353 ;
  assign n9402 = n9323 & ~n9401 ;
  assign n9403 = n9300 | n9355 ;
  assign n9404 = ( x39 & n9402 ) | ( x39 & n9403 ) | ( n9402 & n9403 ) ;
  assign n9405 = n9403 ^ n9402 ^ 1'b0 ;
  assign n9406 = ( x39 & n9404 ) | ( x39 & n9405 ) | ( n9404 & n9405 ) ;
  assign n9407 = n9400 & ~n9406 ;
  assign n9408 = ( n1205 & ~n9382 ) | ( n1205 & n9407 ) | ( ~n9382 & n9407 ) ;
  assign n9409 = ~n9382 & n9408 ;
  assign n9410 = n1205 & ~n9350 ;
  assign n9411 = x87 & ~n9410 ;
  assign n9412 = x228 & ~n9366 ;
  assign n9413 = n9349 & ~n9412 ;
  assign n9414 = ~x43 & n9097 ;
  assign n9415 = x43 & ~n9104 ;
  assign n9416 = ( n9412 & n9414 ) | ( n9412 & ~n9415 ) | ( n9414 & ~n9415 ) ;
  assign n9417 = ~n9414 & n9416 ;
  assign n9418 = ( n2036 & ~n9413 ) | ( n2036 & n9417 ) | ( ~n9413 & n9417 ) ;
  assign n9419 = n9413 | n9418 ;
  assign n9420 = n9411 & n9419 ;
  assign n9421 = ~n9361 & n9420 ;
  assign n9422 = ( x75 & ~n9409 ) | ( x75 & n9421 ) | ( ~n9409 & n9421 ) ;
  assign n9423 = n9409 | n9422 ;
  assign n9424 = n6414 & n9098 ;
  assign n9425 = n9369 & n9424 ;
  assign n9426 = x72 | n9216 ;
  assign n9427 = x43 & ~n9426 ;
  assign n9428 = n9425 | n9427 ;
  assign n9429 = n9367 & n9428 ;
  assign n9430 = ( n6824 & n9368 ) | ( n6824 & ~n9429 ) | ( n9368 & ~n9429 ) ;
  assign n9431 = ~n9368 & n9430 ;
  assign n9432 = ( x39 & n9365 ) | ( x39 & ~n9431 ) | ( n9365 & ~n9431 ) ;
  assign n9433 = n9432 ^ n9365 ^ 1'b0 ;
  assign n9434 = ( x39 & n9432 ) | ( x39 & ~n9433 ) | ( n9432 & ~n9433 ) ;
  assign n9435 = n9350 ^ n2052 ^ 1'b0 ;
  assign n9436 = ( n9350 & n9434 ) | ( n9350 & ~n9435 ) | ( n9434 & ~n9435 ) ;
  assign n9437 = ~n9361 & n9436 ;
  assign n9438 = x75 & ~n9437 ;
  assign n9439 = ( n6782 & n9423 ) | ( n6782 & ~n9438 ) | ( n9423 & ~n9438 ) ;
  assign n9440 = ~n6782 & n9439 ;
  assign n9441 = ( n9233 & n9363 ) | ( n9233 & ~n9440 ) | ( n9363 & ~n9440 ) ;
  assign n9442 = ~n9363 & n9441 ;
  assign n9443 = ~n9242 & n9283 ;
  assign n9444 = n9350 & ~n9443 ;
  assign n9445 = x38 & ~n9444 ;
  assign n9446 = n9378 & ~n9443 ;
  assign n9447 = n5018 & ~n9446 ;
  assign n9448 = ( x87 & ~n9445 ) | ( x87 & n9447 ) | ( ~n9445 & n9447 ) ;
  assign n9449 = n9445 | n9448 ;
  assign n9452 = ~n9249 & n9323 ;
  assign n9450 = n9238 | n9302 ;
  assign n9451 = ~n9300 & n9450 ;
  assign n9453 = n9452 ^ n9451 ^ 1'b0 ;
  assign n9454 = ( x39 & ~n9451 ) | ( x39 & n9452 ) | ( ~n9451 & n9452 ) ;
  assign n9455 = ( x39 & ~n9453 ) | ( x39 & n9454 ) | ( ~n9453 & n9454 ) ;
  assign n9456 = ( n9383 & n9390 ) | ( n9383 & ~n9397 ) | ( n9390 & ~n9397 ) ;
  assign n9457 = ~n9383 & n9456 ;
  assign n9458 = ( x39 & ~n9455 ) | ( x39 & n9457 ) | ( ~n9455 & n9457 ) ;
  assign n9459 = ~n9455 & n9458 ;
  assign n9460 = ( n1205 & ~n9449 ) | ( n1205 & n9459 ) | ( ~n9449 & n9459 ) ;
  assign n9461 = ~n9449 & n9460 ;
  assign n9462 = n9420 & ~n9443 ;
  assign n9463 = ( x75 & ~n9461 ) | ( x75 & n9462 ) | ( ~n9461 & n9462 ) ;
  assign n9464 = n9461 | n9463 ;
  assign n9465 = n9436 & ~n9443 ;
  assign n9466 = x75 & ~n9465 ;
  assign n9467 = ( n6782 & n9464 ) | ( n6782 & ~n9466 ) | ( n9464 & ~n9466 ) ;
  assign n9468 = ~n6782 & n9467 ;
  assign n9469 = n6782 & n9444 ;
  assign n9470 = ( n9233 & ~n9468 ) | ( n9233 & n9469 ) | ( ~n9468 & n9469 ) ;
  assign n9471 = n9468 | n9470 ;
  assign n9472 = n9346 & ~n9471 ;
  assign n9473 = ( n9346 & n9442 ) | ( n9346 & n9472 ) | ( n9442 & n9472 ) ;
  assign n9474 = ~n9360 & n9436 ;
  assign n9475 = x75 & ~n9474 ;
  assign n9476 = x39 & ~n9359 ;
  assign n9477 = ( n9350 & ~n9360 ) | ( n9350 & n9476 ) | ( ~n9360 & n9476 ) ;
  assign n9478 = n2095 & ~n9477 ;
  assign n9479 = n9420 & ~n9478 ;
  assign n9480 = x38 & ~n9477 ;
  assign n9481 = ~n9360 & n9378 ;
  assign n9482 = n5018 & ~n9481 ;
  assign n9483 = ( x87 & ~n9480 ) | ( x87 & n9482 ) | ( ~n9480 & n9482 ) ;
  assign n9484 = n9480 | n9483 ;
  assign n9485 = x232 & ~n9401 ;
  assign n9486 = n9356 | n9485 ;
  assign n9487 = x39 & n9486 ;
  assign n9488 = n9400 & ~n9487 ;
  assign n9489 = ( n1205 & ~n9484 ) | ( n1205 & n9488 ) | ( ~n9484 & n9488 ) ;
  assign n9490 = ~n9484 & n9489 ;
  assign n9491 = ( x75 & ~n9479 ) | ( x75 & n9490 ) | ( ~n9479 & n9490 ) ;
  assign n9492 = n9479 | n9491 ;
  assign n9493 = ( n6782 & ~n9475 ) | ( n6782 & n9492 ) | ( ~n9475 & n9492 ) ;
  assign n9494 = ~n6782 & n9493 ;
  assign n9495 = n6782 & n9477 ;
  assign n9496 = ( n9233 & n9494 ) | ( n9233 & ~n9495 ) | ( n9494 & ~n9495 ) ;
  assign n9497 = ~n9494 & n9496 ;
  assign n9498 = ~n9243 & n9436 ;
  assign n9499 = x75 & ~n9498 ;
  assign n9500 = ~n9243 & n9420 ;
  assign n9501 = ~n9243 & n9350 ;
  assign n9502 = x38 & ~n9501 ;
  assign n9503 = ~n9243 & n9378 ;
  assign n9504 = n5018 & ~n9503 ;
  assign n9505 = ( x87 & ~n9502 ) | ( x87 & n9504 ) | ( ~n9502 & n9504 ) ;
  assign n9506 = n9502 | n9505 ;
  assign n9507 = x232 & ~n9249 ;
  assign n9508 = x39 & ~n9239 ;
  assign n9509 = ( x39 & n9507 ) | ( x39 & n9508 ) | ( n9507 & n9508 ) ;
  assign n9510 = ( x39 & n9457 ) | ( x39 & ~n9509 ) | ( n9457 & ~n9509 ) ;
  assign n9511 = ~n9509 & n9510 ;
  assign n9512 = ( n1205 & ~n9506 ) | ( n1205 & n9511 ) | ( ~n9506 & n9511 ) ;
  assign n9513 = ~n9506 & n9512 ;
  assign n9514 = ( x75 & ~n9500 ) | ( x75 & n9513 ) | ( ~n9500 & n9513 ) ;
  assign n9515 = n9500 | n9514 ;
  assign n9516 = ( n6782 & ~n9499 ) | ( n6782 & n9515 ) | ( ~n9499 & n9515 ) ;
  assign n9517 = ~n6782 & n9516 ;
  assign n9518 = n6782 | n9233 ;
  assign n9519 = ( n9233 & n9501 ) | ( n9233 & n9518 ) | ( n9501 & n9518 ) ;
  assign n9520 = ( ~n9497 & n9517 ) | ( ~n9497 & n9519 ) | ( n9517 & n9519 ) ;
  assign n9521 = ~n9497 & n9520 ;
  assign n9522 = ( ~n7318 & n9346 ) | ( ~n7318 & n9521 ) | ( n9346 & n9521 ) ;
  assign n9523 = ~n7318 & n9522 ;
  assign n9524 = ( n9352 & ~n9473 ) | ( n9352 & n9523 ) | ( ~n9473 & n9523 ) ;
  assign n9525 = n9473 ^ n9352 ^ 1'b0 ;
  assign n9526 = ( n9352 & n9524 ) | ( n9352 & ~n9525 ) | ( n9524 & ~n9525 ) ;
  assign n9527 = x39 & n6412 ;
  assign n9528 = ~x72 & n9527 ;
  assign n9529 = ~x72 & n6412 ;
  assign n9530 = x39 & ~n9529 ;
  assign n9531 = x39 | n8996 ;
  assign n9532 = ( n9528 & ~n9530 ) | ( n9528 & n9531 ) | ( ~n9530 & n9531 ) ;
  assign n9533 = n2052 & n9532 ;
  assign n9534 = n6824 | n8996 ;
  assign n9535 = ~n1615 & n8996 ;
  assign n9536 = n6824 & ~n9535 ;
  assign n9537 = n6416 & ~n9001 ;
  assign n9538 = n6480 & ~n8919 ;
  assign n9539 = n6414 & n9538 ;
  assign n9540 = x44 & ~n8932 ;
  assign n9541 = n9539 | n9540 ;
  assign n9542 = n9536 & ~n9541 ;
  assign n9543 = ( n9536 & ~n9537 ) | ( n9536 & n9542 ) | ( ~n9537 & n9542 ) ;
  assign n9544 = ( x39 & n9534 ) | ( x39 & ~n9543 ) | ( n9534 & ~n9543 ) ;
  assign n9545 = ~x39 & n9544 ;
  assign n9546 = ( ~n2052 & n9528 ) | ( ~n2052 & n9545 ) | ( n9528 & n9545 ) ;
  assign n9547 = ~n2052 & n9546 ;
  assign n9548 = ( x75 & n9533 ) | ( x75 & ~n9547 ) | ( n9533 & ~n9547 ) ;
  assign n9549 = ~n9533 & n9548 ;
  assign n9550 = x228 & ~n1205 ;
  assign n9551 = ~n8948 & n9550 ;
  assign n9552 = n8996 & ~n9551 ;
  assign n9553 = ~n8919 & n9550 ;
  assign n9554 = ( x39 & ~n9552 ) | ( x39 & n9553 ) | ( ~n9552 & n9553 ) ;
  assign n9555 = n9552 | n9554 ;
  assign n9556 = n9555 ^ x75 ^ 1'b0 ;
  assign n9557 = x87 & ~n9530 ;
  assign n9558 = ( n9555 & ~n9556 ) | ( n9555 & n9557 ) | ( ~n9556 & n9557 ) ;
  assign n9559 = ( x75 & n9556 ) | ( x75 & n9558 ) | ( n9556 & n9558 ) ;
  assign n9560 = x38 & ~n9532 ;
  assign n9561 = x87 | n9560 ;
  assign n9565 = n1615 & ~n9046 ;
  assign n9566 = ~n9053 & n9565 ;
  assign n9562 = n1615 | n9012 ;
  assign n9563 = x44 & ~n9024 ;
  assign n9564 = n9562 | n9563 ;
  assign n9567 = n9566 ^ n9564 ^ 1'b0 ;
  assign n9568 = ( x228 & ~n9564 ) | ( x228 & n9566 ) | ( ~n9564 & n9566 ) ;
  assign n9569 = ( x228 & ~n9567 ) | ( x228 & n9568 ) | ( ~n9567 & n9568 ) ;
  assign n9570 = x44 & ~n9000 ;
  assign n9571 = ( x228 & n8993 ) | ( x228 & ~n9570 ) | ( n8993 & ~n9570 ) ;
  assign n9572 = n9570 | n9571 ;
  assign n9573 = ( x39 & ~n9569 ) | ( x39 & n9572 ) | ( ~n9569 & n9572 ) ;
  assign n9574 = ~x39 & n9573 ;
  assign n9575 = x287 & ~n8948 ;
  assign n9576 = x72 | n9575 ;
  assign n9577 = n9527 & ~n9576 ;
  assign n9578 = ( n1205 & ~n9574 ) | ( n1205 & n9577 ) | ( ~n9574 & n9577 ) ;
  assign n9579 = n9574 | n9578 ;
  assign n9580 = ~x39 & n9534 ;
  assign n9581 = ~n9536 & n9580 ;
  assign n9582 = n6480 & ~n8948 ;
  assign n9583 = x44 & ~n9582 ;
  assign n9584 = n9538 | n9583 ;
  assign n9585 = n9537 & n9584 ;
  assign n9586 = ( n9580 & n9581 ) | ( n9580 & n9585 ) | ( n9581 & n9585 ) ;
  assign n9587 = ( n5018 & n9528 ) | ( n5018 & ~n9586 ) | ( n9528 & ~n9586 ) ;
  assign n9588 = ~n9528 & n9587 ;
  assign n9589 = ( n9561 & n9579 ) | ( n9561 & ~n9588 ) | ( n9579 & ~n9588 ) ;
  assign n9590 = ~n9561 & n9589 ;
  assign n9591 = ( ~n9549 & n9559 ) | ( ~n9549 & n9590 ) | ( n9559 & n9590 ) ;
  assign n9592 = ~n9549 & n9591 ;
  assign n9593 = ( x74 & n5015 ) | ( x74 & ~n9592 ) | ( n5015 & ~n9592 ) ;
  assign n9594 = n9592 | n9593 ;
  assign n9595 = ~n1329 & n6411 ;
  assign n9596 = ~x72 & n9595 ;
  assign n9597 = x39 & ~n9596 ;
  assign n9598 = n7318 & ~n9597 ;
  assign n9599 = n9531 & n9598 ;
  assign n9600 = n6782 & ~n9532 ;
  assign n9601 = n7318 | n9600 ;
  assign n9602 = ~n9599 & n9601 ;
  assign n9603 = ( n9594 & n9599 ) | ( n9594 & ~n9602 ) | ( n9599 & ~n9602 ) ;
  assign n9604 = ~x38 & x39 ;
  assign n9605 = ~n8793 & n9604 ;
  assign n9606 = x979 & n9605 ;
  assign n9607 = ~n5362 & n9606 ;
  assign n9608 = ~n1372 & n1840 ;
  assign n9609 = x24 & n9608 ;
  assign n9610 = x49 | x76 ;
  assign n9611 = n7490 | n9610 ;
  assign n9612 = x102 | x104 ;
  assign n9613 = x111 | n9612 ;
  assign n9614 = n8771 | n9613 ;
  assign n9615 = n9611 | n9614 ;
  assign n9616 = x61 & ~x82 ;
  assign n9617 = x83 | x89 ;
  assign n9618 = n9616 & ~n9617 ;
  assign n9619 = n6379 | n7501 ;
  assign n9620 = ( n7487 & n9618 ) | ( n7487 & ~n9619 ) | ( n9618 & ~n9619 ) ;
  assign n9621 = ~n7487 & n9620 ;
  assign n9622 = ( n8797 & ~n8798 ) | ( n8797 & n9621 ) | ( ~n8798 & n9621 ) ;
  assign n9623 = ~n8797 & n9622 ;
  assign n9624 = ( n7511 & ~n9615 ) | ( n7511 & n9623 ) | ( ~n9615 & n9623 ) ;
  assign n9625 = ~n7511 & n9624 ;
  assign n9626 = ~x841 & n9625 ;
  assign n9627 = ( ~n8761 & n9609 ) | ( ~n8761 & n9626 ) | ( n9609 & n9626 ) ;
  assign n9628 = ~n8761 & n9627 ;
  assign n9629 = n1473 | n6379 ;
  assign n9630 = n7500 | n7586 ;
  assign n9631 = x82 | n1239 ;
  assign n9632 = ~x84 & x104 ;
  assign n9633 = ( n1490 & ~n8774 ) | ( n1490 & n9632 ) | ( ~n8774 & n9632 ) ;
  assign n9634 = ~n1490 & n9633 ;
  assign n9635 = n9634 ^ n9631 ^ 1'b0 ;
  assign n9636 = ( n9631 & n9634 ) | ( n9631 & n9635 ) | ( n9634 & n9635 ) ;
  assign n9637 = ( x36 & ~n9631 ) | ( x36 & n9636 ) | ( ~n9631 & n9636 ) ;
  assign n9638 = x67 | x103 ;
  assign n9639 = n1230 | n9638 ;
  assign n9640 = x98 | n9639 ;
  assign n9641 = ( n9630 & n9637 ) | ( n9630 & ~n9640 ) | ( n9637 & ~n9640 ) ;
  assign n9642 = ~n9630 & n9641 ;
  assign n9643 = ~n1528 & n9642 ;
  assign n9644 = x88 | n9643 ;
  assign n9645 = ( n1408 & ~n9629 ) | ( n1408 & n9644 ) | ( ~n9629 & n9644 ) ;
  assign n9646 = ~n1408 & n9645 ;
  assign n9647 = ~n1370 & n9646 ;
  assign n9648 = ( n8754 & ~n8757 ) | ( n8754 & n9647 ) | ( ~n8757 & n9647 ) ;
  assign n9649 = ~n8757 & n9648 ;
  assign n9650 = n6490 & ~n9649 ;
  assign n9651 = n1272 | n8770 ;
  assign n9652 = ~x36 & n9642 ;
  assign n9653 = x88 | n9652 ;
  assign n9654 = ~n9629 & n9653 ;
  assign n9655 = ~n9651 & n9654 ;
  assign n9656 = ~x824 & n5020 ;
  assign n9657 = n9655 & n9656 ;
  assign n9658 = ~n5020 & n9649 ;
  assign n9659 = ( x829 & n9657 ) | ( x829 & ~n9658 ) | ( n9657 & ~n9658 ) ;
  assign n9660 = ~n9657 & n9659 ;
  assign n9661 = ~n1614 & n9660 ;
  assign n9662 = ( x1091 & n9650 ) | ( x1091 & n9661 ) | ( n9650 & n9661 ) ;
  assign n9663 = n9661 ^ n9650 ^ 1'b0 ;
  assign n9664 = ( x1091 & n9662 ) | ( x1091 & n9663 ) | ( n9662 & n9663 ) ;
  assign n9665 = ~n6425 & n9649 ;
  assign n9666 = n6425 & ~n8757 ;
  assign n9667 = n8755 & n9666 ;
  assign n9668 = n5377 & ~n6489 ;
  assign n9669 = n9667 | n9668 ;
  assign n9670 = ( ~n8760 & n9665 ) | ( ~n8760 & n9669 ) | ( n9665 & n9669 ) ;
  assign n9671 = ~n8760 & n9670 ;
  assign n9672 = x829 | n9665 ;
  assign n9673 = ~n9660 & n9672 ;
  assign n9674 = x1093 | n9673 ;
  assign n9675 = ( n9664 & n9671 ) | ( n9664 & n9674 ) | ( n9671 & n9674 ) ;
  assign n9676 = ~n9664 & n9675 ;
  assign n9677 = ~x72 & x841 ;
  assign n9678 = ~n1375 & n9677 ;
  assign n9679 = ~x51 & n9678 ;
  assign n9680 = n8808 & n9679 ;
  assign n9681 = ( n8760 & ~n8770 ) | ( n8760 & n9680 ) | ( ~n8770 & n9680 ) ;
  assign n9682 = ~n8760 & n9681 ;
  assign n9683 = x103 | n1522 ;
  assign n9684 = n8797 | n9683 ;
  assign n9685 = n7490 | n7500 ;
  assign n9686 = n9684 | n9685 ;
  assign n9687 = n1228 | n1230 ;
  assign n9688 = ~x45 & x49 ;
  assign n9689 = ~n9613 & n9688 ;
  assign n9690 = ~n9687 & n9689 ;
  assign n9691 = ( n9631 & ~n9686 ) | ( n9631 & n9690 ) | ( ~n9686 & n9690 ) ;
  assign n9692 = ~n9631 & n9691 ;
  assign n9693 = n1376 | n7511 ;
  assign n9694 = n9692 & ~n9693 ;
  assign n9695 = ~n8756 & n9678 ;
  assign n9696 = n9694 & n9695 ;
  assign n9697 = x74 | n9696 ;
  assign n9698 = ( ~n6336 & n7318 ) | ( ~n6336 & n9697 ) | ( n7318 & n9697 ) ;
  assign n9699 = ~n7318 & n9698 ;
  assign n9700 = ( x74 & n7455 ) | ( x74 & ~n9699 ) | ( n7455 & ~n9699 ) ;
  assign n9701 = n9700 ^ n9699 ^ 1'b0 ;
  assign n9702 = ( n9699 & ~n9700 ) | ( n9699 & n9701 ) | ( ~n9700 & n9701 ) ;
  assign n9703 = n7451 ^ x252 ^ 1'b0 ;
  assign n9704 = ( n7451 & n7457 ) | ( n7451 & ~n9703 ) | ( n7457 & ~n9703 ) ;
  assign n9705 = x24 & ~x94 ;
  assign n9706 = ~n7470 & n9705 ;
  assign n9707 = ( n8757 & n9704 ) | ( n8757 & ~n9706 ) | ( n9704 & ~n9706 ) ;
  assign n9708 = ~n8757 & n9707 ;
  assign n9709 = x24 & ~n7472 ;
  assign n9710 = n9709 ^ n8981 ^ 1'b0 ;
  assign n9711 = ( n8981 & n9709 ) | ( n8981 & ~n9710 ) | ( n9709 & ~n9710 ) ;
  assign n9712 = ( n9708 & n9710 ) | ( n9708 & n9711 ) | ( n9710 & n9711 ) ;
  assign n9713 = n1411 | n6399 ;
  assign n9714 = x24 & ~x90 ;
  assign n9715 = ( n9704 & ~n9713 ) | ( n9704 & n9714 ) | ( ~n9713 & n9714 ) ;
  assign n9716 = ~n9704 & n9715 ;
  assign n9717 = n7474 & n9716 ;
  assign n9718 = ( ~x100 & n9712 ) | ( ~x100 & n9717 ) | ( n9712 & n9717 ) ;
  assign n9719 = ~x100 & n9718 ;
  assign n9720 = n9719 ^ n5421 ^ 1'b0 ;
  assign n9721 = x100 & n5044 ;
  assign n9722 = ( n5421 & ~n9720 ) | ( n5421 & n9721 ) | ( ~n9720 & n9721 ) ;
  assign n9723 = ( n9719 & n9720 ) | ( n9719 & n9722 ) | ( n9720 & n9722 ) ;
  assign n9724 = n5045 & n7461 ;
  assign n9725 = ~n7456 & n9724 ;
  assign n9726 = n1994 | n2044 ;
  assign n9727 = ~n9725 & n9726 ;
  assign n9728 = ( n9723 & n9725 ) | ( n9723 & ~n9727 ) | ( n9725 & ~n9727 ) ;
  assign n9729 = ( n5015 & ~n7448 ) | ( n5015 & n9728 ) | ( ~n7448 & n9728 ) ;
  assign n9730 = ~n5015 & n9729 ;
  assign n9731 = n1370 | n8761 ;
  assign n9732 = n1408 | n9731 ;
  assign n9733 = n7587 | n9687 ;
  assign n9734 = n1232 | n9733 ;
  assign n9735 = x69 | n9734 ;
  assign n9736 = n1522 | n9735 ;
  assign n9737 = n1524 & ~n9736 ;
  assign n9738 = ~n9732 & n9737 ;
  assign n9739 = x52 & ~x72 ;
  assign n9740 = ~x39 & n9739 ;
  assign n9741 = x211 | n9344 ;
  assign n9742 = x219 | n9741 ;
  assign n9743 = x39 & ~n9742 ;
  assign n9744 = ~n9277 & n9743 ;
  assign n9745 = ( n7318 & n9740 ) | ( n7318 & ~n9744 ) | ( n9740 & ~n9744 ) ;
  assign n9746 = ~n9740 & n9745 ;
  assign n9747 = n6782 & ~n9740 ;
  assign n9748 = n9233 & ~n9747 ;
  assign n9749 = n5028 | n5031 ;
  assign n9750 = ~n9739 & n9749 ;
  assign n9751 = ~x52 & n9140 ;
  assign n9752 = n9749 | n9751 ;
  assign n9753 = n9136 & ~n9752 ;
  assign n9754 = ( x52 & n9752 ) | ( x52 & ~n9753 ) | ( n9752 & ~n9753 ) ;
  assign n9755 = ( x228 & ~n9750 ) | ( x228 & n9754 ) | ( ~n9750 & n9754 ) ;
  assign n9756 = ~x228 & n9755 ;
  assign n9757 = ~x52 & n9149 ;
  assign n9758 = x52 & ~n9156 ;
  assign n9759 = ( n9093 & n9757 ) | ( n9093 & ~n9758 ) | ( n9757 & ~n9758 ) ;
  assign n9760 = ~n9757 & n9759 ;
  assign n9761 = x115 | n1615 ;
  assign n9762 = ~x52 & n9163 ;
  assign n9763 = n9761 | n9762 ;
  assign n9764 = x52 & ~n9171 ;
  assign n9765 = ( ~n9760 & n9763 ) | ( ~n9760 & n9764 ) | ( n9763 & n9764 ) ;
  assign n9766 = ~n9760 & n9765 ;
  assign n9767 = ( x114 & n5028 ) | ( x114 & ~n9766 ) | ( n5028 & ~n9766 ) ;
  assign n9768 = n9766 | n9767 ;
  assign n9769 = ( x228 & n9750 ) | ( x228 & n9768 ) | ( n9750 & n9768 ) ;
  assign n9770 = ~n9750 & n9769 ;
  assign n9771 = ( x39 & ~n9756 ) | ( x39 & n9770 ) | ( ~n9756 & n9770 ) ;
  assign n9772 = n9756 | n9771 ;
  assign n9773 = ~n9487 & n9772 ;
  assign n9774 = n1205 | n9773 ;
  assign n9775 = x87 ^ x75 ^ 1'b0 ;
  assign n9776 = n9476 | n9740 ;
  assign n9777 = n1205 & n9776 ;
  assign n9778 = n9097 ^ x52 ^ 1'b0 ;
  assign n9779 = ( n9097 & ~n9104 ) | ( n9097 & n9778 ) | ( ~n9104 & n9778 ) ;
  assign n9780 = x228 & ~n9749 ;
  assign n9781 = n9780 ^ n9779 ^ 1'b0 ;
  assign n9782 = ( n9739 & ~n9779 ) | ( n9739 & n9781 ) | ( ~n9779 & n9781 ) ;
  assign n9783 = x39 | n9782 ;
  assign n9784 = n1205 | n9360 ;
  assign n9785 = n9783 & ~n9784 ;
  assign n9786 = n9777 | n9785 ;
  assign n9787 = ( x87 & ~n9775 ) | ( x87 & n9786 ) | ( ~n9775 & n9786 ) ;
  assign n9788 = ( x75 & n9775 ) | ( x75 & n9787 ) | ( n9775 & n9787 ) ;
  assign n9789 = x38 & ~n9776 ;
  assign n9790 = x87 | n9789 ;
  assign n9791 = x114 | n5028 ;
  assign n9792 = n9109 & ~n9791 ;
  assign n9793 = n6480 & n9792 ;
  assign n9794 = ~n9103 & n9793 ;
  assign n9795 = n9739 & ~n9794 ;
  assign n9796 = x39 | n9795 ;
  assign n9797 = ~n9360 & n9796 ;
  assign n9798 = ~n9790 & n9797 ;
  assign n9799 = ( n5018 & n9790 ) | ( n5018 & ~n9798 ) | ( n9790 & ~n9798 ) ;
  assign n9800 = ~n9788 & n9799 ;
  assign n9801 = ( n9774 & n9788 ) | ( n9774 & ~n9800 ) | ( n9788 & ~n9800 ) ;
  assign n9802 = n2052 | n9360 ;
  assign n9803 = n9216 & n9792 ;
  assign n9804 = n9739 & ~n9803 ;
  assign n9805 = ( x39 & ~n9802 ) | ( x39 & n9804 ) | ( ~n9802 & n9804 ) ;
  assign n9806 = ~n9802 & n9805 ;
  assign n9807 = n2052 & n9776 ;
  assign n9808 = ( x75 & n9806 ) | ( x75 & ~n9807 ) | ( n9806 & ~n9807 ) ;
  assign n9809 = ~n9806 & n9808 ;
  assign n9810 = ( n9518 & n9801 ) | ( n9518 & ~n9809 ) | ( n9801 & ~n9809 ) ;
  assign n9811 = ~n9518 & n9810 ;
  assign n9812 = ~n2052 & n9803 ;
  assign n9813 = n9740 & ~n9812 ;
  assign n9814 = x75 & n9813 ;
  assign n9815 = ~x100 & n9604 ;
  assign n9816 = x87 & ~n9815 ;
  assign n9817 = x100 & ~n9740 ;
  assign n9818 = n9816 & ~n9817 ;
  assign n9819 = x38 & ~n9740 ;
  assign n9820 = x38 | n9782 ;
  assign n9821 = ~n9819 & n9820 ;
  assign n9822 = x100 | n9821 ;
  assign n9823 = n9818 & n9822 ;
  assign n9824 = x100 & ~n9795 ;
  assign n9825 = x39 | n9824 ;
  assign n9826 = x100 | n9772 ;
  assign n9827 = n9826 ^ n9825 ^ 1'b0 ;
  assign n9828 = ( n9825 & n9826 ) | ( n9825 & n9827 ) | ( n9826 & n9827 ) ;
  assign n9829 = ( x38 & ~n9825 ) | ( x38 & n9828 ) | ( ~n9825 & n9828 ) ;
  assign n9830 = ( x87 & ~n9819 ) | ( x87 & n9829 ) | ( ~n9819 & n9829 ) ;
  assign n9831 = ~x87 & n9830 ;
  assign n9832 = ( ~x75 & n9823 ) | ( ~x75 & n9831 ) | ( n9823 & n9831 ) ;
  assign n9833 = ~x75 & n9832 ;
  assign n9834 = ( n6782 & ~n9814 ) | ( n6782 & n9833 ) | ( ~n9814 & n9833 ) ;
  assign n9835 = n9814 | n9834 ;
  assign n9836 = n9811 ^ n9748 ^ 1'b0 ;
  assign n9837 = ( ~n9748 & n9835 ) | ( ~n9748 & n9836 ) | ( n9835 & n9836 ) ;
  assign n9838 = ( n9748 & n9811 ) | ( n9748 & n9837 ) | ( n9811 & n9837 ) ;
  assign n9839 = n9741 ^ x219 ^ 1'b0 ;
  assign n9840 = ( x219 & n9741 ) | ( x219 & ~n9839 ) | ( n9741 & ~n9839 ) ;
  assign n9841 = ( n9838 & n9839 ) | ( n9838 & n9840 ) | ( n9839 & n9840 ) ;
  assign n9842 = ~n9406 & n9772 ;
  assign n9843 = n1205 | n9842 ;
  assign n9844 = ~n9361 & n9796 ;
  assign n9845 = n5018 & ~n9844 ;
  assign n9846 = ~n9283 & n9796 ;
  assign n9847 = n5018 & ~n9846 ;
  assign n9848 = n9740 ^ n9283 ^ x39 ;
  assign n9849 = ~n9847 & n9848 ;
  assign n9850 = ( n9789 & n9845 ) | ( n9789 & ~n9849 ) | ( n9845 & ~n9849 ) ;
  assign n9851 = ( x87 & n9843 ) | ( x87 & ~n9850 ) | ( n9843 & ~n9850 ) ;
  assign n9852 = n9851 ^ n9843 ^ 1'b0 ;
  assign n9853 = ( x87 & n9851 ) | ( x87 & ~n9852 ) | ( n9851 & ~n9852 ) ;
  assign n9854 = n1205 & n9848 ;
  assign n9855 = x87 & ~n9854 ;
  assign n9856 = n1205 | n9361 ;
  assign n9857 = n9783 & ~n9856 ;
  assign n9858 = ( n9777 & n9855 ) | ( n9777 & ~n9857 ) | ( n9855 & ~n9857 ) ;
  assign n9859 = ~n9777 & n9858 ;
  assign n9860 = ( n9233 & n9853 ) | ( n9233 & ~n9859 ) | ( n9853 & ~n9859 ) ;
  assign n9861 = ~n9233 & n9860 ;
  assign n9862 = n1205 | n9283 ;
  assign n9863 = n9783 & ~n9862 ;
  assign n9864 = n9855 & ~n9863 ;
  assign n9865 = ~n9300 & n9302 ;
  assign n9866 = x39 & ~n9865 ;
  assign n9867 = ( n1205 & n9772 ) | ( n1205 & ~n9866 ) | ( n9772 & ~n9866 ) ;
  assign n9868 = n9867 ^ n9772 ^ 1'b0 ;
  assign n9869 = ( n1205 & n9867 ) | ( n1205 & ~n9868 ) | ( n9867 & ~n9868 ) ;
  assign n9870 = ( x38 & n9847 ) | ( x38 & ~n9849 ) | ( n9847 & ~n9849 ) ;
  assign n9871 = ( x87 & n9869 ) | ( x87 & ~n9870 ) | ( n9869 & ~n9870 ) ;
  assign n9872 = n9871 ^ n9869 ^ 1'b0 ;
  assign n9873 = ( x87 & n9871 ) | ( x87 & ~n9872 ) | ( n9871 & ~n9872 ) ;
  assign n9874 = ( n9233 & n9864 ) | ( n9233 & n9873 ) | ( n9864 & n9873 ) ;
  assign n9875 = ~n9864 & n9874 ;
  assign n9876 = ( ~x75 & n9861 ) | ( ~x75 & n9875 ) | ( n9861 & n9875 ) ;
  assign n9877 = ~x75 & n9876 ;
  assign n9878 = ~n9233 & n9361 ;
  assign n9879 = x39 | n9813 ;
  assign n9880 = n9233 & n9283 ;
  assign n9881 = x75 & ~n9880 ;
  assign n9882 = ( n9878 & n9879 ) | ( n9878 & n9881 ) | ( n9879 & n9881 ) ;
  assign n9883 = ~n9878 & n9882 ;
  assign n9884 = ( n6782 & ~n9877 ) | ( n6782 & n9883 ) | ( ~n9877 & n9883 ) ;
  assign n9885 = n9877 | n9884 ;
  assign n9886 = n6782 & ~n9848 ;
  assign n9887 = ( n9742 & n9885 ) | ( n9742 & ~n9886 ) | ( n9885 & ~n9886 ) ;
  assign n9888 = ~n9742 & n9887 ;
  assign n9889 = n6782 & ~n9233 ;
  assign n9890 = n9776 & n9889 ;
  assign n9891 = ( n7318 & ~n9888 ) | ( n7318 & n9890 ) | ( ~n9888 & n9890 ) ;
  assign n9892 = n9888 | n9891 ;
  assign n9893 = ( ~n9746 & n9841 ) | ( ~n9746 & n9892 ) | ( n9841 & n9892 ) ;
  assign n9894 = ~n9746 & n9893 ;
  assign n9895 = x24 & ~n8757 ;
  assign n9896 = x53 & ~n1387 ;
  assign n9897 = ( n1388 & ~n1395 ) | ( n1388 & n9896 ) | ( ~n1395 & n9896 ) ;
  assign n9898 = ~n1388 & n9897 ;
  assign n9899 = n9895 & n9898 ;
  assign n9900 = x39 | n9899 ;
  assign n9901 = x38 | n8793 ;
  assign n9902 = x287 | x979 ;
  assign n9903 = n5066 & ~n9902 ;
  assign n9904 = x39 & ~n9903 ;
  assign n9905 = n9901 | n9904 ;
  assign n9906 = ( n2217 & n9900 ) | ( n2217 & ~n9905 ) | ( n9900 & ~n9905 ) ;
  assign n9907 = ~n2217 & n9906 ;
  assign n9908 = n7472 | n7592 ;
  assign n9909 = x60 | x85 ;
  assign n9910 = x106 & ~n9909 ;
  assign n9911 = n1244 | n7488 ;
  assign n9912 = ( n9611 & n9910 ) | ( n9611 & ~n9911 ) | ( n9910 & ~n9911 ) ;
  assign n9913 = ~n9611 & n9912 ;
  assign n9914 = n7504 | n9684 ;
  assign n9915 = ( n9687 & n9913 ) | ( n9687 & ~n9914 ) | ( n9913 & ~n9914 ) ;
  assign n9916 = ~n9687 & n9915 ;
  assign n9917 = ~n9908 & n9916 ;
  assign n9918 = x841 | n1374 ;
  assign n9919 = n7453 | n9918 ;
  assign n9920 = n1376 | n2056 ;
  assign n9921 = n9919 | n9920 ;
  assign n9922 = n9917 & ~n9921 ;
  assign n9923 = x54 | n9922 ;
  assign n9924 = ~n7448 & n9923 ;
  assign n9925 = ~n2054 & n8766 ;
  assign n9926 = n9925 ^ n9924 ^ 1'b0 ;
  assign n9927 = ( ~x54 & n9925 ) | ( ~x54 & n9926 ) | ( n9925 & n9926 ) ;
  assign n9928 = ( n9924 & ~n9926 ) | ( n9924 & n9927 ) | ( ~n9926 & n9927 ) ;
  assign n9929 = x45 & ~n1244 ;
  assign n9930 = ~n1230 & n9929 ;
  assign n9931 = ( n1241 & ~n9686 ) | ( n1241 & n9930 ) | ( ~n9686 & n9930 ) ;
  assign n9932 = ~n1241 & n9931 ;
  assign n9933 = n5203 | n7908 ;
  assign n9934 = n1229 | n2070 ;
  assign n9935 = n9933 | n9934 ;
  assign n9936 = n9932 & ~n9935 ;
  assign n9937 = x55 | n9936 ;
  assign n9938 = ~x54 & n9925 ;
  assign n9939 = ~x74 & n9938 ;
  assign n9940 = x55 & ~n9939 ;
  assign n9941 = ( n7446 & n9937 ) | ( n7446 & ~n9940 ) | ( n9937 & ~n9940 ) ;
  assign n9942 = ~n7446 & n9941 ;
  assign n9943 = x56 & ~x62 ;
  assign n9944 = x55 & ~n8663 ;
  assign n9945 = n9943 | n9944 ;
  assign n9946 = n1289 | n2099 ;
  assign n9947 = n5162 & ~n9946 ;
  assign n9948 = x56 & ~n9947 ;
  assign n9949 = ( n2120 & n9945 ) | ( n2120 & ~n9948 ) | ( n9945 & ~n9948 ) ;
  assign n9950 = ~n2120 & n9949 ;
  assign n9951 = n5283 | n9946 ;
  assign n9952 = ~x56 & x62 ;
  assign n9953 = x924 & n9952 ;
  assign n9954 = n9953 ^ n9952 ^ n9943 ;
  assign n9955 = n9954 ^ n9951 ^ 1'b0 ;
  assign n9956 = ( n9951 & n9954 ) | ( n9951 & n9955 ) | ( n9954 & n9955 ) ;
  assign n9957 = ( x57 & ~n9951 ) | ( x57 & n9956 ) | ( ~n9951 & n9956 ) ;
  assign n9958 = ~n5192 & n9939 ;
  assign n9959 = x57 & ~n9958 ;
  assign n9960 = ( x59 & n9957 ) | ( x59 & ~n9959 ) | ( n9957 & ~n9959 ) ;
  assign n9961 = ~x59 & n9960 ;
  assign n9962 = x93 | n9713 ;
  assign n9963 = n8760 | n9962 ;
  assign n9964 = n6375 & ~n9963 ;
  assign n9965 = ~n9951 & n9953 ;
  assign n9966 = x59 | n9965 ;
  assign n9967 = x59 & ~n9958 ;
  assign n9968 = ( x57 & n9966 ) | ( x57 & ~n9967 ) | ( n9966 & ~n9967 ) ;
  assign n9969 = ~x57 & n9968 ;
  assign n9970 = ~x39 & n9895 ;
  assign n9971 = n1385 & ~n9908 ;
  assign n9972 = n9970 & n9971 ;
  assign n9973 = x39 & ~x979 ;
  assign n9974 = ~n5066 & n9973 ;
  assign n9975 = ( ~n5067 & n5362 ) | ( ~n5067 & n9974 ) | ( n5362 & n9974 ) ;
  assign n9976 = ~n5362 & n9975 ;
  assign n9977 = ~n9901 & n9976 ;
  assign n9978 = ( ~n9901 & n9972 ) | ( ~n9901 & n9977 ) | ( n9972 & n9977 ) ;
  assign n9979 = ~x24 & n9971 ;
  assign n9980 = x841 & n9625 ;
  assign n9981 = ( ~n8761 & n9979 ) | ( ~n8761 & n9980 ) | ( n9979 & n9980 ) ;
  assign n9982 = ~n8761 & n9981 ;
  assign n9984 = ( x59 & n2120 ) | ( x59 & n8664 ) | ( n2120 & n8664 ) ;
  assign n9983 = n9947 & n9952 ;
  assign n9985 = ( x57 & n9983 ) | ( x57 & ~n9984 ) | ( n9983 & ~n9984 ) ;
  assign n9986 = ~n9984 & n9985 ;
  assign n9987 = n1478 & ~n7511 ;
  assign n9988 = ~n7589 & n9987 ;
  assign n9989 = x999 & n9988 ;
  assign n9990 = ~x24 & n9608 ;
  assign n9991 = ( ~n8761 & n9989 ) | ( ~n8761 & n9990 ) | ( n9989 & n9990 ) ;
  assign n9992 = ~n8761 & n9991 ;
  assign n9993 = ~x63 & x107 ;
  assign n9994 = ~n7589 & n9993 ;
  assign n9995 = x841 | n9994 ;
  assign n9996 = ~n1251 & n9993 ;
  assign n9997 = x64 | n9996 ;
  assign n9998 = ~n1229 & n9997 ;
  assign n9999 = n9998 ^ n8768 ^ 1'b0 ;
  assign n10000 = ( x841 & n8768 ) | ( x841 & ~n9998 ) | ( n8768 & ~n9998 ) ;
  assign n10001 = ( x841 & ~n9999 ) | ( x841 & n10000 ) | ( ~n9999 & n10000 ) ;
  assign n10002 = ( n9732 & n9995 ) | ( n9732 & ~n10001 ) | ( n9995 & ~n10001 ) ;
  assign n10003 = ~n9732 & n10002 ;
  assign n10004 = x39 & n8843 ;
  assign n10005 = ~n9901 & n10004 ;
  assign n10006 = ( n8861 & n8870 ) | ( n8861 & n10005 ) | ( n8870 & n10005 ) ;
  assign n10007 = ~n8861 & n10006 ;
  assign n10008 = x199 & ~x299 ;
  assign n10009 = ~n1206 & n10008 ;
  assign n10010 = x314 & ~n1228 ;
  assign n10011 = ~n9933 & n10010 ;
  assign n10012 = x81 & ~x102 ;
  assign n10013 = ( n1253 & n10011 ) | ( n1253 & n10012 ) | ( n10011 & n10012 ) ;
  assign n10014 = ~n1253 & n10013 ;
  assign n10015 = n1205 | n2068 ;
  assign n10016 = n10014 & ~n10015 ;
  assign n10017 = n10009 & n10016 ;
  assign n10018 = x219 | n10017 ;
  assign n10019 = x199 | x299 ;
  assign n10020 = ~n2070 & n10014 ;
  assign n10021 = n10019 & n10020 ;
  assign n10022 = x219 & ~n10021 ;
  assign n10023 = ( n7318 & n10018 ) | ( n7318 & ~n10022 ) | ( n10018 & ~n10022 ) ;
  assign n10024 = ~n7318 & n10023 ;
  assign n10025 = x83 & ~x103 ;
  assign n10026 = ( n8760 & ~n9733 ) | ( n8760 & n10025 ) | ( ~n9733 & n10025 ) ;
  assign n10027 = ~n8760 & n10026 ;
  assign n10028 = ( n1249 & n10011 ) | ( n1249 & n10027 ) | ( n10011 & n10027 ) ;
  assign n10029 = ~n1249 & n10028 ;
  assign n10030 = n5115 & n5379 ;
  assign n10031 = n2161 & ~n2290 ;
  assign n10032 = n10030 & n10031 ;
  assign n10033 = n5100 & n5379 ;
  assign n10034 = n2125 & n4736 ;
  assign n10035 = n10033 & n10034 ;
  assign n10036 = ( n9605 & n10032 ) | ( n9605 & n10035 ) | ( n10032 & n10035 ) ;
  assign n10037 = n10035 ^ n10032 ^ 1'b0 ;
  assign n10038 = ( n9605 & n10036 ) | ( n9605 & n10037 ) | ( n10036 & n10037 ) ;
  assign n10039 = x71 & x314 ;
  assign n10040 = ~n6379 & n10039 ;
  assign n10041 = ( n1250 & ~n8746 ) | ( n1250 & n10040 ) | ( ~n8746 & n10040 ) ;
  assign n10042 = ~n1250 & n10041 ;
  assign n10043 = x81 | x314 ;
  assign n10044 = ( n1229 & n5226 ) | ( n1229 & ~n10043 ) | ( n5226 & ~n10043 ) ;
  assign n10045 = n10043 | n10044 ;
  assign n10046 = x69 & ~n9683 ;
  assign n10047 = ~n8743 & n10046 ;
  assign n10048 = ( x71 & ~n10045 ) | ( x71 & n10047 ) | ( ~n10045 & n10047 ) ;
  assign n10049 = ~n10045 & n10048 ;
  assign n10050 = ( ~n9732 & n10042 ) | ( ~n9732 & n10049 ) | ( n10042 & n10049 ) ;
  assign n10051 = ~n9732 & n10050 ;
  assign n10052 = x210 & x589 ;
  assign n10053 = ~x221 & n4736 ;
  assign n10054 = ~x216 & n10053 ;
  assign n10055 = n5100 & n10054 ;
  assign n10056 = n10052 & n10055 ;
  assign n10057 = x198 & x589 ;
  assign n10058 = ~n2291 & n5115 ;
  assign n10059 = n10057 & n10058 ;
  assign n10060 = n10056 | n10059 ;
  assign n10061 = n10060 ^ x287 ^ 1'b0 ;
  assign n10062 = ~x593 & n5363 ;
  assign n10063 = n5369 & n10062 ;
  assign n10064 = ( n10060 & ~n10061 ) | ( n10060 & n10063 ) | ( ~n10061 & n10063 ) ;
  assign n10065 = ( x287 & n10061 ) | ( x287 & n10064 ) | ( n10061 & n10064 ) ;
  assign n10066 = x39 & ~n1292 ;
  assign n10067 = n10065 & n10066 ;
  assign n10068 = ~n1269 & n1436 ;
  assign n10069 = ~x96 & n10068 ;
  assign n10070 = n8765 & n10069 ;
  assign n10071 = ( ~n9901 & n10067 ) | ( ~n9901 & n10070 ) | ( n10067 & n10070 ) ;
  assign n10072 = ~n9901 & n10071 ;
  assign n10073 = ~x199 & x200 ;
  assign n10074 = ~x299 & n10073 ;
  assign n10075 = x211 & ~x219 ;
  assign n10076 = x299 & n10075 ;
  assign n10077 = n10074 | n10076 ;
  assign n10078 = n9630 | n10077 ;
  assign n10079 = n1234 | n1246 ;
  assign n10080 = n5210 & ~n10079 ;
  assign n10081 = ~n9639 & n10080 ;
  assign n10082 = ( n10011 & n10078 ) | ( n10011 & n10081 ) | ( n10078 & n10081 ) ;
  assign n10083 = ~n10078 & n10082 ;
  assign n10084 = x50 | n7511 ;
  assign n10085 = x314 & n10077 ;
  assign n10086 = x64 | n7500 ;
  assign n10087 = n10081 & ~n10086 ;
  assign n10088 = x81 | n10087 ;
  assign n10089 = ( n8757 & n10085 ) | ( n8757 & n10088 ) | ( n10085 & n10088 ) ;
  assign n10090 = ~n8757 & n10089 ;
  assign n10091 = ( n5209 & ~n10084 ) | ( n5209 & n10090 ) | ( ~n10084 & n10090 ) ;
  assign n10092 = ~n5209 & n10091 ;
  assign n10093 = ( ~n8760 & n10083 ) | ( ~n8760 & n10092 ) | ( n10083 & n10092 ) ;
  assign n10094 = ~n8760 & n10093 ;
  assign n10095 = x88 & ~n8742 ;
  assign n10096 = n5368 & ~n7786 ;
  assign n10097 = ( n1472 & n10095 ) | ( n1472 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10098 = ~n1472 & n10097 ;
  assign n10099 = x24 & ~n1379 ;
  assign n10100 = n10098 ^ x72 ^ 1'b0 ;
  assign n10101 = ( ~x72 & n10099 ) | ( ~x72 & n10100 ) | ( n10099 & n10100 ) ;
  assign n10102 = ( x72 & n10098 ) | ( x72 & n10101 ) | ( n10098 & n10101 ) ;
  assign n10103 = n10102 ^ n5203 ^ 1'b0 ;
  assign n10104 = ( n5203 & n10102 ) | ( n5203 & n10103 ) | ( n10102 & n10103 ) ;
  assign n10105 = ( x39 & ~n5203 ) | ( x39 & n10104 ) | ( ~n5203 & n10104 ) ;
  assign n10106 = n6463 & n10030 ;
  assign n10107 = n6466 & n10033 ;
  assign n10108 = ( x39 & n10106 ) | ( x39 & ~n10107 ) | ( n10106 & ~n10107 ) ;
  assign n10109 = ~n10106 & n10108 ;
  assign n10110 = ( n9901 & n10105 ) | ( n9901 & ~n10109 ) | ( n10105 & ~n10109 ) ;
  assign n10111 = ~n9901 & n10110 ;
  assign n10112 = n7678 & n10030 ;
  assign n10113 = ~x299 & n10112 ;
  assign n10114 = n7669 & n10033 ;
  assign n10115 = x299 & ~n10114 ;
  assign n10116 = ( n6263 & n10113 ) | ( n6263 & ~n10115 ) | ( n10113 & ~n10115 ) ;
  assign n10117 = x39 & ~n10116 ;
  assign n10118 = ~x314 & x1050 ;
  assign n10119 = n8132 & ~n8757 ;
  assign n10120 = n10118 & n10119 ;
  assign n10121 = x39 | n10120 ;
  assign n10122 = ( n9901 & ~n10117 ) | ( n9901 & n10121 ) | ( ~n10117 & n10121 ) ;
  assign n10123 = ~n9901 & n10122 ;
  assign n10124 = ~n1414 & n6432 ;
  assign n10125 = x96 | n10124 ;
  assign n10126 = x96 | n5165 ;
  assign n10127 = x479 & n10126 ;
  assign n10128 = n2177 | n6782 ;
  assign n10129 = ( x1093 & n9011 ) | ( x1093 & ~n10128 ) | ( n9011 & ~n10128 ) ;
  assign n10130 = ( n6425 & n10128 ) | ( n6425 & ~n10129 ) | ( n10128 & ~n10129 ) ;
  assign n10131 = ( n7451 & ~n10127 ) | ( n7451 & n10130 ) | ( ~n10127 & n10130 ) ;
  assign n10132 = n10127 | n10131 ;
  assign n10133 = ( n6394 & n10125 ) | ( n6394 & ~n10132 ) | ( n10125 & ~n10132 ) ;
  assign n10134 = ~n6394 & n10133 ;
  assign n10135 = x74 & n9938 ;
  assign n10136 = ( ~n7318 & n10134 ) | ( ~n7318 & n10135 ) | ( n10134 & n10135 ) ;
  assign n10137 = ~n7318 & n10136 ;
  assign n10138 = n5015 | n7448 ;
  assign n10139 = n6443 ^ x75 ^ 1'b0 ;
  assign n10140 = ~n1614 & n8670 ;
  assign n10141 = n10125 & n10140 ;
  assign n10142 = ( ~n1207 & n9011 ) | ( ~n1207 & n10141 ) | ( n9011 & n10141 ) ;
  assign n10143 = ~n1207 & n10142 ;
  assign n10144 = ( n6443 & ~n10139 ) | ( n6443 & n10143 ) | ( ~n10139 & n10143 ) ;
  assign n10145 = ( x75 & n10139 ) | ( x75 & n10144 ) | ( n10139 & n10144 ) ;
  assign n10146 = ~n2052 & n8766 ;
  assign n10147 = x75 & ~n10146 ;
  assign n10148 = ( n10138 & n10145 ) | ( n10138 & ~n10147 ) | ( n10145 & ~n10147 ) ;
  assign n10149 = ~n10138 & n10148 ;
  assign n10150 = n1328 | n8898 ;
  assign n10151 = ~x137 & n1615 ;
  assign n10152 = x94 | n7507 ;
  assign n10153 = n7472 & ~n8981 ;
  assign n10154 = ( n8757 & n10152 ) | ( n8757 & ~n10153 ) | ( n10152 & ~n10153 ) ;
  assign n10155 = ~n8757 & n10154 ;
  assign n10156 = n6442 | n10155 ;
  assign n10157 = n7506 & ~n9651 ;
  assign n10158 = x252 & n10157 ;
  assign n10159 = ~x252 & n10155 ;
  assign n10160 = ( n6442 & n10158 ) | ( n6442 & ~n10159 ) | ( n10158 & ~n10159 ) ;
  assign n10161 = ~n10158 & n10160 ;
  assign n10162 = n10156 & ~n10161 ;
  assign n10163 = n10162 ^ x122 ^ 1'b0 ;
  assign n10164 = ~n1290 & n8982 ;
  assign n10165 = x252 & n6442 ;
  assign n10166 = n10164 & ~n10165 ;
  assign n10167 = ( n10162 & ~n10163 ) | ( n10162 & n10166 ) | ( ~n10163 & n10166 ) ;
  assign n10174 = x122 & ~n10162 ;
  assign n10168 = n6425 & ~n10156 ;
  assign n10169 = n5022 | n10164 ;
  assign n10170 = ~n10161 & n10169 ;
  assign n10171 = n10170 ^ n10168 ^ 1'b0 ;
  assign n10172 = ( n10168 & n10170 ) | ( n10168 & n10171 ) | ( n10170 & n10171 ) ;
  assign n10173 = ( x122 & ~n10168 ) | ( x122 & n10172 ) | ( ~n10168 & n10172 ) ;
  assign n10175 = n10174 ^ n10173 ^ 1'b0 ;
  assign n10176 = n10175 ^ x1093 ^ 1'b0 ;
  assign n10177 = ( n10167 & n10175 ) | ( n10167 & n10176 ) | ( n10175 & n10176 ) ;
  assign n10178 = ( x1091 & n1614 ) | ( x1091 & ~n10177 ) | ( n1614 & ~n10177 ) ;
  assign n10179 = ~n1614 & n10178 ;
  assign n10180 = n10151 | n10179 ;
  assign n10181 = ~x137 & n10166 ;
  assign n10182 = n10180 & ~n10181 ;
  assign n10183 = x252 & x1092 ;
  assign n10184 = ~x1093 & n10183 ;
  assign n10185 = n1610 & n10184 ;
  assign n10186 = ( x137 & n10164 ) | ( x137 & ~n10185 ) | ( n10164 & ~n10185 ) ;
  assign n10187 = ~x137 & n10186 ;
  assign n10188 = ( x1093 & n10173 ) | ( x1093 & ~n10174 ) | ( n10173 & ~n10174 ) ;
  assign n10189 = ~x122 & n10164 ;
  assign n10190 = x1093 & ~n10155 ;
  assign n10191 = n6783 | n10190 ;
  assign n10192 = n10188 & ~n10191 ;
  assign n10193 = ( n10188 & n10189 ) | ( n10188 & n10192 ) | ( n10189 & n10192 ) ;
  assign n10194 = n1614 & ~n10193 ;
  assign n10195 = ( x1091 & n10193 ) | ( x1091 & ~n10194 ) | ( n10193 & ~n10194 ) ;
  assign n10196 = x137 | n1615 ;
  assign n10197 = n10195 & n10196 ;
  assign n10198 = ( ~n10182 & n10187 ) | ( ~n10182 & n10197 ) | ( n10187 & n10197 ) ;
  assign n10199 = ~n10182 & n10198 ;
  assign n10200 = ~n10179 & n10195 ;
  assign n10201 = n10199 ^ x210 ^ 1'b0 ;
  assign n10202 = ( n10199 & n10200 ) | ( n10199 & n10201 ) | ( n10200 & n10201 ) ;
  assign n10203 = ( x299 & n10150 ) | ( x299 & n10202 ) | ( n10150 & n10202 ) ;
  assign n10204 = n10202 ^ n10150 ^ 1'b0 ;
  assign n10205 = ( x299 & n10203 ) | ( x299 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10206 = ~x137 & n5035 ;
  assign n10207 = n8686 & n10157 ;
  assign n10208 = n10207 ^ n5035 ^ 1'b0 ;
  assign n10209 = ( n5035 & n10206 ) | ( n5035 & n10208 ) | ( n10206 & n10208 ) ;
  assign n10210 = ( n5035 & n10199 ) | ( n5035 & ~n10209 ) | ( n10199 & ~n10209 ) ;
  assign n10211 = ~n10209 & n10210 ;
  assign n10212 = ( n10200 & n10207 ) | ( n10200 & ~n10208 ) | ( n10207 & ~n10208 ) ;
  assign n10213 = n10211 ^ x210 ^ 1'b0 ;
  assign n10214 = ( n10211 & n10212 ) | ( n10211 & n10213 ) | ( n10212 & n10213 ) ;
  assign n10215 = n10214 ^ n10205 ^ 1'b0 ;
  assign n10216 = ( ~n10150 & n10214 ) | ( ~n10150 & n10215 ) | ( n10214 & n10215 ) ;
  assign n10217 = ( n10205 & ~n10215 ) | ( n10205 & n10216 ) | ( ~n10215 & n10216 ) ;
  assign n10218 = n1283 | n5075 ;
  assign n10219 = n10199 ^ x198 ^ 1'b0 ;
  assign n10220 = ( n10199 & n10200 ) | ( n10199 & n10219 ) | ( n10200 & n10219 ) ;
  assign n10221 = ( ~x299 & n10218 ) | ( ~x299 & n10220 ) | ( n10218 & n10220 ) ;
  assign n10222 = ~x299 & n10221 ;
  assign n10223 = n10211 ^ x198 ^ 1'b0 ;
  assign n10224 = ( n10211 & n10212 ) | ( n10211 & n10223 ) | ( n10212 & n10223 ) ;
  assign n10225 = n10224 ^ n10222 ^ 1'b0 ;
  assign n10226 = ( ~n10218 & n10224 ) | ( ~n10218 & n10225 ) | ( n10224 & n10225 ) ;
  assign n10227 = ( n10222 & ~n10225 ) | ( n10222 & n10226 ) | ( ~n10225 & n10226 ) ;
  assign n10228 = ( x232 & n10217 ) | ( x232 & n10227 ) | ( n10217 & n10227 ) ;
  assign n10229 = n10227 ^ n10217 ^ 1'b0 ;
  assign n10230 = ( x232 & n10228 ) | ( x232 & n10229 ) | ( n10228 & n10229 ) ;
  assign n10231 = x299 | n10224 ;
  assign n10232 = x299 & ~n10214 ;
  assign n10233 = ( x232 & n10231 ) | ( x232 & ~n10232 ) | ( n10231 & ~n10232 ) ;
  assign n10234 = ~x232 & n10233 ;
  assign n10235 = ( ~n6612 & n10230 ) | ( ~n6612 & n10234 ) | ( n10230 & n10234 ) ;
  assign n10236 = ~n6612 & n10235 ;
  assign n10237 = n5035 & n10157 ;
  assign n10238 = ~n8685 & n10237 ;
  assign n10239 = n6442 ^ x252 ^ 1'b0 ;
  assign n10240 = ( ~x252 & n10155 ) | ( ~x252 & n10239 ) | ( n10155 & n10239 ) ;
  assign n10241 = n10240 ^ n10164 ^ 1'b0 ;
  assign n10242 = ( ~n6442 & n10164 ) | ( ~n6442 & n10241 ) | ( n10164 & n10241 ) ;
  assign n10243 = ( n10240 & ~n10241 ) | ( n10240 & n10242 ) | ( ~n10241 & n10242 ) ;
  assign n10244 = n6783 & ~n10243 ;
  assign n10245 = n10174 | n10244 ;
  assign n10246 = n1615 & n10245 ;
  assign n10247 = x1093 | n10162 ;
  assign n10248 = ~n1615 & n10190 ;
  assign n10249 = ( n10246 & n10247 ) | ( n10246 & ~n10248 ) | ( n10247 & ~n10248 ) ;
  assign n10250 = ~n10246 & n10249 ;
  assign n10251 = ~n5035 & n10250 ;
  assign n10252 = n10238 | n10251 ;
  assign n10253 = x137 & ~n10247 ;
  assign n10254 = n10190 | n10253 ;
  assign n10255 = x137 | n10243 ;
  assign n10256 = x1093 | n10255 ;
  assign n10257 = ~n10254 & n10256 ;
  assign n10258 = ~n5035 & n10257 ;
  assign n10259 = n10237 | n10258 ;
  assign n10260 = x137 & ~n6783 ;
  assign n10261 = n6442 & ~n10260 ;
  assign n10262 = n10157 & ~n10261 ;
  assign n10263 = n1615 & ~n5035 ;
  assign n10264 = ( n1615 & n10262 ) | ( n1615 & n10263 ) | ( n10262 & n10263 ) ;
  assign n10265 = ~n10253 & n10255 ;
  assign n10266 = x137 & n10245 ;
  assign n10267 = n10265 & ~n10266 ;
  assign n10268 = n10267 ^ n5035 ^ 1'b0 ;
  assign n10269 = ( n5035 & n10267 ) | ( n5035 & ~n10268 ) | ( n10267 & ~n10268 ) ;
  assign n10270 = ( n10264 & n10268 ) | ( n10264 & n10269 ) | ( n10268 & n10269 ) ;
  assign n10271 = n7450 & n10206 ;
  assign n10272 = n1615 | n10271 ;
  assign n10273 = ~n10270 & n10272 ;
  assign n10274 = ( n10259 & n10270 ) | ( n10259 & ~n10273 ) | ( n10270 & ~n10273 ) ;
  assign n10275 = n10252 ^ x198 ^ 1'b0 ;
  assign n10276 = ( n10252 & n10274 ) | ( n10252 & ~n10275 ) | ( n10274 & ~n10275 ) ;
  assign n10277 = ~x299 & n10276 ;
  assign n10278 = n10252 ^ x210 ^ 1'b0 ;
  assign n10279 = ( n10252 & n10274 ) | ( n10252 & ~n10278 ) | ( n10274 & ~n10278 ) ;
  assign n10280 = x299 & n10279 ;
  assign n10281 = ( x232 & ~n10277 ) | ( x232 & n10280 ) | ( ~n10277 & n10280 ) ;
  assign n10282 = n10277 | n10281 ;
  assign n10294 = x210 & ~n10250 ;
  assign n10295 = n10150 | n10294 ;
  assign n10283 = n10257 ^ n1615 ^ 1'b0 ;
  assign n10284 = ( n10257 & n10267 ) | ( n10257 & n10283 ) | ( n10267 & n10283 ) ;
  assign n10293 = x210 | n10284 ;
  assign n10296 = n10295 ^ n10293 ^ 1'b0 ;
  assign n10297 = ( x299 & ~n10293 ) | ( x299 & n10295 ) | ( ~n10293 & n10295 ) ;
  assign n10298 = ( x299 & ~n10296 ) | ( x299 & n10297 ) | ( ~n10296 & n10297 ) ;
  assign n10299 = ( n10150 & n10279 ) | ( n10150 & ~n10298 ) | ( n10279 & ~n10298 ) ;
  assign n10300 = n10299 ^ n10298 ^ 1'b0 ;
  assign n10301 = ( n10298 & ~n10299 ) | ( n10298 & n10300 ) | ( ~n10299 & n10300 ) ;
  assign n10285 = n10250 ^ x198 ^ 1'b0 ;
  assign n10286 = ( n10250 & n10284 ) | ( n10250 & ~n10285 ) | ( n10284 & ~n10285 ) ;
  assign n10287 = n10286 ^ n10218 ^ 1'b0 ;
  assign n10288 = ( n10218 & n10286 ) | ( n10218 & n10287 ) | ( n10286 & n10287 ) ;
  assign n10289 = ( x299 & ~n10218 ) | ( x299 & n10288 ) | ( ~n10218 & n10288 ) ;
  assign n10290 = n10289 ^ n10218 ^ 1'b0 ;
  assign n10291 = ( ~n10218 & n10276 ) | ( ~n10218 & n10290 ) | ( n10276 & n10290 ) ;
  assign n10292 = ( n10218 & n10289 ) | ( n10218 & n10291 ) | ( n10289 & n10291 ) ;
  assign n10302 = n10301 ^ n10292 ^ 1'b0 ;
  assign n10303 = ( x232 & ~n10292 ) | ( x232 & n10301 ) | ( ~n10292 & n10301 ) ;
  assign n10304 = ( x232 & ~n10302 ) | ( x232 & n10303 ) | ( ~n10302 & n10303 ) ;
  assign n10305 = n6612 & ~n10304 ;
  assign n10306 = n10282 & n10305 ;
  assign n10307 = ( ~n8760 & n10236 ) | ( ~n8760 & n10306 ) | ( n10236 & n10306 ) ;
  assign n10308 = ~n8760 & n10307 ;
  assign n10309 = x86 & ~n7472 ;
  assign n10310 = ~n1464 & n10309 ;
  assign n10311 = x314 & ~n10310 ;
  assign n10312 = n8761 | n10311 ;
  assign n10313 = n1564 | n5207 ;
  assign n10314 = ~n1456 & n1470 ;
  assign n10315 = x86 | n10314 ;
  assign n10316 = ~n10313 & n10315 ;
  assign n10317 = ~n1372 & n10316 ;
  assign n10318 = ( x314 & ~n10312 ) | ( x314 & n10317 ) | ( ~n10312 & n10317 ) ;
  assign n10319 = ~n10312 & n10318 ;
  assign n10320 = x119 & x232 ;
  assign n10321 = ~x468 & n10320 ;
  assign n10322 = x34 | n8653 ;
  assign n10323 = x163 & ~n5075 ;
  assign n10324 = n10323 ^ n8276 ^ n5075 ;
  assign n10325 = x232 & n10324 ;
  assign n10326 = x75 & ~n10325 ;
  assign n10327 = x100 & ~n10325 ;
  assign n10328 = n10326 | n10327 ;
  assign n10329 = x147 & n6411 ;
  assign n10330 = ~n7555 & n10329 ;
  assign n10331 = n10328 | n10330 ;
  assign n10332 = n7555 & n10325 ;
  assign n10333 = x74 & ~n10332 ;
  assign n10334 = n2120 & ~n10333 ;
  assign n10335 = ~n10331 & n10334 ;
  assign n10336 = n10331 ^ x54 ^ 1'b0 ;
  assign n10337 = x38 | x40 ;
  assign n10338 = x38 & ~n10329 ;
  assign n10339 = x100 | n10338 ;
  assign n10340 = n10337 & ~n10339 ;
  assign n10341 = n10327 | n10340 ;
  assign n10342 = ~x75 & n10341 ;
  assign n10343 = n10326 | n10342 ;
  assign n10344 = ( n10331 & ~n10336 ) | ( n10331 & n10343 ) | ( ~n10336 & n10343 ) ;
  assign n10345 = x74 | n10344 ;
  assign n10346 = ( ~x74 & n10333 ) | ( ~x74 & n10345 ) | ( n10333 & n10345 ) ;
  assign n10347 = ( n2109 & ~n7546 ) | ( n2109 & n10346 ) | ( ~n7546 & n10346 ) ;
  assign n10348 = ( n2120 & n7546 ) | ( n2120 & n10347 ) | ( n7546 & n10347 ) ;
  assign n10349 = x54 & n10331 ;
  assign n10350 = n1273 | n8098 ;
  assign n10351 = x163 & x232 ;
  assign n10352 = x92 | n1206 ;
  assign n10353 = n10351 & ~n10352 ;
  assign n10354 = n10353 ^ n10350 ^ 1'b0 ;
  assign n10355 = ( n10350 & n10353 ) | ( n10350 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10356 = ( n10337 & ~n10350 ) | ( n10337 & n10355 ) | ( ~n10350 & n10355 ) ;
  assign n10357 = ( x75 & ~n10339 ) | ( x75 & n10356 ) | ( ~n10339 & n10356 ) ;
  assign n10358 = ~x75 & n10357 ;
  assign n10359 = ( ~x54 & n10328 ) | ( ~x54 & n10358 ) | ( n10328 & n10358 ) ;
  assign n10360 = ~x54 & n10359 ;
  assign n10361 = ( ~x74 & n10349 ) | ( ~x74 & n10360 ) | ( n10349 & n10360 ) ;
  assign n10362 = ~x74 & n10361 ;
  assign n10363 = ( x55 & n10333 ) | ( x55 & ~n10362 ) | ( n10333 & ~n10362 ) ;
  assign n10364 = ~n10333 & n10363 ;
  assign n10365 = x299 ^ x147 ^ 1'b0 ;
  assign n10366 = ( x147 & x187 ) | ( x147 & ~n10365 ) | ( x187 & ~n10365 ) ;
  assign n10367 = n6411 & n10366 ;
  assign n10368 = n7555 | n10367 ;
  assign n10369 = n8304 & n8305 ;
  assign n10370 = ~x184 & n10369 ;
  assign n10371 = x184 & ~n5075 ;
  assign n10372 = ~n10369 & n10371 ;
  assign n10373 = ( x299 & ~n10370 ) | ( x299 & n10372 ) | ( ~n10370 & n10372 ) ;
  assign n10374 = n10370 | n10373 ;
  assign n10375 = x299 & ~n10324 ;
  assign n10376 = x232 & ~n10375 ;
  assign n10377 = n10374 & n10376 ;
  assign n10378 = n7555 & n10377 ;
  assign n10379 = x54 & ~n10378 ;
  assign n10380 = n10368 & n10379 ;
  assign n10381 = ~x147 & x187 ;
  assign n10382 = n7656 & n10381 ;
  assign n10383 = x187 & ~n7659 ;
  assign n10384 = x187 | n7662 ;
  assign n10385 = ( x147 & n10383 ) | ( x147 & n10384 ) | ( n10383 & n10384 ) ;
  assign n10386 = ~n10383 & n10385 ;
  assign n10387 = ( x38 & n10382 ) | ( x38 & n10386 ) | ( n10382 & n10386 ) ;
  assign n10388 = n10386 ^ n10382 ^ 1'b0 ;
  assign n10389 = ( x38 & n10387 ) | ( x38 & n10388 ) | ( n10387 & n10388 ) ;
  assign n10390 = x40 | x232 ;
  assign n10391 = x153 & ~n8098 ;
  assign n10392 = n8105 & n10391 ;
  assign n10393 = x40 | x163 ;
  assign n10394 = n8147 & ~n8898 ;
  assign n10395 = ( ~n10392 & n10393 ) | ( ~n10392 & n10394 ) | ( n10393 & n10394 ) ;
  assign n10396 = n10392 | n10395 ;
  assign n10397 = ~x32 & x95 ;
  assign n10398 = ~x479 & n10397 ;
  assign n10399 = ~n1273 & n10398 ;
  assign n10400 = ~n5075 & n10399 ;
  assign n10401 = n10396 | n10400 ;
  assign n10402 = ~x210 & n8127 ;
  assign n10403 = n8129 | n10402 ;
  assign n10404 = ( x153 & n8163 ) | ( x153 & n10403 ) | ( n8163 & n10403 ) ;
  assign n10405 = ~n8898 & n10404 ;
  assign n10406 = ~x40 & x163 ;
  assign n10407 = x166 & ~n5075 ;
  assign n10408 = x153 & n8117 ;
  assign n10409 = ( n8157 & n10407 ) | ( n8157 & n10408 ) | ( n10407 & n10408 ) ;
  assign n10410 = n10407 & n10409 ;
  assign n10411 = ( n10405 & n10406 ) | ( n10405 & ~n10410 ) | ( n10406 & ~n10410 ) ;
  assign n10412 = ~n10405 & n10411 ;
  assign n10413 = ( x160 & n10396 ) | ( x160 & ~n10412 ) | ( n10396 & ~n10412 ) ;
  assign n10414 = ~x160 & n10413 ;
  assign n10415 = x40 | n10399 ;
  assign n10416 = n8129 | n10415 ;
  assign n10417 = n10402 | n10416 ;
  assign n10418 = ~n8898 & n10417 ;
  assign n10419 = n8157 | n10415 ;
  assign n10420 = n10407 & n10419 ;
  assign n10421 = ( n8117 & n10407 ) | ( n8117 & n10420 ) | ( n10407 & n10420 ) ;
  assign n10422 = ( x153 & n10418 ) | ( x153 & ~n10421 ) | ( n10418 & ~n10421 ) ;
  assign n10423 = ~n10418 & n10422 ;
  assign n10424 = n8163 | n10415 ;
  assign n10425 = ~n8898 & n10424 ;
  assign n10426 = x153 | n10420 ;
  assign n10427 = ( ~n10423 & n10425 ) | ( ~n10423 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10428 = ~n10423 & n10427 ;
  assign n10429 = x40 & n5075 ;
  assign n10430 = ( x163 & n10428 ) | ( x163 & ~n10429 ) | ( n10428 & ~n10429 ) ;
  assign n10431 = ~n10428 & n10430 ;
  assign n10432 = ~n10414 & n10431 ;
  assign n10433 = ( x160 & n10414 ) | ( x160 & ~n10432 ) | ( n10414 & ~n10432 ) ;
  assign n10434 = ( ~x299 & n10401 ) | ( ~x299 & n10433 ) | ( n10401 & n10433 ) ;
  assign n10435 = x299 & n10434 ;
  assign n10436 = x175 | x299 ;
  assign n10437 = x184 | n8147 ;
  assign n10438 = x184 & ~n8143 ;
  assign n10439 = ( x189 & n10437 ) | ( x189 & ~n10438 ) | ( n10437 & ~n10438 ) ;
  assign n10440 = ~x189 & n10439 ;
  assign n10441 = x182 & n10399 ;
  assign n10442 = x184 & x189 ;
  assign n10443 = n8140 & n10442 ;
  assign n10444 = n10441 | n10443 ;
  assign n10445 = ( ~n5075 & n10440 ) | ( ~n5075 & n10444 ) | ( n10440 & n10444 ) ;
  assign n10446 = ~n5075 & n10445 ;
  assign n10447 = x40 | n10446 ;
  assign n10448 = ~n10436 & n10447 ;
  assign n10454 = n8130 & ~n8905 ;
  assign n10455 = ( ~n8905 & n10415 ) | ( ~n8905 & n10454 ) | ( n10415 & n10454 ) ;
  assign n10449 = x189 & ~n5075 ;
  assign n10450 = n8118 | n10415 ;
  assign n10451 = n10449 & n10450 ;
  assign n10452 = x182 & x184 ;
  assign n10453 = ~n10429 & n10452 ;
  assign n10456 = ( ~n10451 & n10453 ) | ( ~n10451 & n10455 ) | ( n10453 & n10455 ) ;
  assign n10457 = ~n10455 & n10456 ;
  assign n10458 = ( x175 & x299 ) | ( x175 & ~n10457 ) | ( x299 & ~n10457 ) ;
  assign n10459 = ~x299 & n10458 ;
  assign n10460 = n10459 ^ n10448 ^ 1'b0 ;
  assign n10461 = x189 & n8119 ;
  assign n10462 = ~x182 & x184 ;
  assign n10463 = ( n10454 & ~n10461 ) | ( n10454 & n10462 ) | ( ~n10461 & n10462 ) ;
  assign n10464 = ~n10454 & n10463 ;
  assign n10465 = x189 & ~n8105 ;
  assign n10466 = n1289 | n10465 ;
  assign n10467 = x189 | n8133 ;
  assign n10468 = n10467 ^ n10466 ^ 1'b0 ;
  assign n10469 = ( n10466 & n10467 ) | ( n10466 & n10468 ) | ( n10467 & n10468 ) ;
  assign n10470 = ( n10441 & ~n10466 ) | ( n10441 & n10469 ) | ( ~n10466 & n10469 ) ;
  assign n10471 = n10470 ^ n5075 ^ 1'b0 ;
  assign n10472 = ( n5075 & n10470 ) | ( n5075 & n10471 ) | ( n10470 & n10471 ) ;
  assign n10473 = ( x184 & ~n5075 ) | ( x184 & n10472 ) | ( ~n5075 & n10472 ) ;
  assign n10474 = n10473 ^ n10464 ^ 1'b0 ;
  assign n10475 = ( n10464 & n10473 ) | ( n10464 & n10474 ) | ( n10473 & n10474 ) ;
  assign n10476 = ( x40 & ~n10464 ) | ( x40 & n10475 ) | ( ~n10464 & n10475 ) ;
  assign n10477 = ( n10459 & ~n10460 ) | ( n10459 & n10476 ) | ( ~n10460 & n10476 ) ;
  assign n10478 = ( n10448 & n10460 ) | ( n10448 & n10477 ) | ( n10460 & n10477 ) ;
  assign n10479 = ( ~x39 & n10435 ) | ( ~x39 & n10478 ) | ( n10435 & n10478 ) ;
  assign n10480 = ~x39 & n10479 ;
  assign n10481 = ~x166 & n7673 ;
  assign n10482 = x156 & n5096 ;
  assign n10483 = n10481 | n10482 ;
  assign n10484 = ( ~n5061 & n7669 ) | ( ~n5061 & n10483 ) | ( n7669 & n10483 ) ;
  assign n10485 = n5061 & n10484 ;
  assign n10486 = ( n1273 & ~n8098 ) | ( n1273 & n10485 ) | ( ~n8098 & n10485 ) ;
  assign n10487 = ~n1273 & n10486 ;
  assign n10488 = ( x40 & x299 ) | ( x40 & ~n10487 ) | ( x299 & ~n10487 ) ;
  assign n10489 = ~x40 & n10488 ;
  assign n10490 = ~x189 & n7673 ;
  assign n10491 = x179 & n5096 ;
  assign n10492 = n10490 | n10491 ;
  assign n10493 = ( ~n5114 & n7678 ) | ( ~n5114 & n10492 ) | ( n7678 & n10492 ) ;
  assign n10494 = n5114 & n10493 ;
  assign n10495 = ( n1273 & ~n8098 ) | ( n1273 & n10494 ) | ( ~n8098 & n10494 ) ;
  assign n10496 = ~n1273 & n10495 ;
  assign n10497 = ( x40 & x299 ) | ( x40 & ~n10496 ) | ( x299 & ~n10496 ) ;
  assign n10498 = n10496 | n10497 ;
  assign n10499 = ( x39 & n10489 ) | ( x39 & n10498 ) | ( n10489 & n10498 ) ;
  assign n10500 = ~n10489 & n10499 ;
  assign n10501 = ( x232 & n10480 ) | ( x232 & ~n10500 ) | ( n10480 & ~n10500 ) ;
  assign n10502 = ~n10480 & n10501 ;
  assign n10503 = ( x38 & n10390 ) | ( x38 & ~n10502 ) | ( n10390 & ~n10502 ) ;
  assign n10504 = ~x38 & n10503 ;
  assign n10505 = ( ~n2051 & n10389 ) | ( ~n2051 & n10504 ) | ( n10389 & n10504 ) ;
  assign n10506 = ~n2051 & n10505 ;
  assign n10507 = x100 & ~n10377 ;
  assign n10508 = x38 & ~n10367 ;
  assign n10509 = x100 | n10508 ;
  assign n10510 = x87 & n10337 ;
  assign n10511 = ~n10509 & n10510 ;
  assign n10512 = n10507 | n10511 ;
  assign n10513 = ( ~n2053 & n10506 ) | ( ~n2053 & n10512 ) | ( n10506 & n10512 ) ;
  assign n10514 = ~n2053 & n10513 ;
  assign n10515 = x299 ^ x156 ^ 1'b0 ;
  assign n10516 = ( x156 & x179 ) | ( x156 & ~n10515 ) | ( x179 & ~n10515 ) ;
  assign n10517 = n6411 & n10516 ;
  assign n10518 = n1206 | n1289 ;
  assign n10519 = ( n1273 & n10517 ) | ( n1273 & ~n10518 ) | ( n10517 & ~n10518 ) ;
  assign n10520 = ~n1273 & n10519 ;
  assign n10521 = ( n10337 & ~n10509 ) | ( n10337 & n10520 ) | ( ~n10509 & n10520 ) ;
  assign n10522 = ~n10509 & n10521 ;
  assign n10523 = ( n7639 & n10507 ) | ( n7639 & n10522 ) | ( n10507 & n10522 ) ;
  assign n10524 = n10522 ^ n10507 ^ 1'b0 ;
  assign n10525 = ( n7639 & n10523 ) | ( n7639 & n10524 ) | ( n10523 & n10524 ) ;
  assign n10526 = n10377 & ~n10525 ;
  assign n10527 = ( x75 & n10525 ) | ( x75 & ~n10526 ) | ( n10525 & ~n10526 ) ;
  assign n10528 = ( ~x54 & n10514 ) | ( ~x54 & n10527 ) | ( n10514 & n10527 ) ;
  assign n10529 = ~x54 & n10528 ;
  assign n10530 = ( ~x74 & n10380 ) | ( ~x74 & n10529 ) | ( n10380 & n10529 ) ;
  assign n10531 = ~x74 & n10530 ;
  assign n10532 = x74 & ~n10378 ;
  assign n10533 = ( x55 & ~n10531 ) | ( x55 & n10532 ) | ( ~n10531 & n10532 ) ;
  assign n10534 = n10531 | n10533 ;
  assign n10535 = ( n2109 & ~n10364 ) | ( n2109 & n10534 ) | ( ~n10364 & n10534 ) ;
  assign n10536 = ~n2109 & n10535 ;
  assign n10537 = ( ~n10335 & n10348 ) | ( ~n10335 & n10536 ) | ( n10348 & n10536 ) ;
  assign n10538 = ~n10335 & n10537 ;
  assign n10539 = x79 & n10538 ;
  assign n10540 = n10322 & ~n10539 ;
  assign n10541 = ~x79 & n8261 ;
  assign n10542 = n10538 & n10541 ;
  assign n10543 = n10322 | n10542 ;
  assign n10544 = ~n7678 & n7812 ;
  assign n10547 = n1230 | n7681 ;
  assign n10548 = ~n7853 & n10547 ;
  assign n10549 = ( x40 & n7598 ) | ( x40 & ~n7812 ) | ( n7598 & ~n7812 ) ;
  assign n10550 = ( n7674 & n7812 ) | ( n7674 & ~n10549 ) | ( n7812 & ~n10549 ) ;
  assign n10551 = n5099 & n10550 ;
  assign n10552 = n5083 & n7812 ;
  assign n10553 = n10551 | n10552 ;
  assign n10554 = n10548 | n10553 ;
  assign n10555 = x189 & n5114 ;
  assign n10556 = ~n10554 & n10555 ;
  assign n10545 = ~x40 & n7677 ;
  assign n10546 = x189 | n10545 ;
  assign n10557 = n10556 ^ n10546 ^ 1'b0 ;
  assign n10558 = ( x179 & ~n10546 ) | ( x179 & n10556 ) | ( ~n10546 & n10556 ) ;
  assign n10559 = ( x179 & ~n10557 ) | ( x179 & n10558 ) | ( ~n10557 & n10558 ) ;
  assign n10560 = n1230 | n7697 ;
  assign n10561 = n7853 | n10560 ;
  assign n10562 = ( ~n7853 & n10553 ) | ( ~n7853 & n10561 ) | ( n10553 & n10561 ) ;
  assign n10563 = ~x189 & n10562 ;
  assign n10564 = ~x179 & n5114 ;
  assign n10565 = n7812 ^ n5083 ^ 1'b0 ;
  assign n10566 = ( n7812 & n10550 ) | ( n7812 & ~n10565 ) | ( n10550 & ~n10565 ) ;
  assign n10567 = x189 & n10566 ;
  assign n10568 = ( n10563 & n10564 ) | ( n10563 & ~n10567 ) | ( n10564 & ~n10567 ) ;
  assign n10569 = ~n10563 & n10568 ;
  assign n10570 = ( n5114 & n10545 ) | ( n5114 & ~n10569 ) | ( n10545 & ~n10569 ) ;
  assign n10571 = ~n10569 & n10570 ;
  assign n10572 = ( n7678 & n10559 ) | ( n7678 & n10571 ) | ( n10559 & n10571 ) ;
  assign n10573 = ~n10559 & n10572 ;
  assign n10574 = ( x299 & ~n10544 ) | ( x299 & n10573 ) | ( ~n10544 & n10573 ) ;
  assign n10575 = n10544 | n10574 ;
  assign n10576 = x166 & n5061 ;
  assign n10577 = ~n10554 & n10576 ;
  assign n10578 = n10545 | n10576 ;
  assign n10579 = ( n7669 & n10577 ) | ( n7669 & n10578 ) | ( n10577 & n10578 ) ;
  assign n10580 = ~n10577 & n10579 ;
  assign n10581 = ~n7669 & n7812 ;
  assign n10582 = x299 & ~n10581 ;
  assign n10583 = n10575 & ~n10582 ;
  assign n10584 = ( n10575 & n10580 ) | ( n10575 & n10583 ) | ( n10580 & n10583 ) ;
  assign n10585 = ( x156 & x232 ) | ( x156 & n10584 ) | ( x232 & n10584 ) ;
  assign n10586 = ~n10584 & n10585 ;
  assign n10587 = ~x166 & n5061 ;
  assign n10588 = ~n10562 & n10587 ;
  assign n10589 = n10545 ^ n5061 ^ 1'b0 ;
  assign n10590 = ( n10545 & n10566 ) | ( n10545 & n10589 ) | ( n10566 & n10589 ) ;
  assign n10591 = n10587 | n10590 ;
  assign n10592 = ( n7669 & n10588 ) | ( n7669 & n10591 ) | ( n10588 & n10591 ) ;
  assign n10593 = ~n10588 & n10592 ;
  assign n10594 = ( n10575 & n10583 ) | ( n10575 & n10593 ) | ( n10583 & n10593 ) ;
  assign n10595 = ( x156 & x232 ) | ( x156 & ~n10594 ) | ( x232 & ~n10594 ) ;
  assign n10596 = ~x156 & n10595 ;
  assign n10597 = n7671 & n10590 ;
  assign n10598 = n7678 | n7812 ;
  assign n10599 = n5114 & ~n10566 ;
  assign n10600 = n5114 | n10545 ;
  assign n10601 = n7678 & ~n10600 ;
  assign n10602 = ( n7678 & n10599 ) | ( n7678 & n10601 ) | ( n10599 & n10601 ) ;
  assign n10603 = ( x299 & n10598 ) | ( x299 & ~n10602 ) | ( n10598 & ~n10602 ) ;
  assign n10604 = ~x299 & n10603 ;
  assign n10605 = ( x232 & ~n10597 ) | ( x232 & n10604 ) | ( ~n10597 & n10604 ) ;
  assign n10606 = n10597 | n10605 ;
  assign n10607 = ( x39 & n10596 ) | ( x39 & n10606 ) | ( n10596 & n10606 ) ;
  assign n10608 = ~n10596 & n10607 ;
  assign n10609 = n10608 ^ n10586 ^ 1'b0 ;
  assign n10610 = ( n10586 & n10608 ) | ( n10586 & n10609 ) | ( n10608 & n10609 ) ;
  assign n10611 = ( x38 & ~n10586 ) | ( x38 & n10610 ) | ( ~n10586 & n10610 ) ;
  assign n10614 = n1224 | n7813 ;
  assign n10615 = ( n7732 & n7734 ) | ( n7732 & n10614 ) | ( n7734 & n10614 ) ;
  assign n10691 = ~x40 & n8032 ;
  assign n10692 = x95 | n10691 ;
  assign n10693 = ~n10615 & n10692 ;
  assign n10694 = n5075 & n10693 ;
  assign n10668 = ~x40 & n7911 ;
  assign n10695 = x95 | n10668 ;
  assign n10696 = ~n10119 & n10695 ;
  assign n10697 = x166 & n10695 ;
  assign n10698 = x153 & ~n10697 ;
  assign n10699 = ~n10696 & n10698 ;
  assign n10700 = x160 | n5075 ;
  assign n10701 = ( n10615 & ~n10699 ) | ( n10615 & n10700 ) | ( ~n10699 & n10700 ) ;
  assign n10702 = n10699 | n10701 ;
  assign n10631 = ~x40 & n7835 ;
  assign n10632 = x95 | n10631 ;
  assign n10633 = ~x40 & n7849 ;
  assign n10703 = x166 & n10633 ;
  assign n10704 = n10632 | n10703 ;
  assign n10705 = ( x153 & ~n10702 ) | ( x153 & n10704 ) | ( ~n10702 & n10704 ) ;
  assign n10706 = ~n10702 & n10705 ;
  assign n10707 = n7812 & ~n8898 ;
  assign n10636 = n5075 | n7813 ;
  assign n10708 = ~n10636 & n10697 ;
  assign n10709 = ( x153 & n10707 ) | ( x153 & ~n10708 ) | ( n10707 & ~n10708 ) ;
  assign n10710 = ~n10707 & n10709 ;
  assign n10711 = ~n10636 & n10704 ;
  assign n10712 = x153 | n10711 ;
  assign n10713 = ( x160 & n10710 ) | ( x160 & n10712 ) | ( n10710 & n10712 ) ;
  assign n10714 = ~n10710 & n10713 ;
  assign n10715 = ( x163 & n10706 ) | ( x163 & ~n10714 ) | ( n10706 & ~n10714 ) ;
  assign n10716 = ~n10706 & n10715 ;
  assign n10717 = x210 & ~n7818 ;
  assign n10619 = n7815 & ~n7894 ;
  assign n10620 = x95 | n10619 ;
  assign n10621 = ~n7813 & n10620 ;
  assign n10718 = x210 | n10621 ;
  assign n10719 = ~n8898 & n10718 ;
  assign n10720 = n10719 ^ n10717 ^ 1'b0 ;
  assign n10721 = ( n10717 & n10719 ) | ( n10717 & n10720 ) | ( n10719 & n10720 ) ;
  assign n10722 = ( x153 & ~n10717 ) | ( x153 & n10721 ) | ( ~n10717 & n10721 ) ;
  assign n10723 = n10722 ^ n10691 ^ 1'b0 ;
  assign n10724 = ( n10407 & ~n10691 ) | ( n10407 & n10723 ) | ( ~n10691 & n10723 ) ;
  assign n10725 = ( n10691 & n10722 ) | ( n10691 & n10724 ) | ( n10722 & n10724 ) ;
  assign n10726 = n10725 ^ x163 ^ 1'b0 ;
  assign n10644 = x95 | n7926 ;
  assign n10645 = ~n7813 & n10644 ;
  assign n10732 = x210 & ~n10645 ;
  assign n10733 = x210 | n7933 ;
  assign n10734 = ( n10407 & n10732 ) | ( n10407 & n10733 ) | ( n10732 & n10733 ) ;
  assign n10735 = ~n10732 & n10734 ;
  assign n10727 = x210 & ~n7892 ;
  assign n10728 = n8898 | n10727 ;
  assign n10729 = x210 | n7897 ;
  assign n10730 = x153 & ~n10729 ;
  assign n10731 = ( x153 & n10728 ) | ( x153 & n10730 ) | ( n10728 & n10730 ) ;
  assign n10736 = n10735 ^ n10731 ^ 1'b0 ;
  assign n10737 = ( x160 & ~n10731 ) | ( x160 & n10735 ) | ( ~n10731 & n10735 ) ;
  assign n10738 = ( x160 & ~n10736 ) | ( x160 & n10737 ) | ( ~n10736 & n10737 ) ;
  assign n10739 = ( n10725 & ~n10726 ) | ( n10725 & n10738 ) | ( ~n10726 & n10738 ) ;
  assign n10740 = ( x163 & n10726 ) | ( x163 & n10739 ) | ( n10726 & n10739 ) ;
  assign n10680 = ~n10615 & n10620 ;
  assign n10741 = x210 | n10680 ;
  assign n10682 = n7817 & ~n10615 ;
  assign n10742 = x210 & ~n10682 ;
  assign n10743 = n8898 | n10742 ;
  assign n10744 = ( x153 & n10741 ) | ( x153 & ~n10743 ) | ( n10741 & ~n10743 ) ;
  assign n10745 = n10744 ^ n10741 ^ 1'b0 ;
  assign n10746 = ( x153 & n10744 ) | ( x153 & ~n10745 ) | ( n10744 & ~n10745 ) ;
  assign n10747 = n10746 ^ x166 ^ 1'b0 ;
  assign n10748 = ( ~x166 & n10693 ) | ( ~x166 & n10747 ) | ( n10693 & n10747 ) ;
  assign n10749 = ( x166 & n10746 ) | ( x166 & n10748 ) | ( n10746 & n10748 ) ;
  assign n10655 = ~n10615 & n10644 ;
  assign n10750 = x210 & ~n10655 ;
  assign n10653 = n7932 & ~n10615 ;
  assign n10751 = x210 | n10653 ;
  assign n10752 = ( n10407 & n10750 ) | ( n10407 & n10751 ) | ( n10750 & n10751 ) ;
  assign n10753 = ~n10750 & n10752 ;
  assign n10754 = n7891 & ~n10615 ;
  assign n10755 = x210 & ~n10754 ;
  assign n10756 = n7896 & ~n10615 ;
  assign n10757 = x210 | n10756 ;
  assign n10758 = ( n8898 & ~n10755 ) | ( n8898 & n10757 ) | ( ~n10755 & n10757 ) ;
  assign n10759 = ~n8898 & n10758 ;
  assign n10760 = ( x153 & n10753 ) | ( x153 & ~n10759 ) | ( n10753 & ~n10759 ) ;
  assign n10761 = ~n10753 & n10760 ;
  assign n10762 = ( x160 & n10749 ) | ( x160 & ~n10761 ) | ( n10749 & ~n10761 ) ;
  assign n10763 = ~x160 & n10762 ;
  assign n10764 = ( ~n10716 & n10740 ) | ( ~n10716 & n10763 ) | ( n10740 & n10763 ) ;
  assign n10765 = ~n10716 & n10764 ;
  assign n10766 = ( x299 & n10694 ) | ( x299 & ~n10765 ) | ( n10694 & ~n10765 ) ;
  assign n10767 = ~n10694 & n10766 ;
  assign n10612 = ~x40 & n7855 ;
  assign n10613 = x95 | n10612 ;
  assign n10616 = n10613 & ~n10615 ;
  assign n10617 = n5075 & n10616 ;
  assign n10618 = x198 & ~n7818 ;
  assign n10622 = x198 | n10621 ;
  assign n10623 = ( n8905 & ~n10618 ) | ( n8905 & n10622 ) | ( ~n10618 & n10622 ) ;
  assign n10624 = ~n8905 & n10623 ;
  assign n10625 = ( x182 & x184 ) | ( x182 & ~n10624 ) | ( x184 & ~n10624 ) ;
  assign n10626 = ~x184 & n10625 ;
  assign n10627 = ( n10449 & n10612 ) | ( n10449 & ~n10626 ) | ( n10612 & ~n10626 ) ;
  assign n10628 = n10627 ^ n10626 ^ 1'b0 ;
  assign n10629 = ( n10626 & ~n10627 ) | ( n10626 & n10628 ) | ( ~n10627 & n10628 ) ;
  assign n10630 = ~x182 & n10615 ;
  assign n10634 = x189 & n10633 ;
  assign n10635 = n10632 | n10634 ;
  assign n10637 = ( x182 & n5075 ) | ( x182 & n10636 ) | ( n5075 & n10636 ) ;
  assign n10638 = ( n10630 & n10635 ) | ( n10630 & ~n10637 ) | ( n10635 & ~n10637 ) ;
  assign n10639 = ~n10630 & n10638 ;
  assign n10640 = ~n10629 & n10639 ;
  assign n10641 = ( x184 & n10629 ) | ( x184 & ~n10640 ) | ( n10629 & ~n10640 ) ;
  assign n10642 = ( x175 & ~x299 ) | ( x175 & n10641 ) | ( ~x299 & n10641 ) ;
  assign n10643 = ~x175 & n10642 ;
  assign n10646 = x198 & ~n10645 ;
  assign n10647 = x198 | n7933 ;
  assign n10648 = ( n10449 & n10646 ) | ( n10449 & n10647 ) | ( n10646 & n10647 ) ;
  assign n10649 = ~n10646 & n10648 ;
  assign n10650 = n7899 & ~n8905 ;
  assign n10651 = ( x182 & n10649 ) | ( x182 & ~n10650 ) | ( n10649 & ~n10650 ) ;
  assign n10652 = ~n10649 & n10651 ;
  assign n10654 = x198 | n10653 ;
  assign n10656 = x198 & ~n10655 ;
  assign n10657 = n10449 & ~n10656 ;
  assign n10658 = n10654 & n10657 ;
  assign n10659 = ( x182 & ~n10652 ) | ( x182 & n10658 ) | ( ~n10652 & n10658 ) ;
  assign n10660 = ~n10652 & n10659 ;
  assign n10661 = n8905 | n10615 ;
  assign n10662 = x95 & ~x182 ;
  assign n10663 = n7899 | n10662 ;
  assign n10664 = ~n10661 & n10663 ;
  assign n10665 = ( ~x184 & n10660 ) | ( ~x184 & n10664 ) | ( n10660 & n10664 ) ;
  assign n10666 = ~x184 & n10665 ;
  assign n10667 = x175 & ~x299 ;
  assign n10669 = ~x95 & x189 ;
  assign n10670 = ( n7812 & n10668 ) | ( n7812 & n10669 ) | ( n10668 & n10669 ) ;
  assign n10671 = x182 & ~n10670 ;
  assign n10672 = ( x95 & n10670 ) | ( x95 & ~n10671 ) | ( n10670 & ~n10671 ) ;
  assign n10673 = n10371 & ~n10630 ;
  assign n10674 = n10672 & n10673 ;
  assign n10675 = ( n10666 & n10667 ) | ( n10666 & ~n10674 ) | ( n10667 & ~n10674 ) ;
  assign n10676 = ~n10666 & n10675 ;
  assign n10677 = ( ~n10617 & n10643 ) | ( ~n10617 & n10676 ) | ( n10643 & n10676 ) ;
  assign n10678 = ~n10617 & n10677 ;
  assign n10679 = n8905 & n10616 ;
  assign n10681 = x198 | n10680 ;
  assign n10683 = x198 & ~n10682 ;
  assign n10684 = ( n8905 & n10681 ) | ( n8905 & ~n10683 ) | ( n10681 & ~n10683 ) ;
  assign n10685 = ~n8905 & n10684 ;
  assign n10686 = x182 | x184 ;
  assign n10687 = ( n10436 & ~n10685 ) | ( n10436 & n10686 ) | ( ~n10685 & n10686 ) ;
  assign n10688 = n10685 | n10687 ;
  assign n10689 = ( ~n10678 & n10679 ) | ( ~n10678 & n10688 ) | ( n10679 & n10688 ) ;
  assign n10690 = ~n10678 & n10689 ;
  assign n10768 = n10767 ^ n10690 ^ 1'b0 ;
  assign n10769 = ( x232 & ~n10690 ) | ( x232 & n10767 ) | ( ~n10690 & n10767 ) ;
  assign n10770 = ( x232 & ~n10768 ) | ( x232 & n10769 ) | ( ~n10768 & n10769 ) ;
  assign n10771 = ~x299 & n10616 ;
  assign n10772 = x299 & n10693 ;
  assign n10773 = ( x232 & ~n10771 ) | ( x232 & n10772 ) | ( ~n10771 & n10772 ) ;
  assign n10774 = n10771 | n10773 ;
  assign n10775 = ( x39 & ~n10770 ) | ( x39 & n10774 ) | ( ~n10770 & n10774 ) ;
  assign n10776 = ~x39 & n10775 ;
  assign n10777 = ( ~n10389 & n10611 ) | ( ~n10389 & n10776 ) | ( n10611 & n10776 ) ;
  assign n10778 = ~n10389 & n10777 ;
  assign n10779 = ( x87 & x100 ) | ( x87 & ~n10778 ) | ( x100 & ~n10778 ) ;
  assign n10780 = n10778 | n10779 ;
  assign n10781 = x87 & n1230 ;
  assign n10782 = ~n10337 & n10781 ;
  assign n10783 = n10509 | n10782 ;
  assign n10784 = x87 & ~n10783 ;
  assign n10785 = ( n10507 & n10780 ) | ( n10507 & ~n10784 ) | ( n10780 & ~n10784 ) ;
  assign n10786 = ~n10507 & n10785 ;
  assign n10787 = ( x75 & x92 ) | ( x75 & ~n10786 ) | ( x92 & ~n10786 ) ;
  assign n10788 = n10786 | n10787 ;
  assign n10789 = x39 & ~n7812 ;
  assign n10790 = n8223 | n10789 ;
  assign n10791 = ~n1230 & n10517 ;
  assign n10792 = ( ~x39 & n10549 ) | ( ~x39 & n10791 ) | ( n10549 & n10791 ) ;
  assign n10793 = ~x39 & n10792 ;
  assign n10794 = ( ~n10783 & n10790 ) | ( ~n10783 & n10793 ) | ( n10790 & n10793 ) ;
  assign n10795 = ~n10783 & n10794 ;
  assign n10796 = ( n7639 & n10507 ) | ( n7639 & n10795 ) | ( n10507 & n10795 ) ;
  assign n10797 = n10795 ^ n10507 ^ 1'b0 ;
  assign n10798 = ( n7639 & n10796 ) | ( n7639 & n10797 ) | ( n10796 & n10797 ) ;
  assign n10799 = n10377 & ~n10798 ;
  assign n10800 = ( x75 & n10798 ) | ( x75 & ~n10799 ) | ( n10798 & ~n10799 ) ;
  assign n10801 = ( x54 & n10788 ) | ( x54 & ~n10800 ) | ( n10788 & ~n10800 ) ;
  assign n10802 = n10801 ^ n10788 ^ 1'b0 ;
  assign n10803 = ( x54 & n10801 ) | ( x54 & ~n10802 ) | ( n10801 & ~n10802 ) ;
  assign n10804 = n10803 ^ n10380 ^ 1'b0 ;
  assign n10805 = ( n10380 & n10803 ) | ( n10380 & n10804 ) | ( n10803 & n10804 ) ;
  assign n10806 = ( x74 & ~n10380 ) | ( x74 & n10805 ) | ( ~n10380 & n10805 ) ;
  assign n10807 = ( x55 & ~n10532 ) | ( x55 & n10806 ) | ( ~n10532 & n10806 ) ;
  assign n10808 = ~x55 & n10807 ;
  assign n10809 = n7643 & ~n10341 ;
  assign n10810 = n7639 & ~n10809 ;
  assign n10811 = n10326 | n10810 ;
  assign n10812 = n5075 & ~n7598 ;
  assign n10813 = n7569 | n10812 ;
  assign n10814 = n10351 & ~n10813 ;
  assign n10815 = n10549 | n10814 ;
  assign n10816 = x39 | n10815 ;
  assign n10817 = ( ~x39 & n10790 ) | ( ~x39 & n10816 ) | ( n10790 & n10816 ) ;
  assign n10818 = ( ~n10339 & n10782 ) | ( ~n10339 & n10817 ) | ( n10782 & n10817 ) ;
  assign n10819 = ~n10782 & n10818 ;
  assign n10820 = ( ~n2053 & n10327 ) | ( ~n2053 & n10819 ) | ( n10327 & n10819 ) ;
  assign n10821 = ~n2053 & n10820 ;
  assign n10822 = ( ~x54 & n10811 ) | ( ~x54 & n10821 ) | ( n10811 & n10821 ) ;
  assign n10823 = ~x54 & n10822 ;
  assign n10824 = ( ~x74 & n10349 ) | ( ~x74 & n10823 ) | ( n10349 & n10823 ) ;
  assign n10825 = ~x74 & n10824 ;
  assign n10826 = ( x55 & n10333 ) | ( x55 & ~n10825 ) | ( n10333 & ~n10825 ) ;
  assign n10827 = ~n10333 & n10826 ;
  assign n10828 = ( n2109 & ~n10808 ) | ( n2109 & n10827 ) | ( ~n10808 & n10827 ) ;
  assign n10829 = n10808 | n10828 ;
  assign n10830 = ( n7573 & ~n10348 ) | ( n7573 & n10829 ) | ( ~n10348 & n10829 ) ;
  assign n10831 = ~n7573 & n10830 ;
  assign n10832 = ( ~n10331 & n10334 ) | ( ~n10331 & n10831 ) | ( n10334 & n10831 ) ;
  assign n10833 = n10831 ^ n10331 ^ 1'b0 ;
  assign n10834 = ( n10831 & n10832 ) | ( n10831 & ~n10833 ) | ( n10832 & ~n10833 ) ;
  assign n10835 = ( n10541 & ~n10543 ) | ( n10541 & n10834 ) | ( ~n10543 & n10834 ) ;
  assign n10836 = ~n10543 & n10835 ;
  assign n10837 = x79 | n10834 ;
  assign n10838 = n10836 ^ n10540 ^ 1'b0 ;
  assign n10839 = ( ~n10540 & n10837 ) | ( ~n10540 & n10838 ) | ( n10837 & n10838 ) ;
  assign n10840 = ( n10540 & n10836 ) | ( n10540 & n10839 ) | ( n10836 & n10839 ) ;
  assign n10841 = x1163 | n7441 ;
  assign n10842 = x98 & x1092 ;
  assign n10843 = x1093 & n10842 ;
  assign n10844 = ~x567 & n1611 ;
  assign n10845 = n10843 | n10844 ;
  assign n10846 = n7276 & ~n10845 ;
  assign n10847 = x588 & ~n10846 ;
  assign n10849 = n6782 & ~n10845 ;
  assign n10850 = n6782 | n10844 ;
  assign n10851 = ( x1093 & n6489 ) | ( x1093 & n10842 ) | ( n6489 & n10842 ) ;
  assign n10852 = n6513 & n10851 ;
  assign n10853 = x1091 & n10843 ;
  assign n10854 = x110 | n1371 ;
  assign n10855 = x88 | n1261 ;
  assign n10856 = n8975 | n10855 ;
  assign n10857 = n10854 | n10856 ;
  assign n10858 = n6381 | n10857 ;
  assign n10859 = n6388 | n10858 ;
  assign n10860 = x824 & x950 ;
  assign n10861 = ~n1291 & n10860 ;
  assign n10862 = ~n10859 & n10861 ;
  assign n10863 = ( x98 & x1092 ) | ( x98 & n10862 ) | ( x1092 & n10862 ) ;
  assign n10864 = x1092 & n10863 ;
  assign n10865 = n10853 | n10864 ;
  assign n10866 = n10852 & n10865 ;
  assign n10867 = n2036 & n10843 ;
  assign n10868 = n10866 | n10867 ;
  assign n10869 = ~n1207 & n10851 ;
  assign n10870 = ~x841 & n1374 ;
  assign n10871 = x90 & x93 ;
  assign n10872 = n10870 & ~n10871 ;
  assign n10873 = ( n1411 & ~n10858 ) | ( n1411 & n10872 ) | ( ~n10858 & n10872 ) ;
  assign n10874 = ~n1411 & n10873 ;
  assign n10875 = n10859 & ~n10874 ;
  assign n10876 = ( x51 & n10874 ) | ( x51 & ~n10875 ) | ( n10874 & ~n10875 ) ;
  assign n10877 = ( n6399 & n10860 ) | ( n6399 & n10876 ) | ( n10860 & n10876 ) ;
  assign n10878 = ~n6399 & n10877 ;
  assign n10879 = ( x98 & x1092 ) | ( x98 & n10878 ) | ( x1092 & n10878 ) ;
  assign n10880 = x1092 & n10879 ;
  assign n10881 = n10853 | n10880 ;
  assign n10882 = n10869 & n10881 ;
  assign n10883 = ( x75 & ~n10868 ) | ( x75 & n10882 ) | ( ~n10868 & n10882 ) ;
  assign n10884 = n10868 | n10883 ;
  assign n10885 = x75 & ~n10843 ;
  assign n10886 = x567 & ~n10885 ;
  assign n10887 = n10884 & n10886 ;
  assign n10888 = ( ~n10849 & n10850 ) | ( ~n10849 & n10887 ) | ( n10850 & n10887 ) ;
  assign n10889 = ~n10849 & n10888 ;
  assign n10890 = x592 & ~n10889 ;
  assign n10891 = x592 | n10845 ;
  assign n10892 = ~n10890 & n10891 ;
  assign n10893 = n10892 ^ n10889 ^ n10845 ;
  assign n10848 = x443 & ~n10845 ;
  assign n10894 = x443 | n10893 ;
  assign n10895 = ~n10848 & n10894 ;
  assign n10896 = n10895 ^ n10893 ^ n10845 ;
  assign n10897 = n10896 ^ n7280 ^ 1'b0 ;
  assign n10898 = ( n10895 & n10896 ) | ( n10895 & n10897 ) | ( n10896 & n10897 ) ;
  assign n10899 = n10898 ^ x435 ^ 1'b0 ;
  assign n10900 = n10898 ^ n10893 ^ n10845 ;
  assign n10901 = ( n10898 & n10899 ) | ( n10898 & n10900 ) | ( n10899 & n10900 ) ;
  assign n10902 = x429 & n10901 ;
  assign n10903 = ( n10898 & ~n10899 ) | ( n10898 & n10900 ) | ( ~n10899 & n10900 ) ;
  assign n10904 = ~x429 & n10903 ;
  assign n10905 = ( n7278 & n10902 ) | ( n7278 & ~n10904 ) | ( n10902 & ~n10904 ) ;
  assign n10906 = ~n10902 & n10905 ;
  assign n10907 = ~x429 & n10901 ;
  assign n10908 = x429 & n10903 ;
  assign n10909 = ( n7278 & ~n10907 ) | ( n7278 & n10908 ) | ( ~n10907 & n10908 ) ;
  assign n10910 = n10907 | n10909 ;
  assign n10911 = ( x1196 & n10906 ) | ( x1196 & n10910 ) | ( n10906 & n10910 ) ;
  assign n10912 = ~n10906 & n10911 ;
  assign n10913 = ~x1196 & n10845 ;
  assign n10914 = ( n7327 & ~n10912 ) | ( n7327 & n10913 ) | ( ~n10912 & n10913 ) ;
  assign n10915 = n10912 | n10914 ;
  assign n10916 = n10915 ^ n10893 ^ 1'b0 ;
  assign n10917 = ( ~n7327 & n10893 ) | ( ~n7327 & n10916 ) | ( n10893 & n10916 ) ;
  assign n10918 = ( n10915 & ~n10916 ) | ( n10915 & n10917 ) | ( ~n10916 & n10917 ) ;
  assign n10919 = n10893 ^ x428 ^ 1'b0 ;
  assign n10920 = ( n10893 & n10918 ) | ( n10893 & ~n10919 ) | ( n10918 & ~n10919 ) ;
  assign n10921 = ( n10893 & n10918 ) | ( n10893 & n10919 ) | ( n10918 & n10919 ) ;
  assign n10922 = n10920 ^ x427 ^ 1'b0 ;
  assign n10923 = ( n10920 & n10921 ) | ( n10920 & n10922 ) | ( n10921 & n10922 ) ;
  assign n10924 = ( n10920 & n10921 ) | ( n10920 & ~n10922 ) | ( n10921 & ~n10922 ) ;
  assign n10925 = n10923 ^ x430 ^ 1'b0 ;
  assign n10926 = ( n10923 & n10924 ) | ( n10923 & ~n10925 ) | ( n10924 & ~n10925 ) ;
  assign n10927 = ( n10923 & n10924 ) | ( n10923 & n10925 ) | ( n10924 & n10925 ) ;
  assign n10928 = n10926 ^ x426 ^ 1'b0 ;
  assign n10929 = ( n10926 & n10927 ) | ( n10926 & ~n10928 ) | ( n10927 & ~n10928 ) ;
  assign n10930 = ( n10926 & n10927 ) | ( n10926 & n10928 ) | ( n10927 & n10928 ) ;
  assign n10931 = n10929 ^ x445 ^ 1'b0 ;
  assign n10932 = ( n10929 & n10930 ) | ( n10929 & ~n10931 ) | ( n10930 & ~n10931 ) ;
  assign n10933 = x448 & n10932 ;
  assign n10934 = ( n10929 & n10930 ) | ( n10929 & n10931 ) | ( n10930 & n10931 ) ;
  assign n10935 = ~x448 & n10934 ;
  assign n10936 = ( n7302 & ~n10933 ) | ( n7302 & n10935 ) | ( ~n10933 & n10935 ) ;
  assign n10937 = n10933 | n10936 ;
  assign n10938 = x448 & n10934 ;
  assign n10939 = ~x448 & n10932 ;
  assign n10940 = ( n7302 & n10938 ) | ( n7302 & ~n10939 ) | ( n10938 & ~n10939 ) ;
  assign n10941 = ~n10938 & n10940 ;
  assign n10942 = x1199 & ~n10941 ;
  assign n10943 = n10937 & n10942 ;
  assign n10944 = ~x1199 & n10918 ;
  assign n10945 = ( n7276 & ~n10943 ) | ( n7276 & n10944 ) | ( ~n10943 & n10944 ) ;
  assign n10946 = n10943 | n10945 ;
  assign n10947 = n10847 & n10946 ;
  assign n10948 = x591 & n10845 ;
  assign n10949 = ~n7179 & n10845 ;
  assign n10950 = n7179 & n10893 ;
  assign n10951 = ( x1198 & n10949 ) | ( x1198 & ~n10950 ) | ( n10949 & ~n10950 ) ;
  assign n10952 = ~n10949 & n10951 ;
  assign n10953 = x1198 | n10913 ;
  assign n10954 = ~n6533 & n10845 ;
  assign n10955 = n6533 & n10893 ;
  assign n10956 = n10954 | n10955 ;
  assign n10957 = n10956 ^ x355 ^ 1'b0 ;
  assign n10958 = n10956 ^ n10893 ^ n10845 ;
  assign n10959 = ( n10956 & n10957 ) | ( n10956 & n10958 ) | ( n10957 & n10958 ) ;
  assign n10960 = x458 & n10959 ;
  assign n10961 = ( n10956 & ~n10957 ) | ( n10956 & n10958 ) | ( ~n10957 & n10958 ) ;
  assign n10962 = ~x458 & n10961 ;
  assign n10963 = ( n6531 & n10960 ) | ( n6531 & ~n10962 ) | ( n10960 & ~n10962 ) ;
  assign n10964 = ~n10960 & n10963 ;
  assign n10965 = ~x458 & n10959 ;
  assign n10966 = x458 & n10961 ;
  assign n10967 = ( n6531 & ~n10965 ) | ( n6531 & n10966 ) | ( ~n10965 & n10966 ) ;
  assign n10968 = n10965 | n10967 ;
  assign n10969 = ( x1196 & n10964 ) | ( x1196 & n10968 ) | ( n10964 & n10968 ) ;
  assign n10970 = ~n10964 & n10969 ;
  assign n10971 = ( ~n10952 & n10953 ) | ( ~n10952 & n10970 ) | ( n10953 & n10970 ) ;
  assign n10972 = ~n10952 & n10971 ;
  assign n10973 = n10893 ^ n6585 ^ 1'b0 ;
  assign n10974 = ( n10893 & n10972 ) | ( n10893 & ~n10973 ) | ( n10972 & ~n10973 ) ;
  assign n10975 = ~n6529 & n10974 ;
  assign n10976 = x1199 & n10893 ;
  assign n10977 = x351 & n10976 ;
  assign n10978 = n10975 | n10977 ;
  assign n10979 = ~n6590 & n10974 ;
  assign n10980 = ~x351 & n10976 ;
  assign n10981 = n10979 | n10980 ;
  assign n10982 = n10978 ^ x461 ^ 1'b0 ;
  assign n10983 = ( n10978 & n10981 ) | ( n10978 & n10982 ) | ( n10981 & n10982 ) ;
  assign n10984 = ( n10978 & n10981 ) | ( n10978 & ~n10982 ) | ( n10981 & ~n10982 ) ;
  assign n10985 = n10983 ^ x357 ^ 1'b0 ;
  assign n10986 = ( n10983 & n10984 ) | ( n10983 & n10985 ) | ( n10984 & n10985 ) ;
  assign n10987 = ( n10983 & n10984 ) | ( n10983 & ~n10985 ) | ( n10984 & ~n10985 ) ;
  assign n10988 = n10986 ^ x356 ^ 1'b0 ;
  assign n10989 = ( n10986 & n10987 ) | ( n10986 & n10988 ) | ( n10987 & n10988 ) ;
  assign n10990 = x354 & n10989 ;
  assign n10991 = ( n10986 & n10987 ) | ( n10986 & ~n10988 ) | ( n10987 & ~n10988 ) ;
  assign n10992 = ~x354 & n10991 ;
  assign n10993 = ( n6507 & n10990 ) | ( n6507 & ~n10992 ) | ( n10990 & ~n10992 ) ;
  assign n10994 = ~n10990 & n10993 ;
  assign n10995 = ~x354 & n10989 ;
  assign n10996 = x354 & n10991 ;
  assign n10997 = ( n6507 & ~n10995 ) | ( n6507 & n10996 ) | ( ~n10995 & n10996 ) ;
  assign n10998 = n10995 | n10997 ;
  assign n10999 = ( x591 & ~n10994 ) | ( x591 & n10998 ) | ( ~n10994 & n10998 ) ;
  assign n11000 = ~x591 & n10999 ;
  assign n11001 = ( x590 & n10948 ) | ( x590 & ~n11000 ) | ( n10948 & ~n11000 ) ;
  assign n11002 = ~n10948 & n11001 ;
  assign n11003 = n7211 | n10845 ;
  assign n11004 = x1199 & n11003 ;
  assign n11005 = n6652 & ~n10892 ;
  assign n11006 = n6623 & ~n10892 ;
  assign n11007 = n6623 | n10845 ;
  assign n11008 = ( x1197 & n11006 ) | ( x1197 & n11007 ) | ( n11006 & n11007 ) ;
  assign n11009 = ~n11006 & n11008 ;
  assign n11010 = ~x1197 & n10845 ;
  assign n11011 = ( n6652 & ~n11009 ) | ( n6652 & n11010 ) | ( ~n11009 & n11010 ) ;
  assign n11012 = n11009 | n11011 ;
  assign n11013 = ( x1199 & ~n11005 ) | ( x1199 & n11012 ) | ( ~n11005 & n11012 ) ;
  assign n11014 = ~x1199 & n11013 ;
  assign n11015 = n7211 & ~n10892 ;
  assign n11016 = ~n11014 & n11015 ;
  assign n11017 = ( n11004 & n11014 ) | ( n11004 & ~n11016 ) | ( n11014 & ~n11016 ) ;
  assign n11018 = n10892 ^ x1198 ^ 1'b0 ;
  assign n11019 = ( n10892 & n11017 ) | ( n10892 & ~n11018 ) | ( n11017 & ~n11018 ) ;
  assign n11020 = n11017 ^ x374 ^ 1'b0 ;
  assign n11021 = ( n11017 & n11019 ) | ( n11017 & n11020 ) | ( n11019 & n11020 ) ;
  assign n11022 = x369 & n11021 ;
  assign n11023 = n7068 ^ x371 ^ x370 ;
  assign n11024 = ( n11017 & n11019 ) | ( n11017 & ~n11020 ) | ( n11019 & ~n11020 ) ;
  assign n11025 = ~x369 & n11024 ;
  assign n11026 = ( n11022 & n11023 ) | ( n11022 & ~n11025 ) | ( n11023 & ~n11025 ) ;
  assign n11027 = ~n11022 & n11026 ;
  assign n11028 = ~x369 & n11021 ;
  assign n11029 = x369 & n11024 ;
  assign n11030 = ( n11023 & ~n11028 ) | ( n11023 & n11029 ) | ( ~n11028 & n11029 ) ;
  assign n11031 = n11028 | n11030 ;
  assign n11032 = ( x591 & ~n11027 ) | ( x591 & n11031 ) | ( ~n11027 & n11031 ) ;
  assign n11033 = ~x591 & n11032 ;
  assign n11034 = n6862 & ~n10849 ;
  assign n11035 = ~x411 & n10842 ;
  assign n11036 = n6693 | n11035 ;
  assign n11037 = x411 & n10880 ;
  assign n11038 = n11036 | n11037 ;
  assign n11039 = x411 & n10842 ;
  assign n11040 = n6693 & ~n11039 ;
  assign n11041 = ~x411 & n10880 ;
  assign n11042 = n11040 & ~n11041 ;
  assign n11043 = n11038 & ~n11042 ;
  assign n11044 = n10853 | n11043 ;
  assign n11045 = n10869 & n11044 ;
  assign n11046 = ~x411 & n10864 ;
  assign n11047 = n11040 & ~n11046 ;
  assign n11048 = x411 & n10864 ;
  assign n11049 = ( n11036 & ~n11047 ) | ( n11036 & n11048 ) | ( ~n11047 & n11048 ) ;
  assign n11050 = ~n11047 & n11049 ;
  assign n11051 = n10853 | n11050 ;
  assign n11052 = n10852 & n11051 ;
  assign n11053 = ( n10867 & ~n11045 ) | ( n10867 & n11052 ) | ( ~n11045 & n11052 ) ;
  assign n11054 = n11045 | n11053 ;
  assign n11055 = x75 | n11054 ;
  assign n11056 = n10886 & n11055 ;
  assign n11057 = ( n10850 & n11034 ) | ( n10850 & n11056 ) | ( n11034 & n11056 ) ;
  assign n11058 = n11034 & n11057 ;
  assign n11059 = x592 & n10845 ;
  assign n11060 = n10913 | n11059 ;
  assign n11061 = ( x1199 & ~n11058 ) | ( x1199 & n11060 ) | ( ~n11058 & n11060 ) ;
  assign n11062 = n11058 | n11061 ;
  assign n11063 = n6702 & n10864 ;
  assign n11064 = ( n10842 & n10864 ) | ( n10842 & n11063 ) | ( n10864 & n11063 ) ;
  assign n11065 = n10866 & n11064 ;
  assign n11066 = ( n6702 & n10842 ) | ( n6702 & n10880 ) | ( n10842 & n10880 ) ;
  assign n11067 = n10882 & n11066 ;
  assign n11068 = ( n10867 & ~n11065 ) | ( n10867 & n11067 ) | ( ~n11065 & n11067 ) ;
  assign n11069 = n11065 | n11068 ;
  assign n11070 = ( n6917 & ~n10849 ) | ( n6917 & n11069 ) | ( ~n10849 & n11069 ) ;
  assign n11071 = ~n6917 & n11070 ;
  assign n11072 = n6702 & n10866 ;
  assign n11073 = ( n11054 & ~n11067 ) | ( n11054 & n11072 ) | ( ~n11067 & n11072 ) ;
  assign n11074 = n11067 | n11073 ;
  assign n11075 = n11071 ^ n11034 ^ 1'b0 ;
  assign n11076 = ( ~n11034 & n11074 ) | ( ~n11034 & n11075 ) | ( n11074 & n11075 ) ;
  assign n11077 = ( n11034 & n11071 ) | ( n11034 & n11076 ) | ( n11071 & n11076 ) ;
  assign n11078 = ( x75 & x567 ) | ( x75 & n11077 ) | ( x567 & n11077 ) ;
  assign n11079 = ~x75 & n11078 ;
  assign n11080 = n6707 | n10850 ;
  assign n11081 = n10845 & n11080 ;
  assign n11082 = ( x1199 & n11079 ) | ( x1199 & ~n11081 ) | ( n11079 & ~n11081 ) ;
  assign n11083 = ~n11079 & n11082 ;
  assign n11084 = ( n6689 & n11062 ) | ( n6689 & ~n11083 ) | ( n11062 & ~n11083 ) ;
  assign n11085 = ~n6689 & n11084 ;
  assign n11086 = ~x1197 & n11085 ;
  assign n11087 = x1197 | n6689 ;
  assign n11088 = n10893 & n11087 ;
  assign n11089 = n11086 | n11088 ;
  assign n11090 = n11089 ^ x333 ^ 1'b0 ;
  assign n11091 = ( n10893 & n11084 ) | ( n10893 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11092 = ( n11089 & n11090 ) | ( n11089 & n11091 ) | ( n11090 & n11091 ) ;
  assign n11093 = ( n11089 & ~n11090 ) | ( n11089 & n11091 ) | ( ~n11090 & n11091 ) ;
  assign n11094 = n11092 ^ x391 ^ 1'b0 ;
  assign n11095 = ( n11092 & n11093 ) | ( n11092 & n11094 ) | ( n11093 & n11094 ) ;
  assign n11096 = ( n11092 & n11093 ) | ( n11092 & ~n11094 ) | ( n11093 & ~n11094 ) ;
  assign n11097 = n11095 ^ x392 ^ 1'b0 ;
  assign n11098 = ( n11095 & n11096 ) | ( n11095 & ~n11097 ) | ( n11096 & ~n11097 ) ;
  assign n11099 = x393 & n11098 ;
  assign n11100 = ( n11095 & n11096 ) | ( n11095 & n11097 ) | ( n11096 & n11097 ) ;
  assign n11101 = ~x393 & n11100 ;
  assign n11102 = ( n6780 & n11099 ) | ( n6780 & ~n11101 ) | ( n11099 & ~n11101 ) ;
  assign n11103 = ~n11099 & n11102 ;
  assign n11104 = ~x393 & n11098 ;
  assign n11105 = x393 & n11100 ;
  assign n11106 = ( n6780 & ~n11104 ) | ( n6780 & n11105 ) | ( ~n11104 & n11105 ) ;
  assign n11107 = n11104 | n11106 ;
  assign n11108 = ( x591 & n11103 ) | ( x591 & n11107 ) | ( n11103 & n11107 ) ;
  assign n11109 = ~n11103 & n11108 ;
  assign n11110 = ( x590 & ~n11033 ) | ( x590 & n11109 ) | ( ~n11033 & n11109 ) ;
  assign n11111 = n11033 | n11110 ;
  assign n11112 = ( x588 & ~n11002 ) | ( x588 & n11111 ) | ( ~n11002 & n11111 ) ;
  assign n11113 = ~x588 & n11112 ;
  assign n11114 = ( n6612 & ~n10947 ) | ( n6612 & n11113 ) | ( ~n10947 & n11113 ) ;
  assign n11115 = n10947 | n11114 ;
  assign n11116 = n7180 | n10845 ;
  assign n11117 = x592 & n7327 ;
  assign n11118 = n6787 & n7298 ;
  assign n11119 = n11118 ^ n11117 ^ 1'b0 ;
  assign n11120 = ( n11117 & n11118 ) | ( n11117 & n11119 ) | ( n11118 & n11119 ) ;
  assign n11121 = ( n10845 & ~n11117 ) | ( n10845 & n11120 ) | ( ~n11117 & n11120 ) ;
  assign n11122 = n11116 ^ x428 ^ 1'b0 ;
  assign n11123 = ( n11116 & n11121 ) | ( n11116 & ~n11122 ) | ( n11121 & ~n11122 ) ;
  assign n11124 = ( n11116 & n11121 ) | ( n11116 & n11122 ) | ( n11121 & n11122 ) ;
  assign n11125 = n11123 ^ x427 ^ 1'b0 ;
  assign n11126 = ( n11123 & n11124 ) | ( n11123 & n11125 ) | ( n11124 & n11125 ) ;
  assign n11127 = ( n11123 & n11124 ) | ( n11123 & ~n11125 ) | ( n11124 & ~n11125 ) ;
  assign n11128 = n11126 ^ x430 ^ 1'b0 ;
  assign n11129 = ( n11126 & n11127 ) | ( n11126 & n11128 ) | ( n11127 & n11128 ) ;
  assign n11130 = ( n11126 & n11127 ) | ( n11126 & ~n11128 ) | ( n11127 & ~n11128 ) ;
  assign n11131 = n11129 ^ x426 ^ 1'b0 ;
  assign n11132 = ( n11129 & n11130 ) | ( n11129 & n11131 ) | ( n11130 & n11131 ) ;
  assign n11133 = ( n11129 & n11130 ) | ( n11129 & ~n11131 ) | ( n11130 & ~n11131 ) ;
  assign n11134 = n11132 ^ x445 ^ 1'b0 ;
  assign n11135 = ( n11132 & n11133 ) | ( n11132 & ~n11134 ) | ( n11133 & ~n11134 ) ;
  assign n11136 = x448 & n11135 ;
  assign n11137 = ( n11132 & n11133 ) | ( n11132 & n11134 ) | ( n11133 & n11134 ) ;
  assign n11138 = ~x448 & n11137 ;
  assign n11139 = ( n7302 & ~n11136 ) | ( n7302 & n11138 ) | ( ~n11136 & n11138 ) ;
  assign n11140 = n11136 | n11139 ;
  assign n11141 = x448 & n11137 ;
  assign n11142 = ~x448 & n11135 ;
  assign n11143 = ( n7302 & n11141 ) | ( n7302 & ~n11142 ) | ( n11141 & ~n11142 ) ;
  assign n11144 = ~n11141 & n11143 ;
  assign n11145 = x1199 & ~n11144 ;
  assign n11146 = n11140 & n11145 ;
  assign n11147 = ~x1199 & n11121 ;
  assign n11148 = ( n7276 & ~n11146 ) | ( n7276 & n11147 ) | ( ~n11146 & n11147 ) ;
  assign n11149 = n11146 | n11148 ;
  assign n11150 = n10847 & n11149 ;
  assign n11151 = n1611 ^ x567 ^ 1'b0 ;
  assign n11152 = x411 ^ x404 ^ x397 ;
  assign n11153 = n11152 ^ x410 ^ x390 ;
  assign n11154 = n6425 & ~n11153 ;
  assign n11155 = n10842 | n11154 ;
  assign n11156 = x412 & n11155 ;
  assign n11157 = n6425 & n11153 ;
  assign n11158 = n10842 | n11157 ;
  assign n11159 = ~x412 & n11158 ;
  assign n11160 = ( n6690 & ~n11156 ) | ( n6690 & n11159 ) | ( ~n11156 & n11159 ) ;
  assign n11161 = n11156 | n11160 ;
  assign n11162 = x412 & n11158 ;
  assign n11163 = ~x412 & n11155 ;
  assign n11164 = ( n6690 & n11162 ) | ( n6690 & ~n11163 ) | ( n11162 & ~n11163 ) ;
  assign n11165 = ~n11162 & n11164 ;
  assign n11166 = ( x122 & n11161 ) | ( x122 & ~n11165 ) | ( n11161 & ~n11165 ) ;
  assign n11167 = ~x122 & n11166 ;
  assign n11168 = n10842 | n11167 ;
  assign n11169 = n6489 & n11168 ;
  assign n11170 = n10853 | n11169 ;
  assign n11171 = ( n1611 & n11151 ) | ( n1611 & n11170 ) | ( n11151 & n11170 ) ;
  assign n11172 = n6862 & n11171 ;
  assign n11173 = n11060 | n11172 ;
  assign n11174 = n6425 & n6702 ;
  assign n11175 = x122 | n10842 ;
  assign n11176 = n11174 | n11175 ;
  assign n11177 = n10851 & n11176 ;
  assign n11178 = n6425 & n6783 ;
  assign n11179 = ~x1091 & n11178 ;
  assign n11180 = n10843 | n11179 ;
  assign n11181 = ( n10843 & n11177 ) | ( n10843 & n11180 ) | ( n11177 & n11180 ) ;
  assign n11182 = ( n1611 & n11151 ) | ( n1611 & n11181 ) | ( n11151 & n11181 ) ;
  assign n11183 = ( x567 & n11171 ) | ( x567 & n11182 ) | ( n11171 & n11182 ) ;
  assign n11184 = n6862 & n11183 ;
  assign n11185 = ~n6917 & n11182 ;
  assign n11186 = ( n11059 & ~n11184 ) | ( n11059 & n11185 ) | ( ~n11184 & n11185 ) ;
  assign n11187 = n11184 | n11186 ;
  assign n11188 = n11173 ^ x1199 ^ 1'b0 ;
  assign n11189 = ( n11173 & n11187 ) | ( n11173 & n11188 ) | ( n11187 & n11188 ) ;
  assign n11190 = n11116 ^ n11087 ^ 1'b0 ;
  assign n11191 = ( n11116 & n11189 ) | ( n11116 & ~n11190 ) | ( n11189 & ~n11190 ) ;
  assign n11192 = n11116 ^ n6689 ^ 1'b0 ;
  assign n11193 = ( n11116 & n11189 ) | ( n11116 & ~n11192 ) | ( n11189 & ~n11192 ) ;
  assign n11194 = n11191 ^ x333 ^ 1'b0 ;
  assign n11195 = ( n11191 & n11193 ) | ( n11191 & n11194 ) | ( n11193 & n11194 ) ;
  assign n11196 = ~x391 & n11195 ;
  assign n11197 = n6781 ^ x392 ^ 1'b0 ;
  assign n11198 = ( n11191 & n11193 ) | ( n11191 & ~n11194 ) | ( n11193 & ~n11194 ) ;
  assign n11199 = x391 & n11198 ;
  assign n11200 = ( n11196 & n11197 ) | ( n11196 & ~n11199 ) | ( n11197 & ~n11199 ) ;
  assign n11201 = ~n11196 & n11200 ;
  assign n11202 = ~x391 & n11198 ;
  assign n11203 = x391 & n11195 ;
  assign n11204 = ( n11197 & ~n11202 ) | ( n11197 & n11203 ) | ( ~n11202 & n11203 ) ;
  assign n11205 = n11202 | n11204 ;
  assign n11206 = ( x591 & n11201 ) | ( x591 & n11205 ) | ( n11201 & n11205 ) ;
  assign n11207 = ~n11201 & n11206 ;
  assign n11208 = ( n7219 & n7223 ) | ( n7219 & n7224 ) | ( n7223 & n7224 ) ;
  assign n11209 = ( ~x591 & n10845 ) | ( ~x591 & n11208 ) | ( n10845 & n11208 ) ;
  assign n11210 = ~x591 & n11209 ;
  assign n11211 = ( x590 & ~n11207 ) | ( x590 & n11210 ) | ( ~n11207 & n11210 ) ;
  assign n11212 = n11207 | n11211 ;
  assign n11213 = n7161 | n10845 ;
  assign n11214 = n7185 | n11213 ;
  assign n11215 = n6529 | n11214 ;
  assign n11216 = n11116 & n11215 ;
  assign n11217 = n6590 | n11214 ;
  assign n11218 = n11116 & n11217 ;
  assign n11219 = n11216 ^ x461 ^ 1'b0 ;
  assign n11220 = ( n11216 & n11218 ) | ( n11216 & ~n11219 ) | ( n11218 & ~n11219 ) ;
  assign n11221 = ( n11216 & n11218 ) | ( n11216 & n11219 ) | ( n11218 & n11219 ) ;
  assign n11222 = n11220 ^ x357 ^ 1'b0 ;
  assign n11223 = ( n11220 & n11221 ) | ( n11220 & ~n11222 ) | ( n11221 & ~n11222 ) ;
  assign n11224 = ( n11220 & n11221 ) | ( n11220 & n11222 ) | ( n11221 & n11222 ) ;
  assign n11225 = n11223 ^ x356 ^ 1'b0 ;
  assign n11226 = ( n11223 & n11224 ) | ( n11223 & ~n11225 ) | ( n11224 & ~n11225 ) ;
  assign n11227 = ~x354 & n11226 ;
  assign n11228 = ( n11223 & n11224 ) | ( n11223 & n11225 ) | ( n11224 & n11225 ) ;
  assign n11229 = x354 & n11228 ;
  assign n11230 = ( n6507 & n11227 ) | ( n6507 & ~n11229 ) | ( n11227 & ~n11229 ) ;
  assign n11231 = ~n11227 & n11230 ;
  assign n11232 = x354 & n11226 ;
  assign n11233 = ~x354 & n11228 ;
  assign n11234 = ( n6507 & ~n11232 ) | ( n6507 & n11233 ) | ( ~n11232 & n11233 ) ;
  assign n11235 = n11232 | n11234 ;
  assign n11236 = ( x591 & ~n11231 ) | ( x591 & n11235 ) | ( ~n11231 & n11235 ) ;
  assign n11237 = ~x591 & n11236 ;
  assign n11238 = ( x590 & n10948 ) | ( x590 & ~n11237 ) | ( n10948 & ~n11237 ) ;
  assign n11239 = ~n10948 & n11238 ;
  assign n11240 = ( x588 & n11212 ) | ( x588 & ~n11239 ) | ( n11212 & ~n11239 ) ;
  assign n11241 = ~x588 & n11240 ;
  assign n11242 = ( n6612 & n11150 ) | ( n6612 & ~n11241 ) | ( n11150 & ~n11241 ) ;
  assign n11243 = ~n11150 & n11242 ;
  assign n11244 = ~x80 & n7318 ;
  assign n11245 = n6612 | n10845 ;
  assign n11246 = n11244 & n11245 ;
  assign n11247 = n11246 ^ n11243 ^ 1'b0 ;
  assign n11248 = ( n11243 & n11246 ) | ( n11243 & n11247 ) | ( n11246 & n11247 ) ;
  assign n11249 = ( x217 & ~n11243 ) | ( x217 & n11248 ) | ( ~n11243 & n11248 ) ;
  assign n11250 = n6369 & ~n11180 ;
  assign n11251 = n2036 | n10853 ;
  assign n11252 = ( n6489 & n11175 ) | ( n6489 & n11179 ) | ( n11175 & n11179 ) ;
  assign n11253 = n11251 | n11252 ;
  assign n11254 = x87 & ~n11251 ;
  assign n11255 = ~n10864 & n11254 ;
  assign n11256 = x87 | n11251 ;
  assign n11257 = n10880 | n11256 ;
  assign n11258 = x122 & ~n11257 ;
  assign n11259 = ( x122 & n11255 ) | ( x122 & n11258 ) | ( n11255 & n11258 ) ;
  assign n11260 = ( x75 & n11253 ) | ( x75 & ~n11259 ) | ( n11253 & ~n11259 ) ;
  assign n11261 = n11260 ^ n11253 ^ 1'b0 ;
  assign n11262 = ( x75 & n11260 ) | ( x75 & ~n11261 ) | ( n11260 & ~n11261 ) ;
  assign n11263 = x567 & ~n6782 ;
  assign n11264 = ( n11250 & n11262 ) | ( n11250 & n11263 ) | ( n11262 & n11263 ) ;
  assign n11265 = ~n11250 & n11264 ;
  assign n11266 = n6782 & n11180 ;
  assign n11267 = ( n10844 & ~n11265 ) | ( n10844 & n11266 ) | ( ~n11265 & n11266 ) ;
  assign n11268 = n11265 | n11267 ;
  assign n11269 = x592 & ~n11268 ;
  assign n11270 = n10891 & ~n11269 ;
  assign n11271 = n11270 ^ n11268 ^ n10845 ;
  assign n11272 = x1199 & n11271 ;
  assign n11273 = x351 & n11272 ;
  assign n11274 = n7179 & n11271 ;
  assign n11275 = ( x1198 & n10949 ) | ( x1198 & ~n11274 ) | ( n10949 & ~n11274 ) ;
  assign n11276 = ~n10949 & n11275 ;
  assign n11277 = n6533 & n11271 ;
  assign n11278 = n10954 | n11277 ;
  assign n11279 = n11278 ^ x355 ^ 1'b0 ;
  assign n11280 = n11278 ^ n11271 ^ n10845 ;
  assign n11281 = ( n11278 & n11279 ) | ( n11278 & n11280 ) | ( n11279 & n11280 ) ;
  assign n11282 = ~x458 & n11281 ;
  assign n11283 = ( n11278 & ~n11279 ) | ( n11278 & n11280 ) | ( ~n11279 & n11280 ) ;
  assign n11284 = x458 & n11283 ;
  assign n11285 = ( n6531 & ~n11282 ) | ( n6531 & n11284 ) | ( ~n11282 & n11284 ) ;
  assign n11286 = n11282 | n11285 ;
  assign n11287 = x458 & n11281 ;
  assign n11288 = ~x458 & n11283 ;
  assign n11289 = ( n6531 & n11287 ) | ( n6531 & ~n11288 ) | ( n11287 & ~n11288 ) ;
  assign n11290 = ~n11287 & n11289 ;
  assign n11291 = x1196 & ~n11290 ;
  assign n11292 = n11286 & n11291 ;
  assign n11293 = n10953 | n11292 ;
  assign n11294 = ~n11276 & n11293 ;
  assign n11295 = n11271 ^ n6585 ^ 1'b0 ;
  assign n11296 = ( n11271 & n11294 ) | ( n11271 & ~n11295 ) | ( n11294 & ~n11295 ) ;
  assign n11297 = ~n6529 & n11296 ;
  assign n11298 = n11273 | n11297 ;
  assign n11299 = ~x351 & n11272 ;
  assign n11300 = ~n6590 & n11296 ;
  assign n11301 = n11299 | n11300 ;
  assign n11302 = n11298 ^ x461 ^ 1'b0 ;
  assign n11303 = ( n11298 & n11301 ) | ( n11298 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11304 = ( n11298 & n11301 ) | ( n11298 & ~n11302 ) | ( n11301 & ~n11302 ) ;
  assign n11305 = n11303 ^ x357 ^ 1'b0 ;
  assign n11306 = ( n11303 & n11304 ) | ( n11303 & n11305 ) | ( n11304 & n11305 ) ;
  assign n11307 = ( n11303 & n11304 ) | ( n11303 & ~n11305 ) | ( n11304 & ~n11305 ) ;
  assign n11308 = n11306 ^ x356 ^ 1'b0 ;
  assign n11309 = ( n11306 & n11307 ) | ( n11306 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11310 = x354 & n11309 ;
  assign n11311 = ( n11306 & n11307 ) | ( n11306 & ~n11308 ) | ( n11307 & ~n11308 ) ;
  assign n11312 = ~x354 & n11311 ;
  assign n11313 = ( n6507 & n11310 ) | ( n6507 & ~n11312 ) | ( n11310 & ~n11312 ) ;
  assign n11314 = ~n11310 & n11313 ;
  assign n11315 = ~x354 & n11309 ;
  assign n11316 = x354 & n11311 ;
  assign n11317 = ( n6507 & ~n11315 ) | ( n6507 & n11316 ) | ( ~n11315 & n11316 ) ;
  assign n11318 = n11315 | n11317 ;
  assign n11319 = ( x591 & ~n11314 ) | ( x591 & n11318 ) | ( ~n11314 & n11318 ) ;
  assign n11320 = ~x591 & n11319 ;
  assign n11321 = ( x590 & n10948 ) | ( x590 & ~n11320 ) | ( n10948 & ~n11320 ) ;
  assign n11322 = ~n10948 & n11321 ;
  assign n11323 = x75 & ~n11170 ;
  assign n11324 = n11256 ^ n6489 ^ 1'b0 ;
  assign n11325 = x122 & n11043 ;
  assign n11326 = n11167 | n11325 ;
  assign n11327 = ( n6489 & ~n11324 ) | ( n6489 & n11326 ) | ( ~n11324 & n11326 ) ;
  assign n11328 = ( n11256 & n11324 ) | ( n11256 & n11327 ) | ( n11324 & n11327 ) ;
  assign n11329 = x122 & n11050 ;
  assign n11330 = n11167 | n11329 ;
  assign n11331 = ( n6489 & ~n11254 ) | ( n6489 & n11330 ) | ( ~n11254 & n11330 ) ;
  assign n11332 = n11254 ^ n6489 ^ 1'b0 ;
  assign n11333 = ( n11254 & ~n11331 ) | ( n11254 & n11332 ) | ( ~n11331 & n11332 ) ;
  assign n11334 = n11170 & ~n11333 ;
  assign n11335 = ( n2036 & n11333 ) | ( n2036 & ~n11334 ) | ( n11333 & ~n11334 ) ;
  assign n11336 = ( x75 & n11328 ) | ( x75 & ~n11335 ) | ( n11328 & ~n11335 ) ;
  assign n11337 = n11336 ^ n11328 ^ 1'b0 ;
  assign n11338 = ( x75 & n11336 ) | ( x75 & ~n11337 ) | ( n11336 & ~n11337 ) ;
  assign n11339 = ( n11263 & n11323 ) | ( n11263 & n11338 ) | ( n11323 & n11338 ) ;
  assign n11340 = ~n11323 & n11339 ;
  assign n11341 = n11340 ^ n10850 ^ 1'b0 ;
  assign n11342 = ( ~n10850 & n11171 ) | ( ~n10850 & n11341 ) | ( n11171 & n11341 ) ;
  assign n11343 = ( n10850 & n11340 ) | ( n10850 & n11342 ) | ( n11340 & n11342 ) ;
  assign n11344 = ( x592 & x1196 ) | ( x592 & n11343 ) | ( x1196 & n11343 ) ;
  assign n11345 = ~x592 & n11344 ;
  assign n11346 = ( ~x1199 & n10913 ) | ( ~x1199 & n11345 ) | ( n10913 & n11345 ) ;
  assign n11347 = ~x1199 & n11346 ;
  assign n11348 = n2036 | n11177 ;
  assign n11349 = ~n11064 & n11254 ;
  assign n11350 = n11066 | n11256 ;
  assign n11351 = x122 & ~n11350 ;
  assign n11352 = ( x122 & n11349 ) | ( x122 & n11351 ) | ( n11349 & n11351 ) ;
  assign n11353 = ( x75 & n11348 ) | ( x75 & ~n11352 ) | ( n11348 & ~n11352 ) ;
  assign n11354 = n11353 ^ n11348 ^ 1'b0 ;
  assign n11355 = ( x75 & n11353 ) | ( x75 & ~n11354 ) | ( n11353 & ~n11354 ) ;
  assign n11356 = n6369 & ~n11181 ;
  assign n11357 = n11263 & ~n11356 ;
  assign n11358 = n11355 & n11357 ;
  assign n11359 = n10850 & n11182 ;
  assign n11360 = ( ~n6917 & n11358 ) | ( ~n6917 & n11359 ) | ( n11358 & n11359 ) ;
  assign n11361 = ~n6917 & n11360 ;
  assign n11362 = ~n11169 & n11356 ;
  assign n11363 = ~x122 & n11174 ;
  assign n11364 = ( n11050 & ~n11063 ) | ( n11050 & n11254 ) | ( ~n11063 & n11254 ) ;
  assign n11365 = ~n11050 & n11364 ;
  assign n11366 = ( n6694 & n11041 ) | ( n6694 & n11043 ) | ( n11041 & n11043 ) ;
  assign n11367 = ( n11350 & ~n11365 ) | ( n11350 & n11366 ) | ( ~n11365 & n11366 ) ;
  assign n11368 = ~n11365 & n11367 ;
  assign n11369 = ( n11167 & ~n11363 ) | ( n11167 & n11368 ) | ( ~n11363 & n11368 ) ;
  assign n11370 = n11363 | n11369 ;
  assign n11371 = n11370 ^ x75 ^ 1'b0 ;
  assign n11372 = n11169 | n11348 ;
  assign n11373 = ( n11370 & ~n11371 ) | ( n11370 & n11372 ) | ( ~n11371 & n11372 ) ;
  assign n11374 = ( x75 & n11371 ) | ( x75 & n11373 ) | ( n11371 & n11373 ) ;
  assign n11375 = ( n11263 & n11362 ) | ( n11263 & n11374 ) | ( n11362 & n11374 ) ;
  assign n11376 = ~n11362 & n11375 ;
  assign n11377 = n11376 ^ n10850 ^ 1'b0 ;
  assign n11378 = ( ~n10850 & n11183 ) | ( ~n10850 & n11377 ) | ( n11183 & n11377 ) ;
  assign n11379 = ( n10850 & n11376 ) | ( n10850 & n11378 ) | ( n11376 & n11378 ) ;
  assign n11380 = ( x592 & x1196 ) | ( x592 & n11379 ) | ( x1196 & n11379 ) ;
  assign n11381 = ~x592 & n11380 ;
  assign n11382 = ( x1199 & n11361 ) | ( x1199 & n11381 ) | ( n11361 & n11381 ) ;
  assign n11383 = n11381 ^ n11361 ^ 1'b0 ;
  assign n11384 = ( x1199 & n11382 ) | ( x1199 & n11383 ) | ( n11382 & n11383 ) ;
  assign n11385 = ( n11059 & ~n11347 ) | ( n11059 & n11384 ) | ( ~n11347 & n11384 ) ;
  assign n11386 = n11347 | n11385 ;
  assign n11387 = n11271 ^ n11087 ^ 1'b0 ;
  assign n11388 = ( n11271 & n11386 ) | ( n11271 & ~n11387 ) | ( n11386 & ~n11387 ) ;
  assign n11389 = n11271 ^ n6689 ^ 1'b0 ;
  assign n11390 = ( n11271 & n11386 ) | ( n11271 & ~n11389 ) | ( n11386 & ~n11389 ) ;
  assign n11391 = n11388 ^ x333 ^ 1'b0 ;
  assign n11392 = ( n11388 & n11390 ) | ( n11388 & ~n11391 ) | ( n11390 & ~n11391 ) ;
  assign n11393 = ( n11388 & n11390 ) | ( n11388 & n11391 ) | ( n11390 & n11391 ) ;
  assign n11394 = n11392 ^ x391 ^ 1'b0 ;
  assign n11395 = ( n11392 & n11393 ) | ( n11392 & ~n11394 ) | ( n11393 & ~n11394 ) ;
  assign n11396 = ( n11392 & n11393 ) | ( n11392 & n11394 ) | ( n11393 & n11394 ) ;
  assign n11397 = n11395 ^ x392 ^ 1'b0 ;
  assign n11398 = ( n11395 & n11396 ) | ( n11395 & n11397 ) | ( n11396 & n11397 ) ;
  assign n11399 = ( n11395 & n11396 ) | ( n11395 & ~n11397 ) | ( n11396 & ~n11397 ) ;
  assign n11400 = n11398 ^ x393 ^ 1'b0 ;
  assign n11401 = ( n11398 & n11399 ) | ( n11398 & n11400 ) | ( n11399 & n11400 ) ;
  assign n11402 = n6780 & ~n11401 ;
  assign n11403 = ( n11398 & n11399 ) | ( n11398 & ~n11400 ) | ( n11399 & ~n11400 ) ;
  assign n11404 = n6780 | n11403 ;
  assign n11405 = ( x591 & n11402 ) | ( x591 & n11404 ) | ( n11402 & n11404 ) ;
  assign n11406 = ~n11402 & n11405 ;
  assign n11407 = n10845 ^ x367 ^ 1'b0 ;
  assign n11408 = ( n10845 & n11270 ) | ( n10845 & ~n11407 ) | ( n11270 & ~n11407 ) ;
  assign n11409 = ( n10845 & n11270 ) | ( n10845 & n11407 ) | ( n11270 & n11407 ) ;
  assign n11410 = n11408 ^ n6622 ^ 1'b0 ;
  assign n11411 = ( n11408 & n11409 ) | ( n11408 & ~n11410 ) | ( n11409 & ~n11410 ) ;
  assign n11412 = ~n6620 & n11411 ;
  assign n11413 = ( n11408 & n11409 ) | ( n11408 & n11410 ) | ( n11409 & n11410 ) ;
  assign n11414 = n6620 & n11413 ;
  assign n11415 = ( n6619 & ~n11412 ) | ( n6619 & n11414 ) | ( ~n11412 & n11414 ) ;
  assign n11416 = n11412 | n11415 ;
  assign n11417 = n6620 & n11411 ;
  assign n11418 = ~n6620 & n11413 ;
  assign n11419 = ( n6619 & n11417 ) | ( n6619 & ~n11418 ) | ( n11417 & ~n11418 ) ;
  assign n11420 = ~n11417 & n11419 ;
  assign n11421 = x1197 & ~n11420 ;
  assign n11422 = n11416 & n11421 ;
  assign n11423 = ( n6652 & n11010 ) | ( n6652 & ~n11422 ) | ( n11010 & ~n11422 ) ;
  assign n11424 = n11422 | n11423 ;
  assign n11425 = n6652 & ~n11270 ;
  assign n11426 = ( x1199 & n11424 ) | ( x1199 & ~n11425 ) | ( n11424 & ~n11425 ) ;
  assign n11427 = ~x1199 & n11426 ;
  assign n11428 = ~x1198 & n11427 ;
  assign n11429 = n10845 ^ n7211 ^ 1'b0 ;
  assign n11430 = ( n10845 & n11270 ) | ( n10845 & n11429 ) | ( n11270 & n11429 ) ;
  assign n11431 = n6658 & n11430 ;
  assign n11432 = x1198 & n11270 ;
  assign n11433 = ( ~n11428 & n11431 ) | ( ~n11428 & n11432 ) | ( n11431 & n11432 ) ;
  assign n11434 = n11428 | n11433 ;
  assign n11435 = n11434 ^ x374 ^ 1'b0 ;
  assign n11436 = ( n11426 & n11427 ) | ( n11426 & n11430 ) | ( n11427 & n11430 ) ;
  assign n11437 = ( n11434 & ~n11435 ) | ( n11434 & n11436 ) | ( ~n11435 & n11436 ) ;
  assign n11438 = ~x369 & n11437 ;
  assign n11439 = ( n11434 & n11435 ) | ( n11434 & n11436 ) | ( n11435 & n11436 ) ;
  assign n11440 = x369 & n11439 ;
  assign n11441 = ( n11023 & ~n11438 ) | ( n11023 & n11440 ) | ( ~n11438 & n11440 ) ;
  assign n11442 = n11438 | n11441 ;
  assign n11443 = ~x369 & n11439 ;
  assign n11444 = x369 & n11437 ;
  assign n11445 = ( n11023 & n11443 ) | ( n11023 & ~n11444 ) | ( n11443 & ~n11444 ) ;
  assign n11446 = ~n11443 & n11445 ;
  assign n11447 = ( x591 & n11442 ) | ( x591 & ~n11446 ) | ( n11442 & ~n11446 ) ;
  assign n11448 = ~x591 & n11447 ;
  assign n11449 = ( x590 & ~n11406 ) | ( x590 & n11448 ) | ( ~n11406 & n11448 ) ;
  assign n11450 = n11406 | n11449 ;
  assign n11451 = ( x588 & ~n11322 ) | ( x588 & n11450 ) | ( ~n11322 & n11450 ) ;
  assign n11452 = ~x588 & n11451 ;
  assign n11453 = x443 | n11271 ;
  assign n11454 = ~n10848 & n11453 ;
  assign n11455 = n11454 ^ n11271 ^ n10845 ;
  assign n11456 = n11455 ^ n7280 ^ 1'b0 ;
  assign n11457 = ( n11454 & n11455 ) | ( n11454 & n11456 ) | ( n11455 & n11456 ) ;
  assign n11458 = n11457 ^ x435 ^ 1'b0 ;
  assign n11459 = n11457 ^ n11271 ^ n10845 ;
  assign n11460 = ( n11457 & n11458 ) | ( n11457 & n11459 ) | ( n11458 & n11459 ) ;
  assign n11461 = x429 & n11460 ;
  assign n11462 = ( n11457 & ~n11458 ) | ( n11457 & n11459 ) | ( ~n11458 & n11459 ) ;
  assign n11463 = ~x429 & n11462 ;
  assign n11464 = ( n7278 & n11461 ) | ( n7278 & ~n11463 ) | ( n11461 & ~n11463 ) ;
  assign n11465 = ~n11461 & n11464 ;
  assign n11466 = ~x429 & n11460 ;
  assign n11467 = x429 & n11462 ;
  assign n11468 = ( n7278 & ~n11466 ) | ( n7278 & n11467 ) | ( ~n11466 & n11467 ) ;
  assign n11469 = n11466 | n11468 ;
  assign n11470 = ( x1196 & n11465 ) | ( x1196 & n11469 ) | ( n11465 & n11469 ) ;
  assign n11471 = ~n11465 & n11470 ;
  assign n11472 = ( n7327 & n10913 ) | ( n7327 & ~n11471 ) | ( n10913 & ~n11471 ) ;
  assign n11473 = n11471 | n11472 ;
  assign n11474 = n11473 ^ n11271 ^ 1'b0 ;
  assign n11475 = ( ~n7327 & n11271 ) | ( ~n7327 & n11474 ) | ( n11271 & n11474 ) ;
  assign n11476 = ( n11473 & ~n11474 ) | ( n11473 & n11475 ) | ( ~n11474 & n11475 ) ;
  assign n11477 = n11271 ^ x428 ^ 1'b0 ;
  assign n11478 = ( n11271 & n11476 ) | ( n11271 & ~n11477 ) | ( n11476 & ~n11477 ) ;
  assign n11479 = ( n11271 & n11476 ) | ( n11271 & n11477 ) | ( n11476 & n11477 ) ;
  assign n11480 = n11478 ^ x427 ^ 1'b0 ;
  assign n11481 = ( n11478 & n11479 ) | ( n11478 & n11480 ) | ( n11479 & n11480 ) ;
  assign n11482 = ( n11478 & n11479 ) | ( n11478 & ~n11480 ) | ( n11479 & ~n11480 ) ;
  assign n11483 = n11481 ^ x430 ^ 1'b0 ;
  assign n11484 = ( n11481 & n11482 ) | ( n11481 & ~n11483 ) | ( n11482 & ~n11483 ) ;
  assign n11485 = ( n11481 & n11482 ) | ( n11481 & n11483 ) | ( n11482 & n11483 ) ;
  assign n11486 = n11484 ^ x426 ^ 1'b0 ;
  assign n11487 = ( n11484 & n11485 ) | ( n11484 & ~n11486 ) | ( n11485 & ~n11486 ) ;
  assign n11488 = ( n11484 & n11485 ) | ( n11484 & n11486 ) | ( n11485 & n11486 ) ;
  assign n11489 = n11487 ^ x445 ^ 1'b0 ;
  assign n11490 = ( n11487 & n11488 ) | ( n11487 & ~n11489 ) | ( n11488 & ~n11489 ) ;
  assign n11491 = ~x448 & n11490 ;
  assign n11492 = ( n11487 & n11488 ) | ( n11487 & n11489 ) | ( n11488 & n11489 ) ;
  assign n11493 = x448 & n11492 ;
  assign n11494 = ( n7302 & n11491 ) | ( n7302 & ~n11493 ) | ( n11491 & ~n11493 ) ;
  assign n11495 = ~n11491 & n11494 ;
  assign n11496 = x448 & n11490 ;
  assign n11497 = ~x448 & n11492 ;
  assign n11498 = ( n7302 & ~n11496 ) | ( n7302 & n11497 ) | ( ~n11496 & n11497 ) ;
  assign n11499 = n11496 | n11498 ;
  assign n11500 = ( x1199 & n11495 ) | ( x1199 & n11499 ) | ( n11495 & n11499 ) ;
  assign n11501 = ~n11495 & n11500 ;
  assign n11502 = ~x1199 & n11476 ;
  assign n11503 = ( n7276 & ~n11501 ) | ( n7276 & n11502 ) | ( ~n11501 & n11502 ) ;
  assign n11504 = n11501 | n11503 ;
  assign n11505 = n10847 & n11504 ;
  assign n11506 = ( n6612 & n11452 ) | ( n6612 & ~n11505 ) | ( n11452 & ~n11505 ) ;
  assign n11507 = ~n11452 & n11506 ;
  assign n11508 = ( x80 & n7318 ) | ( x80 & ~n11507 ) | ( n7318 & ~n11507 ) ;
  assign n11509 = n11507 | n11508 ;
  assign n11510 = ~n11249 & n11509 ;
  assign n11511 = ( n11115 & n11249 ) | ( n11115 & ~n11510 ) | ( n11249 & ~n11510 ) ;
  assign n11512 = ~x80 & n10845 ;
  assign n11513 = x217 & ~n11512 ;
  assign n11514 = ( n10841 & n11511 ) | ( n10841 & ~n11513 ) | ( n11511 & ~n11513 ) ;
  assign n11515 = ~n10841 & n11514 ;
  assign n11516 = x81 & ~x314 ;
  assign n11517 = ~n1253 & n11516 ;
  assign n11518 = x68 & ~x81 ;
  assign n11519 = ~n1245 & n11518 ;
  assign n11520 = ( n9639 & ~n10086 ) | ( n9639 & n11519 ) | ( ~n10086 & n11519 ) ;
  assign n11521 = ~n9639 & n11520 ;
  assign n11522 = n1488 | n11521 ;
  assign n11523 = ( ~n1488 & n11517 ) | ( ~n1488 & n11522 ) | ( n11517 & n11522 ) ;
  assign n11524 = ( n7318 & ~n9935 ) | ( n7318 & n11523 ) | ( ~n9935 & n11523 ) ;
  assign n11525 = ~n7318 & n11524 ;
  assign n11526 = x66 & ~x73 ;
  assign n11527 = ( n1233 & ~n1247 ) | ( n1233 & n11526 ) | ( ~n1247 & n11526 ) ;
  assign n11528 = ~n1233 & n11527 ;
  assign n11529 = x69 & x314 ;
  assign n11530 = ( ~n1481 & n11528 ) | ( ~n1481 & n11529 ) | ( n11528 & n11529 ) ;
  assign n11531 = n11528 ^ n1481 ^ 1'b0 ;
  assign n11532 = ( n11528 & n11530 ) | ( n11528 & ~n11531 ) | ( n11530 & ~n11531 ) ;
  assign n11533 = ( n9732 & ~n9734 ) | ( n9732 & n11532 ) | ( ~n9734 & n11532 ) ;
  assign n11534 = ~n9732 & n11533 ;
  assign n11535 = n1263 | n9733 ;
  assign n11536 = n1372 | n11535 ;
  assign n11537 = n1245 | n1487 ;
  assign n11538 = x84 & ~n7755 ;
  assign n11539 = ~n11537 & n11538 ;
  assign n11540 = ~n1232 & n11539 ;
  assign n11541 = ~n11536 & n11540 ;
  assign n11542 = x314 & ~n11541 ;
  assign n11543 = n8761 | n11542 ;
  assign n11544 = x83 | n11539 ;
  assign n11545 = ( n1483 & ~n11536 ) | ( n1483 & n11544 ) | ( ~n11536 & n11544 ) ;
  assign n11546 = ~n1483 & n11545 ;
  assign n11547 = ( x314 & ~n11543 ) | ( x314 & n11546 ) | ( ~n11543 & n11546 ) ;
  assign n11548 = ~n11543 & n11547 ;
  assign n11549 = x211 & x299 ;
  assign n11550 = x219 & x299 ;
  assign n11551 = n11549 | n11550 ;
  assign n11552 = n9354 | n11551 ;
  assign n11553 = n7318 | n11552 ;
  assign n11554 = n10020 & ~n11553 ;
  assign n11555 = x314 | n9736 ;
  assign n11556 = n10080 & ~n11555 ;
  assign n11557 = n5219 & ~n9735 ;
  assign n11558 = ( ~n9732 & n11556 ) | ( ~n9732 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11559 = ~n9732 & n11558 ;
  assign n11560 = n6461 & n10031 ;
  assign n11561 = n6465 & n10034 ;
  assign n11562 = ( n9605 & n11560 ) | ( n9605 & n11561 ) | ( n11560 & n11561 ) ;
  assign n11563 = n11561 ^ n11560 ^ 1'b0 ;
  assign n11564 = ( n9605 & n11562 ) | ( n9605 & n11563 ) | ( n11562 & n11563 ) ;
  assign n11565 = n1534 & ~n11535 ;
  assign n11566 = x314 & ~n8761 ;
  assign n11567 = ~n1372 & n11566 ;
  assign n11568 = n11565 & n11567 ;
  assign n11569 = ~n1378 & n6425 ;
  assign n11570 = x1093 | n1290 ;
  assign n11571 = n2070 | n11570 ;
  assign n11572 = n11569 & ~n11571 ;
  assign n11573 = ( n1472 & n10095 ) | ( n1472 & n11572 ) | ( n10095 & n11572 ) ;
  assign n11574 = ~n1472 & n11573 ;
  assign n11575 = ( n6612 & n7318 ) | ( n6612 & ~n11574 ) | ( n7318 & ~n11574 ) ;
  assign n11576 = n11575 ^ n6612 ^ 1'b0 ;
  assign n11577 = ( n7318 & n11575 ) | ( n7318 & ~n11576 ) | ( n11575 & ~n11576 ) ;
  assign n11578 = n2070 | n8671 ;
  assign n11579 = n6425 & n9655 ;
  assign n11580 = x1093 | n11579 ;
  assign n11581 = n6380 | n10856 ;
  assign n11582 = n9652 & ~n11581 ;
  assign n11583 = n9666 & ~n10854 ;
  assign n11584 = n11582 & n11583 ;
  assign n11585 = x1093 & ~n11584 ;
  assign n11586 = ( n11578 & n11580 ) | ( n11578 & ~n11585 ) | ( n11580 & ~n11585 ) ;
  assign n11587 = ~n11578 & n11586 ;
  assign n11588 = ( n6612 & ~n11577 ) | ( n6612 & n11587 ) | ( ~n11577 & n11587 ) ;
  assign n11589 = ~n11577 & n11588 ;
  assign n11590 = n1229 | n7496 ;
  assign n11591 = ( n7511 & n8782 ) | ( n7511 & ~n11590 ) | ( n8782 & ~n11590 ) ;
  assign n11592 = ~n7511 & n11591 ;
  assign n11593 = x841 & ~n6387 ;
  assign n11594 = n11592 & n11593 ;
  assign n11595 = x70 | n11594 ;
  assign n11596 = ( n1291 & ~n8760 ) | ( n1291 & n11595 ) | ( ~n8760 & n11595 ) ;
  assign n11597 = ~n1291 & n11596 ;
  assign n11598 = ( x70 & n7452 ) | ( x70 & ~n11597 ) | ( n7452 & ~n11597 ) ;
  assign n11599 = n11598 ^ n11597 ^ 1'b0 ;
  assign n11600 = ( n11597 & ~n11598 ) | ( n11597 & n11599 ) | ( ~n11598 & n11599 ) ;
  assign n11601 = ~x1050 & n8132 ;
  assign n11602 = x90 | n11601 ;
  assign n11603 = ~n9963 & n11602 ;
  assign n11604 = ( n1440 & ~n6375 ) | ( n1440 & n11603 ) | ( ~n6375 & n11603 ) ;
  assign n11605 = ~n1440 & n11604 ;
  assign n11606 = x24 & ~n1412 ;
  assign n11607 = ( n1670 & ~n9713 ) | ( n1670 & n11606 ) | ( ~n9713 & n11606 ) ;
  assign n11608 = ~n1670 & n11607 ;
  assign n11609 = n1443 & n11608 ;
  assign n11610 = ~x58 & n1443 ;
  assign n11611 = n8753 | n11610 ;
  assign n11612 = n1670 & ~n8757 ;
  assign n11613 = n11611 & n11612 ;
  assign n11614 = ( x39 & ~n11609 ) | ( x39 & n11613 ) | ( ~n11609 & n11613 ) ;
  assign n11615 = n11609 | n11614 ;
  assign n11616 = ( n6471 & ~n8793 ) | ( n6471 & n11615 ) | ( ~n8793 & n11615 ) ;
  assign n11617 = ~n6471 & n11616 ;
  assign n11618 = ~n2290 & n5106 ;
  assign n11619 = n6461 & n11618 ;
  assign n11620 = n4736 & n5097 ;
  assign n11621 = n6465 & n11620 ;
  assign n11622 = n11619 | n11621 ;
  assign n11623 = ( n2096 & n9815 ) | ( n2096 & n11622 ) | ( n9815 & n11622 ) ;
  assign n11624 = ~n2096 & n11623 ;
  assign n11625 = x92 & ~n1292 ;
  assign n11626 = ~n2177 & n10118 ;
  assign n11627 = n11625 & n11626 ;
  assign n11628 = ( ~n8758 & n11624 ) | ( ~n8758 & n11627 ) | ( n11624 & n11627 ) ;
  assign n11629 = ~n8758 & n11628 ;
  assign n11630 = x1050 | n1292 ;
  assign n11631 = x92 & n11630 ;
  assign n11632 = x93 & ~n9713 ;
  assign n11633 = n1594 & n11632 ;
  assign n11634 = x92 | n11633 ;
  assign n11635 = ( n8759 & ~n11631 ) | ( n8759 & n11634 ) | ( ~n11631 & n11634 ) ;
  assign n11636 = ~n8759 & n11635 ;
  assign n11637 = n9694 & ~n9919 ;
  assign n11638 = n7457 | n11637 ;
  assign n11639 = n1395 | n8757 ;
  assign n11640 = ~n8815 & n9692 ;
  assign n11641 = n1466 | n11640 ;
  assign n11642 = ( x252 & n11639 ) | ( x252 & n11641 ) | ( n11639 & n11641 ) ;
  assign n11643 = ~n11639 & n11642 ;
  assign n11644 = n1615 & n11637 ;
  assign n11645 = x1093 & ~n11644 ;
  assign n11646 = ~n11643 & n11645 ;
  assign n11647 = ( n6442 & n11643 ) | ( n6442 & ~n11646 ) | ( n11643 & ~n11646 ) ;
  assign n11648 = x252 & ~n11647 ;
  assign n11649 = ~n7451 & n11647 ;
  assign n11650 = n11637 | n11649 ;
  assign n11651 = n7457 & ~n11650 ;
  assign n11652 = ( n7457 & n11648 ) | ( n7457 & n11651 ) | ( n11648 & n11651 ) ;
  assign n11653 = ( n8760 & n11638 ) | ( n8760 & ~n11652 ) | ( n11638 & ~n11652 ) ;
  assign n11654 = ~n8760 & n11653 ;
  assign n11655 = ~n1288 & n10397 ;
  assign n11656 = n10099 & n11655 ;
  assign n11657 = x332 | n8757 ;
  assign n11658 = n9918 | n11657 ;
  assign n11659 = n11592 & ~n11658 ;
  assign n11660 = ( x39 & ~n11656 ) | ( x39 & n11659 ) | ( ~n11656 & n11659 ) ;
  assign n11661 = n11656 | n11660 ;
  assign n11662 = n5115 & n5374 ;
  assign n11663 = n2291 | n10057 ;
  assign n11664 = n11662 & ~n11663 ;
  assign n11665 = ~n10052 & n10055 ;
  assign n11666 = n5374 & n11665 ;
  assign n11667 = ( x39 & n11664 ) | ( x39 & ~n11666 ) | ( n11664 & ~n11666 ) ;
  assign n11668 = ~n11664 & n11667 ;
  assign n11669 = ( n9901 & n11661 ) | ( n9901 & ~n11668 ) | ( n11661 & ~n11668 ) ;
  assign n11670 = ~n9901 & n11669 ;
  assign n11671 = x479 & ~n7451 ;
  assign n11672 = n1791 & n11671 ;
  assign n11673 = x96 & ~n1274 ;
  assign n11674 = ~n1410 & n11673 ;
  assign n11675 = n1596 & ~n11671 ;
  assign n11676 = n11674 & n11675 ;
  assign n11677 = ( ~x95 & n11672 ) | ( ~x95 & n11676 ) | ( n11672 & n11676 ) ;
  assign n11678 = ~x95 & n11677 ;
  assign n11679 = ~n8929 & n11655 ;
  assign n11680 = ( ~n8760 & n11678 ) | ( ~n8760 & n11679 ) | ( n11678 & n11679 ) ;
  assign n11681 = ~n8760 & n11680 ;
  assign n11682 = x96 | n8764 ;
  assign n11683 = n5165 & n11671 ;
  assign n11684 = n5023 | n11683 ;
  assign n11685 = ( n10124 & n11682 ) | ( n10124 & n11684 ) | ( n11682 & n11684 ) ;
  assign n11686 = ~n11682 & n11685 ;
  assign n11687 = x39 & x593 ;
  assign n11688 = ( ~n5374 & n10060 ) | ( ~n5374 & n11687 ) | ( n10060 & n11687 ) ;
  assign n11689 = n5374 & n11688 ;
  assign n11690 = ( ~n9901 & n11686 ) | ( ~n9901 & n11689 ) | ( n11686 & n11689 ) ;
  assign n11691 = ~n9901 & n11690 ;
  assign n11692 = ~x92 & n10119 ;
  assign n11693 = n11625 | n11692 ;
  assign n11694 = x314 & x1050 ;
  assign n11695 = ( n8759 & n11693 ) | ( n8759 & n11694 ) | ( n11693 & n11694 ) ;
  assign n11696 = ~n8759 & n11695 ;
  assign n11697 = ~x72 & x174 ;
  assign n11698 = ( x299 & n8906 ) | ( x299 & n11697 ) | ( n8906 & n11697 ) ;
  assign n11699 = ~x299 & n11698 ;
  assign n11700 = ~x72 & x152 ;
  assign n11701 = n8899 & n11700 ;
  assign n11702 = n11699 ^ x299 ^ 1'b0 ;
  assign n11703 = ( ~x299 & n11701 ) | ( ~x299 & n11702 ) | ( n11701 & n11702 ) ;
  assign n11704 = ( x299 & n11699 ) | ( x299 & n11703 ) | ( n11699 & n11703 ) ;
  assign n11705 = x232 & n11704 ;
  assign n11706 = x39 & ~n11705 ;
  assign n11707 = ~x72 & x99 ;
  assign n11708 = x39 | n11707 ;
  assign n11709 = ~n11706 & n11708 ;
  assign n11710 = n2052 & n11709 ;
  assign n11711 = n6824 | n11707 ;
  assign n11712 = ~n1615 & n11707 ;
  assign n11713 = ~n8934 & n11707 ;
  assign n11714 = ~n5027 & n9539 ;
  assign n11715 = ( n9068 & n11713 ) | ( n9068 & n11714 ) | ( n11713 & n11714 ) ;
  assign n11716 = n11714 ^ n11713 ^ 1'b0 ;
  assign n11717 = ( n9068 & n11715 ) | ( n9068 & n11716 ) | ( n11715 & n11716 ) ;
  assign n11718 = ( n6824 & n11712 ) | ( n6824 & ~n11717 ) | ( n11712 & ~n11717 ) ;
  assign n11719 = ~n11712 & n11718 ;
  assign n11720 = ( x39 & n11711 ) | ( x39 & ~n11719 ) | ( n11711 & ~n11719 ) ;
  assign n11721 = n11720 ^ n11711 ^ 1'b0 ;
  assign n11722 = ( x39 & n11720 ) | ( x39 & ~n11721 ) | ( n11720 & ~n11721 ) ;
  assign n11723 = ( n2052 & ~n11706 ) | ( n2052 & n11722 ) | ( ~n11706 & n11722 ) ;
  assign n11724 = ~n2052 & n11723 ;
  assign n11725 = ( x75 & n11710 ) | ( x75 & ~n11724 ) | ( n11710 & ~n11724 ) ;
  assign n11726 = ~n11710 & n11725 ;
  assign n11727 = x228 & ~n8950 ;
  assign n11728 = n11707 & ~n11727 ;
  assign n11729 = x228 & ~n9096 ;
  assign n11730 = ( n2095 & ~n11728 ) | ( n2095 & n11729 ) | ( ~n11728 & n11729 ) ;
  assign n11731 = n11728 | n11730 ;
  assign n11732 = n11731 ^ x75 ^ 1'b0 ;
  assign n11733 = n2095 & ~n11709 ;
  assign n11734 = x87 & ~n11733 ;
  assign n11735 = ( n11731 & ~n11732 ) | ( n11731 & n11734 ) | ( ~n11732 & n11734 ) ;
  assign n11736 = ( x75 & n11732 ) | ( x75 & n11735 ) | ( n11732 & n11735 ) ;
  assign n11737 = n6824 & ~n11712 ;
  assign n11738 = n11711 & ~n11737 ;
  assign n11739 = ~n5026 & n8921 ;
  assign n11740 = ~n9066 & n11707 ;
  assign n11741 = n11739 | n11740 ;
  assign n11742 = n9068 & n11741 ;
  assign n11743 = ( n11711 & n11738 ) | ( n11711 & n11742 ) | ( n11738 & n11742 ) ;
  assign n11744 = x39 | n11743 ;
  assign n11745 = ~n11706 & n11744 ;
  assign n11746 = ( x38 & x100 ) | ( x38 & ~n11745 ) | ( x100 & ~n11745 ) ;
  assign n11747 = ~x38 & n11746 ;
  assign n11748 = ( x99 & n8924 ) | ( x99 & n11707 ) | ( n8924 & n11707 ) ;
  assign n11751 = ~n9056 & n11748 ;
  assign n11752 = n9384 & ~n11751 ;
  assign n11749 = ~n9027 & n11748 ;
  assign n11750 = n9385 | n11749 ;
  assign n11753 = n11752 ^ n11750 ^ 1'b0 ;
  assign n11754 = ( x228 & ~n11750 ) | ( x228 & n11752 ) | ( ~n11750 & n11752 ) ;
  assign n11755 = ( x228 & ~n11753 ) | ( x228 & n11754 ) | ( ~n11753 & n11754 ) ;
  assign n11756 = ~n9004 & n11748 ;
  assign n11757 = x228 | n9138 ;
  assign n11758 = n11756 | n11757 ;
  assign n11759 = ( x39 & ~n11755 ) | ( x39 & n11758 ) | ( ~n11755 & n11758 ) ;
  assign n11760 = ~x39 & n11759 ;
  assign n11761 = n8901 & n11704 ;
  assign n11762 = ~n9575 & n11761 ;
  assign n11763 = ( n1205 & ~n11760 ) | ( n1205 & n11762 ) | ( ~n11760 & n11762 ) ;
  assign n11764 = n11760 | n11763 ;
  assign n11765 = x38 & ~n11709 ;
  assign n11766 = x87 | n11765 ;
  assign n11767 = ( n11747 & n11764 ) | ( n11747 & ~n11766 ) | ( n11764 & ~n11766 ) ;
  assign n11768 = ~n11747 & n11767 ;
  assign n11769 = ( ~n11726 & n11736 ) | ( ~n11726 & n11768 ) | ( n11736 & n11768 ) ;
  assign n11770 = ~n11726 & n11769 ;
  assign n11771 = ( x74 & n5015 ) | ( x74 & ~n11770 ) | ( n5015 & ~n11770 ) ;
  assign n11772 = n11770 | n11771 ;
  assign n11773 = x232 & n11701 ;
  assign n11774 = x39 & ~n11773 ;
  assign n11775 = ( n7318 & n11708 ) | ( n7318 & n11774 ) | ( n11708 & n11774 ) ;
  assign n11776 = ~n11774 & n11775 ;
  assign n11777 = n6782 & ~n11709 ;
  assign n11778 = n7318 | n11777 ;
  assign n11779 = ~n11776 & n11778 ;
  assign n11780 = ( n11772 & n11776 ) | ( n11772 & ~n11779 ) | ( n11776 & ~n11779 ) ;
  assign n11781 = ~x24 & n7461 ;
  assign n11782 = n7451 & ~n7458 ;
  assign n11783 = n11781 & n11782 ;
  assign n11784 = n5037 & n5044 ;
  assign n11785 = x129 & ~n8675 ;
  assign n11786 = ~n11784 & n11785 ;
  assign n11787 = ( n5043 & n11784 ) | ( n5043 & ~n11786 ) | ( n11784 & ~n11786 ) ;
  assign n11788 = ( x129 & n6411 ) | ( x129 & n11785 ) | ( n6411 & n11785 ) ;
  assign n11789 = ( n5040 & ~n11787 ) | ( n5040 & n11788 ) | ( ~n11787 & n11788 ) ;
  assign n11790 = ~n11787 & n11789 ;
  assign n11791 = x75 | n1206 ;
  assign n11792 = n5018 & ~n11791 ;
  assign n11793 = ( n11783 & ~n11790 ) | ( n11783 & n11792 ) | ( ~n11790 & n11792 ) ;
  assign n11794 = n11790 ^ n11783 ^ 1'b0 ;
  assign n11795 = ( n11783 & n11793 ) | ( n11783 & ~n11794 ) | ( n11793 & ~n11794 ) ;
  assign n11796 = ( n1292 & ~n10138 ) | ( n1292 & n11795 ) | ( ~n10138 & n11795 ) ;
  assign n11797 = ~n1292 & n11796 ;
  assign n11798 = n10218 ^ n8906 ^ n8905 ;
  assign n11799 = ~x72 & n11798 ;
  assign n11800 = x299 | n11799 ;
  assign n11801 = n10150 ^ n8899 ^ n8898 ;
  assign n11802 = ~x72 & n11801 ;
  assign n11803 = ( x232 & n9323 ) | ( x232 & n11802 ) | ( n9323 & n11802 ) ;
  assign n11804 = x39 & ~n11803 ;
  assign n11805 = ( x39 & ~n11800 ) | ( x39 & n11804 ) | ( ~n11800 & n11804 ) ;
  assign n11806 = x39 | n8927 ;
  assign n11807 = ~n11805 & n11806 ;
  assign n11808 = n2052 & n11807 ;
  assign n11809 = n6824 | n8927 ;
  assign n11810 = ~n1615 & n8927 ;
  assign n11811 = n6824 & ~n11810 ;
  assign n11812 = n1615 & n5034 ;
  assign n11813 = n8927 & ~n8933 ;
  assign n11814 = n8922 | n11813 ;
  assign n11815 = n11811 & ~n11814 ;
  assign n11816 = ( n11811 & ~n11812 ) | ( n11811 & n11815 ) | ( ~n11812 & n11815 ) ;
  assign n11817 = ( x39 & n11809 ) | ( x39 & ~n11816 ) | ( n11809 & ~n11816 ) ;
  assign n11818 = n11817 ^ n11809 ^ 1'b0 ;
  assign n11819 = ( x39 & n11817 ) | ( x39 & ~n11818 ) | ( n11817 & ~n11818 ) ;
  assign n11820 = ( n2052 & ~n11805 ) | ( n2052 & n11819 ) | ( ~n11805 & n11819 ) ;
  assign n11821 = ~n2052 & n11820 ;
  assign n11822 = ( x75 & n11808 ) | ( x75 & ~n11821 ) | ( n11808 & ~n11821 ) ;
  assign n11823 = ~n11808 & n11822 ;
  assign n11824 = ~x101 & n9553 ;
  assign n11825 = ~n8949 & n9550 ;
  assign n11826 = n8927 & ~n11825 ;
  assign n11827 = ( x39 & ~n11824 ) | ( x39 & n11826 ) | ( ~n11824 & n11826 ) ;
  assign n11828 = n11824 | n11827 ;
  assign n11829 = n11828 ^ x75 ^ 1'b0 ;
  assign n11830 = x87 & ~n11805 ;
  assign n11831 = ( n11828 & ~n11829 ) | ( n11828 & n11830 ) | ( ~n11829 & n11830 ) ;
  assign n11832 = ( x75 & n11829 ) | ( x75 & n11831 ) | ( n11829 & n11831 ) ;
  assign n11833 = x38 & ~n11807 ;
  assign n11834 = x87 | n11833 ;
  assign n11837 = n1615 & ~n9047 ;
  assign n11838 = ~n9055 & n11837 ;
  assign n11835 = n1615 | n9013 ;
  assign n11836 = n9026 | n11835 ;
  assign n11839 = n11838 ^ n11836 ^ 1'b0 ;
  assign n11840 = ( x228 & ~n11836 ) | ( x228 & n11838 ) | ( ~n11836 & n11838 ) ;
  assign n11841 = ( x228 & ~n11839 ) | ( x228 & n11840 ) | ( ~n11839 & n11840 ) ;
  assign n11842 = x228 | n8994 ;
  assign n11843 = n9003 | n11842 ;
  assign n11844 = ( x39 & ~n11841 ) | ( x39 & n11843 ) | ( ~n11841 & n11843 ) ;
  assign n11845 = ~x39 & n11844 ;
  assign n11846 = ~n9576 & n11801 ;
  assign n11847 = x299 & ~n11846 ;
  assign n11848 = ~n9576 & n11798 ;
  assign n11849 = x299 | n11848 ;
  assign n11850 = ( n8901 & n11847 ) | ( n8901 & n11849 ) | ( n11847 & n11849 ) ;
  assign n11851 = ~n11847 & n11850 ;
  assign n11852 = ( n1205 & ~n11845 ) | ( n1205 & n11851 ) | ( ~n11845 & n11851 ) ;
  assign n11853 = n11845 | n11852 ;
  assign n11854 = n11809 & ~n11811 ;
  assign n11855 = ~x44 & n9582 ;
  assign n11856 = n8927 & ~n11855 ;
  assign n11857 = ( n8921 & n11812 ) | ( n8921 & n11856 ) | ( n11812 & n11856 ) ;
  assign n11858 = n11812 & n11857 ;
  assign n11859 = ( n11809 & n11854 ) | ( n11809 & n11858 ) | ( n11854 & n11858 ) ;
  assign n11860 = x39 | n11859 ;
  assign n11861 = ~n11805 & n11860 ;
  assign n11862 = ( x38 & x100 ) | ( x38 & ~n11861 ) | ( x100 & ~n11861 ) ;
  assign n11863 = ~x38 & n11862 ;
  assign n11864 = ( n11834 & n11853 ) | ( n11834 & ~n11863 ) | ( n11853 & ~n11863 ) ;
  assign n11865 = ~n11834 & n11864 ;
  assign n11866 = ( ~n11823 & n11832 ) | ( ~n11823 & n11865 ) | ( n11832 & n11865 ) ;
  assign n11867 = ~n11823 & n11866 ;
  assign n11868 = ( x74 & n5015 ) | ( x74 & ~n11867 ) | ( n5015 & ~n11867 ) ;
  assign n11869 = n11867 | n11868 ;
  assign n11870 = x232 & n11802 ;
  assign n11871 = x39 & ~n11870 ;
  assign n11872 = ( n7318 & n11806 ) | ( n7318 & n11871 ) | ( n11806 & n11871 ) ;
  assign n11873 = ~n11871 & n11872 ;
  assign n11874 = n6782 & ~n11807 ;
  assign n11875 = n7318 | n11874 ;
  assign n11876 = ~n11873 & n11875 ;
  assign n11877 = ( n11869 & n11873 ) | ( n11869 & ~n11876 ) | ( n11873 & ~n11876 ) ;
  assign n11878 = n7318 | n9935 ;
  assign n11879 = n1546 & ~n7497 ;
  assign n11880 = ~n11878 & n11879 ;
  assign n11881 = x109 & ~n1452 ;
  assign n11882 = ~n1369 & n11881 ;
  assign n11883 = ( x314 & n9731 ) | ( x314 & ~n11882 ) | ( n9731 & ~n11882 ) ;
  assign n11884 = n11882 ^ n9731 ^ 1'b0 ;
  assign n11885 = ( n9731 & n11883 ) | ( n9731 & ~n11884 ) | ( n11883 & ~n11884 ) ;
  assign n11886 = ( ~n5206 & n11565 ) | ( ~n5206 & n11882 ) | ( n11565 & n11882 ) ;
  assign n11887 = ( x314 & ~n11885 ) | ( x314 & n11886 ) | ( ~n11885 & n11886 ) ;
  assign n11888 = ~n11885 & n11887 ;
  assign n11889 = n6612 | n7457 ;
  assign n11890 = n8967 & ~n11889 ;
  assign n11891 = ( ~n8672 & n8967 ) | ( ~n8672 & n11890 ) | ( n8967 & n11890 ) ;
  assign n11892 = n6611 ^ x288 ^ 1'b0 ;
  assign n11893 = ( x288 & n6611 ) | ( x288 & ~n11892 ) | ( n6611 & ~n11892 ) ;
  assign n11894 = n6412 | n8671 ;
  assign n11895 = ~x47 & n9666 ;
  assign n11896 = x110 | n11582 ;
  assign n11897 = ( n8972 & n11895 ) | ( n8972 & n11896 ) | ( n11895 & n11896 ) ;
  assign n11898 = ~n8972 & n11897 ;
  assign n11899 = n5035 | n11898 ;
  assign n11900 = n5035 & ~n11584 ;
  assign n11901 = ( n11894 & n11899 ) | ( n11894 & ~n11900 ) | ( n11899 & ~n11900 ) ;
  assign n11902 = ~n11894 & n11901 ;
  assign n11903 = n11902 ^ n11898 ^ 1'b0 ;
  assign n11904 = n6412 & ~n8671 ;
  assign n11905 = ( n11898 & ~n11903 ) | ( n11898 & n11904 ) | ( ~n11903 & n11904 ) ;
  assign n11906 = ( n11902 & n11903 ) | ( n11902 & n11905 ) | ( n11903 & n11905 ) ;
  assign n11907 = ( n11892 & n11893 ) | ( n11892 & n11906 ) | ( n11893 & n11906 ) ;
  assign n11908 = ( ~n8760 & n11891 ) | ( ~n8760 & n11907 ) | ( n11891 & n11907 ) ;
  assign n11909 = ~n8760 & n11908 ;
  assign n11910 = x24 & n9917 ;
  assign n11911 = x53 | n9916 ;
  assign n11912 = ~n1390 & n11911 ;
  assign n11913 = x24 | n1395 ;
  assign n11914 = n11912 & ~n11913 ;
  assign n11915 = ( x841 & n11910 ) | ( x841 & n11914 ) | ( n11910 & n11914 ) ;
  assign n11916 = n11914 ^ n11910 ^ 1'b0 ;
  assign n11917 = ( x841 & n11915 ) | ( x841 & n11916 ) | ( n11915 & n11916 ) ;
  assign n11918 = ~n7477 & n9898 ;
  assign n11919 = ( ~n8761 & n11917 ) | ( ~n8761 & n11918 ) | ( n11917 & n11918 ) ;
  assign n11920 = ~n8761 & n11919 ;
  assign n11921 = x999 | n8761 ;
  assign n11922 = n9988 & ~n11921 ;
  assign n11923 = n2036 | n6423 ;
  assign n11924 = ( ~x97 & x108 ) | ( ~x97 & n6385 ) | ( x108 & n6385 ) ;
  assign n11925 = ( n1371 & ~n8813 ) | ( n1371 & n11924 ) | ( ~n8813 & n11924 ) ;
  assign n11926 = ~n1371 & n11925 ;
  assign n11927 = ~n6388 & n8824 ;
  assign n11928 = n11926 & n11927 ;
  assign n11929 = n6388 | n8824 ;
  assign n11930 = x314 & ~n6386 ;
  assign n11931 = n11929 | n11930 ;
  assign n11932 = ( x314 & n11926 ) | ( x314 & ~n11931 ) | ( n11926 & ~n11931 ) ;
  assign n11933 = ~n11931 & n11932 ;
  assign n11934 = ( x51 & ~n11928 ) | ( x51 & n11933 ) | ( ~n11928 & n11933 ) ;
  assign n11935 = n11928 | n11934 ;
  assign n11936 = n11935 ^ n11923 ^ 1'b0 ;
  assign n11937 = ( n11923 & n11935 ) | ( n11923 & n11936 ) | ( n11935 & n11936 ) ;
  assign n11938 = ( x87 & ~n11923 ) | ( x87 & n11937 ) | ( ~n11923 & n11937 ) ;
  assign n11939 = ( n5014 & ~n10138 ) | ( n5014 & n11938 ) | ( ~n10138 & n11938 ) ;
  assign n11940 = ~n5014 & n11939 ;
  assign n11941 = n1470 & ~n10084 ;
  assign n11942 = n11566 & n11941 ;
  assign n11943 = n7457 & n8672 ;
  assign n11944 = n8966 & n11943 ;
  assign n11945 = x82 | x109 ;
  assign n11946 = x111 & ~n11945 ;
  assign n11947 = ( n1263 & ~n10854 ) | ( n1263 & n11946 ) | ( ~n10854 & n11946 ) ;
  assign n11948 = ~n1263 & n11947 ;
  assign n11949 = ( n1518 & ~n9736 ) | ( n1518 & n11948 ) | ( ~n9736 & n11948 ) ;
  assign n11950 = ~n1518 & n11949 ;
  assign n11951 = x314 & n11950 ;
  assign n11952 = ( ~n8761 & n11944 ) | ( ~n8761 & n11951 ) | ( n11944 & n11951 ) ;
  assign n11953 = ~n8761 & n11952 ;
  assign n11954 = ~x314 & n11950 ;
  assign n11955 = ~n7786 & n11954 ;
  assign n11956 = x72 & ~n8929 ;
  assign n11957 = n11955 | n11956 ;
  assign n11958 = ( n5203 & ~n8760 ) | ( n5203 & n11957 ) | ( ~n8760 & n11957 ) ;
  assign n11959 = ~n5203 & n11958 ;
  assign n11960 = x124 & ~x468 ;
  assign n11961 = ~x39 & n9132 ;
  assign n11962 = n2052 & n11961 ;
  assign n11963 = n1615 & n6824 ;
  assign n11964 = n9132 & ~n11963 ;
  assign n11965 = n5033 & ~n9214 ;
  assign n11966 = ( n9132 & n11964 ) | ( n9132 & n11965 ) | ( n11964 & n11965 ) ;
  assign n11967 = n5033 & n11963 ;
  assign n11968 = ~x113 & n11967 ;
  assign n11969 = n11739 & n11968 ;
  assign n11970 = n6414 & n11969 ;
  assign n11971 = ( ~n1207 & n11966 ) | ( ~n1207 & n11970 ) | ( n11966 & n11970 ) ;
  assign n11972 = ~n1207 & n11971 ;
  assign n11973 = ( x75 & n11962 ) | ( x75 & ~n11972 ) | ( n11962 & ~n11972 ) ;
  assign n11974 = ~n11962 & n11973 ;
  assign n11975 = n1205 & n11961 ;
  assign n11976 = n9132 & ~n9202 ;
  assign n11977 = ~x113 & n11729 ;
  assign n11978 = ( ~n2095 & n11976 ) | ( ~n2095 & n11977 ) | ( n11976 & n11977 ) ;
  assign n11979 = ~n2095 & n11978 ;
  assign n11980 = ( x87 & n11975 ) | ( x87 & ~n11979 ) | ( n11975 & ~n11979 ) ;
  assign n11981 = ~n11975 & n11980 ;
  assign n11982 = n6480 & ~n9102 ;
  assign n11983 = n5033 & ~n11982 ;
  assign n11984 = ( n9132 & n11964 ) | ( n9132 & n11983 ) | ( n11964 & n11983 ) ;
  assign n11985 = ( ~x39 & n11969 ) | ( ~x39 & n11984 ) | ( n11969 & n11984 ) ;
  assign n11986 = ~x39 & n11985 ;
  assign n11987 = ( x38 & x100 ) | ( x38 & ~n11986 ) | ( x100 & ~n11986 ) ;
  assign n11988 = ~x38 & n11987 ;
  assign n11989 = n11961 & ~n11988 ;
  assign n11990 = ( x38 & n11988 ) | ( x38 & ~n11989 ) | ( n11988 & ~n11989 ) ;
  assign n11991 = x228 | n9139 ;
  assign n11992 = n9131 | n11991 ;
  assign n11993 = n1615 | n9027 ;
  assign n11994 = ( x99 & ~n9057 ) | ( x99 & n11993 ) | ( ~n9057 & n11993 ) ;
  assign n11995 = ~x99 & n11994 ;
  assign n11996 = ( x113 & n9128 ) | ( x113 & ~n11995 ) | ( n9128 & ~n11995 ) ;
  assign n11997 = ~n9128 & n11996 ;
  assign n11998 = ~x113 & n9386 ;
  assign n11999 = ( x228 & n11997 ) | ( x228 & ~n11998 ) | ( n11997 & ~n11998 ) ;
  assign n12000 = ~n11997 & n11999 ;
  assign n12001 = ( x39 & n11992 ) | ( x39 & ~n12000 ) | ( n11992 & ~n12000 ) ;
  assign n12002 = ~x39 & n12001 ;
  assign n12003 = ( n1205 & ~n11990 ) | ( n1205 & n12002 ) | ( ~n11990 & n12002 ) ;
  assign n12004 = ~n11990 & n12003 ;
  assign n12005 = ( x87 & ~n11981 ) | ( x87 & n12004 ) | ( ~n11981 & n12004 ) ;
  assign n12006 = ~n11981 & n12005 ;
  assign n12007 = ( x75 & ~n11974 ) | ( x75 & n12006 ) | ( ~n11974 & n12006 ) ;
  assign n12008 = ~n11974 & n12007 ;
  assign n12009 = n11961 ^ n10138 ^ 1'b0 ;
  assign n12010 = ( n11961 & n12008 ) | ( n11961 & ~n12009 ) | ( n12008 & ~n12009 ) ;
  assign n12011 = ~x72 & x114 ;
  assign n12012 = ~x39 & n12011 ;
  assign n12013 = n9109 | n12011 ;
  assign n12014 = x114 & ~n9426 ;
  assign n12015 = ( n9109 & n9218 ) | ( n9109 & ~n12014 ) | ( n9218 & ~n12014 ) ;
  assign n12016 = ~n9218 & n12015 ;
  assign n12017 = ( n1207 & n12013 ) | ( n1207 & ~n12016 ) | ( n12013 & ~n12016 ) ;
  assign n12018 = ~n1207 & n12017 ;
  assign n12019 = n2052 & n12012 ;
  assign n12020 = ( x75 & n12018 ) | ( x75 & ~n12019 ) | ( n12018 & ~n12019 ) ;
  assign n12021 = ~n12018 & n12020 ;
  assign n12022 = x114 & ~n9105 ;
  assign n12023 = ( n9100 & n9109 ) | ( n9100 & ~n12022 ) | ( n9109 & ~n12022 ) ;
  assign n12024 = ~n9100 & n12023 ;
  assign n12025 = ~x39 & n12013 ;
  assign n12026 = n5018 & ~n12025 ;
  assign n12027 = ( n5018 & n12024 ) | ( n5018 & n12026 ) | ( n12024 & n12026 ) ;
  assign n12028 = x38 & ~n12012 ;
  assign n12029 = ( x87 & ~n12027 ) | ( x87 & n12028 ) | ( ~n12027 & n12028 ) ;
  assign n12030 = n12027 | n12029 ;
  assign n12031 = x115 & ~n12011 ;
  assign n12032 = x39 | n12031 ;
  assign n12033 = n9389 ^ x114 ^ 1'b0 ;
  assign n12034 = ( n9389 & ~n9395 ) | ( n9389 & n12033 ) | ( ~n9395 & n12033 ) ;
  assign n12035 = ( x115 & ~n12032 ) | ( x115 & n12034 ) | ( ~n12032 & n12034 ) ;
  assign n12036 = ~n12032 & n12035 ;
  assign n12037 = ( n1205 & ~n12030 ) | ( n1205 & n12036 ) | ( ~n12030 & n12036 ) ;
  assign n12038 = ~n12030 & n12037 ;
  assign n12039 = x228 & ~n9103 ;
  assign n12040 = ~x115 & n12039 ;
  assign n12041 = n12011 & ~n12040 ;
  assign n12042 = ( n1205 & n9200 ) | ( n1205 & ~n12041 ) | ( n9200 & ~n12041 ) ;
  assign n12043 = n12041 | n12042 ;
  assign n12044 = n12043 ^ x75 ^ 1'b0 ;
  assign n12045 = n1205 & ~n12012 ;
  assign n12046 = n9816 & ~n12045 ;
  assign n12047 = ( n12043 & ~n12044 ) | ( n12043 & n12046 ) | ( ~n12044 & n12046 ) ;
  assign n12048 = ( x75 & n12044 ) | ( x75 & n12047 ) | ( n12044 & n12047 ) ;
  assign n12049 = ( ~n12021 & n12038 ) | ( ~n12021 & n12048 ) | ( n12038 & n12048 ) ;
  assign n12050 = ~n12021 & n12049 ;
  assign n12051 = n12012 ^ n10138 ^ 1'b0 ;
  assign n12052 = ( n12012 & n12050 ) | ( n12012 & ~n12051 ) | ( n12050 & ~n12051 ) ;
  assign n12053 = ~x72 & x115 ;
  assign n12054 = ~x39 & n12053 ;
  assign n12055 = n2052 & n12054 ;
  assign n12056 = x52 | n9791 ;
  assign n12057 = ( x115 & n9098 ) | ( x115 & n12056 ) | ( n9098 & n12056 ) ;
  assign n12058 = ~x115 & n12057 ;
  assign n12059 = n6414 & n12058 ;
  assign n12060 = x115 & ~n9426 ;
  assign n12061 = ( n11963 & n12059 ) | ( n11963 & ~n12060 ) | ( n12059 & ~n12060 ) ;
  assign n12062 = ~n12059 & n12061 ;
  assign n12063 = n11963 | n12053 ;
  assign n12064 = ( n1207 & ~n12062 ) | ( n1207 & n12063 ) | ( ~n12062 & n12063 ) ;
  assign n12065 = ~n1207 & n12064 ;
  assign n12066 = ( x75 & n12055 ) | ( x75 & ~n12065 ) | ( n12055 & ~n12065 ) ;
  assign n12067 = ~n12055 & n12066 ;
  assign n12068 = x115 & ~n9105 ;
  assign n12069 = ( n11963 & n12058 ) | ( n11963 & ~n12068 ) | ( n12058 & ~n12068 ) ;
  assign n12070 = ~n12058 & n12069 ;
  assign n12071 = ~x39 & n12063 ;
  assign n12072 = n5018 & ~n12071 ;
  assign n12073 = ( n5018 & n12070 ) | ( n5018 & n12072 ) | ( n12070 & n12072 ) ;
  assign n12074 = x38 & ~n12054 ;
  assign n12075 = ( x87 & ~n12073 ) | ( x87 & n12074 ) | ( ~n12073 & n12074 ) ;
  assign n12076 = n12073 | n12075 ;
  assign n12077 = x115 | n9389 ;
  assign n12078 = x115 & n9395 ;
  assign n12079 = ( x39 & n12077 ) | ( x39 & ~n12078 ) | ( n12077 & ~n12078 ) ;
  assign n12080 = ~x39 & n12079 ;
  assign n12081 = ( n1205 & ~n12076 ) | ( n1205 & n12080 ) | ( ~n12076 & n12080 ) ;
  assign n12082 = ~n12076 & n12081 ;
  assign n12083 = ~n12039 & n12053 ;
  assign n12084 = ( n1205 & n9199 ) | ( n1205 & ~n12083 ) | ( n9199 & ~n12083 ) ;
  assign n12085 = n12083 | n12084 ;
  assign n12086 = n12085 ^ x75 ^ 1'b0 ;
  assign n12087 = n1205 & ~n12054 ;
  assign n12088 = n9816 & ~n12087 ;
  assign n12089 = ( n12085 & ~n12086 ) | ( n12085 & n12088 ) | ( ~n12086 & n12088 ) ;
  assign n12090 = ( x75 & n12086 ) | ( x75 & n12089 ) | ( n12086 & n12089 ) ;
  assign n12091 = ( ~n12067 & n12082 ) | ( ~n12067 & n12090 ) | ( n12082 & n12090 ) ;
  assign n12092 = ~n12067 & n12091 ;
  assign n12093 = n12054 ^ n10138 ^ 1'b0 ;
  assign n12094 = ( n12054 & n12092 ) | ( n12054 & ~n12093 ) | ( n12092 & ~n12093 ) ;
  assign n12095 = ~x39 & n9135 ;
  assign n12096 = n2052 & n12095 ;
  assign n12097 = n9135 & ~n11963 ;
  assign n12098 = n9135 & ~n9215 ;
  assign n12099 = ( n9424 & n11967 ) | ( n9424 & n12098 ) | ( n11967 & n12098 ) ;
  assign n12100 = n11967 & n12099 ;
  assign n12101 = ( ~n1207 & n12097 ) | ( ~n1207 & n12100 ) | ( n12097 & n12100 ) ;
  assign n12102 = ~n1207 & n12101 ;
  assign n12103 = ( x75 & n12096 ) | ( x75 & ~n12102 ) | ( n12096 & ~n12102 ) ;
  assign n12104 = ~n12096 & n12103 ;
  assign n12105 = x38 & ~n12095 ;
  assign n12106 = x87 | n12105 ;
  assign n12107 = ~x113 & n11982 ;
  assign n12108 = n9135 & ~n12107 ;
  assign n12109 = ( n9098 & n11967 ) | ( n9098 & n12108 ) | ( n11967 & n12108 ) ;
  assign n12110 = n11967 & n12109 ;
  assign n12111 = ( ~x39 & n12097 ) | ( ~x39 & n12110 ) | ( n12097 & n12110 ) ;
  assign n12112 = ~x39 & n12111 ;
  assign n12113 = ~n12106 & n12112 ;
  assign n12114 = ( n5018 & n12106 ) | ( n5018 & ~n12113 ) | ( n12106 & ~n12113 ) ;
  assign n12115 = x228 | n9140 ;
  assign n12116 = n9134 | n12115 ;
  assign n12117 = n1615 & n9154 ;
  assign n12118 = x116 & ~n12117 ;
  assign n12119 = n9149 | n12118 ;
  assign n12120 = n9170 ^ n1615 ^ 1'b0 ;
  assign n12121 = ( n1615 & n9170 ) | ( n1615 & ~n12120 ) | ( n9170 & ~n12120 ) ;
  assign n12122 = ( n12119 & n12120 ) | ( n12119 & n12121 ) | ( n12120 & n12121 ) ;
  assign n12123 = ~n1615 & n9163 ;
  assign n12124 = ( x228 & n12122 ) | ( x228 & ~n12123 ) | ( n12122 & ~n12123 ) ;
  assign n12125 = ~n12122 & n12124 ;
  assign n12126 = ( x39 & n12116 ) | ( x39 & ~n12125 ) | ( n12116 & ~n12125 ) ;
  assign n12127 = ~x39 & n12126 ;
  assign n12128 = ( n1205 & ~n12114 ) | ( n1205 & n12127 ) | ( ~n12114 & n12127 ) ;
  assign n12129 = ~n12114 & n12128 ;
  assign n12130 = ~x113 & n9202 ;
  assign n12131 = n9135 & ~n12130 ;
  assign n12132 = ( x38 & n9198 ) | ( x38 & ~n12131 ) | ( n9198 & ~n12131 ) ;
  assign n12133 = n12131 | n12132 ;
  assign n12134 = n12133 ^ n12105 ^ 1'b0 ;
  assign n12135 = ( n12105 & n12133 ) | ( n12105 & n12134 ) | ( n12133 & n12134 ) ;
  assign n12136 = ( x100 & ~n12105 ) | ( x100 & n12135 ) | ( ~n12105 & n12135 ) ;
  assign n12137 = n12136 ^ x75 ^ 1'b0 ;
  assign n12138 = x100 & ~n12095 ;
  assign n12139 = n9816 & ~n12138 ;
  assign n12140 = ( n12136 & ~n12137 ) | ( n12136 & n12139 ) | ( ~n12137 & n12139 ) ;
  assign n12141 = ( x75 & n12137 ) | ( x75 & n12140 ) | ( n12137 & n12140 ) ;
  assign n12142 = ( ~n12104 & n12129 ) | ( ~n12104 & n12141 ) | ( n12129 & n12141 ) ;
  assign n12143 = ~n12104 & n12142 ;
  assign n12144 = n12095 ^ n10138 ^ 1'b0 ;
  assign n12145 = ( n12095 & n12143 ) | ( n12095 & ~n12144 ) | ( n12143 & ~n12144 ) ;
  assign n12146 = x54 | n6257 ;
  assign n12147 = x74 | n12146 ;
  assign n12148 = n2509 & ~n6312 ;
  assign n12149 = n2508 | n12148 ;
  assign n12150 = x38 | n12149 ;
  assign n12151 = ( ~x38 & x87 ) | ( ~x38 & n12150 ) | ( x87 & n12150 ) ;
  assign n12152 = n12151 ^ n5014 ^ 1'b0 ;
  assign n12153 = ( n5014 & n12151 ) | ( n5014 & n12152 ) | ( n12151 & n12152 ) ;
  assign n12154 = ( x92 & ~n5014 ) | ( x92 & n12153 ) | ( ~n5014 & n12153 ) ;
  assign n12155 = n12154 ^ n12147 ^ 1'b0 ;
  assign n12156 = ( n12147 & n12154 ) | ( n12147 & n12155 ) | ( n12154 & n12155 ) ;
  assign n12157 = ( x55 & ~n12147 ) | ( x55 & n12156 ) | ( ~n12147 & n12156 ) ;
  assign n12158 = n12157 ^ n6249 ^ 1'b0 ;
  assign n12159 = ( n6249 & n12157 ) | ( n6249 & n12158 ) | ( n12157 & n12158 ) ;
  assign n12160 = ( x56 & ~n6249 ) | ( x56 & n12159 ) | ( ~n6249 & n12159 ) ;
  assign n12161 = n12160 ^ n5008 ^ 1'b0 ;
  assign n12162 = ( n5008 & n12160 ) | ( n5008 & n12161 ) | ( n12160 & n12161 ) ;
  assign n12163 = ( x62 & ~n5008 ) | ( x62 & n12162 ) | ( ~n5008 & n12162 ) ;
  assign n12164 = ( x57 & ~n5006 ) | ( x57 & n12163 ) | ( ~n5006 & n12163 ) ;
  assign n12165 = ~x57 & n12164 ;
  assign n12166 = x79 | n10322 ;
  assign n12167 = x163 | n8272 ;
  assign n12168 = n10323 | n10324 ;
  assign n12169 = ~x150 & n12168 ;
  assign n12170 = x150 & ~n8275 ;
  assign n12171 = n12167 | n12170 ;
  assign n12172 = ( ~n12167 & n12169 ) | ( ~n12167 & n12171 ) | ( n12169 & n12171 ) ;
  assign n12173 = x232 & n12172 ;
  assign n12174 = n7555 & n12173 ;
  assign n12175 = x74 & ~n12174 ;
  assign n12176 = x165 & n6411 ;
  assign n12177 = x38 | x54 ;
  assign n12178 = ~n12176 & n12177 ;
  assign n12179 = ~n7555 & n12178 ;
  assign n12180 = x74 | n12174 ;
  assign n12181 = n12179 | n12180 ;
  assign n12182 = ~n12175 & n12181 ;
  assign n12183 = n2109 & ~n12182 ;
  assign n12184 = n2120 | n12183 ;
  assign n12185 = ~n7555 & n12176 ;
  assign n12186 = n2120 & ~n12185 ;
  assign n12187 = n7555 & ~n12173 ;
  assign n12188 = ( n12175 & n12186 ) | ( n12175 & ~n12187 ) | ( n12186 & ~n12187 ) ;
  assign n12189 = ~n12175 & n12188 ;
  assign n12190 = x184 | n10369 ;
  assign n12191 = x185 & n12190 ;
  assign n12192 = n5075 | n12191 ;
  assign n12193 = ( x185 & n12190 ) | ( x185 & ~n12192 ) | ( n12190 & ~n12192 ) ;
  assign n12194 = ~n12192 & n12193 ;
  assign n12195 = ( x232 & x299 ) | ( x232 & n12194 ) | ( x299 & n12194 ) ;
  assign n12196 = n12194 ^ x299 ^ 1'b0 ;
  assign n12197 = ( x232 & n12195 ) | ( x232 & n12196 ) | ( n12195 & n12196 ) ;
  assign n12198 = n12197 ^ n12172 ^ 1'b0 ;
  assign n12199 = ( ~x299 & n12172 ) | ( ~x299 & n12198 ) | ( n12172 & n12198 ) ;
  assign n12200 = ( n12197 & ~n12198 ) | ( n12197 & n12199 ) | ( ~n12198 & n12199 ) ;
  assign n12201 = n7555 & n12200 ;
  assign n12202 = x74 & ~n12201 ;
  assign n12203 = x299 ^ x165 ^ 1'b0 ;
  assign n12204 = ( x143 & x165 ) | ( x143 & ~n12203 ) | ( x165 & ~n12203 ) ;
  assign n12205 = n6411 & n12204 ;
  assign n12206 = n7555 | n12205 ;
  assign n12207 = x54 & ~n12201 ;
  assign n12208 = n12206 & n12207 ;
  assign n12209 = x100 & ~n12200 ;
  assign n12210 = x38 & ~n12205 ;
  assign n12211 = n6512 & ~n12210 ;
  assign n12212 = ~n5165 & n8127 ;
  assign n12213 = x232 | n8129 ;
  assign n12214 = n12212 | n12213 ;
  assign n12215 = x168 & ~n8105 ;
  assign n12216 = x151 | n12215 ;
  assign n12217 = ( x168 & n8133 ) | ( x168 & ~n12216 ) | ( n8133 & ~n12216 ) ;
  assign n12218 = ~n12216 & n12217 ;
  assign n12219 = x151 & ~x168 ;
  assign n12220 = n12218 ^ n8146 ^ 1'b0 ;
  assign n12221 = ( ~n8146 & n12219 ) | ( ~n8146 & n12220 ) | ( n12219 & n12220 ) ;
  assign n12222 = ( n8146 & n12218 ) | ( n8146 & n12221 ) | ( n12218 & n12221 ) ;
  assign n12223 = n12222 ^ n8099 ^ 1'b0 ;
  assign n12224 = ( x150 & n8099 ) | ( x150 & ~n12222 ) | ( n8099 & ~n12222 ) ;
  assign n12225 = ( x150 & ~n12223 ) | ( x150 & n12224 ) | ( ~n12223 & n12224 ) ;
  assign n12226 = ~x151 & n8129 ;
  assign n12227 = ( ~x168 & n8163 ) | ( ~x168 & n12226 ) | ( n8163 & n12226 ) ;
  assign n12228 = ~x168 & n12227 ;
  assign n12229 = x168 & ~n5075 ;
  assign n12230 = ~x151 & n8117 ;
  assign n12231 = ( n8157 & n12229 ) | ( n8157 & n12230 ) | ( n12229 & n12230 ) ;
  assign n12232 = n12229 & n12231 ;
  assign n12233 = x150 | n12232 ;
  assign n12234 = ( ~n12225 & n12228 ) | ( ~n12225 & n12233 ) | ( n12228 & n12233 ) ;
  assign n12235 = ~n12225 & n12234 ;
  assign n12236 = n5075 & n10403 ;
  assign n12237 = ( x299 & n12235 ) | ( x299 & ~n12236 ) | ( n12235 & ~n12236 ) ;
  assign n12238 = ~n12235 & n12237 ;
  assign n12239 = n5075 & n8130 ;
  assign n12240 = ~x173 & x190 ;
  assign n12241 = n8106 & n12240 ;
  assign n12242 = ~n5203 & n8146 ;
  assign n12243 = x173 & n12242 ;
  assign n12244 = x173 | n5203 ;
  assign n12245 = ~n12243 & n12244 ;
  assign n12246 = ( n8133 & n12243 ) | ( n8133 & ~n12245 ) | ( n12243 & ~n12245 ) ;
  assign n12247 = ( x190 & ~n5075 ) | ( x190 & n12246 ) | ( ~n5075 & n12246 ) ;
  assign n12248 = ~x190 & n12247 ;
  assign n12249 = ( x185 & n12241 ) | ( x185 & ~n12248 ) | ( n12241 & ~n12248 ) ;
  assign n12250 = ~n12241 & n12249 ;
  assign n12251 = ~x173 & n8129 ;
  assign n12252 = ( ~x190 & n8143 ) | ( ~x190 & n12251 ) | ( n8143 & n12251 ) ;
  assign n12253 = ~x190 & n12252 ;
  assign n12254 = x173 & ~n8140 ;
  assign n12255 = x190 & n8119 ;
  assign n12256 = n12255 ^ n12254 ^ 1'b0 ;
  assign n12257 = ( n12254 & n12255 ) | ( n12254 & n12256 ) | ( n12255 & n12256 ) ;
  assign n12258 = ( x185 & ~n12254 ) | ( x185 & n12257 ) | ( ~n12254 & n12257 ) ;
  assign n12259 = ( ~n12250 & n12253 ) | ( ~n12250 & n12258 ) | ( n12253 & n12258 ) ;
  assign n12260 = ~n12250 & n12259 ;
  assign n12261 = ( x299 & ~n12239 ) | ( x299 & n12260 ) | ( ~n12239 & n12260 ) ;
  assign n12262 = n12239 | n12261 ;
  assign n12263 = x232 & ~n12262 ;
  assign n12264 = ( x232 & n12238 ) | ( x232 & n12263 ) | ( n12238 & n12263 ) ;
  assign n12265 = ( x39 & n12214 ) | ( x39 & ~n12264 ) | ( n12214 & ~n12264 ) ;
  assign n12266 = ~x39 & n12265 ;
  assign n12267 = n6261 & n8201 ;
  assign n12268 = n5100 & n11620 ;
  assign n12269 = n5374 & n12268 ;
  assign n12270 = ( x232 & ~n12267 ) | ( x232 & n12269 ) | ( ~n12267 & n12269 ) ;
  assign n12271 = n12267 | n12270 ;
  assign n12272 = n5099 & n5374 ;
  assign n12273 = x178 & ~n8196 ;
  assign n12274 = ~n12272 & n12273 ;
  assign n12275 = x190 | n12274 ;
  assign n12276 = ( x178 & n11662 ) | ( x178 & ~n12275 ) | ( n11662 & ~n12275 ) ;
  assign n12277 = ~n12275 & n12276 ;
  assign n12278 = ~x178 & n5114 ;
  assign n12279 = n8188 & n12278 ;
  assign n12280 = n12272 | n12279 ;
  assign n12281 = n12277 ^ x190 ^ 1'b0 ;
  assign n12282 = ( ~x190 & n12280 ) | ( ~x190 & n12281 ) | ( n12280 & n12281 ) ;
  assign n12283 = ( x190 & n12277 ) | ( x190 & n12282 ) | ( n12277 & n12282 ) ;
  assign n12284 = ( n2290 & n5106 ) | ( n2290 & n12283 ) | ( n5106 & n12283 ) ;
  assign n12285 = ~n2290 & n12284 ;
  assign n12286 = ~x157 & n8189 ;
  assign n12287 = x168 & ~n12286 ;
  assign n12288 = x157 | x168 ;
  assign n12289 = n8184 | n12288 ;
  assign n12290 = x157 & ~n8182 ;
  assign n12291 = ( n12287 & n12289 ) | ( n12287 & ~n12290 ) | ( n12289 & ~n12290 ) ;
  assign n12292 = ~n12287 & n12291 ;
  assign n12293 = ( n11620 & n12272 ) | ( n11620 & n12292 ) | ( n12272 & n12292 ) ;
  assign n12294 = n12292 ^ n12272 ^ 1'b0 ;
  assign n12295 = ( n11620 & n12293 ) | ( n11620 & n12294 ) | ( n12293 & n12294 ) ;
  assign n12296 = ( x232 & n12285 ) | ( x232 & ~n12295 ) | ( n12285 & ~n12295 ) ;
  assign n12297 = ~n12285 & n12296 ;
  assign n12298 = x39 & ~n12297 ;
  assign n12299 = n12271 & n12298 ;
  assign n12300 = ( ~x38 & n12266 ) | ( ~x38 & n12299 ) | ( n12266 & n12299 ) ;
  assign n12301 = ~x38 & n12300 ;
  assign n12302 = x143 & ~n7659 ;
  assign n12303 = x165 & ~n12302 ;
  assign n12304 = x143 | n7662 ;
  assign n12305 = n12303 & n12304 ;
  assign n12306 = x143 & ~x165 ;
  assign n12307 = n7656 & n12306 ;
  assign n12308 = ( x38 & n12305 ) | ( x38 & ~n12307 ) | ( n12305 & ~n12307 ) ;
  assign n12309 = ~n12305 & n12308 ;
  assign n12310 = ( n2051 & ~n12301 ) | ( n2051 & n12309 ) | ( ~n12301 & n12309 ) ;
  assign n12311 = n12301 | n12310 ;
  assign n12312 = ( n12209 & ~n12211 ) | ( n12209 & n12311 ) | ( ~n12211 & n12311 ) ;
  assign n12313 = ~n12209 & n12312 ;
  assign n12314 = ( x75 & x92 ) | ( x75 & ~n12313 ) | ( x92 & ~n12313 ) ;
  assign n12315 = n12313 | n12314 ;
  assign n12316 = x75 & ~n12200 ;
  assign n12317 = n12316 ^ n7639 ^ 1'b0 ;
  assign n12318 = x100 | n12210 ;
  assign n12319 = x178 | x299 ;
  assign n12320 = ~x157 & x299 ;
  assign n12321 = n6411 & ~n12320 ;
  assign n12322 = n12319 & n12321 ;
  assign n12323 = n7459 | n12322 ;
  assign n12324 = n1292 | n12323 ;
  assign n12325 = n12324 ^ n12318 ^ 1'b0 ;
  assign n12326 = ( n12318 & n12324 ) | ( n12318 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12327 = ( n12209 & ~n12318 ) | ( n12209 & n12326 ) | ( ~n12318 & n12326 ) ;
  assign n12328 = ( n7639 & ~n12317 ) | ( n7639 & n12327 ) | ( ~n12317 & n12327 ) ;
  assign n12329 = ( n12316 & n12317 ) | ( n12316 & n12328 ) | ( n12317 & n12328 ) ;
  assign n12330 = ( x54 & n12315 ) | ( x54 & ~n12329 ) | ( n12315 & ~n12329 ) ;
  assign n12331 = n12330 ^ n12315 ^ 1'b0 ;
  assign n12332 = ( x54 & n12330 ) | ( x54 & ~n12331 ) | ( n12330 & ~n12331 ) ;
  assign n12333 = n12332 ^ n12208 ^ 1'b0 ;
  assign n12334 = ( n12208 & n12332 ) | ( n12208 & n12333 ) | ( n12332 & n12333 ) ;
  assign n12335 = ( x74 & ~n12208 ) | ( x74 & n12334 ) | ( ~n12208 & n12334 ) ;
  assign n12336 = ( x55 & ~n12202 ) | ( x55 & n12335 ) | ( ~n12202 & n12335 ) ;
  assign n12337 = ~x55 & n12336 ;
  assign n12338 = x92 | n7555 ;
  assign n12339 = x150 & n6411 ;
  assign n12340 = ( n7459 & ~n12338 ) | ( n7459 & n12339 ) | ( ~n12338 & n12339 ) ;
  assign n12341 = n12338 | n12340 ;
  assign n12342 = n12341 ^ x54 ^ 1'b0 ;
  assign n12343 = ( ~x54 & n12176 ) | ( ~x54 & n12342 ) | ( n12176 & n12342 ) ;
  assign n12344 = ( x54 & n12341 ) | ( x54 & n12343 ) | ( n12341 & n12343 ) ;
  assign n12345 = n1292 | n12344 ;
  assign n12346 = ~n12181 & n12345 ;
  assign n12347 = ( x55 & n12175 ) | ( x55 & ~n12346 ) | ( n12175 & ~n12346 ) ;
  assign n12348 = ~n12175 & n12347 ;
  assign n12349 = ( n2109 & ~n12337 ) | ( n2109 & n12348 ) | ( ~n12337 & n12348 ) ;
  assign n12350 = n12337 | n12349 ;
  assign n12351 = n12184 | n12350 ;
  assign n12352 = ( ~n12184 & n12189 ) | ( ~n12184 & n12351 ) | ( n12189 & n12351 ) ;
  assign n12353 = x118 | n12352 ;
  assign n12354 = n12166 & n12353 ;
  assign n12355 = ~x118 & n8260 ;
  assign n12356 = n12352 | n12355 ;
  assign n12357 = n8298 & n12184 ;
  assign n12358 = n7569 | n12177 ;
  assign n12359 = x92 | n7648 ;
  assign n12360 = n12339 & ~n12359 ;
  assign n12361 = ( ~n12178 & n12358 ) | ( ~n12178 & n12360 ) | ( n12358 & n12360 ) ;
  assign n12362 = ~n12178 & n12361 ;
  assign n12363 = n7555 | n12362 ;
  assign n12364 = ~n12180 & n12363 ;
  assign n12365 = ( x55 & n12175 ) | ( x55 & ~n12364 ) | ( n12175 & ~n12364 ) ;
  assign n12366 = ~n12175 & n12365 ;
  assign n12367 = x178 & ~n7726 ;
  assign n12368 = x190 | n12367 ;
  assign n12369 = ~x299 & n12368 ;
  assign n12370 = x157 & n7697 ;
  assign n12371 = x168 & n7681 ;
  assign n12372 = n12370 | n12371 ;
  assign n12373 = n5061 & n7669 ;
  assign n12374 = ~n5075 & n12373 ;
  assign n12375 = ( ~x299 & n12372 ) | ( ~x299 & n12374 ) | ( n12372 & n12374 ) ;
  assign n12376 = x299 & n12375 ;
  assign n12377 = x299 & ~n12376 ;
  assign n12378 = ( x178 & n12376 ) | ( x178 & ~n12377 ) | ( n12376 & ~n12377 ) ;
  assign n12379 = ( n7569 & ~n12369 ) | ( n7569 & n12378 ) | ( ~n12369 & n12378 ) ;
  assign n12380 = ~n12369 & n12379 ;
  assign n12381 = ( n5114 & n7678 ) | ( n5114 & n7722 ) | ( n7678 & n7722 ) ;
  assign n12382 = x178 & n12381 ;
  assign n12383 = ~n7715 & n12382 ;
  assign n12384 = ~x299 & n7679 ;
  assign n12385 = x190 & n12384 ;
  assign n12386 = ~x178 & n12381 ;
  assign n12387 = ~n7684 & n12386 ;
  assign n12388 = ( n12383 & n12385 ) | ( n12383 & ~n12387 ) | ( n12385 & ~n12387 ) ;
  assign n12389 = ~n12383 & n12388 ;
  assign n12390 = ( x232 & n12380 ) | ( x232 & ~n12389 ) | ( n12380 & ~n12389 ) ;
  assign n12391 = ~n12380 & n12390 ;
  assign n12392 = x232 | n7569 ;
  assign n12393 = ( x39 & n12391 ) | ( x39 & n12392 ) | ( n12391 & n12392 ) ;
  assign n12394 = ~n12391 & n12393 ;
  assign n12395 = x232 | n7944 ;
  assign n12396 = n5075 & ~n7944 ;
  assign n12397 = n8051 & n12219 ;
  assign n12398 = x168 & ~n8044 ;
  assign n12399 = x168 | n8041 ;
  assign n12400 = ( x151 & ~n12398 ) | ( x151 & n12399 ) | ( ~n12398 & n12399 ) ;
  assign n12401 = ~x151 & n12400 ;
  assign n12402 = ( ~n12396 & n12397 ) | ( ~n12396 & n12401 ) | ( n12397 & n12401 ) ;
  assign n12403 = ~n12396 & n12402 ;
  assign n12404 = n7978 ^ n7976 ^ n7944 ;
  assign n12405 = ( ~x151 & x168 ) | ( ~x151 & n12404 ) | ( x168 & n12404 ) ;
  assign n12406 = x151 & n12405 ;
  assign n12407 = ( x150 & n12403 ) | ( x150 & ~n12406 ) | ( n12403 & ~n12406 ) ;
  assign n12408 = ~n12403 & n12407 ;
  assign n12409 = x168 & ~n7958 ;
  assign n12410 = n7944 | n12229 ;
  assign n12411 = ( x151 & ~n12409 ) | ( x151 & n12410 ) | ( ~n12409 & n12410 ) ;
  assign n12412 = ~x151 & n12411 ;
  assign n12413 = n7984 & ~n12396 ;
  assign n12414 = x168 | n12413 ;
  assign n12415 = n5075 & n7944 ;
  assign n12416 = n7866 | n12415 ;
  assign n12417 = ( x151 & n12219 ) | ( x151 & n12416 ) | ( n12219 & n12416 ) ;
  assign n12418 = n12414 & n12417 ;
  assign n12419 = ( x150 & ~n12412 ) | ( x150 & n12418 ) | ( ~n12412 & n12418 ) ;
  assign n12420 = n12412 | n12419 ;
  assign n12421 = ( x299 & n12408 ) | ( x299 & n12420 ) | ( n12408 & n12420 ) ;
  assign n12422 = ~n12408 & n12421 ;
  assign n12423 = x173 & ~n12416 ;
  assign n12424 = x173 & ~n12415 ;
  assign n12425 = ( n7958 & ~n12396 ) | ( n7958 & n12424 ) | ( ~n12396 & n12424 ) ;
  assign n12426 = ( x185 & ~n12423 ) | ( x185 & n12425 ) | ( ~n12423 & n12425 ) ;
  assign n12427 = ~x185 & n12426 ;
  assign n12428 = ~n5075 & n7795 ;
  assign n12429 = n12424 & ~n12428 ;
  assign n12430 = ( n7965 & ~n12396 ) | ( n7965 & n12424 ) | ( ~n12396 & n12424 ) ;
  assign n12431 = ( x185 & n12429 ) | ( x185 & n12430 ) | ( n12429 & n12430 ) ;
  assign n12432 = ~n12429 & n12431 ;
  assign n12433 = ( x190 & n12427 ) | ( x190 & ~n12432 ) | ( n12427 & ~n12432 ) ;
  assign n12434 = ~n12427 & n12433 ;
  assign n12435 = x173 | n7944 ;
  assign n12436 = x173 & ~n12413 ;
  assign n12437 = ( x185 & n12435 ) | ( x185 & ~n12436 ) | ( n12435 & ~n12436 ) ;
  assign n12438 = ~x185 & n12437 ;
  assign n12439 = x185 & ~n12396 ;
  assign n12440 = ~x173 & n7951 ;
  assign n12441 = x173 & n8367 ;
  assign n12442 = ( n5075 & ~n12440 ) | ( n5075 & n12441 ) | ( ~n12440 & n12441 ) ;
  assign n12443 = n12440 | n12442 ;
  assign n12444 = n12439 & n12443 ;
  assign n12445 = ( x190 & ~n12438 ) | ( x190 & n12444 ) | ( ~n12438 & n12444 ) ;
  assign n12446 = n12438 | n12445 ;
  assign n12447 = ( x299 & ~n12434 ) | ( x299 & n12446 ) | ( ~n12434 & n12446 ) ;
  assign n12448 = ~x299 & n12447 ;
  assign n12449 = ( x232 & n12422 ) | ( x232 & ~n12448 ) | ( n12422 & ~n12448 ) ;
  assign n12450 = ~n12422 & n12449 ;
  assign n12451 = ( x39 & n12395 ) | ( x39 & ~n12450 ) | ( n12395 & ~n12450 ) ;
  assign n12452 = ~x39 & n12451 ;
  assign n12453 = ( x38 & ~n12394 ) | ( x38 & n12452 ) | ( ~n12394 & n12452 ) ;
  assign n12454 = n12394 | n12453 ;
  assign n12455 = ( n2051 & ~n12309 ) | ( n2051 & n12454 ) | ( ~n12309 & n12454 ) ;
  assign n12456 = ~n2051 & n12455 ;
  assign n12457 = n7570 & n12211 ;
  assign n12458 = n12209 | n12457 ;
  assign n12459 = ( ~n2053 & n12456 ) | ( ~n2053 & n12458 ) | ( n12456 & n12458 ) ;
  assign n12460 = ~n2053 & n12459 ;
  assign n12461 = ~n7648 & n12322 ;
  assign n12462 = n7570 | n12461 ;
  assign n12463 = n12462 ^ n12318 ^ 1'b0 ;
  assign n12464 = ( n12318 & n12462 ) | ( n12318 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = ( n12209 & ~n12318 ) | ( n12209 & n12464 ) | ( ~n12318 & n12464 ) ;
  assign n12466 = ( x75 & x92 ) | ( x75 & n12465 ) | ( x92 & n12465 ) ;
  assign n12467 = ~x75 & n12466 ;
  assign n12468 = n12200 & ~n12467 ;
  assign n12469 = ( x75 & n12467 ) | ( x75 & ~n12468 ) | ( n12467 & ~n12468 ) ;
  assign n12470 = ( ~x54 & n12460 ) | ( ~x54 & n12469 ) | ( n12460 & n12469 ) ;
  assign n12471 = ~x54 & n12470 ;
  assign n12472 = ( ~x74 & n12208 ) | ( ~x74 & n12471 ) | ( n12208 & n12471 ) ;
  assign n12473 = ~x74 & n12472 ;
  assign n12474 = ( x55 & n12202 ) | ( x55 & ~n12473 ) | ( n12202 & ~n12473 ) ;
  assign n12475 = n12473 | n12474 ;
  assign n12476 = ( n2109 & ~n12366 ) | ( n2109 & n12475 ) | ( ~n12366 & n12475 ) ;
  assign n12477 = ~n2109 & n12476 ;
  assign n12478 = ( ~n12189 & n12357 ) | ( ~n12189 & n12477 ) | ( n12357 & n12477 ) ;
  assign n12479 = ~n12189 & n12478 ;
  assign n12480 = n12355 & n12479 ;
  assign n12481 = ( n12166 & n12356 ) | ( n12166 & ~n12480 ) | ( n12356 & ~n12480 ) ;
  assign n12482 = ~n12166 & n12481 ;
  assign n12483 = x118 & n12479 ;
  assign n12484 = ~n12482 & n12483 ;
  assign n12485 = ( n12354 & n12482 ) | ( n12354 & ~n12484 ) | ( n12482 & ~n12484 ) ;
  assign n12486 = x128 & x228 ;
  assign n12487 = ~n1457 & n8752 ;
  assign n12488 = ( ~n1564 & n10315 ) | ( ~n1564 & n12487 ) | ( n10315 & n12487 ) ;
  assign n12489 = ~n1564 & n12488 ;
  assign n12490 = x97 | n12489 ;
  assign n12491 = ~x46 & n1670 ;
  assign n12492 = ( n1622 & n12490 ) | ( n1622 & n12491 ) | ( n12490 & n12491 ) ;
  assign n12493 = ~n1622 & n12492 ;
  assign n12494 = x299 & n5304 ;
  assign n12495 = ( n5355 & n6411 ) | ( n5355 & n12494 ) | ( n6411 & n12494 ) ;
  assign n12496 = n6411 & n12495 ;
  assign n12497 = x109 & ~n12496 ;
  assign n12498 = ~n1670 & n10316 ;
  assign n12499 = ( ~n12493 & n12497 ) | ( ~n12493 & n12498 ) | ( n12497 & n12498 ) ;
  assign n12500 = n12493 | n12499 ;
  assign n12501 = n12496 ^ n5306 ^ 1'b0 ;
  assign n12502 = ( n5206 & n5306 ) | ( n5206 & ~n12501 ) | ( n5306 & ~n12501 ) ;
  assign n12503 = ( x91 & n12500 ) | ( x91 & ~n12502 ) | ( n12500 & ~n12502 ) ;
  assign n12504 = n12503 ^ n12500 ^ 1'b0 ;
  assign n12505 = ( x91 & n12503 ) | ( x91 & ~n12504 ) | ( n12503 & ~n12504 ) ;
  assign n12506 = ( ~n1412 & n5261 ) | ( ~n1412 & n12505 ) | ( n5261 & n12505 ) ;
  assign n12507 = ~n5261 & n12506 ;
  assign n12508 = n1267 & ~n12507 ;
  assign n12509 = ( x93 & n12507 ) | ( x93 & ~n12508 ) | ( n12507 & ~n12508 ) ;
  assign n12510 = ( x39 & ~n9713 ) | ( x39 & n12509 ) | ( ~n9713 & n12509 ) ;
  assign n12511 = ~x39 & n12510 ;
  assign n12512 = n2263 & n4736 ;
  assign n12513 = n6465 & n12512 ;
  assign n12514 = n1359 & ~n2290 ;
  assign n12515 = n6461 & n12514 ;
  assign n12516 = ( x39 & n12513 ) | ( x39 & n12515 ) | ( n12513 & n12515 ) ;
  assign n12517 = n12515 ^ n12513 ^ 1'b0 ;
  assign n12518 = ( x39 & n12516 ) | ( x39 & n12517 ) | ( n12516 & n12517 ) ;
  assign n12519 = ( ~x38 & n12511 ) | ( ~x38 & n12518 ) | ( n12511 & n12518 ) ;
  assign n12520 = ~x38 & n12519 ;
  assign n12521 = ~x228 & n12520 ;
  assign n12522 = ( ~x100 & n12486 ) | ( ~x100 & n12521 ) | ( n12486 & n12521 ) ;
  assign n12523 = ~x100 & n12522 ;
  assign n12524 = n1994 | n2142 ;
  assign n12525 = ~n12486 & n12524 ;
  assign n12526 = x100 & ~n12525 ;
  assign n12527 = ( x87 & ~n12523 ) | ( x87 & n12526 ) | ( ~n12523 & n12526 ) ;
  assign n12528 = n12523 | n12527 ;
  assign n12529 = x87 & ~n12486 ;
  assign n12530 = ( x75 & n12528 ) | ( x75 & ~n12529 ) | ( n12528 & ~n12529 ) ;
  assign n12531 = ~x75 & n12530 ;
  assign n12532 = n6317 | n7459 ;
  assign n12533 = ~n12486 & n12532 ;
  assign n12534 = x75 & ~n12533 ;
  assign n12535 = ( x92 & ~n12531 ) | ( x92 & n12534 ) | ( ~n12531 & n12534 ) ;
  assign n12536 = n12531 | n12535 ;
  assign n12537 = x92 & ~n12486 ;
  assign n12538 = n6331 & n12537 ;
  assign n12539 = ( n8758 & n12536 ) | ( n8758 & ~n12538 ) | ( n12536 & ~n12538 ) ;
  assign n12540 = ~n8758 & n12539 ;
  assign n12541 = n12540 ^ n8758 ^ 1'b0 ;
  assign n12542 = ( ~n8758 & n12486 ) | ( ~n8758 & n12541 ) | ( n12486 & n12541 ) ;
  assign n12543 = ( n8758 & n12540 ) | ( n8758 & n12542 ) | ( n12540 & n12542 ) ;
  assign n12544 = x31 | x80 ;
  assign n12545 = x818 & ~n12544 ;
  assign n12546 = n12545 ^ n7318 ^ 1'b0 ;
  assign n12547 = n6782 & n11179 ;
  assign n12548 = n6612 & ~n12547 ;
  assign n12549 = ~x120 & n6782 ;
  assign n12550 = ~x1093 & n12549 ;
  assign n12551 = n12548 & ~n12550 ;
  assign n12552 = x120 | x1093 ;
  assign n12553 = n6421 & n12552 ;
  assign n12554 = x87 & ~n6499 ;
  assign n12555 = n12552 & n12554 ;
  assign n12556 = x38 & ~n12552 ;
  assign n12557 = x100 | n12556 ;
  assign n12558 = x1093 & ~n5099 ;
  assign n12559 = ~n5114 & n12558 ;
  assign n12560 = n5083 & n5114 ;
  assign n12561 = n6801 & ~n12560 ;
  assign n12562 = ( n6460 & n12559 ) | ( n6460 & n12561 ) | ( n12559 & n12561 ) ;
  assign n12563 = ~n12559 & n12562 ;
  assign n12564 = ( x299 & n12552 ) | ( x299 & ~n12563 ) | ( n12552 & ~n12563 ) ;
  assign n12565 = ~x299 & n12564 ;
  assign n12566 = ~n5061 & n12558 ;
  assign n12567 = n5061 & n5083 ;
  assign n12568 = n6810 & ~n12567 ;
  assign n12569 = ( n6460 & n12566 ) | ( n6460 & n12568 ) | ( n12566 & n12568 ) ;
  assign n12570 = ~n12566 & n12569 ;
  assign n12571 = ( x299 & n12552 ) | ( x299 & n12570 ) | ( n12552 & n12570 ) ;
  assign n12572 = ~n12570 & n12571 ;
  assign n12573 = ( x39 & n12565 ) | ( x39 & ~n12572 ) | ( n12565 & ~n12572 ) ;
  assign n12574 = ~n12565 & n12573 ;
  assign n12575 = x1093 | n6403 ;
  assign n12576 = x120 & ~n12575 ;
  assign n12577 = x39 | n12576 ;
  assign n12578 = n6400 & n6425 ;
  assign n12579 = n6489 & ~n12578 ;
  assign n12580 = x122 & ~n6401 ;
  assign n12581 = ~x829 & n12578 ;
  assign n12582 = n6443 & n9041 ;
  assign n12583 = ( x122 & ~n12581 ) | ( x122 & n12582 ) | ( ~n12581 & n12582 ) ;
  assign n12584 = n12581 | n12583 ;
  assign n12585 = ( n1614 & ~n12580 ) | ( n1614 & n12584 ) | ( ~n12580 & n12584 ) ;
  assign n12586 = ~n1614 & n12585 ;
  assign n12587 = ( x1091 & x1093 ) | ( x1091 & n12586 ) | ( x1093 & n12586 ) ;
  assign n12588 = ~n12586 & n12587 ;
  assign n12589 = n12579 | n12588 ;
  assign n12590 = ( ~n12574 & n12577 ) | ( ~n12574 & n12589 ) | ( n12577 & n12589 ) ;
  assign n12591 = ~n12574 & n12590 ;
  assign n12592 = x38 | n12591 ;
  assign n12593 = ~n12557 & n12592 ;
  assign n12594 = ~n1292 & n6417 ;
  assign n12595 = n6483 ^ x120 ^ 1'b0 ;
  assign n12596 = ( n6483 & n12594 ) | ( n6483 & ~n12595 ) | ( n12594 & ~n12595 ) ;
  assign n12597 = ( n1994 & n6824 ) | ( n1994 & n12596 ) | ( n6824 & n12596 ) ;
  assign n12598 = ~n1994 & n12597 ;
  assign n12599 = ( x100 & n12552 ) | ( x100 & n12598 ) | ( n12552 & n12598 ) ;
  assign n12600 = ~n12598 & n12599 ;
  assign n12601 = ( ~x87 & n12593 ) | ( ~x87 & n12600 ) | ( n12593 & n12600 ) ;
  assign n12602 = ~x87 & n12601 ;
  assign n12603 = ( ~x75 & n12555 ) | ( ~x75 & n12602 ) | ( n12555 & n12602 ) ;
  assign n12604 = ~x75 & n12603 ;
  assign n12605 = ( n6782 & ~n12553 ) | ( n6782 & n12604 ) | ( ~n12553 & n12604 ) ;
  assign n12606 = n12553 | n12605 ;
  assign n12607 = ( n6612 & ~n12550 ) | ( n6612 & n12606 ) | ( ~n12550 & n12606 ) ;
  assign n12608 = ~n6612 & n12607 ;
  assign n12609 = n2036 & n11179 ;
  assign n12610 = x87 & ~n12609 ;
  assign n12611 = ~x122 & n6425 ;
  assign n12612 = ( n6494 & n6499 ) | ( n6494 & n12611 ) | ( n6499 & n12611 ) ;
  assign n12613 = n12610 & ~n12612 ;
  assign n12614 = n12555 & n12613 ;
  assign n12615 = ~x120 & x1093 ;
  assign n12616 = n6483 & ~n12615 ;
  assign n12617 = x120 & ~n11179 ;
  assign n12618 = ~n6483 & n12617 ;
  assign n12619 = n12594 & ~n12618 ;
  assign n12620 = n12616 | n12619 ;
  assign n12621 = ( n1994 & n6824 ) | ( n1994 & n12620 ) | ( n6824 & n12620 ) ;
  assign n12622 = ~n1994 & n12621 ;
  assign n12623 = n6489 & ~n12611 ;
  assign n12624 = ( n8670 & n12615 ) | ( n8670 & n12623 ) | ( n12615 & n12623 ) ;
  assign n12625 = n12617 | n12624 ;
  assign n12626 = ( x100 & n12622 ) | ( x100 & n12625 ) | ( n12622 & n12625 ) ;
  assign n12627 = ~n12622 & n12626 ;
  assign n12628 = n12579 & ~n12611 ;
  assign n12629 = n12588 | n12628 ;
  assign n12630 = n12577 | n12629 ;
  assign n12631 = n6810 | n12625 ;
  assign n12632 = ~n6460 & n12617 ;
  assign n12633 = x1091 & x1092 ;
  assign n12634 = n6458 & n12633 ;
  assign n12635 = n12624 & ~n12634 ;
  assign n12636 = n12632 | n12635 ;
  assign n12637 = ( n5083 & n12625 ) | ( n5083 & n12636 ) | ( n12625 & n12636 ) ;
  assign n12638 = n5061 & n12637 ;
  assign n12639 = n12625 ^ n5099 ^ 1'b0 ;
  assign n12640 = ( n12625 & n12636 ) | ( n12625 & n12639 ) | ( n12636 & n12639 ) ;
  assign n12641 = ~n5061 & n12640 ;
  assign n12642 = ( n6810 & n12638 ) | ( n6810 & ~n12641 ) | ( n12638 & ~n12641 ) ;
  assign n12643 = ~n12638 & n12642 ;
  assign n12644 = x299 & ~n12643 ;
  assign n12645 = n12631 & n12644 ;
  assign n12646 = n5114 & n12637 ;
  assign n12647 = ~n5114 & n12640 ;
  assign n12648 = ( n6801 & n12646 ) | ( n6801 & ~n12647 ) | ( n12646 & ~n12647 ) ;
  assign n12649 = ~n12646 & n12648 ;
  assign n12650 = n6801 | n12625 ;
  assign n12651 = ( x299 & ~n12649 ) | ( x299 & n12650 ) | ( ~n12649 & n12650 ) ;
  assign n12652 = ~x299 & n12651 ;
  assign n12653 = ( x39 & n12645 ) | ( x39 & ~n12652 ) | ( n12645 & ~n12652 ) ;
  assign n12654 = ~n12645 & n12653 ;
  assign n12655 = ( x38 & n12630 ) | ( x38 & ~n12654 ) | ( n12630 & ~n12654 ) ;
  assign n12656 = n12655 ^ n12630 ^ 1'b0 ;
  assign n12657 = ( x38 & n12655 ) | ( x38 & ~n12656 ) | ( n12655 & ~n12656 ) ;
  assign n12658 = x38 & n11179 ;
  assign n12659 = ( n12557 & n12657 ) | ( n12557 & ~n12658 ) | ( n12657 & ~n12658 ) ;
  assign n12660 = ~n12557 & n12659 ;
  assign n12661 = ( ~x87 & n12627 ) | ( ~x87 & n12660 ) | ( n12627 & n12660 ) ;
  assign n12662 = ~x87 & n12661 ;
  assign n12663 = ( ~x75 & n12614 ) | ( ~x75 & n12662 ) | ( n12614 & n12662 ) ;
  assign n12664 = ~x75 & n12663 ;
  assign n12665 = n1207 & ~n12625 ;
  assign n12666 = n6412 & ~n12625 ;
  assign n12667 = n11179 ^ n6846 ^ x1091 ;
  assign n12668 = x120 & ~n12667 ;
  assign n12669 = n6412 | n12668 ;
  assign n12670 = ~n6418 & n12624 ;
  assign n12671 = ( ~n12666 & n12669 ) | ( ~n12666 & n12670 ) | ( n12669 & n12670 ) ;
  assign n12672 = ~n12666 & n12671 ;
  assign n12673 = ( n1205 & n1206 ) | ( n1205 & ~n12672 ) | ( n1206 & ~n12672 ) ;
  assign n12674 = n12672 | n12673 ;
  assign n12675 = ( x75 & n12665 ) | ( x75 & n12674 ) | ( n12665 & n12674 ) ;
  assign n12676 = ~n12665 & n12675 ;
  assign n12677 = ( n6782 & ~n12664 ) | ( n6782 & n12676 ) | ( ~n12664 & n12676 ) ;
  assign n12678 = n12664 | n12677 ;
  assign n12679 = n12608 ^ n12551 ^ 1'b0 ;
  assign n12680 = ( ~n12551 & n12678 ) | ( ~n12551 & n12679 ) | ( n12678 & n12679 ) ;
  assign n12681 = ( n12551 & n12608 ) | ( n12551 & n12680 ) | ( n12608 & n12680 ) ;
  assign n12682 = ( n12545 & ~n12546 ) | ( n12545 & n12681 ) | ( ~n12546 & n12681 ) ;
  assign n12683 = ( n7318 & n12546 ) | ( n7318 & n12682 ) | ( n12546 & n12682 ) ;
  assign n12684 = n6612 & ~n12625 ;
  assign n12685 = n6782 & ~n12684 ;
  assign n12686 = n6413 & n11179 ;
  assign n12687 = ~n6413 & n12667 ;
  assign n12688 = ( x75 & n12686 ) | ( x75 & ~n12687 ) | ( n12686 & ~n12687 ) ;
  assign n12689 = ~n12686 & n12688 ;
  assign n12690 = n6486 & ~n11179 ;
  assign n12691 = ~n6810 & n11179 ;
  assign n12692 = n6460 | n11179 ;
  assign n12693 = ( n6798 & n11179 ) | ( n6798 & n12692 ) | ( n11179 & n12692 ) ;
  assign n12694 = n5061 & ~n12693 ;
  assign n12695 = ( n5099 & n11179 ) | ( n5099 & n12692 ) | ( n11179 & n12692 ) ;
  assign n12696 = n5061 | n12695 ;
  assign n12697 = ( n6810 & n12694 ) | ( n6810 & n12696 ) | ( n12694 & n12696 ) ;
  assign n12698 = ~n12694 & n12697 ;
  assign n12699 = ( x299 & n12691 ) | ( x299 & ~n12698 ) | ( n12691 & ~n12698 ) ;
  assign n12700 = ~n12691 & n12699 ;
  assign n12701 = n5114 & ~n12693 ;
  assign n12702 = n5114 | n12695 ;
  assign n12703 = ( n6801 & n12701 ) | ( n6801 & n12702 ) | ( n12701 & n12702 ) ;
  assign n12704 = ~n12701 & n12703 ;
  assign n12705 = ~n6801 & n11179 ;
  assign n12706 = x299 | n12705 ;
  assign n12707 = ( ~n12700 & n12704 ) | ( ~n12700 & n12706 ) | ( n12704 & n12706 ) ;
  assign n12708 = ~n12700 & n12707 ;
  assign n12709 = ( x38 & x39 ) | ( x38 & ~n12708 ) | ( x39 & ~n12708 ) ;
  assign n12710 = n12709 ^ x39 ^ 1'b0 ;
  assign n12711 = ( x38 & n12709 ) | ( x38 & ~n12710 ) | ( n12709 & ~n12710 ) ;
  assign n12712 = n12575 & ~n12629 ;
  assign n12713 = ( x39 & ~n12711 ) | ( x39 & n12712 ) | ( ~n12711 & n12712 ) ;
  assign n12714 = ~n12711 & n12713 ;
  assign n12715 = x100 | n12658 ;
  assign n12716 = ( ~n12690 & n12714 ) | ( ~n12690 & n12715 ) | ( n12714 & n12715 ) ;
  assign n12717 = ~n12690 & n12716 ;
  assign n12718 = x87 | n12717 ;
  assign n12719 = ~n12613 & n12718 ;
  assign n12720 = ( x75 & ~n12689 ) | ( x75 & n12719 ) | ( ~n12689 & n12719 ) ;
  assign n12721 = ~n12689 & n12720 ;
  assign n12722 = n12548 & ~n12721 ;
  assign n12723 = n12685 | n12722 ;
  assign n12724 = n12575 & ~n12589 ;
  assign n12725 = x39 | n12724 ;
  assign n12726 = ~n6471 & n12725 ;
  assign n12727 = x100 | n12726 ;
  assign n12728 = ~n6486 & n12727 ;
  assign n12729 = x87 | n12728 ;
  assign n12730 = ~n12554 & n12729 ;
  assign n12731 = x75 | n12730 ;
  assign n12732 = ~n6421 & n12731 ;
  assign n12733 = n6612 | n12549 ;
  assign n12734 = ( ~n12723 & n12732 ) | ( ~n12723 & n12733 ) | ( n12732 & n12733 ) ;
  assign n12735 = ~n12723 & n12734 ;
  assign n12736 = x120 & ~n12684 ;
  assign n12737 = n12545 & n12552 ;
  assign n12738 = ~n12684 & n12737 ;
  assign n12739 = n7318 & ~n12738 ;
  assign n12740 = ~n12736 & n12739 ;
  assign n12741 = n10841 & ~n12740 ;
  assign n12742 = ( x120 & n12735 ) | ( x120 & n12741 ) | ( n12735 & n12741 ) ;
  assign n12743 = ~n12735 & n12742 ;
  assign n12744 = x951 & x982 ;
  assign n12745 = x1092 & n12744 ;
  assign n12746 = x1093 & n12745 ;
  assign n12747 = x120 | n12746 ;
  assign n12748 = ~n12684 & n12747 ;
  assign n12749 = n12739 & ~n12748 ;
  assign n12750 = n10841 | n12749 ;
  assign n12751 = n6412 & ~n12747 ;
  assign n12752 = x120 & n6419 ;
  assign n12753 = ~x1091 & n12746 ;
  assign n12754 = x120 | n12753 ;
  assign n12755 = x93 | x122 ;
  assign n12756 = n1270 | n12755 ;
  assign n12757 = n1610 & ~n7467 ;
  assign n12758 = ( n1411 & ~n12756 ) | ( n1411 & n12757 ) | ( ~n12756 & n12757 ) ;
  assign n12759 = ~n1411 & n12758 ;
  assign n12760 = n8930 & n12759 ;
  assign n12761 = ( n1373 & n6415 ) | ( n1373 & n12760 ) | ( n6415 & n12760 ) ;
  assign n12762 = ~n1373 & n12761 ;
  assign n12763 = ( n8670 & n12745 ) | ( n8670 & n12762 ) | ( n12745 & n12762 ) ;
  assign n12764 = ~n12762 & n12763 ;
  assign n12765 = n12754 | n12764 ;
  assign n12766 = n12765 ^ n12752 ^ 1'b0 ;
  assign n12767 = ( n12752 & n12765 ) | ( n12752 & n12766 ) | ( n12765 & n12766 ) ;
  assign n12768 = ( n6412 & ~n12752 ) | ( n6412 & n12767 ) | ( ~n12752 & n12767 ) ;
  assign n12769 = ( n1207 & ~n12751 ) | ( n1207 & n12768 ) | ( ~n12751 & n12768 ) ;
  assign n12770 = ~n1207 & n12769 ;
  assign n12771 = n1207 & n12747 ;
  assign n12772 = ( x75 & n12770 ) | ( x75 & ~n12771 ) | ( n12770 & ~n12771 ) ;
  assign n12773 = ~n12770 & n12772 ;
  assign n12774 = n2036 & ~n12747 ;
  assign n12775 = x87 & ~n12774 ;
  assign n12776 = n8670 & n12745 ;
  assign n12777 = x950 & ~n1292 ;
  assign n12778 = ~n1614 & n5021 ;
  assign n12779 = n12777 & n12778 ;
  assign n12780 = n12776 & ~n12779 ;
  assign n12781 = x824 & n12777 ;
  assign n12782 = n12753 & ~n12781 ;
  assign n12783 = ( ~x120 & n12780 ) | ( ~x120 & n12782 ) | ( n12780 & n12782 ) ;
  assign n12784 = ~x120 & n12783 ;
  assign n12785 = ( x120 & n2036 ) | ( x120 & ~n6497 ) | ( n2036 & ~n6497 ) ;
  assign n12786 = ( n2036 & ~n6498 ) | ( n2036 & n12785 ) | ( ~n6498 & n12785 ) ;
  assign n12787 = n12784 | n12786 ;
  assign n12788 = n12775 & n12787 ;
  assign n12789 = x75 | n12788 ;
  assign n12790 = n6395 & n6415 ;
  assign n12791 = n12777 & n12790 ;
  assign n12792 = n12776 & ~n12791 ;
  assign n12793 = n12754 | n12792 ;
  assign n12794 = x120 & n6483 ;
  assign n12795 = n12793 & ~n12794 ;
  assign n12796 = ( x39 & n6824 ) | ( x39 & ~n12795 ) | ( n6824 & ~n12795 ) ;
  assign n12797 = ~x39 & n12796 ;
  assign n12798 = ( x38 & x100 ) | ( x38 & ~n12797 ) | ( x100 & ~n12797 ) ;
  assign n12799 = n12798 ^ x100 ^ 1'b0 ;
  assign n12800 = ( x38 & n12798 ) | ( x38 & ~n12799 ) | ( n12798 & ~n12799 ) ;
  assign n12801 = ~n1994 & n6824 ;
  assign n12802 = n12801 ^ n12747 ^ 1'b0 ;
  assign n12803 = ( n12747 & n12801 ) | ( n12747 & ~n12802 ) | ( n12801 & ~n12802 ) ;
  assign n12804 = ( n12800 & n12802 ) | ( n12800 & n12803 ) | ( n12802 & n12803 ) ;
  assign n12805 = x120 & n12724 ;
  assign n12806 = ~n1458 & n6382 ;
  assign n12807 = ~n1454 & n12806 ;
  assign n12808 = ~n8111 & n12807 ;
  assign n12809 = n6373 | n12808 ;
  assign n12810 = ( ~n6373 & n6378 ) | ( ~n6373 & n12809 ) | ( n6378 & n12809 ) ;
  assign n12811 = x950 & ~n6423 ;
  assign n12812 = n12810 & n12811 ;
  assign n12813 = x824 & n12812 ;
  assign n12814 = n12745 & ~n12813 ;
  assign n12815 = ~x829 & n12814 ;
  assign n12816 = x97 | n12807 ;
  assign n12817 = ~n1625 & n12816 ;
  assign n12818 = n1623 | n12817 ;
  assign n12819 = ( ~n1623 & n6428 ) | ( ~n1623 & n12818 ) | ( n6428 & n12818 ) ;
  assign n12820 = n1225 | n12819 ;
  assign n12821 = ( ~n1225 & n6376 ) | ( ~n1225 & n12820 ) | ( n6376 & n12820 ) ;
  assign n12822 = n12821 ^ n6373 ^ 1'b0 ;
  assign n12823 = ( n6373 & n12821 ) | ( n6373 & n12822 ) | ( n12821 & n12822 ) ;
  assign n12824 = ( x51 & ~n6373 ) | ( x51 & n12823 ) | ( ~n6373 & n12823 ) ;
  assign n12825 = n12824 ^ n1434 ^ 1'b0 ;
  assign n12826 = ( n1434 & n12824 ) | ( n1434 & n12825 ) | ( n12824 & n12825 ) ;
  assign n12827 = ( x96 & ~n1434 ) | ( x96 & n12826 ) | ( ~n1434 & n12826 ) ;
  assign n12828 = ~x72 & x950 ;
  assign n12829 = ( n9018 & n12827 ) | ( n9018 & n12828 ) | ( n12827 & n12828 ) ;
  assign n12830 = ~n9018 & n12829 ;
  assign n12831 = ( n6395 & n12745 ) | ( n6395 & n12830 ) | ( n12745 & n12830 ) ;
  assign n12832 = ~n12830 & n12831 ;
  assign n12833 = x829 & x1092 ;
  assign n12834 = x122 & n12744 ;
  assign n12835 = ( n12812 & n12833 ) | ( n12812 & n12834 ) | ( n12833 & n12834 ) ;
  assign n12836 = ~n12812 & n12835 ;
  assign n12837 = ( ~n12815 & n12832 ) | ( ~n12815 & n12836 ) | ( n12832 & n12836 ) ;
  assign n12838 = n12815 | n12837 ;
  assign n12839 = n6422 & n12838 ;
  assign n12840 = n1614 & n12746 ;
  assign n12841 = ( x1091 & n12839 ) | ( x1091 & n12840 ) | ( n12839 & n12840 ) ;
  assign n12842 = n12840 ^ n12839 ^ 1'b0 ;
  assign n12843 = ( x1091 & n12841 ) | ( x1091 & n12842 ) | ( n12841 & n12842 ) ;
  assign n12844 = n12753 & ~n12813 ;
  assign n12845 = x120 | n12844 ;
  assign n12846 = n12843 | n12845 ;
  assign n12847 = ( x39 & ~n12805 ) | ( x39 & n12846 ) | ( ~n12805 & n12846 ) ;
  assign n12848 = ~x39 & n12847 ;
  assign n12849 = ~n6798 & n12747 ;
  assign n12850 = n5061 & n12849 ;
  assign n12851 = ~n6867 & n12747 ;
  assign n12852 = ~n5061 & n12851 ;
  assign n12853 = ( n6810 & n12850 ) | ( n6810 & ~n12852 ) | ( n12850 & ~n12852 ) ;
  assign n12854 = ~n12850 & n12853 ;
  assign n12855 = n6810 | n12747 ;
  assign n12856 = ( x299 & n12854 ) | ( x299 & n12855 ) | ( n12854 & n12855 ) ;
  assign n12857 = ~n12854 & n12856 ;
  assign n12858 = n6801 | n12747 ;
  assign n12859 = n5114 & n12849 ;
  assign n12860 = ~n5114 & n12851 ;
  assign n12861 = ( n6801 & n12859 ) | ( n6801 & ~n12860 ) | ( n12859 & ~n12860 ) ;
  assign n12862 = ~n12859 & n12861 ;
  assign n12863 = ( x299 & n12858 ) | ( x299 & ~n12862 ) | ( n12858 & ~n12862 ) ;
  assign n12864 = ~x299 & n12863 ;
  assign n12865 = ( x39 & n12857 ) | ( x39 & n12864 ) | ( n12857 & n12864 ) ;
  assign n12866 = n12864 ^ n12857 ^ 1'b0 ;
  assign n12867 = ( x39 & n12865 ) | ( x39 & n12866 ) | ( n12865 & n12866 ) ;
  assign n12868 = ( ~n1205 & n12848 ) | ( ~n1205 & n12867 ) | ( n12848 & n12867 ) ;
  assign n12869 = ~n1205 & n12868 ;
  assign n12870 = ( ~x87 & n12804 ) | ( ~x87 & n12869 ) | ( n12804 & n12869 ) ;
  assign n12871 = ~x87 & n12870 ;
  assign n12872 = ( ~n12773 & n12789 ) | ( ~n12773 & n12871 ) | ( n12789 & n12871 ) ;
  assign n12873 = ~n12773 & n12872 ;
  assign n12874 = n6782 | n12873 ;
  assign n12875 = ~n6612 & n12874 ;
  assign n12876 = ~n12612 & n12786 ;
  assign n12877 = ~n12611 & n12753 ;
  assign n12878 = n12780 | n12877 ;
  assign n12879 = n12784 & n12878 ;
  assign n12880 = n12876 | n12879 ;
  assign n12881 = ( n12609 & n12775 ) | ( n12609 & n12880 ) | ( n12775 & n12880 ) ;
  assign n12882 = ~n12609 & n12881 ;
  assign n12883 = n12625 & n12747 ;
  assign n12884 = n1994 & ~n12883 ;
  assign n12885 = x100 & ~n12884 ;
  assign n12886 = ~n6824 & n12883 ;
  assign n12887 = n12792 | n12877 ;
  assign n12888 = x120 | n12887 ;
  assign n12889 = ( ~x120 & n12618 ) | ( ~x120 & n12888 ) | ( n12618 & n12888 ) ;
  assign n12890 = n6824 & n12889 ;
  assign n12891 = ( n1994 & ~n12886 ) | ( n1994 & n12890 ) | ( ~n12886 & n12890 ) ;
  assign n12892 = n12886 | n12891 ;
  assign n12893 = n12885 & n12892 ;
  assign n12894 = n12623 & n12814 ;
  assign n12895 = ( x120 & n12843 ) | ( x120 & ~n12894 ) | ( n12843 & ~n12894 ) ;
  assign n12896 = n12894 | n12895 ;
  assign n12897 = x120 & n12712 ;
  assign n12898 = ( x39 & n12896 ) | ( x39 & ~n12897 ) | ( n12896 & ~n12897 ) ;
  assign n12899 = n12898 ^ n12896 ^ 1'b0 ;
  assign n12900 = ( x39 & n12898 ) | ( x39 & ~n12899 ) | ( n12898 & ~n12899 ) ;
  assign n12901 = ~n6458 & n12776 ;
  assign n12902 = n12877 | n12901 ;
  assign n12903 = x120 | n12902 ;
  assign n12904 = ( ~x120 & n12632 ) | ( ~x120 & n12903 ) | ( n12632 & n12903 ) ;
  assign n12905 = n12883 ^ n5083 ^ 1'b0 ;
  assign n12906 = ( n12883 & n12904 ) | ( n12883 & ~n12905 ) | ( n12904 & ~n12905 ) ;
  assign n12907 = n5114 & n12906 ;
  assign n12908 = n12883 ^ n5099 ^ 1'b0 ;
  assign n12909 = ( n12883 & n12904 ) | ( n12883 & n12908 ) | ( n12904 & n12908 ) ;
  assign n12910 = ~n5114 & n12909 ;
  assign n12911 = ( n6801 & n12907 ) | ( n6801 & ~n12910 ) | ( n12907 & ~n12910 ) ;
  assign n12912 = ~n12907 & n12911 ;
  assign n12913 = ~x299 & n12858 ;
  assign n12914 = ( n12650 & n12912 ) | ( n12650 & n12913 ) | ( n12912 & n12913 ) ;
  assign n12915 = ~n12912 & n12914 ;
  assign n12916 = n5061 & n12906 ;
  assign n12917 = ~n5061 & n12909 ;
  assign n12918 = ( n6810 & n12916 ) | ( n6810 & ~n12917 ) | ( n12916 & ~n12917 ) ;
  assign n12919 = ~n12916 & n12918 ;
  assign n12920 = x299 & n12855 ;
  assign n12921 = ( ~n12691 & n12919 ) | ( ~n12691 & n12920 ) | ( n12919 & n12920 ) ;
  assign n12922 = ~n12919 & n12921 ;
  assign n12923 = ( x39 & n12915 ) | ( x39 & ~n12922 ) | ( n12915 & ~n12922 ) ;
  assign n12924 = ~n12915 & n12923 ;
  assign n12925 = ( x38 & n12900 ) | ( x38 & ~n12924 ) | ( n12900 & ~n12924 ) ;
  assign n12926 = n12925 ^ n12900 ^ 1'b0 ;
  assign n12927 = ( x38 & n12925 ) | ( x38 & ~n12926 ) | ( n12925 & ~n12926 ) ;
  assign n12928 = x38 & ~n12883 ;
  assign n12929 = ( x100 & n12927 ) | ( x100 & ~n12928 ) | ( n12927 & ~n12928 ) ;
  assign n12930 = ~x100 & n12929 ;
  assign n12931 = ( ~x87 & n12893 ) | ( ~x87 & n12930 ) | ( n12893 & n12930 ) ;
  assign n12932 = ~x87 & n12931 ;
  assign n12933 = ( ~x75 & n12882 ) | ( ~x75 & n12932 ) | ( n12882 & n12932 ) ;
  assign n12934 = ~x75 & n12933 ;
  assign n12935 = n1207 & ~n12883 ;
  assign n12936 = x75 & ~n12935 ;
  assign n12937 = n12764 | n12877 ;
  assign n12938 = x120 | n12937 ;
  assign n12939 = ( ~x120 & n12669 ) | ( ~x120 & n12938 ) | ( n12669 & n12938 ) ;
  assign n12940 = n12939 ^ n12883 ^ 1'b0 ;
  assign n12941 = ( ~n6412 & n12883 ) | ( ~n6412 & n12940 ) | ( n12883 & n12940 ) ;
  assign n12942 = ( n12939 & ~n12940 ) | ( n12939 & n12941 ) | ( ~n12940 & n12941 ) ;
  assign n12943 = ( n1205 & n1206 ) | ( n1205 & ~n12942 ) | ( n1206 & ~n12942 ) ;
  assign n12944 = n12942 | n12943 ;
  assign n12945 = n12936 & n12944 ;
  assign n12946 = ( n6782 & ~n12934 ) | ( n6782 & n12945 ) | ( ~n12934 & n12945 ) ;
  assign n12947 = n12934 | n12946 ;
  assign n12948 = n12875 ^ n12551 ^ 1'b0 ;
  assign n12949 = ( ~n12551 & n12947 ) | ( ~n12551 & n12948 ) | ( n12947 & n12948 ) ;
  assign n12950 = ( n12551 & n12875 ) | ( n12551 & n12949 ) | ( n12875 & n12949 ) ;
  assign n12951 = n12549 & ~n12746 ;
  assign n12952 = ( n12750 & n12950 ) | ( n12750 & ~n12951 ) | ( n12950 & ~n12951 ) ;
  assign n12953 = ~n12750 & n12952 ;
  assign n12954 = ( ~n12545 & n12743 ) | ( ~n12545 & n12953 ) | ( n12743 & n12953 ) ;
  assign n12955 = ~n12545 & n12954 ;
  assign n12956 = ~n12741 & n12750 ;
  assign n12957 = ~n12955 & n12956 ;
  assign n12958 = ( n12683 & n12955 ) | ( n12683 & ~n12957 ) | ( n12955 & ~n12957 ) ;
  assign n12959 = n1243 | n8748 ;
  assign n12960 = x51 | n12959 ;
  assign n12961 = x100 & ~n12960 ;
  assign n12962 = n2097 | n12961 ;
  assign n12963 = ~n5075 & n12960 ;
  assign n12964 = x51 & x146 ;
  assign n12965 = x51 & ~n5075 ;
  assign n12966 = ~x146 & n12965 ;
  assign n12967 = x161 & ~n12966 ;
  assign n12968 = n12964 | n12967 ;
  assign n12969 = n12963 & ~n12968 ;
  assign n12970 = x299 & ~n12969 ;
  assign n12971 = ~x142 & n12965 ;
  assign n12972 = x144 & ~n12971 ;
  assign n12973 = x51 & x142 ;
  assign n12974 = n12963 & ~n12973 ;
  assign n12975 = ~n12972 & n12974 ;
  assign n12976 = x299 | n12975 ;
  assign n12977 = x232 & n12976 ;
  assign n12978 = ~n12970 & n12977 ;
  assign n12979 = x38 & ~n12978 ;
  assign n12980 = x100 | n12979 ;
  assign n12981 = x38 & n12960 ;
  assign n12982 = x100 | n12981 ;
  assign n12983 = n12980 & n12982 ;
  assign n12984 = n1232 | n8747 ;
  assign n12985 = n11537 | n12984 ;
  assign n12986 = ~x50 & x77 ;
  assign n12987 = ~n1261 & n12986 ;
  assign n12988 = ~n12985 & n12987 ;
  assign n12989 = n1375 | n6387 ;
  assign n12990 = ~x24 & x314 ;
  assign n12991 = ~n12989 & n12990 ;
  assign n12992 = ~n7472 & n12991 ;
  assign n12993 = n12988 & n12992 ;
  assign n12994 = ~n1290 & n12993 ;
  assign n12995 = n1457 | n12985 ;
  assign n12996 = x58 | n12989 ;
  assign n12997 = n7591 | n12996 ;
  assign n12998 = n12995 | n12997 ;
  assign n12999 = x72 & ~n5203 ;
  assign n13000 = ~n12998 & n12999 ;
  assign n13001 = x86 & ~n12995 ;
  assign n13002 = n12988 | n13001 ;
  assign n13003 = n9709 & n13002 ;
  assign n13004 = ~x24 & n10309 ;
  assign n13005 = ~n12995 & n13004 ;
  assign n13006 = ( n12959 & ~n13003 ) | ( n12959 & n13005 ) | ( ~n13003 & n13005 ) ;
  assign n13007 = n13003 | n13006 ;
  assign n13008 = ~x51 & n12959 ;
  assign n13009 = ( x51 & n12989 ) | ( x51 & ~n13008 ) | ( n12989 & ~n13008 ) ;
  assign n13010 = n13007 & ~n13009 ;
  assign n13011 = ~n1290 & n13010 ;
  assign n13012 = n12960 | n13011 ;
  assign n13013 = n13000 | n13012 ;
  assign n13014 = n12994 | n13013 ;
  assign n13015 = n1290 | n12998 ;
  assign n13016 = n5525 | n6462 ;
  assign n13017 = ~n13015 & n13016 ;
  assign n13018 = ( x232 & n12960 ) | ( x232 & ~n13017 ) | ( n12960 & ~n13017 ) ;
  assign n13019 = n13017 | n13018 ;
  assign n13020 = ( n5376 & n12960 ) | ( n5376 & ~n12971 ) | ( n12960 & ~n12971 ) ;
  assign n13021 = x144 & n13020 ;
  assign n13022 = ~n12960 & n13015 ;
  assign n13023 = x51 | n13022 ;
  assign n13024 = ( ~x51 & n12965 ) | ( ~x51 & n13023 ) | ( n12965 & n13023 ) ;
  assign n13025 = n5376 & ~n12973 ;
  assign n13026 = n13021 & ~n13025 ;
  assign n13027 = ( n13021 & ~n13024 ) | ( n13021 & n13026 ) | ( ~n13024 & n13026 ) ;
  assign n13028 = ~x287 & n13023 ;
  assign n13029 = ~n5075 & n13008 ;
  assign n13030 = x287 | n5075 ;
  assign n13031 = ~n13029 & n13030 ;
  assign n13032 = n13028 | n13031 ;
  assign n13033 = ~n12974 & n13032 ;
  assign n13034 = n7678 & ~n13033 ;
  assign n13035 = ~n12959 & n13034 ;
  assign n13036 = n13027 & ~n13035 ;
  assign n13037 = x51 | n13030 ;
  assign n13038 = n1286 | n6399 ;
  assign n13039 = ~x51 & n13038 ;
  assign n13040 = ~n5075 & n13022 ;
  assign n13041 = n5075 | n13022 ;
  assign n13042 = ( n13039 & n13040 ) | ( n13039 & n13041 ) | ( n13040 & n13041 ) ;
  assign n13043 = n13042 ^ n13039 ^ n13022 ;
  assign n13044 = n13037 & ~n13043 ;
  assign n13045 = x224 & ~n12971 ;
  assign n13046 = n13044 & n13045 ;
  assign n13047 = x142 & ~n13043 ;
  assign n13048 = n5075 & ~n13022 ;
  assign n13049 = n5088 & ~n13048 ;
  assign n13050 = x142 | n13049 ;
  assign n13051 = ( n5376 & n13047 ) | ( n5376 & n13050 ) | ( n13047 & n13050 ) ;
  assign n13052 = ~n13047 & n13051 ;
  assign n13053 = ( n7678 & ~n13046 ) | ( n7678 & n13052 ) | ( ~n13046 & n13052 ) ;
  assign n13054 = ~n13046 & n13053 ;
  assign n13055 = ~n5376 & n13029 ;
  assign n13056 = n13020 & ~n13055 ;
  assign n13057 = ( ~n13021 & n13054 ) | ( ~n13021 & n13056 ) | ( n13054 & n13056 ) ;
  assign n13058 = ~n13054 & n13057 ;
  assign n13059 = ( x181 & n13036 ) | ( x181 & ~n13058 ) | ( n13036 & ~n13058 ) ;
  assign n13060 = ~n13036 & n13059 ;
  assign n13061 = ~n13021 & n13056 ;
  assign n13062 = ~n13052 & n13061 ;
  assign n13063 = x181 | n13027 ;
  assign n13064 = n13062 | n13063 ;
  assign n13065 = ( x299 & ~n13060 ) | ( x299 & n13064 ) | ( ~n13060 & n13064 ) ;
  assign n13066 = ~x299 & n13065 ;
  assign n13067 = x146 | n13049 ;
  assign n13068 = x146 & ~n13043 ;
  assign n13069 = ( x161 & n13067 ) | ( x161 & ~n13068 ) | ( n13067 & ~n13068 ) ;
  assign n13070 = ~x161 & n13069 ;
  assign n13071 = n12966 | n13022 ;
  assign n13072 = ( ~x161 & n13069 ) | ( ~x161 & n13071 ) | ( n13069 & n13071 ) ;
  assign n13073 = ( x161 & n13070 ) | ( x161 & n13072 ) | ( n13070 & n13072 ) ;
  assign n13074 = ( x215 & x221 ) | ( x215 & n13073 ) | ( x221 & n13073 ) ;
  assign n13075 = ~x215 & n13074 ;
  assign n13076 = ~x159 & x299 ;
  assign n13077 = n12960 & ~n12969 ;
  assign n13078 = n5390 | n13077 ;
  assign n13079 = n13076 & n13078 ;
  assign n13080 = ~n13075 & n13079 ;
  assign n13081 = x232 & ~n13080 ;
  assign n13082 = x159 & x299 ;
  assign n13083 = ~n13015 & n13030 ;
  assign n13084 = n12960 | n13083 ;
  assign n13085 = n12967 & n13084 ;
  assign n13086 = x161 | n12966 ;
  assign n13087 = n13044 & ~n13086 ;
  assign n13088 = ( x216 & n13085 ) | ( x216 & n13087 ) | ( n13085 & n13087 ) ;
  assign n13089 = n13087 ^ n13085 ^ 1'b0 ;
  assign n13090 = ( x216 & n13088 ) | ( x216 & n13089 ) | ( n13088 & n13089 ) ;
  assign n13091 = ( n7669 & n13075 ) | ( n7669 & ~n13090 ) | ( n13075 & ~n13090 ) ;
  assign n13092 = ~n13090 & n13091 ;
  assign n13093 = n13082 & ~n13092 ;
  assign n13094 = n13078 & n13093 ;
  assign n13095 = ( n13066 & n13081 ) | ( n13066 & ~n13094 ) | ( n13081 & ~n13094 ) ;
  assign n13096 = ~n13066 & n13095 ;
  assign n13097 = x39 & ~n13096 ;
  assign n13098 = n13019 & n13097 ;
  assign n13099 = x39 | x232 ;
  assign n13100 = ~n13098 & n13099 ;
  assign n13101 = ( n13014 & n13098 ) | ( n13014 & ~n13100 ) | ( n13098 & ~n13100 ) ;
  assign n13102 = n5075 | n12960 ;
  assign n13103 = n12960 | n12994 ;
  assign n13104 = n13011 | n13103 ;
  assign n13105 = n5075 & ~n13104 ;
  assign n13106 = n13102 & ~n13105 ;
  assign n13107 = n13000 | n13106 ;
  assign n13108 = n12994 | n13107 ;
  assign n13109 = n12972 & n13108 ;
  assign n13110 = n5075 & n13014 ;
  assign n13111 = x72 & ~n8948 ;
  assign n13112 = n12965 | n13111 ;
  assign n13113 = ~n5075 & n13112 ;
  assign n13114 = n13110 | n13113 ;
  assign n13115 = ~x51 & n12991 ;
  assign n13116 = n11941 & n13115 ;
  assign n13117 = n1290 | n5075 ;
  assign n13118 = n13116 & ~n13117 ;
  assign n13119 = n13114 | n13118 ;
  assign n13120 = x142 & ~n13119 ;
  assign n13121 = n1432 | n5203 ;
  assign n13122 = ( n13111 & n13116 ) | ( n13111 & ~n13121 ) | ( n13116 & ~n13121 ) ;
  assign n13123 = ~n5075 & n13122 ;
  assign n13124 = n13110 | n13123 ;
  assign n13125 = x142 | n13124 ;
  assign n13126 = ( x144 & ~n13120 ) | ( x144 & n13125 ) | ( ~n13120 & n13125 ) ;
  assign n13127 = ~x144 & n13126 ;
  assign n13128 = ( x180 & ~n13109 ) | ( x180 & n13127 ) | ( ~n13109 & n13127 ) ;
  assign n13129 = n13109 | n13128 ;
  assign n13130 = n13114 ^ x144 ^ 1'b0 ;
  assign n13131 = ( n13107 & n13114 ) | ( n13107 & n13130 ) | ( n13114 & n13130 ) ;
  assign n13132 = n13131 ^ n12971 ^ 1'b0 ;
  assign n13133 = ( x180 & n12971 ) | ( x180 & ~n13131 ) | ( n12971 & ~n13131 ) ;
  assign n13134 = ( x180 & ~n13132 ) | ( x180 & n13133 ) | ( ~n13132 & n13133 ) ;
  assign n13135 = x179 & ~n13134 ;
  assign n13136 = n13129 & n13135 ;
  assign n13137 = n10317 ^ x24 ^ 1'b0 ;
  assign n13138 = ( n10310 & n10317 ) | ( n10310 & ~n13137 ) | ( n10317 & ~n13137 ) ;
  assign n13139 = n10317 ^ x314 ^ 1'b0 ;
  assign n13140 = ( n10317 & n13138 ) | ( n10317 & ~n13139 ) | ( n13138 & ~n13139 ) ;
  assign n13141 = ~n1378 & n13140 ;
  assign n13142 = x72 | n13141 ;
  assign n13143 = ~n13121 & n13142 ;
  assign n13144 = ~n5075 & n13143 ;
  assign n13145 = n13110 | n13144 ;
  assign n13146 = x142 | n13145 ;
  assign n13147 = n6387 | n7453 ;
  assign n13148 = n13140 & ~n13147 ;
  assign n13149 = x51 | n13148 ;
  assign n13150 = n13111 | n13149 ;
  assign n13151 = n5075 & ~n13111 ;
  assign n13152 = n13150 & ~n13151 ;
  assign n13153 = n13152 ^ n13114 ^ n13112 ;
  assign n13154 = x142 & ~n13153 ;
  assign n13155 = ( x144 & n13146 ) | ( x144 & ~n13154 ) | ( n13146 & ~n13154 ) ;
  assign n13156 = ~x144 & n13155 ;
  assign n13157 = n12972 & n13014 ;
  assign n13158 = ( x180 & ~n13156 ) | ( x180 & n13157 ) | ( ~n13156 & n13157 ) ;
  assign n13159 = n13156 | n13158 ;
  assign n13160 = ~n1378 & n13138 ;
  assign n13161 = ~n13117 & n13160 ;
  assign n13162 = n13113 | n13161 ;
  assign n13163 = n13110 | n13162 ;
  assign n13164 = x142 & ~n13163 ;
  assign n13165 = x144 | n13164 ;
  assign n13166 = x72 | n13160 ;
  assign n13167 = ~n13121 & n13166 ;
  assign n13168 = ~n5075 & n13167 ;
  assign n13169 = n13110 | n13168 ;
  assign n13170 = ( x142 & ~n13165 ) | ( x142 & n13169 ) | ( ~n13165 & n13169 ) ;
  assign n13171 = ~n13165 & n13170 ;
  assign n13172 = x51 | n5075 ;
  assign n13173 = n13013 & ~n13172 ;
  assign n13174 = n13110 | n13173 ;
  assign n13175 = ~n5075 & n13012 ;
  assign n13176 = n13175 ^ x142 ^ 1'b0 ;
  assign n13177 = ~n13029 & n13117 ;
  assign n13178 = ( n1290 & n13011 ) | ( n1290 & ~n13177 ) | ( n13011 & ~n13177 ) ;
  assign n13179 = ( n13175 & n13176 ) | ( n13175 & n13178 ) | ( n13176 & n13178 ) ;
  assign n13180 = n13106 & ~n13179 ;
  assign n13181 = n13174 | n13180 ;
  assign n13182 = x144 & n13181 ;
  assign n13183 = ( x180 & n13171 ) | ( x180 & ~n13182 ) | ( n13171 & ~n13182 ) ;
  assign n13184 = ~n13171 & n13183 ;
  assign n13185 = ( x179 & n13159 ) | ( x179 & ~n13184 ) | ( n13159 & ~n13184 ) ;
  assign n13186 = ~x179 & n13185 ;
  assign n13187 = ( ~x299 & n13136 ) | ( ~x299 & n13186 ) | ( n13136 & n13186 ) ;
  assign n13188 = ~x299 & n13187 ;
  assign n13189 = x146 | n13145 ;
  assign n13190 = x146 & ~n13153 ;
  assign n13191 = n8048 & ~n13190 ;
  assign n13192 = n13189 & n13191 ;
  assign n13193 = x146 & ~n13163 ;
  assign n13194 = x158 & x299 ;
  assign n13195 = x146 | n13169 ;
  assign n13196 = ( n13193 & n13194 ) | ( n13193 & n13195 ) | ( n13194 & n13195 ) ;
  assign n13197 = ~n13193 & n13196 ;
  assign n13198 = ( x161 & ~n13192 ) | ( x161 & n13197 ) | ( ~n13192 & n13197 ) ;
  assign n13199 = n13192 | n13198 ;
  assign n13200 = n13175 ^ x146 ^ 1'b0 ;
  assign n13201 = ( n13175 & n13178 ) | ( n13175 & n13200 ) | ( n13178 & n13200 ) ;
  assign n13202 = n13106 & ~n13201 ;
  assign n13203 = n13174 | n13202 ;
  assign n13204 = n13194 & n13203 ;
  assign n13205 = n8048 & ~n12966 ;
  assign n13206 = n13014 & n13205 ;
  assign n13207 = ( x161 & n13204 ) | ( x161 & ~n13206 ) | ( n13204 & ~n13206 ) ;
  assign n13208 = ~n13204 & n13207 ;
  assign n13209 = ( x156 & n13199 ) | ( x156 & ~n13208 ) | ( n13199 & ~n13208 ) ;
  assign n13210 = ~x156 & n13209 ;
  assign n13211 = n5075 & ~n13014 ;
  assign n13212 = x146 | n13124 ;
  assign n13213 = x146 & ~n13119 ;
  assign n13214 = ( x161 & n13212 ) | ( x161 & ~n13213 ) | ( n13212 & ~n13213 ) ;
  assign n13215 = ~x161 & n13214 ;
  assign n13216 = n12959 | n13000 ;
  assign n13217 = n13172 | n13216 ;
  assign n13218 = n12994 | n13217 ;
  assign n13219 = ~n12965 & n13218 ;
  assign n13220 = x146 & n12960 ;
  assign n13221 = ( x161 & n13219 ) | ( x161 & n13220 ) | ( n13219 & n13220 ) ;
  assign n13222 = n13220 ^ n13219 ^ 1'b0 ;
  assign n13223 = ( x161 & n13221 ) | ( x161 & n13222 ) | ( n13221 & n13222 ) ;
  assign n13224 = n13211 | n13223 ;
  assign n13225 = ( ~n13211 & n13215 ) | ( ~n13211 & n13224 ) | ( n13215 & n13224 ) ;
  assign n13226 = ( x158 & x299 ) | ( x158 & n13225 ) | ( x299 & n13225 ) ;
  assign n13227 = ~x158 & n13226 ;
  assign n13228 = ~n13172 & n13216 ;
  assign n13229 = x146 | n13228 ;
  assign n13230 = n13110 | n13229 ;
  assign n13231 = ( x161 & n8431 ) | ( x161 & n13107 ) | ( n8431 & n13107 ) ;
  assign n13232 = n13230 & n13231 ;
  assign n13233 = n13086 & ~n13232 ;
  assign n13234 = ( n13114 & n13232 ) | ( n13114 & ~n13233 ) | ( n13232 & ~n13233 ) ;
  assign n13235 = ( ~x158 & x299 ) | ( ~x158 & n13234 ) | ( x299 & n13234 ) ;
  assign n13236 = x158 & n13235 ;
  assign n13237 = ( x156 & n13227 ) | ( x156 & n13236 ) | ( n13227 & n13236 ) ;
  assign n13238 = n13236 ^ n13227 ^ 1'b0 ;
  assign n13239 = ( x156 & n13237 ) | ( x156 & n13238 ) | ( n13237 & n13238 ) ;
  assign n13240 = ( ~n13188 & n13210 ) | ( ~n13188 & n13239 ) | ( n13210 & n13239 ) ;
  assign n13241 = n13188 | n13240 ;
  assign n13242 = n13101 ^ n8156 ^ 1'b0 ;
  assign n13243 = ( ~n8156 & n13241 ) | ( ~n8156 & n13242 ) | ( n13241 & n13242 ) ;
  assign n13244 = ( n8156 & n13101 ) | ( n8156 & n13243 ) | ( n13101 & n13243 ) ;
  assign n13245 = x38 | n13244 ;
  assign n13246 = ( ~x38 & n12983 ) | ( ~x38 & n13245 ) | ( n12983 & n13245 ) ;
  assign n13247 = x100 & n12978 ;
  assign n13248 = ( n12962 & n13246 ) | ( n12962 & ~n13247 ) | ( n13246 & ~n13247 ) ;
  assign n13249 = ~n12962 & n13248 ;
  assign n13250 = x134 | x135 ;
  assign n13251 = x136 | n13250 ;
  assign n13252 = x130 | n13251 ;
  assign n13253 = x132 | n13252 ;
  assign n13254 = x126 | n13253 ;
  assign n13255 = x121 | n13254 ;
  assign n13256 = x125 | x133 ;
  assign n13257 = n13256 ^ x121 ^ 1'b0 ;
  assign n13258 = n13255 & ~n13257 ;
  assign n13259 = ~x163 & x299 ;
  assign n13260 = x184 | x299 ;
  assign n13261 = ~n13259 & n13260 ;
  assign n13262 = x87 & ~n13261 ;
  assign n13263 = ( x87 & ~n6411 ) | ( x87 & n13262 ) | ( ~n6411 & n13262 ) ;
  assign n13264 = n13258 | n13263 ;
  assign n13265 = ~x87 & n2068 ;
  assign n13266 = n12960 & n13265 ;
  assign n13267 = ~n12978 & n13266 ;
  assign n13268 = ( ~n13249 & n13264 ) | ( ~n13249 & n13267 ) | ( n13264 & n13267 ) ;
  assign n13269 = n13249 | n13268 ;
  assign n13270 = x87 | n12960 ;
  assign n13271 = n13258 | n13270 ;
  assign n13272 = x87 & ~n10323 ;
  assign n13273 = x232 & ~n13272 ;
  assign n13274 = x87 | n12969 ;
  assign n13275 = n13273 & n13274 ;
  assign n13276 = n7318 & ~n13275 ;
  assign n13277 = n13271 & n13276 ;
  assign n13278 = ~n12978 & n13265 ;
  assign n13279 = n12972 & ~n13161 ;
  assign n13280 = x144 | n13179 ;
  assign n13281 = ( x180 & ~n13279 ) | ( x180 & n13280 ) | ( ~n13279 & n13280 ) ;
  assign n13282 = ~x180 & n13281 ;
  assign n13283 = ~n5075 & n13104 ;
  assign n13284 = ~x142 & n13283 ;
  assign n13285 = n12959 | n12993 ;
  assign n13286 = ~x51 & n13285 ;
  assign n13287 = ( ~n13009 & n13010 ) | ( ~n13009 & n13286 ) | ( n13010 & n13286 ) ;
  assign n13288 = n1290 | n13287 ;
  assign n13289 = ~n13177 & n13288 ;
  assign n13290 = x142 & n13289 ;
  assign n13291 = ( x144 & ~n13284 ) | ( x144 & n13290 ) | ( ~n13284 & n13290 ) ;
  assign n13292 = n13284 | n13291 ;
  assign n13293 = ~n5075 & n13149 ;
  assign n13294 = ~n12973 & n13293 ;
  assign n13295 = x144 & ~n13294 ;
  assign n13296 = x180 & ~n13295 ;
  assign n13297 = n13292 & n13296 ;
  assign n13298 = ( x179 & n13282 ) | ( x179 & ~n13297 ) | ( n13282 & ~n13297 ) ;
  assign n13299 = ~n13282 & n13298 ;
  assign n13300 = ~n5075 & n13103 ;
  assign n13301 = ~x142 & n13300 ;
  assign n13302 = n1290 | n13286 ;
  assign n13303 = ~n13177 & n13302 ;
  assign n13304 = x142 & n13303 ;
  assign n13305 = ( x144 & ~n13301 ) | ( x144 & n13304 ) | ( ~n13301 & n13304 ) ;
  assign n13306 = n13301 | n13305 ;
  assign n13307 = n12972 & ~n13118 ;
  assign n13308 = x180 & ~n13307 ;
  assign n13309 = n13306 & n13308 ;
  assign n13310 = ~x180 & n12975 ;
  assign n13311 = ( x179 & ~n13309 ) | ( x179 & n13310 ) | ( ~n13309 & n13310 ) ;
  assign n13312 = n13309 | n13311 ;
  assign n13313 = n13312 ^ n13299 ^ 1'b0 ;
  assign n13314 = ( n13299 & n13312 ) | ( n13299 & n13313 ) | ( n13312 & n13313 ) ;
  assign n13315 = ( x299 & ~n13299 ) | ( x299 & n13314 ) | ( ~n13299 & n13314 ) ;
  assign n13316 = x144 | n12974 ;
  assign n13317 = n13034 | n13316 ;
  assign n13318 = ~x142 & n13038 ;
  assign n13319 = n7678 & ~n13030 ;
  assign n13320 = x142 & n1292 ;
  assign n13321 = ( n13318 & n13319 ) | ( n13318 & ~n13320 ) | ( n13319 & ~n13320 ) ;
  assign n13322 = ~n13318 & n13321 ;
  assign n13323 = ( x144 & n12971 ) | ( x144 & ~n13322 ) | ( n12971 & ~n13322 ) ;
  assign n13324 = ~n12971 & n13323 ;
  assign n13325 = x181 & ~n13324 ;
  assign n13326 = n13317 & n13325 ;
  assign n13327 = ~x181 & n12975 ;
  assign n13328 = ( x299 & ~n13326 ) | ( x299 & n13327 ) | ( ~n13326 & n13327 ) ;
  assign n13329 = n13326 | n13328 ;
  assign n13330 = n13329 ^ x38 ^ 1'b0 ;
  assign n13331 = ~x159 & n12970 ;
  assign n13332 = n13032 & ~n13086 ;
  assign n13333 = n5075 | n5362 ;
  assign n13334 = n12967 & n13333 ;
  assign n13335 = ( n7669 & n13332 ) | ( n7669 & ~n13334 ) | ( n13332 & ~n13334 ) ;
  assign n13336 = ~n13332 & n13335 ;
  assign n13337 = ~n7669 & n12969 ;
  assign n13338 = ( n13082 & n13336 ) | ( n13082 & ~n13337 ) | ( n13336 & ~n13337 ) ;
  assign n13339 = ~n13336 & n13338 ;
  assign n13340 = ( n8901 & n13331 ) | ( n8901 & ~n13339 ) | ( n13331 & ~n13339 ) ;
  assign n13341 = ~n13331 & n13340 ;
  assign n13342 = ( n13329 & ~n13330 ) | ( n13329 & n13341 ) | ( ~n13330 & n13341 ) ;
  assign n13343 = ( x38 & n13330 ) | ( x38 & n13342 ) | ( n13330 & n13342 ) ;
  assign n13344 = ~n12964 & n13293 ;
  assign n13345 = x161 & ~n13344 ;
  assign n13346 = x146 & n13289 ;
  assign n13347 = ~x146 & n13283 ;
  assign n13348 = x161 | n13347 ;
  assign n13349 = ( ~n13345 & n13346 ) | ( ~n13345 & n13348 ) | ( n13346 & n13348 ) ;
  assign n13350 = ~n13345 & n13349 ;
  assign n13351 = ( x158 & x299 ) | ( x158 & n13350 ) | ( x299 & n13350 ) ;
  assign n13352 = ~n13350 & n13351 ;
  assign n13353 = n12967 & ~n13161 ;
  assign n13354 = x161 | n13201 ;
  assign n13355 = n8048 & ~n13354 ;
  assign n13356 = ( n8048 & n13353 ) | ( n8048 & n13355 ) | ( n13353 & n13355 ) ;
  assign n13357 = ( x232 & n13352 ) | ( x232 & ~n13356 ) | ( n13352 & ~n13356 ) ;
  assign n13358 = ~n13352 & n13357 ;
  assign n13359 = ( x39 & x156 ) | ( x39 & ~n13358 ) | ( x156 & ~n13358 ) ;
  assign n13360 = n13359 ^ x156 ^ 1'b0 ;
  assign n13361 = ( x39 & n13359 ) | ( x39 & ~n13360 ) | ( n13359 & ~n13360 ) ;
  assign n13362 = ~n13343 & n13361 ;
  assign n13363 = ( n13315 & n13343 ) | ( n13315 & ~n13362 ) | ( n13343 & ~n13362 ) ;
  assign n13364 = ~x158 & n12970 ;
  assign n13365 = n12967 & ~n13118 ;
  assign n13366 = x146 & n13303 ;
  assign n13367 = ~x146 & n13300 ;
  assign n13368 = ( x161 & ~n13366 ) | ( x161 & n13367 ) | ( ~n13366 & n13367 ) ;
  assign n13369 = n13366 | n13368 ;
  assign n13370 = n13194 & ~n13369 ;
  assign n13371 = ( n13194 & n13365 ) | ( n13194 & n13370 ) | ( n13365 & n13370 ) ;
  assign n13372 = ( x232 & n13364 ) | ( x232 & ~n13371 ) | ( n13364 & ~n13371 ) ;
  assign n13373 = ~n13364 & n13372 ;
  assign n13374 = ( x156 & n1994 ) | ( x156 & ~n13373 ) | ( n1994 & ~n13373 ) ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = ( n12980 & n13363 ) | ( n12980 & n13375 ) | ( n13363 & n13375 ) ;
  assign n13377 = ~n12980 & n13376 ;
  assign n13378 = ( n2097 & n13247 ) | ( n2097 & ~n13377 ) | ( n13247 & ~n13377 ) ;
  assign n13379 = n13377 | n13378 ;
  assign n13380 = n13258 & ~n13263 ;
  assign n13381 = ( n13278 & n13379 ) | ( n13278 & n13380 ) | ( n13379 & n13380 ) ;
  assign n13382 = ~n13278 & n13381 ;
  assign n13383 = ( x57 & n5193 ) | ( x57 & ~n13382 ) | ( n5193 & ~n13382 ) ;
  assign n13384 = n13382 | n13383 ;
  assign n13385 = ~n13277 & n13384 ;
  assign n13386 = ( n13269 & n13277 ) | ( n13269 & ~n13385 ) | ( n13277 & ~n13385 ) ;
  assign n13387 = ~n6782 & n12732 ;
  assign n13388 = n6612 | n13387 ;
  assign n13389 = ( n6782 & n12548 ) | ( n6782 & n12722 ) | ( n12548 & n12722 ) ;
  assign n13390 = ( n7318 & n13388 ) | ( n7318 & ~n13389 ) | ( n13388 & ~n13389 ) ;
  assign n13391 = ~n7318 & n13390 ;
  assign n13392 = n13391 ^ n11179 ^ 1'b0 ;
  assign n13393 = ( n7437 & ~n11179 ) | ( n7437 & n13392 ) | ( ~n11179 & n13392 ) ;
  assign n13394 = ( n11179 & n13391 ) | ( n11179 & n13393 ) | ( n13391 & n13393 ) ;
  assign n13395 = x110 & n8672 ;
  assign n13396 = n5035 & ~n9595 ;
  assign n13397 = n13395 & n13396 ;
  assign n13398 = ( x39 & n7318 ) | ( x39 & n13397 ) | ( n7318 & n13397 ) ;
  assign n13399 = n7318 & n13398 ;
  assign n13400 = ~x110 & n7673 ;
  assign n13401 = n5115 & n6462 ;
  assign n13402 = x39 & ~n13401 ;
  assign n13403 = ( x39 & ~n13400 ) | ( x39 & n13402 ) | ( ~n13400 & n13402 ) ;
  assign n13404 = n5100 & n5390 ;
  assign n13405 = n13400 & n13404 ;
  assign n13406 = ( x299 & ~n13403 ) | ( x299 & n13405 ) | ( ~n13403 & n13405 ) ;
  assign n13407 = n13406 ^ n13403 ^ 1'b0 ;
  assign n13408 = ( n13403 & ~n13406 ) | ( n13403 & n13407 ) | ( ~n13406 & n13407 ) ;
  assign n13409 = n5209 | n10084 ;
  assign n13410 = x36 | n1519 ;
  assign n13411 = x111 | n5215 ;
  assign n13412 = n13411 ^ n13410 ^ 1'b0 ;
  assign n13413 = ( n13410 & n13411 ) | ( n13410 & n13412 ) | ( n13411 & n13412 ) ;
  assign n13414 = ( n1233 & ~n13410 ) | ( n1233 & n13413 ) | ( ~n13410 & n13413 ) ;
  assign n13415 = ( n1482 & ~n1486 ) | ( n1482 & n13414 ) | ( ~n1486 & n13414 ) ;
  assign n13416 = ~n1482 & n13415 ;
  assign n13417 = x83 | n13416 ;
  assign n13418 = ~n1483 & n13417 ;
  assign n13419 = x71 | n13418 ;
  assign n13420 = ~n5226 & n13419 ;
  assign n13421 = x81 | n13420 ;
  assign n13422 = ~n13409 & n13421 ;
  assign n13423 = x90 | n13422 ;
  assign n13424 = ~n1377 & n13423 ;
  assign n13425 = ~n1441 & n13424 ;
  assign n13426 = x72 | n13425 ;
  assign n13427 = n11943 | n13121 ;
  assign n13428 = ( x39 & n13426 ) | ( x39 & ~n13427 ) | ( n13426 & ~n13427 ) ;
  assign n13429 = n13428 ^ n13426 ^ 1'b0 ;
  assign n13430 = ( x39 & n13428 ) | ( x39 & ~n13429 ) | ( n13428 & ~n13429 ) ;
  assign n13431 = x72 & ~n1378 ;
  assign n13432 = ~n8965 & n13431 ;
  assign n13433 = x90 & n8965 ;
  assign n13434 = n8101 | n13433 ;
  assign n13435 = n13424 & ~n13434 ;
  assign n13436 = ( ~n5203 & n13432 ) | ( ~n5203 & n13435 ) | ( n13432 & n13435 ) ;
  assign n13437 = ~n5203 & n13436 ;
  assign n13438 = ( x110 & n11943 ) | ( x110 & n13437 ) | ( n11943 & n13437 ) ;
  assign n13439 = n11943 & n13438 ;
  assign n13440 = ( ~n13408 & n13430 ) | ( ~n13408 & n13439 ) | ( n13430 & n13439 ) ;
  assign n13441 = ~n13408 & n13440 ;
  assign n13442 = ( x38 & n2069 ) | ( x38 & ~n13441 ) | ( n2069 & ~n13441 ) ;
  assign n13443 = n13441 | n13442 ;
  assign n13444 = x110 & n11943 ;
  assign n13445 = x39 | n13444 ;
  assign n13446 = ~n13408 & n13445 ;
  assign n13447 = ( x38 & n2069 ) | ( x38 & ~n13446 ) | ( n2069 & ~n13446 ) ;
  assign n13448 = ~n13446 & n13447 ;
  assign n13449 = ( n7318 & n13443 ) | ( n7318 & ~n13448 ) | ( n13443 & ~n13448 ) ;
  assign n13450 = ~n7318 & n13449 ;
  assign n13451 = x39 & ~n13405 ;
  assign n13452 = ~n13450 & n13451 ;
  assign n13453 = ( n13399 & n13450 ) | ( n13399 & ~n13452 ) | ( n13450 & ~n13452 ) ;
  assign n13454 = x87 & n6411 ;
  assign n13455 = x162 & n13454 ;
  assign n13456 = n7318 & ~n13455 ;
  assign n13457 = x125 | n13255 ;
  assign n13458 = x133 ^ x125 ^ 1'b0 ;
  assign n13459 = n13457 & ~n13458 ;
  assign n13460 = x162 & x299 ;
  assign n13461 = x140 & ~x299 ;
  assign n13462 = n13460 | n13461 ;
  assign n13463 = x87 & ~n13462 ;
  assign n13464 = ( x87 & ~n6411 ) | ( x87 & n13463 ) | ( ~n6411 & n13463 ) ;
  assign n13465 = n13459 & ~n13464 ;
  assign n13466 = x193 & n12965 ;
  assign n13467 = x299 | n13466 ;
  assign n13468 = ~x174 & n13029 ;
  assign n13469 = ( x232 & n13467 ) | ( x232 & n13468 ) | ( n13467 & n13468 ) ;
  assign n13470 = n13468 ^ n13467 ^ 1'b0 ;
  assign n13471 = ( x232 & n13469 ) | ( x232 & n13470 ) | ( n13469 & n13470 ) ;
  assign n13472 = x172 & n12965 ;
  assign n13473 = ~x152 & n13029 ;
  assign n13474 = n13472 | n13473 ;
  assign n13475 = n13474 ^ n13471 ^ 1'b0 ;
  assign n13476 = ( ~x299 & n13474 ) | ( ~x299 & n13475 ) | ( n13474 & n13475 ) ;
  assign n13477 = ( n13471 & ~n13475 ) | ( n13471 & n13476 ) | ( ~n13475 & n13476 ) ;
  assign n13478 = n13265 & ~n13477 ;
  assign n13479 = n13465 & ~n13478 ;
  assign n13480 = x100 & n13477 ;
  assign n13481 = x38 & ~n13477 ;
  assign n13482 = x100 | n13481 ;
  assign n13483 = ~n5390 & n13474 ;
  assign n13484 = x51 & ~x172 ;
  assign n13489 = x152 | n5075 ;
  assign n13490 = ~n13022 & n13489 ;
  assign n13485 = n5075 | n13039 ;
  assign n13488 = x152 | n13485 ;
  assign n13491 = n13490 ^ n13488 ^ 1'b0 ;
  assign n13486 = n1292 & n5075 ;
  assign n13487 = n13486 ^ n13485 ^ n5075 ;
  assign n13492 = n13491 ^ n13487 ^ n13022 ;
  assign n13493 = ( ~x216 & n13484 ) | ( ~x216 & n13492 ) | ( n13484 & n13492 ) ;
  assign n13494 = ~x216 & n13493 ;
  assign n13495 = n13015 | n13030 ;
  assign n13496 = ~n12963 & n13495 ;
  assign n13497 = ~x152 & n13496 ;
  assign n13498 = n13030 | n13038 ;
  assign n13499 = ~n12965 & n13498 ;
  assign n13500 = x152 & n13499 ;
  assign n13501 = ( x172 & n13497 ) | ( x172 & ~n13500 ) | ( n13497 & ~n13500 ) ;
  assign n13502 = ~n13497 & n13501 ;
  assign n13503 = x152 & n13333 ;
  assign n13504 = ~x152 & n13032 ;
  assign n13505 = ( x172 & ~n13503 ) | ( x172 & n13504 ) | ( ~n13503 & n13504 ) ;
  assign n13506 = n13503 | n13505 ;
  assign n13507 = ( x216 & n13502 ) | ( x216 & n13506 ) | ( n13502 & n13506 ) ;
  assign n13508 = ~n13502 & n13507 ;
  assign n13509 = ( n5390 & n13494 ) | ( n5390 & ~n13508 ) | ( n13494 & ~n13508 ) ;
  assign n13510 = ~n13494 & n13509 ;
  assign n13511 = ( n13194 & n13483 ) | ( n13194 & ~n13510 ) | ( n13483 & ~n13510 ) ;
  assign n13512 = ~n13483 & n13511 ;
  assign n13513 = n5390 & n13494 ;
  assign n13514 = n6810 | n13474 ;
  assign n13515 = ~n13513 & n13514 ;
  assign n13516 = ~n13512 & n13515 ;
  assign n13517 = ( n8048 & n13512 ) | ( n8048 & ~n13516 ) | ( n13512 & ~n13516 ) ;
  assign n13518 = n6801 | n13319 ;
  assign n13519 = ~n1292 & n13518 ;
  assign n13520 = x174 & n13519 ;
  assign n13521 = x224 & n13032 ;
  assign n13522 = n5376 & ~n13521 ;
  assign n13523 = ~n5075 & n13023 ;
  assign n13524 = n13486 | n13523 ;
  assign n13525 = ~x224 & n13524 ;
  assign n13526 = ( n13055 & n13522 ) | ( n13055 & ~n13525 ) | ( n13522 & ~n13525 ) ;
  assign n13527 = n13526 ^ n13522 ^ 1'b0 ;
  assign n13528 = ( n13055 & n13526 ) | ( n13055 & ~n13527 ) | ( n13526 & ~n13527 ) ;
  assign n13529 = ~x174 & n13528 ;
  assign n13530 = ( x193 & ~n13520 ) | ( x193 & n13529 ) | ( ~n13520 & n13529 ) ;
  assign n13531 = n13520 | n13530 ;
  assign n13532 = n13040 | n13486 ;
  assign n13533 = n6801 & n13532 ;
  assign n13534 = x224 & n13495 ;
  assign n13535 = n5376 & ~n13534 ;
  assign n13536 = ( n12963 & ~n13533 ) | ( n12963 & n13535 ) | ( ~n13533 & n13535 ) ;
  assign n13537 = ~n13533 & n13536 ;
  assign n13538 = ~x174 & n13537 ;
  assign n13539 = x224 & n13499 ;
  assign n13540 = n5376 & ~n13539 ;
  assign n13541 = n6801 & n13487 ;
  assign n13542 = n13540 & ~n13541 ;
  assign n13543 = n12965 | n13542 ;
  assign n13544 = x174 & n13543 ;
  assign n13545 = ( x193 & n13538 ) | ( x193 & ~n13544 ) | ( n13538 & ~n13544 ) ;
  assign n13546 = ~n13538 & n13545 ;
  assign n13547 = x180 & ~n13546 ;
  assign n13548 = n13531 & n13547 ;
  assign n13549 = ~n1292 & n6801 ;
  assign n13550 = x174 & n13549 ;
  assign n13551 = n13466 | n13550 ;
  assign n13552 = n6801 | n12963 ;
  assign n13553 = ~n13524 & n13552 ;
  assign n13554 = ~x174 & n13553 ;
  assign n13555 = ( ~x180 & n13551 ) | ( ~x180 & n13554 ) | ( n13551 & n13554 ) ;
  assign n13556 = ~x180 & n13555 ;
  assign n13557 = ( x299 & ~n13548 ) | ( x299 & n13556 ) | ( ~n13548 & n13556 ) ;
  assign n13558 = n13548 | n13557 ;
  assign n13559 = x232 & ~n13558 ;
  assign n13560 = ( x232 & n13517 ) | ( x232 & n13559 ) | ( n13517 & n13559 ) ;
  assign n13561 = ( n6463 & n6466 ) | ( n6463 & n13016 ) | ( n6466 & n13016 ) ;
  assign n13562 = ~n1292 & n13561 ;
  assign n13563 = x232 | n13562 ;
  assign n13564 = ( x39 & n13560 ) | ( x39 & n13563 ) | ( n13560 & n13563 ) ;
  assign n13565 = ~n13560 & n13564 ;
  assign n13566 = x232 | n13111 ;
  assign n13567 = ~x39 & n13566 ;
  assign n13568 = ( x38 & ~n13565 ) | ( x38 & n13567 ) | ( ~n13565 & n13567 ) ;
  assign n13569 = n13565 | n13568 ;
  assign n13574 = n5075 & n13111 ;
  assign n13593 = n13173 | n13574 ;
  assign n13594 = ~x152 & n13593 ;
  assign n13595 = n13168 | n13574 ;
  assign n13596 = x152 & n13595 ;
  assign n13597 = ( x172 & ~n13594 ) | ( x172 & n13596 ) | ( ~n13594 & n13596 ) ;
  assign n13598 = n13594 | n13597 ;
  assign n13599 = n13112 | n13161 ;
  assign n13600 = x152 & n13599 ;
  assign n13601 = n13013 | n13217 ;
  assign n13602 = ~n13151 & n13601 ;
  assign n13603 = ~x152 & n13602 ;
  assign n13604 = ( x172 & n13600 ) | ( x172 & ~n13603 ) | ( n13600 & ~n13603 ) ;
  assign n13605 = ~n13600 & n13604 ;
  assign n13606 = ( x197 & n13598 ) | ( x197 & ~n13605 ) | ( n13598 & ~n13605 ) ;
  assign n13607 = ~x197 & n13606 ;
  assign n13584 = n13172 & ~n13574 ;
  assign n13608 = n5075 | n13014 ;
  assign n13609 = ~n13584 & n13608 ;
  assign n13610 = x152 | n13472 ;
  assign n13611 = n13609 | n13610 ;
  assign n13612 = x172 & n13152 ;
  assign n13613 = n13144 | n13574 ;
  assign n13614 = ~x172 & n13613 ;
  assign n13615 = ( x152 & n13612 ) | ( x152 & ~n13614 ) | ( n13612 & ~n13614 ) ;
  assign n13616 = ~n13612 & n13615 ;
  assign n13617 = x197 & ~n13616 ;
  assign n13618 = n13611 & n13617 ;
  assign n13619 = ( n8465 & n13607 ) | ( n8465 & ~n13618 ) | ( n13607 & ~n13618 ) ;
  assign n13620 = ~n13607 & n13619 ;
  assign n13570 = n12965 | n13118 ;
  assign n13571 = n13111 | n13570 ;
  assign n13572 = x172 & n13571 ;
  assign n13573 = x152 & x197 ;
  assign n13575 = n13123 | n13574 ;
  assign n13576 = ~x172 & n13575 ;
  assign n13577 = ( n13572 & n13573 ) | ( n13572 & ~n13576 ) | ( n13573 & ~n13576 ) ;
  assign n13578 = ~n13572 & n13577 ;
  assign n13579 = n13111 & n13489 ;
  assign n13580 = ~x152 & n13228 ;
  assign n13581 = ( x197 & ~n13579 ) | ( x197 & n13580 ) | ( ~n13579 & n13580 ) ;
  assign n13582 = n13579 | n13581 ;
  assign n13585 = n13218 & ~n13584 ;
  assign n13583 = ~x152 & x197 ;
  assign n13586 = n13585 ^ n13583 ^ 1'b0 ;
  assign n13587 = ( n13582 & ~n13583 ) | ( n13582 & n13585 ) | ( ~n13583 & n13585 ) ;
  assign n13588 = ( n13582 & ~n13586 ) | ( n13582 & n13587 ) | ( ~n13586 & n13587 ) ;
  assign n13589 = ( n13472 & ~n13578 ) | ( n13472 & n13588 ) | ( ~n13578 & n13588 ) ;
  assign n13590 = ~n13578 & n13589 ;
  assign n13591 = ( x38 & x155 ) | ( x38 & ~n13590 ) | ( x155 & ~n13590 ) ;
  assign n13592 = n13590 | n13591 ;
  assign n13621 = n13620 ^ n13592 ^ 1'b0 ;
  assign n13622 = ( x299 & ~n13592 ) | ( x299 & n13620 ) | ( ~n13592 & n13620 ) ;
  assign n13623 = ( x299 & ~n13621 ) | ( x299 & n13622 ) | ( ~n13621 & n13622 ) ;
  assign n13624 = ~x193 & n13593 ;
  assign n13625 = x193 & n13602 ;
  assign n13626 = ( x145 & ~n13624 ) | ( x145 & n13625 ) | ( ~n13624 & n13625 ) ;
  assign n13627 = n13624 | n13626 ;
  assign n13628 = x145 & ~n13466 ;
  assign n13629 = ~n13609 & n13628 ;
  assign n13630 = ( x174 & n13627 ) | ( x174 & ~n13629 ) | ( n13627 & ~n13629 ) ;
  assign n13631 = ~x174 & n13630 ;
  assign n13632 = ~x145 & n13599 ;
  assign n13633 = x145 & n13152 ;
  assign n13634 = ( x193 & n13632 ) | ( x193 & ~n13633 ) | ( n13632 & ~n13633 ) ;
  assign n13635 = ~n13632 & n13634 ;
  assign n13636 = x145 & n13613 ;
  assign n13637 = ~x145 & n13595 ;
  assign n13638 = ( x193 & ~n13636 ) | ( x193 & n13637 ) | ( ~n13636 & n13637 ) ;
  assign n13639 = n13636 | n13638 ;
  assign n13640 = ( x174 & n13635 ) | ( x174 & n13639 ) | ( n13635 & n13639 ) ;
  assign n13641 = ~n13635 & n13640 ;
  assign n13642 = ( n8456 & n13631 ) | ( n8456 & ~n13641 ) | ( n13631 & ~n13641 ) ;
  assign n13643 = ~n13631 & n13642 ;
  assign n13644 = n13118 ^ x145 ^ 1'b0 ;
  assign n13645 = ( x145 & n12965 ) | ( x145 & ~n13644 ) | ( n12965 & ~n13644 ) ;
  assign n13646 = ( x174 & n13111 ) | ( x174 & n13645 ) | ( n13111 & n13645 ) ;
  assign n13647 = n13645 ^ n13111 ^ 1'b0 ;
  assign n13648 = ( x174 & n13646 ) | ( x174 & n13647 ) | ( n13646 & n13647 ) ;
  assign n13649 = n12965 | n12994 ;
  assign n13650 = x145 & n13649 ;
  assign n13651 = n13217 | n13650 ;
  assign n13652 = ( x174 & ~n13151 ) | ( x174 & n13651 ) | ( ~n13151 & n13651 ) ;
  assign n13653 = ~x174 & n13652 ;
  assign n13654 = ( x193 & n13648 ) | ( x193 & ~n13653 ) | ( n13648 & ~n13653 ) ;
  assign n13655 = ~n13648 & n13654 ;
  assign n13656 = x145 & n13575 ;
  assign n13657 = ~x145 & n13111 ;
  assign n13658 = ( x174 & n13656 ) | ( x174 & ~n13657 ) | ( n13656 & ~n13657 ) ;
  assign n13659 = ~n13656 & n13658 ;
  assign n13660 = n13228 | n13574 ;
  assign n13661 = ~x145 & n13660 ;
  assign n13662 = x174 | n13661 ;
  assign n13663 = x145 & n13585 ;
  assign n13664 = ( ~n13659 & n13662 ) | ( ~n13659 & n13663 ) | ( n13662 & n13663 ) ;
  assign n13665 = ~n13659 & n13664 ;
  assign n13666 = ( x193 & ~n13655 ) | ( x193 & n13665 ) | ( ~n13655 & n13665 ) ;
  assign n13667 = ~n13655 & n13666 ;
  assign n13668 = ( x177 & x299 ) | ( x177 & ~n13667 ) | ( x299 & ~n13667 ) ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = n13669 ^ n13643 ^ 1'b0 ;
  assign n13671 = ( n13643 & n13669 ) | ( n13643 & n13670 ) | ( n13669 & n13670 ) ;
  assign n13672 = ( x38 & ~n13643 ) | ( x38 & n13671 ) | ( ~n13643 & n13671 ) ;
  assign n13673 = n8156 & ~n13672 ;
  assign n13674 = ( n8156 & n13623 ) | ( n8156 & n13673 ) | ( n13623 & n13673 ) ;
  assign n13675 = ( n13482 & n13569 ) | ( n13482 & ~n13674 ) | ( n13569 & ~n13674 ) ;
  assign n13676 = ~n13482 & n13675 ;
  assign n13677 = ( n2097 & ~n13480 ) | ( n2097 & n13676 ) | ( ~n13480 & n13676 ) ;
  assign n13678 = n13480 | n13677 ;
  assign n13679 = n13479 & n13678 ;
  assign n13680 = n13266 & ~n13477 ;
  assign n13681 = n12982 & n13482 ;
  assign n13682 = n5075 & n13104 ;
  assign n13683 = n13161 | n13682 ;
  assign n13684 = ~x152 & n13683 ;
  assign n13685 = n13178 | n13682 ;
  assign n13686 = x172 & ~n13685 ;
  assign n13687 = ( n12960 & n13102 ) | ( n12960 & n13103 ) | ( n13102 & n13103 ) ;
  assign n13688 = n13011 | n13687 ;
  assign n13689 = x172 | n13688 ;
  assign n13690 = ( x152 & n13686 ) | ( x152 & n13689 ) | ( n13686 & n13689 ) ;
  assign n13691 = ~n13686 & n13690 ;
  assign n13692 = ~x172 & n12965 ;
  assign n13693 = x197 & ~n13692 ;
  assign n13694 = ( n13684 & ~n13691 ) | ( n13684 & n13693 ) | ( ~n13691 & n13693 ) ;
  assign n13695 = ~n13684 & n13694 ;
  assign n13696 = n13289 | n13682 ;
  assign n13697 = x152 & n13696 ;
  assign n13698 = ~n13117 & n13141 ;
  assign n13699 = n13682 | n13698 ;
  assign n13700 = ~x152 & n13699 ;
  assign n13701 = ( x172 & n13697 ) | ( x172 & ~n13700 ) | ( n13697 & ~n13700 ) ;
  assign n13702 = ~n13697 & n13701 ;
  assign n13703 = ~x152 & n13293 ;
  assign n13704 = n13104 & n13489 ;
  assign n13705 = ( x172 & ~n13703 ) | ( x172 & n13704 ) | ( ~n13703 & n13704 ) ;
  assign n13706 = n13703 | n13705 ;
  assign n13707 = n13706 ^ n13702 ^ 1'b0 ;
  assign n13708 = ( n13702 & n13706 ) | ( n13702 & n13707 ) | ( n13706 & n13707 ) ;
  assign n13709 = ( x197 & ~n13702 ) | ( x197 & n13708 ) | ( ~n13702 & n13708 ) ;
  assign n13710 = x299 & ~n8474 ;
  assign n13711 = ( n13695 & n13709 ) | ( n13695 & n13710 ) | ( n13709 & n13710 ) ;
  assign n13712 = ~n13695 & n13711 ;
  assign n13713 = x145 | n13699 ;
  assign n13714 = x145 & ~n13683 ;
  assign n13715 = x174 | n13714 ;
  assign n13716 = n13713 & ~n13715 ;
  assign n13717 = ~x145 & n13103 ;
  assign n13718 = n13688 | n13717 ;
  assign n13719 = n1290 | n13718 ;
  assign n13720 = x174 & n13696 ;
  assign n13721 = n13719 & n13720 ;
  assign n13722 = ( x193 & n13716 ) | ( x193 & ~n13721 ) | ( n13716 & ~n13721 ) ;
  assign n13723 = ~n13716 & n13722 ;
  assign n13724 = x174 & n13718 ;
  assign n13725 = ~x51 & n13714 ;
  assign n13726 = x174 | n13725 ;
  assign n13727 = x145 | n13682 ;
  assign n13728 = ( n13293 & ~n13726 ) | ( n13293 & n13727 ) | ( ~n13726 & n13727 ) ;
  assign n13729 = ~n13726 & n13728 ;
  assign n13730 = ( x193 & ~n13724 ) | ( x193 & n13729 ) | ( ~n13724 & n13729 ) ;
  assign n13731 = n13724 | n13730 ;
  assign n13732 = ( n8450 & ~n13723 ) | ( n8450 & n13731 ) | ( ~n13723 & n13731 ) ;
  assign n13733 = ~n8450 & n13732 ;
  assign n13734 = ( n13103 & n13104 ) | ( n13103 & n13682 ) | ( n13104 & n13682 ) ;
  assign n13735 = x174 & ~n13734 ;
  assign n13736 = ~n13105 & n13172 ;
  assign n13737 = ~x145 & n13118 ;
  assign n13738 = x174 | n13737 ;
  assign n13739 = x145 & ~n12959 ;
  assign n13740 = n13738 & ~n13739 ;
  assign n13741 = n13736 | n13740 ;
  assign n13742 = n13741 ^ n13735 ^ 1'b0 ;
  assign n13743 = ( n13735 & n13741 ) | ( n13735 & n13742 ) | ( n13741 & n13742 ) ;
  assign n13744 = ( x193 & ~n13735 ) | ( x193 & n13743 ) | ( ~n13735 & n13743 ) ;
  assign n13745 = ~x145 & x174 ;
  assign n13746 = ~n13303 & n13745 ;
  assign n13747 = x145 & ~n13029 ;
  assign n13748 = ( n13738 & n13746 ) | ( n13738 & ~n13747 ) | ( n13746 & ~n13747 ) ;
  assign n13749 = ~n13746 & n13748 ;
  assign n13750 = ( x193 & n13682 ) | ( x193 & ~n13749 ) | ( n13682 & ~n13749 ) ;
  assign n13751 = ~n13682 & n13750 ;
  assign n13752 = n8456 & ~n13751 ;
  assign n13753 = n13744 & n13752 ;
  assign n13754 = ( ~x38 & n13733 ) | ( ~x38 & n13753 ) | ( n13733 & n13753 ) ;
  assign n13755 = ~x38 & n13754 ;
  assign n13756 = n13303 | n13682 ;
  assign n13757 = x152 & ~n13756 ;
  assign n13758 = n13118 | n13682 ;
  assign n13759 = x152 | n13758 ;
  assign n13760 = ( x172 & n13757 ) | ( x172 & n13759 ) | ( n13757 & n13759 ) ;
  assign n13761 = ~n13757 & n13760 ;
  assign n13762 = x152 & ~n13734 ;
  assign n13763 = x172 | n13762 ;
  assign n13764 = ( n12965 & n13759 ) | ( n12965 & ~n13763 ) | ( n13759 & ~n13763 ) ;
  assign n13765 = ~n13763 & n13764 ;
  assign n13766 = ( x197 & ~n13761 ) | ( x197 & n13765 ) | ( ~n13761 & n13765 ) ;
  assign n13767 = n13761 | n13766 ;
  assign n13768 = x299 & n8465 ;
  assign n13769 = x172 | n13473 ;
  assign n13770 = n13106 & ~n13769 ;
  assign n13771 = x152 & n13029 ;
  assign n13772 = n13682 | n13771 ;
  assign n13773 = x172 & n13772 ;
  assign n13774 = ( x197 & n13770 ) | ( x197 & ~n13773 ) | ( n13770 & ~n13773 ) ;
  assign n13775 = ~n13770 & n13774 ;
  assign n13776 = n13768 & ~n13775 ;
  assign n13777 = n13767 & n13776 ;
  assign n13778 = ( ~n13712 & n13755 ) | ( ~n13712 & n13777 ) | ( n13755 & n13777 ) ;
  assign n13779 = n13712 | n13778 ;
  assign n13780 = ( x39 & x232 ) | ( x39 & n13779 ) | ( x232 & n13779 ) ;
  assign n13781 = ~x39 & n13780 ;
  assign n13782 = n7678 & ~n13015 ;
  assign n13783 = n12960 | n13782 ;
  assign n13784 = n7669 & ~n13015 ;
  assign n13785 = n12960 | n13784 ;
  assign n13786 = n13783 ^ x299 ^ 1'b0 ;
  assign n13787 = ( n13783 & n13785 ) | ( n13783 & n13786 ) | ( n13785 & n13786 ) ;
  assign n13788 = ~x232 & n13787 ;
  assign n13789 = n5075 & n12959 ;
  assign n13790 = n7678 | n13789 ;
  assign n13791 = x51 | n13790 ;
  assign n13792 = n7678 & n13043 ;
  assign n13793 = n13791 & ~n13792 ;
  assign n13794 = x180 & ~n13084 ;
  assign n13795 = x174 & n13783 ;
  assign n13796 = n13795 ^ n13794 ^ 1'b0 ;
  assign n13797 = ( n13794 & n13795 ) | ( n13794 & n13796 ) | ( n13795 & n13796 ) ;
  assign n13798 = ( x193 & ~n13794 ) | ( x193 & n13797 ) | ( ~n13794 & n13797 ) ;
  assign n13799 = x180 & ~n13037 ;
  assign n13800 = x174 | n13799 ;
  assign n13801 = ~n13798 & n13800 ;
  assign n13802 = ( n13793 & n13798 ) | ( n13793 & ~n13801 ) | ( n13798 & ~n13801 ) ;
  assign n13803 = ~n12965 & n13783 ;
  assign n13804 = x174 & ~n13803 ;
  assign n13805 = x180 | n13804 ;
  assign n13806 = x51 & n5075 ;
  assign n13807 = n13790 | n13806 ;
  assign n13808 = n7678 & n13049 ;
  assign n13809 = n13807 & ~n13808 ;
  assign n13810 = ( x174 & ~n13805 ) | ( x174 & n13809 ) | ( ~n13805 & n13809 ) ;
  assign n13811 = ~n13805 & n13810 ;
  assign n13812 = ~x51 & n13084 ;
  assign n13813 = n5075 | n13812 ;
  assign n13814 = n13783 & n13813 ;
  assign n13815 = x174 & ~n13814 ;
  assign n13816 = n7678 & ~n13048 ;
  assign n13817 = ~n9182 & n13816 ;
  assign n13818 = n13807 & ~n13817 ;
  assign n13819 = x174 | n13818 ;
  assign n13820 = ( x180 & n13815 ) | ( x180 & n13819 ) | ( n13815 & n13819 ) ;
  assign n13821 = ~n13815 & n13820 ;
  assign n13822 = ( x193 & n13811 ) | ( x193 & ~n13821 ) | ( n13811 & ~n13821 ) ;
  assign n13823 = ~n13811 & n13822 ;
  assign n13824 = ( x299 & n13802 ) | ( x299 & ~n13823 ) | ( n13802 & ~n13823 ) ;
  assign n13825 = ~x299 & n13824 ;
  assign n13826 = n13044 & ~n13610 ;
  assign n13827 = x152 & ~n13472 ;
  assign n13828 = n7669 & ~n13827 ;
  assign n13829 = ( n7669 & ~n13084 ) | ( n7669 & n13828 ) | ( ~n13084 & n13828 ) ;
  assign n13830 = n13194 & ~n13829 ;
  assign n13831 = ( n13194 & n13826 ) | ( n13194 & n13830 ) | ( n13826 & n13830 ) ;
  assign n13832 = ( n13488 & n13490 ) | ( n13488 & n13491 ) | ( n13490 & n13491 ) ;
  assign n13833 = ( x172 & ~n13490 ) | ( x172 & n13832 ) | ( ~n13490 & n13832 ) ;
  assign n13834 = x152 & n13024 ;
  assign n13835 = ~x152 & n13049 ;
  assign n13836 = ( x172 & n13834 ) | ( x172 & ~n13835 ) | ( n13834 & ~n13835 ) ;
  assign n13837 = ~n13834 & n13836 ;
  assign n13838 = n7669 & ~n13837 ;
  assign n13839 = n13833 & n13838 ;
  assign n13840 = ~n13831 & n13839 ;
  assign n13841 = ( n8048 & n13831 ) | ( n8048 & ~n13840 ) | ( n13831 & ~n13840 ) ;
  assign n13842 = n12960 & ~n13474 ;
  assign n13843 = n13842 ^ n7669 ^ 1'b0 ;
  assign n13844 = ( n7669 & n13842 ) | ( n7669 & ~n13843 ) | ( n13842 & ~n13843 ) ;
  assign n13845 = ( n13841 & n13843 ) | ( n13841 & n13844 ) | ( n13843 & n13844 ) ;
  assign n13846 = ( x232 & n13825 ) | ( x232 & n13845 ) | ( n13825 & n13845 ) ;
  assign n13847 = n13845 ^ n13825 ^ 1'b0 ;
  assign n13848 = ( x232 & n13846 ) | ( x232 & n13847 ) | ( n13846 & n13847 ) ;
  assign n13849 = ( x39 & n13788 ) | ( x39 & ~n13848 ) | ( n13788 & ~n13848 ) ;
  assign n13850 = ~n13788 & n13849 ;
  assign n13851 = ~x232 & n13104 ;
  assign n13852 = x39 | n13851 ;
  assign n13853 = ( x38 & ~n13850 ) | ( x38 & n13852 ) | ( ~n13850 & n13852 ) ;
  assign n13854 = ~x38 & n13853 ;
  assign n13855 = ( ~n13681 & n13781 ) | ( ~n13681 & n13854 ) | ( n13781 & n13854 ) ;
  assign n13856 = n13681 | n13855 ;
  assign n13857 = ( n12962 & ~n13480 ) | ( n12962 & n13856 ) | ( ~n13480 & n13856 ) ;
  assign n13858 = ~n12962 & n13857 ;
  assign n13859 = n13459 | n13464 ;
  assign n13860 = ( ~n13680 & n13858 ) | ( ~n13680 & n13859 ) | ( n13858 & n13859 ) ;
  assign n13861 = n13680 | n13860 ;
  assign n13862 = ( n7318 & ~n13679 ) | ( n7318 & n13861 ) | ( ~n13679 & n13861 ) ;
  assign n13863 = ~n7318 & n13862 ;
  assign n13864 = n12960 | n13459 ;
  assign n13865 = x232 & n13474 ;
  assign n13866 = ( x87 & n13864 ) | ( x87 & ~n13865 ) | ( n13864 & ~n13865 ) ;
  assign n13867 = n13866 ^ n13864 ^ 1'b0 ;
  assign n13868 = ( x87 & n13866 ) | ( x87 & ~n13867 ) | ( n13866 & ~n13867 ) ;
  assign n13869 = n13863 ^ n13456 ^ 1'b0 ;
  assign n13870 = ( ~n13456 & n13868 ) | ( ~n13456 & n13869 ) | ( n13868 & n13869 ) ;
  assign n13871 = ( n13456 & n13863 ) | ( n13456 & n13870 ) | ( n13863 & n13870 ) ;
  assign n13872 = x121 | n13256 ;
  assign n13873 = n13872 ^ x126 ^ 1'b0 ;
  assign n13874 = n13254 & ~n13873 ;
  assign n13875 = x51 | n13029 ;
  assign n13876 = x232 & n13875 ;
  assign n13877 = n13874 & ~n13876 ;
  assign n13878 = x153 & n12965 ;
  assign n13879 = ( n10407 & n12960 ) | ( n10407 & n13172 ) | ( n12960 & n13172 ) ;
  assign n13880 = ~n13878 & n13879 ;
  assign n13881 = ~x232 & n12960 ;
  assign n13882 = n13880 | n13881 ;
  assign n13883 = ( ~x87 & n13877 ) | ( ~x87 & n13882 ) | ( n13877 & n13882 ) ;
  assign n13884 = ~x87 & n13883 ;
  assign n13885 = x87 & ~n12339 ;
  assign n13886 = ( n7318 & n13884 ) | ( n7318 & ~n13885 ) | ( n13884 & ~n13885 ) ;
  assign n13887 = ~n13884 & n13886 ;
  assign n13888 = ~x189 & n13029 ;
  assign n13889 = x175 & n12965 ;
  assign n13890 = ( x299 & ~n13888 ) | ( x299 & n13889 ) | ( ~n13888 & n13889 ) ;
  assign n13891 = n13888 | n13890 ;
  assign n13892 = n13875 & ~n13880 ;
  assign n13893 = x299 & ~n13892 ;
  assign n13894 = x232 & ~n13893 ;
  assign n13895 = n13891 & n13894 ;
  assign n13896 = n1205 & n13895 ;
  assign n13897 = n1205 & ~n12960 ;
  assign n13898 = ~n13874 & n13897 ;
  assign n13899 = ( n2097 & ~n13896 ) | ( n2097 & n13898 ) | ( ~n13896 & n13898 ) ;
  assign n13900 = n13896 | n13899 ;
  assign n13920 = ( x160 & n5390 ) | ( x160 & n6810 ) | ( n5390 & n6810 ) ;
  assign n13921 = n13892 & ~n13920 ;
  assign n13922 = n13487 ^ x166 ^ 1'b0 ;
  assign n13923 = ( n13487 & n13532 ) | ( n13487 & ~n13922 ) | ( n13532 & ~n13922 ) ;
  assign n13924 = x51 & ~x153 ;
  assign n13925 = ( ~x216 & n13923 ) | ( ~x216 & n13924 ) | ( n13923 & n13924 ) ;
  assign n13926 = ~x216 & n13925 ;
  assign n13932 = x166 & ~n13499 ;
  assign n13933 = x166 | n13496 ;
  assign n13934 = ( x153 & n13932 ) | ( x153 & n13933 ) | ( n13932 & n13933 ) ;
  assign n13935 = ~n13932 & n13934 ;
  assign n13927 = x166 & ~n13333 ;
  assign n13928 = x166 | n13032 ;
  assign n13929 = ~x153 & n13928 ;
  assign n13930 = x160 & ~n13929 ;
  assign n13931 = ( x160 & n13927 ) | ( x160 & n13930 ) | ( n13927 & n13930 ) ;
  assign n13936 = n13935 ^ n13931 ^ 1'b0 ;
  assign n13937 = ( x216 & ~n13931 ) | ( x216 & n13935 ) | ( ~n13931 & n13935 ) ;
  assign n13938 = ( x216 & ~n13936 ) | ( x216 & n13937 ) | ( ~n13936 & n13937 ) ;
  assign n13939 = ( n5390 & n13926 ) | ( n5390 & ~n13938 ) | ( n13926 & ~n13938 ) ;
  assign n13940 = ~n13926 & n13939 ;
  assign n13941 = ( x299 & n13921 ) | ( x299 & ~n13940 ) | ( n13921 & ~n13940 ) ;
  assign n13942 = ~n13921 & n13941 ;
  assign n13901 = x189 & n13543 ;
  assign n13902 = ~x189 & n13537 ;
  assign n13903 = ( x182 & n13901 ) | ( x182 & ~n13902 ) | ( n13901 & ~n13902 ) ;
  assign n13904 = ~n13901 & n13903 ;
  assign n13905 = ~x189 & n13553 ;
  assign n13906 = x189 & n13549 ;
  assign n13907 = ( x182 & ~n13905 ) | ( x182 & n13906 ) | ( ~n13905 & n13906 ) ;
  assign n13908 = n13905 | n13907 ;
  assign n13909 = ( n12965 & ~n13904 ) | ( n12965 & n13908 ) | ( ~n13904 & n13908 ) ;
  assign n13910 = ~n13904 & n13909 ;
  assign n13911 = ( x175 & x299 ) | ( x175 & ~n13910 ) | ( x299 & ~n13910 ) ;
  assign n13912 = ~x299 & n13911 ;
  assign n13913 = ~x189 & n13528 ;
  assign n13914 = x189 & n13519 ;
  assign n13915 = x182 & ~n13914 ;
  assign n13916 = n13908 & ~n13915 ;
  assign n13917 = ( n13908 & n13913 ) | ( n13908 & n13916 ) | ( n13913 & n13916 ) ;
  assign n13918 = ( n10436 & ~n13912 ) | ( n10436 & n13917 ) | ( ~n13912 & n13917 ) ;
  assign n13919 = ~n13912 & n13918 ;
  assign n13943 = n13942 ^ n13919 ^ 1'b0 ;
  assign n13944 = ( x232 & ~n13919 ) | ( x232 & n13942 ) | ( ~n13919 & n13942 ) ;
  assign n13945 = ( x232 & ~n13943 ) | ( x232 & n13944 ) | ( ~n13943 & n13944 ) ;
  assign n13946 = ( x39 & n13563 ) | ( x39 & n13945 ) | ( n13563 & n13945 ) ;
  assign n13947 = ~n13945 & n13946 ;
  assign n13948 = ( n13254 & n13873 ) | ( n13254 & ~n13947 ) | ( n13873 & ~n13947 ) ;
  assign n13949 = ~n13873 & n13948 ;
  assign n13950 = ~x189 & n13660 ;
  assign n13951 = x189 & n13111 ;
  assign n13952 = x178 | n13951 ;
  assign n13953 = n12965 | n13952 ;
  assign n13954 = ( ~x181 & n13950 ) | ( ~x181 & n13953 ) | ( n13950 & n13953 ) ;
  assign n13955 = ~x181 & n13954 ;
  assign n13956 = x189 & n13599 ;
  assign n13957 = ~x189 & n13602 ;
  assign n13958 = x178 & ~n13957 ;
  assign n13959 = n13955 & ~n13958 ;
  assign n13960 = ( n13955 & n13956 ) | ( n13955 & n13959 ) | ( n13956 & n13959 ) ;
  assign n13961 = x189 & ~n13571 ;
  assign n13962 = x189 | n13585 ;
  assign n13963 = n12965 | n13962 ;
  assign n13964 = n13963 ^ n13961 ^ 1'b0 ;
  assign n13965 = ( n13961 & n13963 ) | ( n13961 & n13964 ) | ( n13963 & n13964 ) ;
  assign n13966 = ( x178 & ~n13961 ) | ( x178 & n13965 ) | ( ~n13961 & n13965 ) ;
  assign n13967 = ~x189 & n13609 ;
  assign n13968 = x178 & ~n13967 ;
  assign n13969 = x189 | n13736 ;
  assign n13970 = n13152 & n13969 ;
  assign n13971 = n13968 & ~n13970 ;
  assign n13972 = x181 & ~n13971 ;
  assign n13973 = n13966 & n13972 ;
  assign n13974 = ( n10667 & n13960 ) | ( n10667 & ~n13973 ) | ( n13960 & ~n13973 ) ;
  assign n13975 = ~n13960 & n13974 ;
  assign n13980 = ~x166 & n13602 ;
  assign n13981 = x166 & n13599 ;
  assign n13982 = ( x153 & n13980 ) | ( x153 & ~n13981 ) | ( n13980 & ~n13981 ) ;
  assign n13983 = ~n13980 & n13982 ;
  assign n13976 = x166 & n13595 ;
  assign n13977 = ~x166 & n13593 ;
  assign n13978 = ( x153 & ~n13976 ) | ( x153 & n13977 ) | ( ~n13976 & n13977 ) ;
  assign n13979 = n13976 | n13978 ;
  assign n13984 = n13983 ^ n13979 ^ 1'b0 ;
  assign n13985 = ( x157 & ~n13979 ) | ( x157 & n13983 ) | ( ~n13979 & n13983 ) ;
  assign n13986 = ( x157 & ~n13984 ) | ( x157 & n13985 ) | ( ~n13984 & n13985 ) ;
  assign n13987 = x157 | n13878 ;
  assign n13988 = x166 & n13111 ;
  assign n13989 = n13987 | n13988 ;
  assign n13990 = ~x166 & n13660 ;
  assign n13991 = ( ~n13986 & n13989 ) | ( ~n13986 & n13990 ) | ( n13989 & n13990 ) ;
  assign n13992 = ~n13986 & n13991 ;
  assign n13993 = ~n13975 & n13992 ;
  assign n13994 = ( n13076 & n13975 ) | ( n13076 & ~n13993 ) | ( n13975 & ~n13993 ) ;
  assign n13999 = x153 & n13152 ;
  assign n14000 = ~x153 & n13613 ;
  assign n14001 = ( x157 & n13999 ) | ( x157 & ~n14000 ) | ( n13999 & ~n14000 ) ;
  assign n14002 = ~n13999 & n14001 ;
  assign n13995 = ~x153 & n13575 ;
  assign n13996 = x153 & n13571 ;
  assign n13997 = ( x157 & ~n13995 ) | ( x157 & n13996 ) | ( ~n13995 & n13996 ) ;
  assign n13998 = n13995 | n13997 ;
  assign n14003 = n14002 ^ n13998 ^ 1'b0 ;
  assign n14004 = ( x166 & ~n13998 ) | ( x166 & n14002 ) | ( ~n13998 & n14002 ) ;
  assign n14005 = ( x166 & ~n14003 ) | ( x166 & n14004 ) | ( ~n14003 & n14004 ) ;
  assign n14006 = x166 | n13878 ;
  assign n14007 = x157 & n13609 ;
  assign n14008 = n14006 | n14007 ;
  assign n14009 = ~x157 & n13585 ;
  assign n14010 = ( ~n14005 & n14008 ) | ( ~n14005 & n14009 ) | ( n14008 & n14009 ) ;
  assign n14011 = ~n14005 & n14010 ;
  assign n14012 = ~n13994 & n14011 ;
  assign n14013 = ( n13082 & n13994 ) | ( n13082 & ~n14012 ) | ( n13994 & ~n14012 ) ;
  assign n14014 = ~x178 & n13962 ;
  assign n14015 = x189 & ~n13575 ;
  assign n14016 = n14014 & ~n14015 ;
  assign n14017 = x189 & n13613 ;
  assign n14018 = n13967 | n14017 ;
  assign n14019 = x178 & n14018 ;
  assign n14020 = ( x181 & n14016 ) | ( x181 & n14019 ) | ( n14016 & n14019 ) ;
  assign n14021 = n14019 ^ n14016 ^ 1'b0 ;
  assign n14022 = ( x181 & n14020 ) | ( x181 & n14021 ) | ( n14020 & n14021 ) ;
  assign n14023 = ~x189 & n13593 ;
  assign n14024 = x189 & n13595 ;
  assign n14025 = ( x178 & n14023 ) | ( x178 & ~n14024 ) | ( n14023 & ~n14024 ) ;
  assign n14026 = ~n14023 & n14025 ;
  assign n14027 = n13660 | n13952 ;
  assign n14028 = ( n13955 & n14026 ) | ( n13955 & n14027 ) | ( n14026 & n14027 ) ;
  assign n14029 = ~n14026 & n14028 ;
  assign n14030 = ( n10436 & ~n14022 ) | ( n10436 & n14029 ) | ( ~n14022 & n14029 ) ;
  assign n14031 = n14022 | n14030 ;
  assign n14032 = x232 & ~n14031 ;
  assign n14033 = ( x232 & n14013 ) | ( x232 & n14032 ) | ( n14013 & n14032 ) ;
  assign n14034 = n14033 ^ n13949 ^ 1'b0 ;
  assign n14035 = ( ~n13567 & n14033 ) | ( ~n13567 & n14034 ) | ( n14033 & n14034 ) ;
  assign n14036 = ( n13949 & ~n14034 ) | ( n13949 & n14035 ) | ( ~n14034 & n14035 ) ;
  assign n14037 = n13044 ^ x166 ^ 1'b0 ;
  assign n14038 = ( n13044 & n13084 ) | ( n13044 & n14037 ) | ( n13084 & n14037 ) ;
  assign n14039 = x160 & ~n13878 ;
  assign n14040 = n14038 & n14039 ;
  assign n14041 = x166 | n13485 ;
  assign n14042 = n8898 & ~n13022 ;
  assign n14043 = ( x153 & n14041 ) | ( x153 & ~n14042 ) | ( n14041 & ~n14042 ) ;
  assign n14044 = n14043 ^ n14041 ^ 1'b0 ;
  assign n14045 = ( x153 & n14043 ) | ( x153 & ~n14044 ) | ( n14043 & ~n14044 ) ;
  assign n14046 = x166 & n13024 ;
  assign n14047 = ~x166 & n13049 ;
  assign n14048 = ( x153 & n14046 ) | ( x153 & ~n14047 ) | ( n14046 & ~n14047 ) ;
  assign n14049 = ~n14046 & n14048 ;
  assign n14050 = ( x160 & n14045 ) | ( x160 & ~n14049 ) | ( n14045 & ~n14049 ) ;
  assign n14051 = n14050 ^ n14045 ^ 1'b0 ;
  assign n14052 = ( x160 & n14050 ) | ( x160 & ~n14051 ) | ( n14050 & ~n14051 ) ;
  assign n14053 = ( n7669 & n14040 ) | ( n7669 & n14052 ) | ( n14040 & n14052 ) ;
  assign n14054 = ~n14040 & n14053 ;
  assign n14055 = n7669 | n13880 ;
  assign n14056 = ( x299 & n14054 ) | ( x299 & n14055 ) | ( n14054 & n14055 ) ;
  assign n14057 = ~n14054 & n14056 ;
  assign n14058 = x189 & n13783 ;
  assign n14059 = x182 & ~n13084 ;
  assign n14060 = n14058 & ~n14059 ;
  assign n14061 = x182 & ~n13037 ;
  assign n14062 = ( x189 & n13793 ) | ( x189 & ~n14061 ) | ( n13793 & ~n14061 ) ;
  assign n14063 = ~x189 & n14062 ;
  assign n14064 = ( ~n10436 & n14060 ) | ( ~n10436 & n14063 ) | ( n14060 & n14063 ) ;
  assign n14065 = ~n10436 & n14064 ;
  assign n14066 = x189 & ~n13803 ;
  assign n14067 = x182 | n14066 ;
  assign n14068 = ( x189 & n13809 ) | ( x189 & ~n14067 ) | ( n13809 & ~n14067 ) ;
  assign n14069 = ~n14067 & n14068 ;
  assign n14070 = x189 & ~n13814 ;
  assign n14071 = x182 & ~n14070 ;
  assign n14072 = n14071 ^ n14069 ^ 1'b0 ;
  assign n14073 = x189 | n13818 ;
  assign n14074 = ( n14071 & ~n14072 ) | ( n14071 & n14073 ) | ( ~n14072 & n14073 ) ;
  assign n14075 = ( n14069 & n14072 ) | ( n14069 & n14074 ) | ( n14072 & n14074 ) ;
  assign n14076 = n14065 ^ n10667 ^ 1'b0 ;
  assign n14077 = ( ~n10667 & n14075 ) | ( ~n10667 & n14076 ) | ( n14075 & n14076 ) ;
  assign n14078 = ( n10667 & n14065 ) | ( n10667 & n14077 ) | ( n14065 & n14077 ) ;
  assign n14079 = ( x232 & n14057 ) | ( x232 & n14078 ) | ( n14057 & n14078 ) ;
  assign n14080 = n14078 ^ n14057 ^ 1'b0 ;
  assign n14081 = ( x232 & n14079 ) | ( x232 & n14080 ) | ( n14079 & n14080 ) ;
  assign n14082 = ( x39 & n13788 ) | ( x39 & ~n14081 ) | ( n13788 & ~n14081 ) ;
  assign n14083 = ~n13788 & n14082 ;
  assign n14084 = n13873 & ~n14083 ;
  assign n14085 = ( n13254 & n14083 ) | ( n13254 & ~n14084 ) | ( n14083 & ~n14084 ) ;
  assign n14086 = ~x189 & n13293 ;
  assign n14087 = n8905 & n13104 ;
  assign n14088 = ( ~x178 & n14086 ) | ( ~x178 & n14087 ) | ( n14086 & n14087 ) ;
  assign n14089 = ~x178 & n14088 ;
  assign n14090 = x178 & n13969 ;
  assign n14091 = x189 | n13758 ;
  assign n14092 = x178 & n14091 ;
  assign n14093 = n14090 | n14092 ;
  assign n14094 = x189 & ~n13734 ;
  assign n14095 = n14093 & ~n14094 ;
  assign n14096 = ( x181 & ~n14089 ) | ( x181 & n14095 ) | ( ~n14089 & n14095 ) ;
  assign n14097 = n14089 | n14096 ;
  assign n14098 = x189 & ~n13756 ;
  assign n14099 = n14092 & ~n14098 ;
  assign n14100 = x189 & ~n13696 ;
  assign n14101 = x178 | n14100 ;
  assign n14102 = ( x189 & n13699 ) | ( x189 & ~n14101 ) | ( n13699 & ~n14101 ) ;
  assign n14103 = ~n14101 & n14102 ;
  assign n14104 = ( x181 & ~n14099 ) | ( x181 & n14103 ) | ( ~n14099 & n14103 ) ;
  assign n14105 = n14099 | n14104 ;
  assign n14106 = x189 & ~n13178 ;
  assign n14107 = x178 | n14106 ;
  assign n14108 = ( x189 & n13161 ) | ( x189 & ~n14107 ) | ( n13161 & ~n14107 ) ;
  assign n14109 = ~n14107 & n14108 ;
  assign n14110 = x178 & n10449 ;
  assign n14111 = x181 & ~n14110 ;
  assign n14112 = ( x181 & ~n13008 ) | ( x181 & n14111 ) | ( ~n13008 & n14111 ) ;
  assign n14113 = ( n13682 & ~n14109 ) | ( n13682 & n14112 ) | ( ~n14109 & n14112 ) ;
  assign n14114 = ~n13682 & n14113 ;
  assign n14115 = n10667 & ~n14114 ;
  assign n14116 = n14105 & n14115 ;
  assign n14117 = x51 & ~n8898 ;
  assign n14118 = x166 & n13688 ;
  assign n14119 = ( ~x153 & n14117 ) | ( ~x153 & n14118 ) | ( n14117 & n14118 ) ;
  assign n14120 = ~x153 & n14119 ;
  assign n14121 = x153 & x166 ;
  assign n14122 = n13685 & n14121 ;
  assign n14123 = ( x157 & ~n14120 ) | ( x157 & n14122 ) | ( ~n14120 & n14122 ) ;
  assign n14124 = n14120 | n14123 ;
  assign n14125 = ( ~x166 & n13683 ) | ( ~x166 & n14124 ) | ( n13683 & n14124 ) ;
  assign n14126 = n14124 ^ x166 ^ 1'b0 ;
  assign n14127 = ( n14124 & n14125 ) | ( n14124 & ~n14126 ) | ( n14125 & ~n14126 ) ;
  assign n14128 = n14127 ^ n14116 ^ 1'b0 ;
  assign n14129 = x153 | n13892 ;
  assign n14130 = n13106 & ~n14129 ;
  assign n14131 = x166 & n13029 ;
  assign n14132 = n13682 | n14131 ;
  assign n14133 = x153 & n14132 ;
  assign n14134 = ( x157 & n14130 ) | ( x157 & ~n14133 ) | ( n14130 & ~n14133 ) ;
  assign n14135 = ~n14130 & n14134 ;
  assign n14136 = ( x159 & x299 ) | ( x159 & n14135 ) | ( x299 & n14135 ) ;
  assign n14137 = ~n14135 & n14136 ;
  assign n14138 = ( n14127 & ~n14128 ) | ( n14127 & n14137 ) | ( ~n14128 & n14137 ) ;
  assign n14139 = ( n14116 & n14128 ) | ( n14116 & n14138 ) | ( n14128 & n14138 ) ;
  assign n14140 = x189 & ~n13688 ;
  assign n14141 = x178 | n14140 ;
  assign n14142 = ( n13161 & n13969 ) | ( n13161 & ~n14141 ) | ( n13969 & ~n14141 ) ;
  assign n14143 = ~n14141 & n14142 ;
  assign n14144 = ( n12963 & n13682 ) | ( n12963 & n14090 ) | ( n13682 & n14090 ) ;
  assign n14145 = ( x181 & n14143 ) | ( x181 & ~n14144 ) | ( n14143 & ~n14144 ) ;
  assign n14146 = ~n14143 & n14145 ;
  assign n14147 = ( x175 & x299 ) | ( x175 & ~n14146 ) | ( x299 & ~n14146 ) ;
  assign n14148 = n14146 | n14147 ;
  assign n14149 = ~n14139 & n14148 ;
  assign n14150 = ( n14097 & n14139 ) | ( n14097 & ~n14149 ) | ( n14139 & ~n14149 ) ;
  assign n14151 = x166 & n13734 ;
  assign n14152 = ( ~x153 & n14117 ) | ( ~x153 & n14151 ) | ( n14117 & n14151 ) ;
  assign n14153 = ~x153 & n14152 ;
  assign n14154 = n13756 & n14121 ;
  assign n14155 = x157 & ~n14154 ;
  assign n14156 = ~x166 & n13758 ;
  assign n14157 = ( n14153 & n14155 ) | ( n14153 & ~n14156 ) | ( n14155 & ~n14156 ) ;
  assign n14158 = ~n14153 & n14157 ;
  assign n14159 = x166 & n13696 ;
  assign n14160 = ~x166 & n13699 ;
  assign n14161 = ( x153 & n14159 ) | ( x153 & ~n14160 ) | ( n14159 & ~n14160 ) ;
  assign n14162 = ~n14159 & n14161 ;
  assign n14163 = ~x166 & n13293 ;
  assign n14164 = n8898 & n13104 ;
  assign n14165 = ( x153 & ~n14163 ) | ( x153 & n14164 ) | ( ~n14163 & n14164 ) ;
  assign n14166 = n14163 | n14165 ;
  assign n14167 = n14166 ^ n14162 ^ 1'b0 ;
  assign n14168 = ( n14162 & n14166 ) | ( n14162 & n14167 ) | ( n14166 & n14167 ) ;
  assign n14169 = ( x157 & ~n14162 ) | ( x157 & n14168 ) | ( ~n14162 & n14168 ) ;
  assign n14170 = ( n13076 & n14158 ) | ( n13076 & n14169 ) | ( n14158 & n14169 ) ;
  assign n14171 = ~n14158 & n14170 ;
  assign n14172 = ( x232 & n14150 ) | ( x232 & n14171 ) | ( n14150 & n14171 ) ;
  assign n14173 = n14171 ^ n14150 ^ 1'b0 ;
  assign n14174 = ( x232 & n14172 ) | ( x232 & n14173 ) | ( n14172 & n14173 ) ;
  assign n14175 = ( n13852 & ~n14085 ) | ( n13852 & n14174 ) | ( ~n14085 & n14174 ) ;
  assign n14176 = ~n14085 & n14175 ;
  assign n14177 = ( x38 & x100 ) | ( x38 & ~n14176 ) | ( x100 & ~n14176 ) ;
  assign n14178 = n14176 | n14177 ;
  assign n14179 = ( ~n13900 & n14036 ) | ( ~n13900 & n14178 ) | ( n14036 & n14178 ) ;
  assign n14180 = ~n13900 & n14179 ;
  assign n14181 = ~x150 & x299 ;
  assign n14182 = x185 | x299 ;
  assign n14183 = ~n14181 & n14182 ;
  assign n14184 = x87 & ~n14183 ;
  assign n14185 = ( x87 & ~n6411 ) | ( x87 & n14184 ) | ( ~n6411 & n14184 ) ;
  assign n14186 = n13895 & ~n14185 ;
  assign n14187 = ( n13265 & n14185 ) | ( n13265 & ~n14186 ) | ( n14185 & ~n14186 ) ;
  assign n14188 = n13874 ^ n13270 ^ 1'b0 ;
  assign n14189 = ( n13270 & n13874 ) | ( n13270 & ~n14188 ) | ( n13874 & ~n14188 ) ;
  assign n14190 = ( n14187 & n14188 ) | ( n14187 & n14189 ) | ( n14188 & n14189 ) ;
  assign n14191 = ( x57 & n5193 ) | ( x57 & ~n14190 ) | ( n5193 & ~n14190 ) ;
  assign n14192 = n14190 | n14191 ;
  assign n14193 = ( ~n13887 & n14180 ) | ( ~n13887 & n14192 ) | ( n14180 & n14192 ) ;
  assign n14194 = ~n13887 & n14193 ;
  assign n14195 = ~n2099 & n7528 ;
  assign n14196 = ~n2109 & n14195 ;
  assign n14197 = ( x57 & x59 ) | ( x57 & ~n14196 ) | ( x59 & ~n14196 ) ;
  assign n14198 = x129 & ~n6255 ;
  assign n14199 = ~n5459 & n14198 ;
  assign n14200 = x74 & ~n14199 ;
  assign n14201 = x54 & ~n2056 ;
  assign n14202 = n7528 & n14201 ;
  assign n14203 = x92 & ~x129 ;
  assign n14204 = x75 & n14198 ;
  assign n14205 = n2036 & n7459 ;
  assign n14206 = n2051 & ~n7528 ;
  assign n14207 = ( n2051 & n14205 ) | ( n2051 & n14206 ) | ( n14205 & n14206 ) ;
  assign n14208 = x75 | n14207 ;
  assign n14209 = x129 & ~n5052 ;
  assign n14210 = x38 & ~n14209 ;
  assign n14211 = ~x39 & x129 ;
  assign n14212 = n1400 | n1701 ;
  assign n14213 = n1473 | n1556 ;
  assign n14214 = n1226 | n1552 ;
  assign n14215 = ~n14213 & n14214 ;
  assign n14216 = ( ~n1469 & n1471 ) | ( ~n1469 & n14215 ) | ( n1471 & n14215 ) ;
  assign n14217 = ~n1469 & n14216 ;
  assign n14218 = ( n1386 & ~n1389 ) | ( n1386 & n14217 ) | ( ~n1389 & n14217 ) ;
  assign n14219 = ~n1389 & n14218 ;
  assign n14220 = x86 | n14219 ;
  assign n14221 = ~n1564 & n14220 ;
  assign n14222 = n1467 | n14221 ;
  assign n14223 = ~n1462 & n14222 ;
  assign n14224 = x108 | n14223 ;
  assign n14225 = ~n1704 & n14224 ;
  assign n14226 = ( ~n1703 & n1841 ) | ( ~n1703 & n14225 ) | ( n1841 & n14225 ) ;
  assign n14227 = ~n1703 & n14226 ;
  assign n14228 = n1452 | n14227 ;
  assign n14229 = ~n1451 & n14228 ;
  assign n14230 = ~n5023 & n14229 ;
  assign n14231 = n14221 ^ x97 ^ 1'b0 ;
  assign n14232 = ( ~n1459 & n14221 ) | ( ~n1459 & n14231 ) | ( n14221 & n14231 ) ;
  assign n14233 = x108 | n14232 ;
  assign n14234 = ~n1704 & n14233 ;
  assign n14235 = ( ~n1703 & n1841 ) | ( ~n1703 & n14234 ) | ( n1841 & n14234 ) ;
  assign n14236 = ~n1703 & n14235 ;
  assign n14237 = n1452 | n14236 ;
  assign n14238 = ~n1451 & n14237 ;
  assign n14239 = n5023 & n14238 ;
  assign n14240 = n7457 & n8969 ;
  assign n14241 = n14240 ^ n7458 ^ x252 ;
  assign n14242 = ( n14230 & ~n14239 ) | ( n14230 & n14241 ) | ( ~n14239 & n14241 ) ;
  assign n14243 = ~n14230 & n14242 ;
  assign n14244 = x127 & n14229 ;
  assign n14245 = ~x127 & n14238 ;
  assign n14246 = n14241 | n14245 ;
  assign n14247 = ( ~n14243 & n14244 ) | ( ~n14243 & n14246 ) | ( n14244 & n14246 ) ;
  assign n14248 = ~n14243 & n14247 ;
  assign n14249 = n1444 | n14248 ;
  assign n14250 = ~n1702 & n14249 ;
  assign n14251 = n1268 | n14250 ;
  assign n14252 = ~n14212 & n14251 ;
  assign n14253 = x70 | n14252 ;
  assign n14254 = ~n1693 & n14253 ;
  assign n14255 = x51 | n14254 ;
  assign n14256 = ~n1435 & n14255 ;
  assign n14257 = ( ~n1432 & n1773 ) | ( ~n1432 & n14256 ) | ( n1773 & n14256 ) ;
  assign n14258 = ~n1432 & n14257 ;
  assign n14259 = ( x32 & x40 ) | ( x32 & ~n14258 ) | ( x40 & ~n14258 ) ;
  assign n14260 = n14258 | n14259 ;
  assign n14261 = n14260 ^ n2219 ^ 1'b0 ;
  assign n14262 = ( n2219 & n14260 ) | ( n2219 & n14261 ) | ( n14260 & n14261 ) ;
  assign n14263 = ( x95 & ~n2219 ) | ( x95 & n14262 ) | ( ~n2219 & n14262 ) ;
  assign n14264 = ( n1422 & n14211 ) | ( n1422 & n14263 ) | ( n14211 & n14263 ) ;
  assign n14265 = ~n1422 & n14264 ;
  assign n14266 = ( x38 & n6259 ) | ( x38 & n7528 ) | ( n6259 & n7528 ) ;
  assign n14267 = ( ~n14210 & n14265 ) | ( ~n14210 & n14266 ) | ( n14265 & n14266 ) ;
  assign n14268 = ~n14210 & n14267 ;
  assign n14269 = ( n2051 & ~n14208 ) | ( n2051 & n14268 ) | ( ~n14208 & n14268 ) ;
  assign n14270 = ~n14208 & n14269 ;
  assign n14271 = ( x92 & ~n14204 ) | ( x92 & n14270 ) | ( ~n14204 & n14270 ) ;
  assign n14272 = n14204 | n14271 ;
  assign n14273 = ( n12146 & ~n14203 ) | ( n12146 & n14272 ) | ( ~n14203 & n14272 ) ;
  assign n14274 = ~n12146 & n14273 ;
  assign n14275 = ( x74 & ~n14202 ) | ( x74 & n14274 ) | ( ~n14202 & n14274 ) ;
  assign n14276 = n14202 | n14275 ;
  assign n14277 = ( x55 & ~n14200 ) | ( x55 & n14276 ) | ( ~n14200 & n14276 ) ;
  assign n14278 = ~x55 & n14277 ;
  assign n14279 = x55 & ~n2068 ;
  assign n14280 = n14198 & n14279 ;
  assign n14281 = ( ~x56 & n14278 ) | ( ~x56 & n14280 ) | ( n14278 & n14280 ) ;
  assign n14282 = ~x56 & n14281 ;
  assign n14283 = ( n9943 & n9952 ) | ( n9943 & ~n14282 ) | ( n9952 & ~n14282 ) ;
  assign n14284 = n14282 | n14283 ;
  assign n14285 = n14284 ^ n14195 ^ 1'b0 ;
  assign n14286 = ( ~n2109 & n14195 ) | ( ~n2109 & n14285 ) | ( n14195 & n14285 ) ;
  assign n14287 = ( n14284 & ~n14285 ) | ( n14284 & n14286 ) | ( ~n14285 & n14286 ) ;
  assign n14288 = ( n2120 & ~n14197 ) | ( n2120 & n14287 ) | ( ~n14197 & n14287 ) ;
  assign n14289 = ~n14197 & n14288 ;
  assign n14290 = n5011 | n6249 ;
  assign n14291 = n5023 & n14240 ;
  assign n14292 = n7461 & ~n14291 ;
  assign n14293 = x129 | n14240 ;
  assign n14294 = ( n1292 & n14292 ) | ( n1292 & n14293 ) | ( n14292 & n14293 ) ;
  assign n14295 = ~n1292 & n14294 ;
  assign n14296 = x38 | n2232 ;
  assign n14297 = ~n5054 & n14296 ;
  assign n14298 = n5019 & ~n5025 ;
  assign n14299 = x87 | n14298 ;
  assign n14300 = ( ~n5014 & n14297 ) | ( ~n5014 & n14299 ) | ( n14297 & n14299 ) ;
  assign n14301 = ~n5014 & n14300 ;
  assign n14302 = ( n5015 & ~n14295 ) | ( n5015 & n14301 ) | ( ~n14295 & n14301 ) ;
  assign n14303 = n14295 | n14302 ;
  assign n14304 = ( ~n6254 & n6257 ) | ( ~n6254 & n14303 ) | ( n6257 & n14303 ) ;
  assign n14305 = ~n6257 & n14304 ;
  assign n14306 = n7447 | n14305 ;
  assign n14307 = ~n14290 & n14306 ;
  assign n14308 = x56 | n14307 ;
  assign n14309 = ~n5008 & n14308 ;
  assign n14310 = x62 | n14309 ;
  assign n14311 = ~n5005 & n14310 ;
  assign n14312 = n2120 | n14311 ;
  assign n14313 = ~n5190 & n14312 ;
  assign n14314 = ~x87 & n13008 ;
  assign n14315 = x169 & n6411 ;
  assign n14316 = n14314 & ~n14315 ;
  assign n14317 = x87 & ~n8284 ;
  assign n14318 = ( n7318 & n14316 ) | ( n7318 & ~n14317 ) | ( n14316 & ~n14317 ) ;
  assign n14319 = ~n14316 & n14318 ;
  assign n14320 = x169 & n13029 ;
  assign n14321 = x51 | x87 ;
  assign n14322 = n14320 | n14321 ;
  assign n14323 = n14322 ^ n14319 ^ 1'b0 ;
  assign n14324 = x126 | n13872 ;
  assign n14325 = x132 | n14324 ;
  assign n14326 = n14325 ^ x130 ^ 1'b0 ;
  assign n14327 = n13252 & ~n14326 ;
  assign n14328 = ( n14322 & n14323 ) | ( n14322 & ~n14327 ) | ( n14323 & ~n14327 ) ;
  assign n14329 = ( n14319 & ~n14323 ) | ( n14319 & n14328 ) | ( ~n14323 & n14328 ) ;
  assign n14330 = x87 & ~n8328 ;
  assign n14331 = n6411 & n7629 ;
  assign n14332 = n13008 & ~n14331 ;
  assign n14333 = n13875 & ~n14332 ;
  assign n14334 = n13265 & ~n14333 ;
  assign n14335 = n14330 | n14334 ;
  assign n14336 = x38 & ~n14333 ;
  assign n14337 = n7629 | n13150 ;
  assign n14338 = ( n13149 & n13608 ) | ( n13149 & n13609 ) | ( n13608 & n13609 ) ;
  assign n14339 = n7629 & ~n14338 ;
  assign n14340 = x232 & ~n14339 ;
  assign n14341 = n14337 & n14340 ;
  assign n14342 = ~x232 & n13150 ;
  assign n14343 = ( x39 & ~n14341 ) | ( x39 & n14342 ) | ( ~n14341 & n14342 ) ;
  assign n14344 = n14341 | n14343 ;
  assign n14345 = n13496 & ~n13806 ;
  assign n14346 = n14345 ^ x224 ^ 1'b0 ;
  assign n14347 = ( n13042 & n14345 ) | ( n13042 & ~n14346 ) | ( n14345 & ~n14346 ) ;
  assign n14348 = n13875 ^ n5376 ^ 1'b0 ;
  assign n14349 = ( n13875 & ~n14347 ) | ( n13875 & n14348 ) | ( ~n14347 & n14348 ) ;
  assign n14350 = x140 & ~n14349 ;
  assign n14351 = n13875 ^ n6801 ^ 1'b0 ;
  assign n14352 = ( ~n13042 & n13875 ) | ( ~n13042 & n14351 ) | ( n13875 & n14351 ) ;
  assign n14353 = x140 | n14352 ;
  assign n14354 = ( n7627 & n14350 ) | ( n7627 & n14353 ) | ( n14350 & n14353 ) ;
  assign n14355 = ~n14350 & n14354 ;
  assign n14356 = x191 | x299 ;
  assign n14357 = n6801 & ~n13038 ;
  assign n14358 = x51 | n14357 ;
  assign n14359 = x140 | n14358 ;
  assign n14360 = ~n14356 & n14359 ;
  assign n14361 = x162 & n7669 ;
  assign n14362 = n6810 | n14361 ;
  assign n14363 = x51 | n14320 ;
  assign n14364 = ~n14362 & n14363 ;
  assign n14365 = x169 & n14345 ;
  assign n14366 = x162 & x216 ;
  assign n14367 = ~x51 & n13498 ;
  assign n14368 = ~x169 & n14367 ;
  assign n14369 = ( n14365 & n14366 ) | ( n14365 & ~n14368 ) | ( n14366 & ~n14368 ) ;
  assign n14370 = ~n14365 & n14369 ;
  assign n14371 = x169 & ~n5075 ;
  assign n14372 = n13039 | n14371 ;
  assign n14373 = x169 & ~n13041 ;
  assign n14374 = n14372 & ~n14373 ;
  assign n14375 = ( x216 & ~n14370 ) | ( x216 & n14374 ) | ( ~n14370 & n14374 ) ;
  assign n14376 = ~n14370 & n14375 ;
  assign n14377 = ( x215 & x221 ) | ( x215 & ~n14376 ) | ( x221 & ~n14376 ) ;
  assign n14378 = ~x215 & n14377 ;
  assign n14379 = ( x299 & n14364 ) | ( x299 & n14378 ) | ( n14364 & n14378 ) ;
  assign n14380 = n14378 ^ n14364 ^ 1'b0 ;
  assign n14381 = ( x299 & n14379 ) | ( x299 & n14380 ) | ( n14379 & n14380 ) ;
  assign n14382 = ~n13038 & n13540 ;
  assign n14383 = x51 | n14382 ;
  assign n14384 = x140 & ~n14383 ;
  assign n14385 = ~n14381 & n14384 ;
  assign n14386 = ( n14360 & n14381 ) | ( n14360 & ~n14385 ) | ( n14381 & ~n14385 ) ;
  assign n14387 = ( x232 & n14355 ) | ( x232 & n14386 ) | ( n14355 & n14386 ) ;
  assign n14388 = n14386 ^ n14355 ^ 1'b0 ;
  assign n14389 = ( x232 & n14387 ) | ( x232 & n14388 ) | ( n14387 & n14388 ) ;
  assign n14390 = ~n13038 & n13561 ;
  assign n14391 = x51 | n14390 ;
  assign n14392 = ~x232 & n14391 ;
  assign n14393 = ( x39 & n14389 ) | ( x39 & ~n14392 ) | ( n14389 & ~n14392 ) ;
  assign n14394 = ~n14389 & n14393 ;
  assign n14395 = ( x38 & n14344 ) | ( x38 & ~n14394 ) | ( n14344 & ~n14394 ) ;
  assign n14396 = n14395 ^ n14344 ^ 1'b0 ;
  assign n14397 = ( x38 & n14395 ) | ( x38 & ~n14396 ) | ( n14395 & ~n14396 ) ;
  assign n14398 = ( x100 & ~n14336 ) | ( x100 & n14397 ) | ( ~n14336 & n14397 ) ;
  assign n14399 = ~x100 & n14398 ;
  assign n14400 = x100 & n14333 ;
  assign n14401 = ( n2097 & ~n14399 ) | ( n2097 & n14400 ) | ( ~n14399 & n14400 ) ;
  assign n14402 = n14399 | n14401 ;
  assign n14403 = ( n14327 & n14335 ) | ( n14327 & n14402 ) | ( n14335 & n14402 ) ;
  assign n14404 = ~n14335 & n14403 ;
  assign n14405 = n2097 | n14400 ;
  assign n14406 = ~n9604 & n14332 ;
  assign n14407 = x51 | n13043 ;
  assign n14408 = n13030 & ~n14407 ;
  assign n14409 = x169 & ~n14408 ;
  assign n14410 = x169 | n13812 ;
  assign n14411 = ( n14361 & n14409 ) | ( n14361 & n14410 ) | ( n14409 & n14410 ) ;
  assign n14412 = ~n14409 & n14411 ;
  assign n14413 = ~n7669 & n13008 ;
  assign n14414 = ~n14371 & n14413 ;
  assign n14415 = x299 & ~n14414 ;
  assign n14416 = n1292 & n14371 ;
  assign n14417 = ~x162 & n7669 ;
  assign n14418 = n13023 & ~n14371 ;
  assign n14419 = ( n14416 & n14417 ) | ( n14416 & ~n14418 ) | ( n14417 & ~n14418 ) ;
  assign n14420 = ~n14416 & n14419 ;
  assign n14421 = ( n14412 & n14415 ) | ( n14412 & ~n14420 ) | ( n14415 & ~n14420 ) ;
  assign n14422 = ~n14412 & n14421 ;
  assign n14423 = x140 & ~n13030 ;
  assign n14424 = ~x51 & n13793 ;
  assign n14425 = n7627 & ~n14424 ;
  assign n14426 = ( n7627 & n14423 ) | ( n7627 & n14425 ) | ( n14423 & n14425 ) ;
  assign n14427 = ~x51 & n13783 ;
  assign n14428 = x140 & ~n13813 ;
  assign n14429 = n14427 & ~n14428 ;
  assign n14430 = ( n14356 & ~n14426 ) | ( n14356 & n14429 ) | ( ~n14426 & n14429 ) ;
  assign n14431 = ~n14426 & n14430 ;
  assign n14432 = x232 & ~n14431 ;
  assign n14433 = ( x232 & n14422 ) | ( x232 & n14432 ) | ( n14422 & n14432 ) ;
  assign n14434 = ~x51 & n13787 ;
  assign n14435 = x232 | n14434 ;
  assign n14436 = ( n9604 & n14433 ) | ( n9604 & n14435 ) | ( n14433 & n14435 ) ;
  assign n14437 = ~n14433 & n14436 ;
  assign n14438 = ( x100 & ~n14406 ) | ( x100 & n14437 ) | ( ~n14406 & n14437 ) ;
  assign n14439 = n14406 | n14438 ;
  assign n14440 = ( n12961 & ~n14405 ) | ( n12961 & n14439 ) | ( ~n14405 & n14439 ) ;
  assign n14441 = ~n12961 & n14440 ;
  assign n14442 = n13270 & n14335 ;
  assign n14443 = n14327 | n14442 ;
  assign n14444 = ( ~n14404 & n14441 ) | ( ~n14404 & n14443 ) | ( n14441 & n14443 ) ;
  assign n14445 = ~n14404 & n14444 ;
  assign n14446 = ( n7318 & ~n14329 ) | ( n7318 & n14445 ) | ( ~n14329 & n14445 ) ;
  assign n14447 = ~n14329 & n14446 ;
  assign n14448 = x87 | n6260 ;
  assign n14449 = x100 | n12520 ;
  assign n14450 = n14449 ^ n14448 ^ 1'b0 ;
  assign n14451 = ( n14448 & n14449 ) | ( n14448 & n14450 ) | ( n14449 & n14450 ) ;
  assign n14452 = ( x75 & ~n14448 ) | ( x75 & n14451 ) | ( ~n14448 & n14451 ) ;
  assign n14453 = n14452 ^ n6256 ^ 1'b0 ;
  assign n14454 = ( n6256 & n14452 ) | ( n6256 & n14453 ) | ( n14452 & n14453 ) ;
  assign n14455 = ( x92 & ~n6256 ) | ( x92 & n14454 ) | ( ~n6256 & n14454 ) ;
  assign n14456 = ( n7448 & ~n12146 ) | ( n7448 & n14455 ) | ( ~n12146 & n14455 ) ;
  assign n14457 = ~n7448 & n14456 ;
  assign n14458 = x164 & n13454 ;
  assign n14459 = n7318 & ~n14458 ;
  assign n14460 = x173 & n12965 ;
  assign n14461 = x299 | n14460 ;
  assign n14462 = x190 & n13029 ;
  assign n14463 = n14461 | n14462 ;
  assign n14464 = x51 & ~x151 ;
  assign n14465 = n12229 | n12965 ;
  assign n14466 = ~n14464 & n14465 ;
  assign n14467 = n12963 & n14466 ;
  assign n14468 = x299 & ~n14467 ;
  assign n14469 = x232 & ~n14468 ;
  assign n14470 = n14463 & n14469 ;
  assign n14471 = n13266 & ~n14470 ;
  assign n14472 = n1205 & n14470 ;
  assign n14473 = n2097 | n13897 ;
  assign n14474 = x232 | n13103 ;
  assign n14475 = n5075 & n13103 ;
  assign n14476 = ~x151 & n12965 ;
  assign n14477 = ( x168 & n13118 ) | ( x168 & ~n14476 ) | ( n13118 & ~n14476 ) ;
  assign n14478 = ~n13118 & n14477 ;
  assign n14479 = ~x151 & n13103 ;
  assign n14480 = x168 | n14479 ;
  assign n14481 = x151 & n13303 ;
  assign n14482 = ( ~n14478 & n14480 ) | ( ~n14478 & n14481 ) | ( n14480 & n14481 ) ;
  assign n14483 = ~n14478 & n14482 ;
  assign n14484 = ( x160 & ~n14475 ) | ( x160 & n14483 ) | ( ~n14475 & n14483 ) ;
  assign n14485 = n14475 | n14484 ;
  assign n14486 = x151 | n14467 ;
  assign n14487 = n13687 & ~n14486 ;
  assign n14488 = ~x168 & n13029 ;
  assign n14489 = n14475 | n14488 ;
  assign n14490 = x151 & n14489 ;
  assign n14491 = ( x160 & n14487 ) | ( x160 & ~n14490 ) | ( n14487 & ~n14490 ) ;
  assign n14492 = ~n14487 & n14491 ;
  assign n14493 = x299 & ~n14492 ;
  assign n14494 = n14485 & n14493 ;
  assign n14495 = x182 & ~n13687 ;
  assign n14496 = x190 | x299 ;
  assign n14497 = n14460 | n14496 ;
  assign n14498 = n13103 & ~n14497 ;
  assign n14499 = x232 & ~n14498 ;
  assign n14500 = ( x232 & n14495 ) | ( x232 & n14499 ) | ( n14495 & n14499 ) ;
  assign n14501 = x190 & ~x299 ;
  assign n14502 = x51 & ~x173 ;
  assign n14503 = n14475 | n14502 ;
  assign n14504 = ~x182 & n13118 ;
  assign n14505 = n14503 | n14504 ;
  assign n14506 = n14501 & n14505 ;
  assign n14507 = ( n14494 & n14500 ) | ( n14494 & ~n14506 ) | ( n14500 & ~n14506 ) ;
  assign n14508 = ~n14494 & n14507 ;
  assign n14509 = ( x39 & n14474 ) | ( x39 & ~n14508 ) | ( n14474 & ~n14508 ) ;
  assign n14510 = ~x39 & n14509 ;
  assign n14511 = x183 & ~n13818 ;
  assign n14512 = x183 | n13809 ;
  assign n14513 = ( x173 & n14511 ) | ( x173 & n14512 ) | ( n14511 & n14512 ) ;
  assign n14514 = ~n14511 & n14513 ;
  assign n14515 = x183 & ~n13037 ;
  assign n14516 = x173 | n14515 ;
  assign n14517 = ~n14514 & n14516 ;
  assign n14518 = ( n13793 & n14514 ) | ( n13793 & ~n14517 ) | ( n14514 & ~n14517 ) ;
  assign n14519 = n14501 & n14518 ;
  assign n14520 = n12229 | n13022 ;
  assign n14521 = x168 & ~n13485 ;
  assign n14522 = ( x151 & n14520 ) | ( x151 & ~n14521 ) | ( n14520 & ~n14521 ) ;
  assign n14523 = ~x151 & n14522 ;
  assign n14524 = x168 & ~n13049 ;
  assign n14525 = x168 | n13024 ;
  assign n14526 = ( x151 & n14524 ) | ( x151 & n14525 ) | ( n14524 & n14525 ) ;
  assign n14527 = ~n14524 & n14526 ;
  assign n14528 = ( x149 & ~n14523 ) | ( x149 & n14527 ) | ( ~n14523 & n14527 ) ;
  assign n14529 = n14523 | n14528 ;
  assign n14530 = ( n13044 & n13499 ) | ( n13044 & n14476 ) | ( n13499 & n14476 ) ;
  assign n14531 = x168 & ~n14530 ;
  assign n14532 = n13084 & ~n14466 ;
  assign n14533 = x168 | n14532 ;
  assign n14534 = ( x149 & n14531 ) | ( x149 & n14533 ) | ( n14531 & n14533 ) ;
  assign n14535 = ~n14531 & n14534 ;
  assign n14536 = n7669 & ~n14535 ;
  assign n14537 = n14529 & n14536 ;
  assign n14538 = n12960 & n14468 ;
  assign n14539 = ( n11620 & ~n14537 ) | ( n11620 & n14538 ) | ( ~n14537 & n14538 ) ;
  assign n14540 = ~n14537 & n14539 ;
  assign n14541 = n13783 & ~n14497 ;
  assign n14542 = x183 & ~n13084 ;
  assign n14543 = ( n14540 & n14541 ) | ( n14540 & ~n14542 ) | ( n14541 & ~n14542 ) ;
  assign n14544 = n14543 ^ n14541 ^ 1'b0 ;
  assign n14545 = ( n14540 & n14543 ) | ( n14540 & ~n14544 ) | ( n14543 & ~n14544 ) ;
  assign n14546 = ( x232 & n14519 ) | ( x232 & n14545 ) | ( n14519 & n14545 ) ;
  assign n14547 = n14545 ^ n14519 ^ 1'b0 ;
  assign n14548 = ( x232 & n14546 ) | ( x232 & n14547 ) | ( n14546 & n14547 ) ;
  assign n14549 = ( x39 & n13788 ) | ( x39 & n14548 ) | ( n13788 & n14548 ) ;
  assign n14550 = n14548 ^ n13788 ^ 1'b0 ;
  assign n14551 = ( x39 & n14549 ) | ( x39 & n14550 ) | ( n14549 & n14550 ) ;
  assign n14552 = ( n1205 & ~n14510 ) | ( n1205 & n14551 ) | ( ~n14510 & n14551 ) ;
  assign n14553 = n14510 | n14552 ;
  assign n14554 = ( n14472 & ~n14473 ) | ( n14472 & n14553 ) | ( ~n14473 & n14553 ) ;
  assign n14555 = ~n14472 & n14554 ;
  assign n14556 = n14324 ^ x132 ^ 1'b0 ;
  assign n14557 = n13253 & ~n14556 ;
  assign n14558 = x87 & ~n7636 ;
  assign n14559 = n14557 | n14558 ;
  assign n14560 = ( ~n14471 & n14555 ) | ( ~n14471 & n14559 ) | ( n14555 & n14559 ) ;
  assign n14561 = n14471 | n14560 ;
  assign n14562 = n14557 & ~n14558 ;
  assign n14587 = ( x149 & n5390 ) | ( x149 & n6810 ) | ( n5390 & n6810 ) ;
  assign n14588 = n14467 & ~n14587 ;
  assign n14589 = n13487 ^ x168 ^ 1'b0 ;
  assign n14590 = ( n13487 & n13532 ) | ( n13487 & n14589 ) | ( n13532 & n14589 ) ;
  assign n14591 = ( ~x216 & n14464 ) | ( ~x216 & n14590 ) | ( n14464 & n14590 ) ;
  assign n14592 = ~x216 & n14591 ;
  assign n14599 = ( x151 & n12219 ) | ( x151 & n13496 ) | ( n12219 & n13496 ) ;
  assign n14600 = x168 | n13499 ;
  assign n14601 = n14599 & n14600 ;
  assign n14594 = x168 & ~n13032 ;
  assign n14595 = x151 | n14594 ;
  assign n14593 = x168 | n13333 ;
  assign n14596 = n14595 ^ n14593 ^ 1'b0 ;
  assign n14597 = ( x149 & ~n14593 ) | ( x149 & n14595 ) | ( ~n14593 & n14595 ) ;
  assign n14598 = ( x149 & ~n14596 ) | ( x149 & n14597 ) | ( ~n14596 & n14597 ) ;
  assign n14602 = n14601 ^ n14598 ^ 1'b0 ;
  assign n14603 = ( x216 & ~n14598 ) | ( x216 & n14601 ) | ( ~n14598 & n14601 ) ;
  assign n14604 = ( x216 & ~n14602 ) | ( x216 & n14603 ) | ( ~n14602 & n14603 ) ;
  assign n14605 = ( n5390 & n14592 ) | ( n5390 & ~n14604 ) | ( n14592 & ~n14604 ) ;
  assign n14606 = ~n14592 & n14605 ;
  assign n14607 = ( x299 & n14588 ) | ( x299 & ~n14606 ) | ( n14588 & ~n14606 ) ;
  assign n14608 = ~n14588 & n14607 ;
  assign n14563 = x183 & n13528 ;
  assign n14564 = x183 | n13524 ;
  assign n14565 = ( x173 & ~n14563 ) | ( x173 & n14564 ) | ( ~n14563 & n14564 ) ;
  assign n14566 = ~x173 & n14565 ;
  assign n14567 = x183 | n13552 ;
  assign n14568 = x183 | n13533 ;
  assign n14569 = x173 & ~n13537 ;
  assign n14570 = n14568 & n14569 ;
  assign n14571 = ( n14566 & n14567 ) | ( n14566 & ~n14570 ) | ( n14567 & ~n14570 ) ;
  assign n14572 = ~n14566 & n14571 ;
  assign n14573 = ( x190 & x299 ) | ( x190 & ~n14572 ) | ( x299 & ~n14572 ) ;
  assign n14574 = ~x299 & n14573 ;
  assign n14575 = x183 | n12965 ;
  assign n14576 = n13549 | n14575 ;
  assign n14577 = x183 & ~n13543 ;
  assign n14578 = x173 & ~n14577 ;
  assign n14579 = n14576 & n14578 ;
  assign n14580 = x183 | n6801 ;
  assign n14581 = ( x173 & n13519 ) | ( x173 & n14580 ) | ( n13519 & n14580 ) ;
  assign n14582 = ~x173 & n14581 ;
  assign n14583 = ( x190 & x299 ) | ( x190 & ~n14582 ) | ( x299 & ~n14582 ) ;
  assign n14584 = n14582 | n14583 ;
  assign n14585 = ( ~n14574 & n14579 ) | ( ~n14574 & n14584 ) | ( n14579 & n14584 ) ;
  assign n14586 = ~n14574 & n14585 ;
  assign n14609 = n14608 ^ n14586 ^ 1'b0 ;
  assign n14610 = ( x232 & ~n14586 ) | ( x232 & n14608 ) | ( ~n14586 & n14608 ) ;
  assign n14611 = ( x232 & ~n14609 ) | ( x232 & n14610 ) | ( ~n14609 & n14610 ) ;
  assign n14612 = ( x39 & n13563 ) | ( x39 & n14611 ) | ( n13563 & n14611 ) ;
  assign n14613 = ~n14611 & n14612 ;
  assign n14614 = n5075 & ~n13167 ;
  assign n14615 = x160 & ~n14614 ;
  assign n14616 = x168 & ~n14464 ;
  assign n14617 = n13014 & n14616 ;
  assign n14618 = x151 & ~n13150 ;
  assign n14619 = x168 | n14618 ;
  assign n14620 = ( x151 & n13143 ) | ( x151 & ~n14619 ) | ( n13143 & ~n14619 ) ;
  assign n14621 = ~n14619 & n14620 ;
  assign n14622 = ( n5075 & ~n14617 ) | ( n5075 & n14621 ) | ( ~n14617 & n14621 ) ;
  assign n14623 = n14617 | n14622 ;
  assign n14624 = n14615 & n14623 ;
  assign n14625 = x168 & n13601 ;
  assign n14626 = ~n14614 & n14625 ;
  assign n14627 = n5075 & n13167 ;
  assign n14628 = n13162 | n14627 ;
  assign n14629 = ~x168 & n14628 ;
  assign n14630 = ( x151 & n14626 ) | ( x151 & ~n14629 ) | ( n14626 & ~n14629 ) ;
  assign n14631 = ~n14626 & n14630 ;
  assign n14632 = ~n12229 & n13167 ;
  assign n14633 = x168 & n13173 ;
  assign n14634 = ( x151 & ~n14632 ) | ( x151 & n14633 ) | ( ~n14632 & n14633 ) ;
  assign n14635 = n14632 | n14634 ;
  assign n14636 = ( x160 & ~n14631 ) | ( x160 & n14635 ) | ( ~n14631 & n14635 ) ;
  assign n14637 = ~x160 & n14636 ;
  assign n14638 = ( x299 & n14624 ) | ( x299 & ~n14637 ) | ( n14624 & ~n14637 ) ;
  assign n14639 = ~n14624 & n14638 ;
  assign n14641 = x182 & ~n14614 ;
  assign n14642 = ( n13144 & n14627 ) | ( n13144 & n14641 ) | ( n14627 & n14641 ) ;
  assign n14640 = ~x182 & n13167 ;
  assign n14643 = ( x173 & n14640 ) | ( x173 & ~n14642 ) | ( n14640 & ~n14642 ) ;
  assign n14644 = n14642 | n14643 ;
  assign n14645 = ~x182 & n14628 ;
  assign n14646 = x173 & ~n14645 ;
  assign n14647 = n14644 & ~n14646 ;
  assign n14648 = ( n13151 & n13152 ) | ( n13151 & n14641 ) | ( n13152 & n14641 ) ;
  assign n14649 = ( n14644 & n14647 ) | ( n14644 & n14648 ) | ( n14647 & n14648 ) ;
  assign n14650 = ( x190 & x299 ) | ( x190 & ~n14649 ) | ( x299 & ~n14649 ) ;
  assign n14651 = n14649 | n14650 ;
  assign n14652 = x182 & n12994 ;
  assign n14653 = n13013 | n14652 ;
  assign n14654 = ( n5075 & ~n14502 ) | ( n5075 & n14653 ) | ( ~n14502 & n14653 ) ;
  assign n14655 = ~n5075 & n14654 ;
  assign n14656 = ( x190 & x299 ) | ( x190 & ~n14655 ) | ( x299 & ~n14655 ) ;
  assign n14657 = ~x299 & n14656 ;
  assign n14658 = n14657 ^ n14627 ^ 1'b0 ;
  assign n14659 = ( x232 & n14627 ) | ( x232 & ~n14657 ) | ( n14627 & ~n14657 ) ;
  assign n14660 = ( x232 & ~n14658 ) | ( x232 & n14659 ) | ( ~n14658 & n14659 ) ;
  assign n14661 = ( n14639 & n14651 ) | ( n14639 & n14660 ) | ( n14651 & n14660 ) ;
  assign n14662 = ~n14639 & n14661 ;
  assign n14663 = ~x232 & n13167 ;
  assign n14664 = ( ~x39 & n14662 ) | ( ~x39 & n14663 ) | ( n14662 & n14663 ) ;
  assign n14665 = ~x39 & n14664 ;
  assign n14666 = ( ~n1205 & n14613 ) | ( ~n1205 & n14665 ) | ( n14613 & n14665 ) ;
  assign n14667 = ~n1205 & n14666 ;
  assign n14668 = ( n2097 & n14472 ) | ( n2097 & ~n14667 ) | ( n14472 & ~n14667 ) ;
  assign n14669 = n14667 | n14668 ;
  assign n14670 = n13265 & ~n14470 ;
  assign n14671 = n14669 & ~n14670 ;
  assign n14672 = n14562 & n14671 ;
  assign n14673 = ( n7318 & n14561 ) | ( n7318 & ~n14672 ) | ( n14561 & ~n14672 ) ;
  assign n14674 = ~n7318 & n14673 ;
  assign n14675 = n12960 | n14557 ;
  assign n14676 = x232 & n14467 ;
  assign n14677 = ( x87 & n14675 ) | ( x87 & ~n14676 ) | ( n14675 & ~n14676 ) ;
  assign n14678 = n14677 ^ n14675 ^ 1'b0 ;
  assign n14679 = ( x87 & n14677 ) | ( x87 & ~n14678 ) | ( n14677 & ~n14678 ) ;
  assign n14680 = n14674 ^ n14459 ^ 1'b0 ;
  assign n14681 = ( ~n14459 & n14679 ) | ( ~n14459 & n14680 ) | ( n14679 & n14680 ) ;
  assign n14682 = ( n14459 & n14674 ) | ( n14459 & n14681 ) | ( n14674 & n14681 ) ;
  assign n14683 = ~x133 & n13457 ;
  assign n14684 = ~n7644 & n13122 ;
  assign n14685 = ~x39 & x176 ;
  assign n14686 = n13613 ^ n13575 ^ n13122 ;
  assign n14687 = n7644 & n14686 ;
  assign n14688 = ( n14684 & n14685 ) | ( n14684 & ~n14687 ) | ( n14685 & ~n14687 ) ;
  assign n14689 = ~n14684 & n14688 ;
  assign n14690 = x154 & x232 ;
  assign n14691 = x299 & n14690 ;
  assign n14692 = n14686 & n14691 ;
  assign n14693 = x39 | x176 ;
  assign n14694 = n13122 & ~n14691 ;
  assign n14695 = ( ~n14692 & n14693 ) | ( ~n14692 & n14694 ) | ( n14693 & n14694 ) ;
  assign n14696 = n14692 | n14695 ;
  assign n14697 = x145 | n6801 ;
  assign n14698 = ( x299 & n13518 ) | ( x299 & n14697 ) | ( n13518 & n14697 ) ;
  assign n14699 = ~x299 & n14698 ;
  assign n14700 = x197 & ~n13030 ;
  assign n14701 = n4652 | n14700 ;
  assign n14702 = n14699 ^ n5525 ^ 1'b0 ;
  assign n14703 = ( ~n5525 & n14701 ) | ( ~n5525 & n14702 ) | ( n14701 & n14702 ) ;
  assign n14704 = ( n5525 & n14699 ) | ( n5525 & n14703 ) | ( n14699 & n14703 ) ;
  assign n14705 = n14704 ^ n1292 ^ 1'b0 ;
  assign n14706 = ( x232 & n1292 ) | ( x232 & ~n14704 ) | ( n1292 & ~n14704 ) ;
  assign n14707 = ( x232 & ~n14705 ) | ( x232 & n14706 ) | ( ~n14705 & n14706 ) ;
  assign n14708 = x39 & ~n13563 ;
  assign n14709 = ( x39 & n14707 ) | ( x39 & n14708 ) | ( n14707 & n14708 ) ;
  assign n14710 = ( n1205 & n2068 ) | ( n1205 & ~n14709 ) | ( n2068 & ~n14709 ) ;
  assign n14711 = n14709 | n14710 ;
  assign n14712 = ( n14689 & n14696 ) | ( n14689 & ~n14711 ) | ( n14696 & ~n14711 ) ;
  assign n14713 = ~n14689 & n14712 ;
  assign n14714 = ( x87 & n14683 ) | ( x87 & ~n14713 ) | ( n14683 & ~n14713 ) ;
  assign n14715 = ~x87 & n14714 ;
  assign n14716 = n13784 & ~n14700 ;
  assign n14717 = n12960 | n14716 ;
  assign n14718 = x299 & n14717 ;
  assign n14719 = ~x299 & n13783 ;
  assign n14720 = x145 & ~n13084 ;
  assign n14721 = n14719 & ~n14720 ;
  assign n14722 = ( x232 & n14718 ) | ( x232 & n14721 ) | ( n14718 & n14721 ) ;
  assign n14723 = n14721 ^ n14718 ^ 1'b0 ;
  assign n14724 = ( x232 & n14722 ) | ( x232 & n14723 ) | ( n14722 & n14723 ) ;
  assign n14725 = ( x39 & n13788 ) | ( x39 & ~n14724 ) | ( n13788 & ~n14724 ) ;
  assign n14726 = ~n13788 & n14725 ;
  assign n14727 = x39 | n12960 ;
  assign n14728 = ~n7647 & n13011 ;
  assign n14729 = n14727 | n14728 ;
  assign n14730 = ( x38 & ~n14726 ) | ( x38 & n14729 ) | ( ~n14726 & n14729 ) ;
  assign n14731 = ~x38 & n14730 ;
  assign n14732 = n12982 | n14731 ;
  assign n14733 = ~n12962 & n14732 ;
  assign n14734 = n13266 | n14733 ;
  assign n14735 = ~n14683 & n14734 ;
  assign n14736 = x299 ^ x149 ^ 1'b0 ;
  assign n14737 = ( x149 & x183 ) | ( x149 & ~n14736 ) | ( x183 & ~n14736 ) ;
  assign n14738 = n6411 & n14737 ;
  assign n14739 = ~n14735 & n14738 ;
  assign n14740 = ( x87 & n14735 ) | ( x87 & ~n14739 ) | ( n14735 & ~n14739 ) ;
  assign n14741 = ( ~n7318 & n14715 ) | ( ~n7318 & n14740 ) | ( n14715 & n14740 ) ;
  assign n14742 = ~n7318 & n14741 ;
  assign n14743 = x149 & n13454 ;
  assign n14744 = n7318 & ~n14743 ;
  assign n14745 = n14744 ^ n14742 ^ 1'b0 ;
  assign n14746 = n13270 | n14683 ;
  assign n14747 = ( n14744 & ~n14745 ) | ( n14744 & n14746 ) | ( ~n14745 & n14746 ) ;
  assign n14748 = ( n14742 & n14745 ) | ( n14742 & n14747 ) | ( n14745 & n14747 ) ;
  assign n14749 = n7318 & ~n14321 ;
  assign n14750 = x171 & ~n5075 ;
  assign n14751 = n12959 & n14750 ;
  assign n14752 = x232 & n14751 ;
  assign n14753 = n14749 & ~n14752 ;
  assign n14754 = x192 & ~x299 ;
  assign n14755 = n13030 & n14424 ;
  assign n14756 = n14754 & ~n14755 ;
  assign n14757 = x192 | x299 ;
  assign n14758 = n13813 & n14427 ;
  assign n14759 = ( ~n14756 & n14757 ) | ( ~n14756 & n14758 ) | ( n14757 & n14758 ) ;
  assign n14760 = ~n14756 & n14759 ;
  assign n14761 = n14413 & ~n14750 ;
  assign n14762 = x171 | n13812 ;
  assign n14763 = x171 & ~n14408 ;
  assign n14764 = n7669 & ~n14763 ;
  assign n14765 = n14762 & n14764 ;
  assign n14766 = ( x299 & n14761 ) | ( x299 & ~n14765 ) | ( n14761 & ~n14765 ) ;
  assign n14767 = ~n14761 & n14766 ;
  assign n14768 = n14760 & ~n14767 ;
  assign n14769 = n14434 ^ x232 ^ 1'b0 ;
  assign n14770 = ( n14434 & n14768 ) | ( n14434 & n14769 ) | ( n14768 & n14769 ) ;
  assign n14771 = ( x39 & x186 ) | ( x39 & n14770 ) | ( x186 & n14770 ) ;
  assign n14772 = ~n14770 & n14771 ;
  assign n14773 = n14427 | n14757 ;
  assign n14774 = ~n14424 & n14754 ;
  assign n14775 = n14773 & ~n14774 ;
  assign n14776 = ~n14767 & n14775 ;
  assign n14777 = ( n14434 & n14769 ) | ( n14434 & n14776 ) | ( n14769 & n14776 ) ;
  assign n14778 = ( x39 & x186 ) | ( x39 & ~n14777 ) | ( x186 & ~n14777 ) ;
  assign n14779 = ~x186 & n14778 ;
  assign n14780 = x171 & x299 ;
  assign n14781 = n14754 | n14780 ;
  assign n14782 = n6411 & n14781 ;
  assign n14783 = n13008 & ~n14782 ;
  assign n14784 = x39 | n14783 ;
  assign n14785 = x164 & n14784 ;
  assign n14786 = ( n14772 & ~n14779 ) | ( n14772 & n14785 ) | ( ~n14779 & n14785 ) ;
  assign n14787 = ~n14772 & n14786 ;
  assign n14788 = n13023 & ~n14750 ;
  assign n14789 = n3094 & ~n5075 ;
  assign n14790 = ( n7669 & n14788 ) | ( n7669 & ~n14789 ) | ( n14788 & ~n14789 ) ;
  assign n14791 = ~n14788 & n14790 ;
  assign n14792 = ( x299 & n14761 ) | ( x299 & ~n14791 ) | ( n14761 & ~n14791 ) ;
  assign n14793 = ~n14761 & n14792 ;
  assign n14794 = n14760 & ~n14793 ;
  assign n14795 = ( n14434 & n14769 ) | ( n14434 & n14794 ) | ( n14769 & n14794 ) ;
  assign n14796 = ( x39 & x186 ) | ( x39 & n14795 ) | ( x186 & n14795 ) ;
  assign n14797 = ~n14795 & n14796 ;
  assign n14798 = n14775 & ~n14793 ;
  assign n14799 = ( n14434 & n14769 ) | ( n14434 & n14798 ) | ( n14769 & n14798 ) ;
  assign n14800 = ( x39 & x186 ) | ( x39 & ~n14799 ) | ( x186 & ~n14799 ) ;
  assign n14801 = ~x186 & n14800 ;
  assign n14802 = ~x164 & n14784 ;
  assign n14803 = ( n14797 & ~n14801 ) | ( n14797 & n14802 ) | ( ~n14801 & n14802 ) ;
  assign n14804 = ~n14797 & n14803 ;
  assign n14805 = ( n1205 & ~n14787 ) | ( n1205 & n14804 ) | ( ~n14787 & n14804 ) ;
  assign n14806 = n14787 | n14805 ;
  assign n14807 = n13875 & ~n14783 ;
  assign n14808 = n1205 & n14807 ;
  assign n14809 = n2097 | n14808 ;
  assign n14810 = ( n13897 & n14806 ) | ( n13897 & ~n14809 ) | ( n14806 & ~n14809 ) ;
  assign n14811 = ~n13897 & n14810 ;
  assign n14812 = x130 | n14325 ;
  assign n14813 = x136 | n14812 ;
  assign n14814 = x135 | n14813 ;
  assign n14815 = x134 & n14814 ;
  assign n14816 = n13265 & n14783 ;
  assign n14817 = ( ~n14811 & n14815 ) | ( ~n14811 & n14816 ) | ( n14815 & n14816 ) ;
  assign n14818 = n14811 | n14817 ;
  assign n14819 = n13265 & ~n14807 ;
  assign n14820 = x232 & n14781 ;
  assign n14821 = n14338 & n14820 ;
  assign n14822 = n13150 & ~n14820 ;
  assign n14823 = ( x39 & ~n14821 ) | ( x39 & n14822 ) | ( ~n14821 & n14822 ) ;
  assign n14824 = n14821 | n14823 ;
  assign n14825 = ( x164 & n5390 ) | ( x164 & n6810 ) | ( n5390 & n6810 ) ;
  assign n14826 = ( x51 & n14751 ) | ( x51 & ~n14825 ) | ( n14751 & ~n14825 ) ;
  assign n14827 = ~n14825 & n14826 ;
  assign n14828 = x171 & n14345 ;
  assign n14829 = x164 & x216 ;
  assign n14830 = ~x171 & n14367 ;
  assign n14831 = ( n14828 & n14829 ) | ( n14828 & ~n14830 ) | ( n14829 & ~n14830 ) ;
  assign n14832 = ~n14828 & n14831 ;
  assign n14833 = n13039 | n14750 ;
  assign n14834 = x171 & ~n13041 ;
  assign n14835 = ( x216 & n14833 ) | ( x216 & ~n14834 ) | ( n14833 & ~n14834 ) ;
  assign n14836 = n14835 ^ n14833 ^ 1'b0 ;
  assign n14837 = ( x216 & n14835 ) | ( x216 & ~n14836 ) | ( n14835 & ~n14836 ) ;
  assign n14838 = n5390 & ~n14837 ;
  assign n14839 = ( n5390 & n14832 ) | ( n5390 & n14838 ) | ( n14832 & n14838 ) ;
  assign n14840 = ( x299 & n14827 ) | ( x299 & n14839 ) | ( n14827 & n14839 ) ;
  assign n14841 = n14839 ^ n14827 ^ 1'b0 ;
  assign n14842 = ( x299 & n14840 ) | ( x299 & n14841 ) | ( n14840 & n14841 ) ;
  assign n14843 = n14349 & n14754 ;
  assign n14844 = n14383 & ~n14757 ;
  assign n14845 = ( x186 & n14843 ) | ( x186 & ~n14844 ) | ( n14843 & ~n14844 ) ;
  assign n14846 = ~n14843 & n14845 ;
  assign n14847 = x39 & x186 ;
  assign n14848 = n14358 & ~n14757 ;
  assign n14849 = n14847 | n14848 ;
  assign n14850 = n14352 & n14754 ;
  assign n14851 = ( ~n14846 & n14849 ) | ( ~n14846 & n14850 ) | ( n14849 & n14850 ) ;
  assign n14852 = ~n14846 & n14851 ;
  assign n14853 = ( x232 & n14842 ) | ( x232 & n14852 ) | ( n14842 & n14852 ) ;
  assign n14854 = n14852 ^ n14842 ^ 1'b0 ;
  assign n14855 = ( x232 & n14853 ) | ( x232 & n14854 ) | ( n14853 & n14854 ) ;
  assign n14856 = ( x39 & n14392 ) | ( x39 & ~n14855 ) | ( n14392 & ~n14855 ) ;
  assign n14857 = ~n14392 & n14856 ;
  assign n14858 = ( n1205 & n14824 ) | ( n1205 & ~n14857 ) | ( n14824 & ~n14857 ) ;
  assign n14859 = ~n1205 & n14858 ;
  assign n14860 = ( n2097 & n14808 ) | ( n2097 & ~n14859 ) | ( n14808 & ~n14859 ) ;
  assign n14861 = n14859 | n14860 ;
  assign n14862 = ( n14815 & n14819 ) | ( n14815 & n14861 ) | ( n14819 & n14861 ) ;
  assign n14863 = ~n14819 & n14862 ;
  assign n14864 = ( n7318 & n14818 ) | ( n7318 & ~n14863 ) | ( n14818 & ~n14863 ) ;
  assign n14865 = ~n7318 & n14864 ;
  assign n14866 = n12959 | n14815 ;
  assign n14867 = n14865 ^ n14753 ^ 1'b0 ;
  assign n14868 = ( ~n14753 & n14866 ) | ( ~n14753 & n14867 ) | ( n14866 & n14867 ) ;
  assign n14869 = ( n14753 & n14865 ) | ( n14753 & n14868 ) | ( n14865 & n14868 ) ;
  assign n14870 = x170 & n6411 ;
  assign n14871 = n12959 & n14870 ;
  assign n14872 = n14749 & ~n14871 ;
  assign n14873 = x135 & n14813 ;
  assign n14874 = x134 & ~n14814 ;
  assign n14875 = n14873 | n14874 ;
  assign n14876 = x170 & ~n5075 ;
  assign n14877 = n9297 & n14876 ;
  assign n14878 = n13008 & ~n14877 ;
  assign n14879 = x194 & n7655 ;
  assign n14880 = n14878 & ~n14879 ;
  assign n14881 = n13875 & ~n14880 ;
  assign n14882 = n13265 & ~n14881 ;
  assign n14883 = n14875 & ~n14882 ;
  assign n14884 = n13875 & ~n14878 ;
  assign n14885 = x38 & ~n14884 ;
  assign n14886 = ~x299 & n13150 ;
  assign n14887 = x170 & ~n14338 ;
  assign n14888 = x170 | n13150 ;
  assign n14889 = ( n9297 & n14887 ) | ( n9297 & n14888 ) | ( n14887 & n14888 ) ;
  assign n14890 = ~n14887 & n14889 ;
  assign n14891 = ( x39 & n14342 ) | ( x39 & ~n14890 ) | ( n14342 & ~n14890 ) ;
  assign n14892 = n14890 | n14891 ;
  assign n14893 = n14886 | n14892 ;
  assign n14894 = ( x51 & x170 ) | ( x51 & n13875 ) | ( x170 & n13875 ) ;
  assign n14895 = n6810 | n14894 ;
  assign n14896 = x170 & ~n13041 ;
  assign n14897 = n6810 & ~n14896 ;
  assign n14898 = n13039 | n14876 ;
  assign n14899 = n14897 & n14898 ;
  assign n14900 = n14181 & ~n14899 ;
  assign n14901 = n14895 & n14900 ;
  assign n14902 = ~x170 & n14367 ;
  assign n14903 = x170 & n14345 ;
  assign n14904 = ( x216 & n14902 ) | ( x216 & ~n14903 ) | ( n14902 & ~n14903 ) ;
  assign n14905 = ~n14902 & n14904 ;
  assign n14906 = ( n7669 & n14899 ) | ( n7669 & ~n14905 ) | ( n14899 & ~n14905 ) ;
  assign n14907 = ~n14905 & n14906 ;
  assign n14908 = x150 & x299 ;
  assign n14909 = n5390 | n14894 ;
  assign n14910 = n14908 & n14909 ;
  assign n14911 = ( n14901 & ~n14907 ) | ( n14901 & n14910 ) | ( ~n14907 & n14910 ) ;
  assign n14912 = n14907 ^ n14901 ^ 1'b0 ;
  assign n14913 = ( n14901 & n14911 ) | ( n14901 & ~n14912 ) | ( n14911 & ~n14912 ) ;
  assign n14914 = x185 | n14358 ;
  assign n14915 = x185 & ~n14383 ;
  assign n14916 = ( x299 & n14914 ) | ( x299 & ~n14915 ) | ( n14914 & ~n14915 ) ;
  assign n14917 = ~x299 & n14916 ;
  assign n14918 = ( x232 & n14913 ) | ( x232 & n14917 ) | ( n14913 & n14917 ) ;
  assign n14919 = n14917 ^ n14913 ^ 1'b0 ;
  assign n14920 = ( x232 & n14918 ) | ( x232 & n14919 ) | ( n14918 & n14919 ) ;
  assign n14921 = ( x39 & n14392 ) | ( x39 & ~n14920 ) | ( n14392 & ~n14920 ) ;
  assign n14922 = ~n14392 & n14921 ;
  assign n14923 = ( x38 & n14893 ) | ( x38 & ~n14922 ) | ( n14893 & ~n14922 ) ;
  assign n14924 = n14923 ^ n14893 ^ 1'b0 ;
  assign n14925 = ( x38 & n14923 ) | ( x38 & ~n14924 ) | ( n14923 & ~n14924 ) ;
  assign n14926 = ( x194 & ~n14885 ) | ( x194 & n14925 ) | ( ~n14885 & n14925 ) ;
  assign n14927 = ~x194 & n14926 ;
  assign n14928 = n7655 | n14870 ;
  assign n14929 = n13008 & ~n14928 ;
  assign n14930 = n13875 & ~n14929 ;
  assign n14931 = x38 & ~n14930 ;
  assign n14932 = x194 & ~n14931 ;
  assign n14933 = n9323 & n14338 ;
  assign n14934 = n14892 | n14933 ;
  assign n14935 = x185 | n14352 ;
  assign n14936 = x185 & ~n14349 ;
  assign n14937 = ( x299 & n14935 ) | ( x299 & ~n14936 ) | ( n14935 & ~n14936 ) ;
  assign n14938 = ~x299 & n14937 ;
  assign n14939 = ( x232 & n14913 ) | ( x232 & n14938 ) | ( n14913 & n14938 ) ;
  assign n14940 = n14938 ^ n14913 ^ 1'b0 ;
  assign n14941 = ( x232 & n14939 ) | ( x232 & n14940 ) | ( n14939 & n14940 ) ;
  assign n14942 = ( x39 & n14392 ) | ( x39 & ~n14941 ) | ( n14392 & ~n14941 ) ;
  assign n14943 = ~n14392 & n14942 ;
  assign n14944 = ( x38 & n14934 ) | ( x38 & ~n14943 ) | ( n14934 & ~n14943 ) ;
  assign n14945 = n14944 ^ n14934 ^ 1'b0 ;
  assign n14946 = ( x38 & n14944 ) | ( x38 & ~n14945 ) | ( n14944 & ~n14945 ) ;
  assign n14947 = n14932 & n14946 ;
  assign n14948 = ( ~x100 & n14927 ) | ( ~x100 & n14947 ) | ( n14927 & n14947 ) ;
  assign n14949 = ~x100 & n14948 ;
  assign n14950 = x100 & n14881 ;
  assign n14951 = ( n2097 & ~n14949 ) | ( n2097 & n14950 ) | ( ~n14949 & n14950 ) ;
  assign n14952 = n14949 | n14951 ;
  assign n14953 = n14883 & n14952 ;
  assign n14954 = n13265 & n14880 ;
  assign n14955 = n2097 | n14950 ;
  assign n14957 = ~n9604 & n14929 ;
  assign n14958 = x194 & ~n14957 ;
  assign n14961 = ~n9604 & n14878 ;
  assign n14962 = x194 | n14961 ;
  assign n14969 = ~n14958 & n14962 ;
  assign n14970 = n3326 & ~n5075 ;
  assign n14971 = n13023 & ~n14876 ;
  assign n14972 = n7669 & ~n14971 ;
  assign n14973 = n14181 & ~n14972 ;
  assign n14974 = ( n14181 & n14970 ) | ( n14181 & n14973 ) | ( n14970 & n14973 ) ;
  assign n14975 = x170 | n13812 ;
  assign n14976 = x170 & ~n14408 ;
  assign n14977 = n7669 & ~n14976 ;
  assign n14978 = n14975 & n14977 ;
  assign n14979 = ~n14974 & n14978 ;
  assign n14980 = ( n14908 & n14974 ) | ( n14908 & ~n14979 ) | ( n14974 & ~n14979 ) ;
  assign n14981 = n14413 & ~n14876 ;
  assign n14982 = ( n14969 & n14980 ) | ( n14969 & ~n14981 ) | ( n14980 & ~n14981 ) ;
  assign n14983 = ~n14969 & n14982 ;
  assign n14956 = ~x185 & n14424 ;
  assign n14959 = ~n14755 & n14958 ;
  assign n14960 = ~n14956 & n14959 ;
  assign n14963 = x185 & ~n13813 ;
  assign n14964 = n14427 & ~n14963 ;
  assign n14965 = n14962 | n14964 ;
  assign n14966 = n14965 ^ n14960 ^ 1'b0 ;
  assign n14967 = ( n14960 & n14965 ) | ( n14960 & n14966 ) | ( n14965 & n14966 ) ;
  assign n14968 = ( x299 & ~n14960 ) | ( x299 & n14967 ) | ( ~n14960 & n14967 ) ;
  assign n14984 = n14983 ^ n14968 ^ 1'b0 ;
  assign n14985 = ( x232 & ~n14968 ) | ( x232 & n14983 ) | ( ~n14968 & n14983 ) ;
  assign n14986 = ( x232 & ~n14984 ) | ( x232 & n14985 ) | ( ~n14984 & n14985 ) ;
  assign n14987 = n9604 & n14435 ;
  assign n14988 = n14969 | n14987 ;
  assign n14989 = n14988 ^ n14986 ^ 1'b0 ;
  assign n14990 = ( n14986 & n14988 ) | ( n14986 & n14989 ) | ( n14988 & n14989 ) ;
  assign n14991 = ( x100 & ~n14986 ) | ( x100 & n14990 ) | ( ~n14986 & n14990 ) ;
  assign n14992 = ( n12961 & ~n14955 ) | ( n12961 & n14991 ) | ( ~n14955 & n14991 ) ;
  assign n14993 = ~n12961 & n14992 ;
  assign n14994 = ( n14875 & ~n14954 ) | ( n14875 & n14993 ) | ( ~n14954 & n14993 ) ;
  assign n14995 = n14954 | n14994 ;
  assign n14996 = ( n7318 & ~n14953 ) | ( n7318 & n14995 ) | ( ~n14953 & n14995 ) ;
  assign n14997 = ~n7318 & n14996 ;
  assign n14998 = n12959 | n14875 ;
  assign n14999 = n14997 ^ n14872 ^ 1'b0 ;
  assign n15000 = ( ~n14872 & n14998 ) | ( ~n14872 & n14999 ) | ( n14998 & n14999 ) ;
  assign n15001 = ( n14872 & n14997 ) | ( n14872 & n15000 ) | ( n14997 & n15000 ) ;
  assign n15002 = n14812 ^ x136 ^ 1'b0 ;
  assign n15003 = n13251 & ~n15002 ;
  assign n15004 = ( x51 & n8320 ) | ( x51 & n13875 ) | ( n8320 & n13875 ) ;
  assign n15005 = n13265 & ~n15004 ;
  assign n15006 = n15003 & ~n15005 ;
  assign n15007 = n1205 & n15004 ;
  assign n15008 = x184 & ~n14349 ;
  assign n15009 = x184 | n14352 ;
  assign n15010 = ( n8317 & n15008 ) | ( n8317 & n15009 ) | ( n15008 & n15009 ) ;
  assign n15011 = ~n15008 & n15010 ;
  assign n15012 = x141 | x299 ;
  assign n15013 = x184 | n14358 ;
  assign n15014 = ~n15012 & n15013 ;
  assign n15015 = ~x287 & n10323 ;
  assign n15016 = x216 & ~n15015 ;
  assign n15017 = ( n5390 & n13038 ) | ( n5390 & ~n15016 ) | ( n13038 & ~n15016 ) ;
  assign n15018 = ~n13038 & n15017 ;
  assign n15019 = ( x51 & x148 ) | ( x51 & ~n15018 ) | ( x148 & ~n15018 ) ;
  assign n15020 = n15018 | n15019 ;
  assign n15021 = n6810 & ~n13042 ;
  assign n15022 = x163 & n5390 ;
  assign n15023 = n14345 & n15022 ;
  assign n15024 = ~n6810 & n13875 ;
  assign n15025 = x163 | n15024 ;
  assign n15026 = n5390 | n13875 ;
  assign n15027 = ( n15023 & n15025 ) | ( n15023 & n15026 ) | ( n15025 & n15026 ) ;
  assign n15028 = ~n15023 & n15027 ;
  assign n15029 = ( x148 & n15021 ) | ( x148 & ~n15028 ) | ( n15021 & ~n15028 ) ;
  assign n15030 = ~n15021 & n15029 ;
  assign n15031 = x299 & ~n15030 ;
  assign n15032 = n15020 & n15031 ;
  assign n15033 = x184 & ~n14383 ;
  assign n15034 = ~n15032 & n15033 ;
  assign n15035 = ( n15014 & n15032 ) | ( n15014 & ~n15034 ) | ( n15032 & ~n15034 ) ;
  assign n15036 = ( x232 & n15011 ) | ( x232 & n15035 ) | ( n15011 & n15035 ) ;
  assign n15037 = n15035 ^ n15011 ^ 1'b0 ;
  assign n15038 = ( x232 & n15036 ) | ( x232 & n15037 ) | ( n15036 & n15037 ) ;
  assign n15039 = ( x39 & n14392 ) | ( x39 & ~n15038 ) | ( n14392 & ~n15038 ) ;
  assign n15040 = ~n14392 & n15039 ;
  assign n15041 = ( x38 & x100 ) | ( x38 & ~n15040 ) | ( x100 & ~n15040 ) ;
  assign n15042 = n15040 | n15041 ;
  assign n15043 = x39 | n14342 ;
  assign n15044 = n8319 | n13150 ;
  assign n15045 = n8319 & ~n14338 ;
  assign n15046 = x232 & ~n15045 ;
  assign n15047 = n15044 & n15046 ;
  assign n15048 = ( ~n15042 & n15043 ) | ( ~n15042 & n15047 ) | ( n15043 & n15047 ) ;
  assign n15049 = ~n15042 & n15048 ;
  assign n15050 = ( n2097 & ~n15007 ) | ( n2097 & n15049 ) | ( ~n15007 & n15049 ) ;
  assign n15051 = n15007 | n15050 ;
  assign n15052 = n15006 & n15051 ;
  assign n15066 = n5075 & n14413 ;
  assign n15067 = n7669 & ~n14407 ;
  assign n15068 = ( x148 & n15066 ) | ( x148 & ~n15067 ) | ( n15066 & ~n15067 ) ;
  assign n15069 = ~n15066 & n15068 ;
  assign n15060 = ~x51 & n13784 ;
  assign n15061 = x148 | n15060 ;
  assign n15062 = ~n15015 & n15061 ;
  assign n15063 = ( ~x148 & n13008 ) | ( ~x148 & n15062 ) | ( n13008 & n15062 ) ;
  assign n15064 = n15062 ^ x148 ^ 1'b0 ;
  assign n15065 = ( n15062 & n15063 ) | ( n15062 & ~n15064 ) | ( n15063 & ~n15064 ) ;
  assign n15070 = n15069 ^ n15065 ^ 1'b0 ;
  assign n15071 = ( x299 & ~n15065 ) | ( x299 & n15069 ) | ( ~n15065 & n15069 ) ;
  assign n15072 = ( x299 & ~n15070 ) | ( x299 & n15071 ) | ( ~n15070 & n15071 ) ;
  assign n15053 = x184 & ~n13030 ;
  assign n15054 = n8317 & ~n14424 ;
  assign n15055 = ( n8317 & n15053 ) | ( n8317 & n15054 ) | ( n15053 & n15054 ) ;
  assign n15056 = x184 & ~n13813 ;
  assign n15057 = n14427 & ~n15056 ;
  assign n15058 = ( n15012 & ~n15055 ) | ( n15012 & n15057 ) | ( ~n15055 & n15057 ) ;
  assign n15059 = ~n15055 & n15058 ;
  assign n15073 = n15072 ^ n15059 ^ 1'b0 ;
  assign n15074 = ( x232 & ~n15059 ) | ( x232 & n15072 ) | ( ~n15059 & n15072 ) ;
  assign n15075 = ( x232 & ~n15073 ) | ( x232 & n15074 ) | ( ~n15073 & n15074 ) ;
  assign n15076 = ( x100 & n14987 ) | ( x100 & ~n15075 ) | ( n14987 & ~n15075 ) ;
  assign n15077 = ~x100 & n15076 ;
  assign n15078 = ~n9815 & n12959 ;
  assign n15079 = ~n15004 & n15078 ;
  assign n15080 = ( ~n2097 & n15077 ) | ( ~n2097 & n15079 ) | ( n15077 & n15079 ) ;
  assign n15081 = ~n2097 & n15080 ;
  assign n15082 = n12959 & n15005 ;
  assign n15083 = ( n15003 & ~n15081 ) | ( n15003 & n15082 ) | ( ~n15081 & n15082 ) ;
  assign n15084 = n15081 | n15083 ;
  assign n15085 = ( n7318 & ~n15052 ) | ( n7318 & n15084 ) | ( ~n15052 & n15084 ) ;
  assign n15086 = ~n7318 & n15085 ;
  assign n15087 = ~n13008 & n15003 ;
  assign n15088 = x148 & n6411 ;
  assign n15089 = ~n15087 & n15088 ;
  assign n15090 = ( n12959 & n15087 ) | ( n12959 & ~n15089 ) | ( n15087 & ~n15089 ) ;
  assign n15091 = n15086 ^ n14749 ^ 1'b0 ;
  assign n15092 = ( ~n14749 & n15090 ) | ( ~n14749 & n15091 ) | ( n15090 & n15091 ) ;
  assign n15093 = ( n14749 & n15086 ) | ( n14749 & n15092 ) | ( n15086 & n15092 ) ;
  assign n15094 = x210 | n10150 ;
  assign n15095 = n7318 & ~n15094 ;
  assign n15096 = ~x210 & x299 ;
  assign n15097 = ~n10150 & n15096 ;
  assign n15098 = x299 | n7318 ;
  assign n15099 = x198 | n10218 ;
  assign n15100 = ( ~n15097 & n15098 ) | ( ~n15097 & n15099 ) | ( n15098 & n15099 ) ;
  assign n15101 = ~n15097 & n15100 ;
  assign n15102 = x38 | n2069 ;
  assign n15103 = ~n15101 & n15102 ;
  assign n15104 = ( n8962 & n15101 ) | ( n8962 & ~n15103 ) | ( n15101 & ~n15103 ) ;
  assign n15105 = n8901 & ~n15104 ;
  assign n15106 = ( n8901 & n15095 ) | ( n8901 & n15105 ) | ( n15095 & n15105 ) ;
  assign n15107 = ( ~x39 & x137 ) | ( ~x39 & n15106 ) | ( x137 & n15106 ) ;
  assign n15108 = n15106 ^ x39 ^ 1'b0 ;
  assign n15109 = ( n15106 & n15107 ) | ( n15106 & ~n15108 ) | ( n15107 & ~n15108 ) ;
  assign n15110 = ~n7571 & n7648 ;
  assign n15111 = x92 & ~n15110 ;
  assign n15112 = n2067 | n15111 ;
  assign n15113 = x75 | n7653 ;
  assign n15114 = n7699 & n10813 ;
  assign n15115 = n7725 & ~n15114 ;
  assign n15116 = n12384 & ~n15115 ;
  assign n15118 = n5061 & n7699 ;
  assign n15117 = n7669 & ~n15114 ;
  assign n15119 = n15118 ^ n15117 ^ 1'b0 ;
  assign n15120 = ( n7671 & ~n15117 ) | ( n7671 & n15118 ) | ( ~n15117 & n15118 ) ;
  assign n15121 = ( n7671 & ~n15119 ) | ( n7671 & n15120 ) | ( ~n15119 & n15120 ) ;
  assign n15122 = n15116 | n15121 ;
  assign n15123 = ~x232 & n15122 ;
  assign n15124 = n7704 | n15114 ;
  assign n15125 = n7670 & n15124 ;
  assign n15126 = x148 & ~n15125 ;
  assign n15127 = ( n8318 & n15121 ) | ( n8318 & ~n15126 ) | ( n15121 & ~n15126 ) ;
  assign n15128 = ~n15126 & n15127 ;
  assign n15129 = ( n7715 & n12384 ) | ( n7715 & n15116 ) | ( n12384 & n15116 ) ;
  assign n15130 = ( x141 & n15116 ) | ( x141 & n15129 ) | ( n15116 & n15129 ) ;
  assign n15131 = ( x232 & n15128 ) | ( x232 & n15130 ) | ( n15128 & n15130 ) ;
  assign n15132 = n15130 ^ n15128 ^ 1'b0 ;
  assign n15133 = ( x232 & n15131 ) | ( x232 & n15132 ) | ( n15131 & n15132 ) ;
  assign n15134 = ( x39 & n15123 ) | ( x39 & n15133 ) | ( n15123 & n15133 ) ;
  assign n15135 = n15133 ^ n15123 ^ 1'b0 ;
  assign n15136 = ( x39 & n15134 ) | ( x39 & n15135 ) | ( n15134 & n15135 ) ;
  assign n15137 = ( x38 & x100 ) | ( x38 & ~n15136 ) | ( x100 & ~n15136 ) ;
  assign n15138 = n15136 | n15137 ;
  assign n15139 = ~x299 & n8367 ;
  assign n15140 = x299 & n8050 ;
  assign n15141 = x232 | n15140 ;
  assign n15142 = n15139 | n15141 ;
  assign n15143 = x148 & ~n5075 ;
  assign n15144 = n8050 & ~n15143 ;
  assign n15145 = x148 & n7980 ;
  assign n15146 = ( x299 & n15144 ) | ( x299 & n15145 ) | ( n15144 & n15145 ) ;
  assign n15147 = n15145 ^ n15144 ^ 1'b0 ;
  assign n15148 = ( x299 & n15146 ) | ( x299 & n15147 ) | ( n15146 & n15147 ) ;
  assign n15149 = ~x141 & n15139 ;
  assign n15150 = x232 & ~n15149 ;
  assign n15151 = ( n7795 & n7952 ) | ( n7795 & n8367 ) | ( n7952 & n8367 ) ;
  assign n15152 = ~x299 & n15151 ;
  assign n15153 = x141 & n15152 ;
  assign n15154 = ( n15148 & n15150 ) | ( n15148 & ~n15153 ) | ( n15150 & ~n15153 ) ;
  assign n15155 = ~n15148 & n15154 ;
  assign n15156 = ( x39 & n15142 ) | ( x39 & ~n15155 ) | ( n15142 & ~n15155 ) ;
  assign n15157 = ~x39 & n15156 ;
  assign n15158 = ( ~x87 & n15138 ) | ( ~x87 & n15157 ) | ( n15138 & n15157 ) ;
  assign n15159 = ~x87 & n15158 ;
  assign n15160 = ( ~x92 & n15113 ) | ( ~x92 & n15159 ) | ( n15113 & n15159 ) ;
  assign n15161 = ~x92 & n15160 ;
  assign n15162 = ( ~x55 & n15112 ) | ( ~x55 & n15161 ) | ( n15112 & n15161 ) ;
  assign n15163 = ~x55 & n15162 ;
  assign n15164 = ~n7572 & n12359 ;
  assign n15165 = ~n15163 & n15164 ;
  assign n15166 = ( x55 & n15163 ) | ( x55 & ~n15165 ) | ( n15163 & ~n15165 ) ;
  assign n15167 = n2109 | n15166 ;
  assign n15168 = ( ~n2109 & n8298 ) | ( ~n2109 & n15167 ) | ( n8298 & n15167 ) ;
  assign n15169 = x138 & ~n15168 ;
  assign n15170 = ~n8320 & n12242 ;
  assign n15171 = x39 | n15170 ;
  assign n15172 = n5099 & n5379 ;
  assign n15173 = n7678 & n15172 ;
  assign n15174 = n8317 & ~n15173 ;
  assign n15175 = ~n5099 & n8318 ;
  assign n15176 = n15174 | n15175 ;
  assign n15177 = n8317 | n10116 ;
  assign n15178 = ( x232 & n15176 ) | ( x232 & n15177 ) | ( n15176 & n15177 ) ;
  assign n15179 = ~n15176 & n15178 ;
  assign n15180 = ~x232 & n10116 ;
  assign n15181 = ( x39 & n15179 ) | ( x39 & ~n15180 ) | ( n15179 & ~n15180 ) ;
  assign n15182 = ~n15179 & n15181 ;
  assign n15183 = ( n9901 & n15171 ) | ( n9901 & ~n15182 ) | ( n15171 & ~n15182 ) ;
  assign n15184 = ~n9901 & n15183 ;
  assign n15185 = ~x138 & n15184 ;
  assign n15186 = x118 | n12166 ;
  assign n15187 = x139 | n15186 ;
  assign n15188 = ( n15169 & ~n15185 ) | ( n15169 & n15187 ) | ( ~n15185 & n15187 ) ;
  assign n15189 = ~n15169 & n15188 ;
  assign n15190 = ~x138 & n8258 ;
  assign n15191 = ~n15168 & n15190 ;
  assign n15192 = n15184 & ~n15190 ;
  assign n15193 = n15187 | n15192 ;
  assign n15194 = ( ~n15189 & n15191 ) | ( ~n15189 & n15193 ) | ( n15191 & n15193 ) ;
  assign n15195 = ~n15189 & n15194 ;
  assign n15196 = x55 & ~n15164 ;
  assign n15197 = ~x191 & n15116 ;
  assign n15198 = x169 | n7699 ;
  assign n15199 = n7669 & ~n15198 ;
  assign n15200 = ( n7669 & ~n15124 ) | ( n7669 & n15199 ) | ( ~n15124 & n15199 ) ;
  assign n15201 = ~n15197 & n15200 ;
  assign n15202 = ( n7671 & n15197 ) | ( n7671 & ~n15201 ) | ( n15197 & ~n15201 ) ;
  assign n15203 = x191 & n15129 ;
  assign n15204 = ( x232 & n15202 ) | ( x232 & n15203 ) | ( n15202 & n15203 ) ;
  assign n15205 = n15203 ^ n15202 ^ 1'b0 ;
  assign n15206 = ( x232 & n15204 ) | ( x232 & n15205 ) | ( n15204 & n15205 ) ;
  assign n15207 = ( x39 & n15123 ) | ( x39 & n15206 ) | ( n15123 & n15206 ) ;
  assign n15208 = n15206 ^ n15123 ^ 1'b0 ;
  assign n15209 = ( x39 & n15207 ) | ( x39 & n15208 ) | ( n15207 & n15208 ) ;
  assign n15210 = n8050 & ~n14371 ;
  assign n15211 = x169 & n7980 ;
  assign n15212 = ( x299 & n15210 ) | ( x299 & n15211 ) | ( n15210 & n15211 ) ;
  assign n15213 = n15211 ^ n15210 ^ 1'b0 ;
  assign n15214 = ( x299 & n15212 ) | ( x299 & n15213 ) | ( n15212 & n15213 ) ;
  assign n15215 = ~x191 & n15139 ;
  assign n15216 = x232 & ~n15215 ;
  assign n15217 = x191 & n15152 ;
  assign n15218 = ( n15214 & n15216 ) | ( n15214 & ~n15217 ) | ( n15216 & ~n15217 ) ;
  assign n15219 = ~n15214 & n15218 ;
  assign n15220 = ( x39 & n15142 ) | ( x39 & ~n15219 ) | ( n15142 & ~n15219 ) ;
  assign n15221 = ~x39 & n15220 ;
  assign n15222 = ( n1205 & ~n15209 ) | ( n1205 & n15221 ) | ( ~n15209 & n15221 ) ;
  assign n15223 = n15209 | n15222 ;
  assign n15224 = x87 | n15223 ;
  assign n15225 = ( ~x87 & n15113 ) | ( ~x87 & n15224 ) | ( n15113 & n15224 ) ;
  assign n15226 = x92 | n15225 ;
  assign n15227 = ( ~x92 & n15112 ) | ( ~x92 & n15226 ) | ( n15112 & n15226 ) ;
  assign n15228 = x55 | n15227 ;
  assign n15229 = ( ~x55 & n15196 ) | ( ~x55 & n15228 ) | ( n15196 & n15228 ) ;
  assign n15230 = n2109 | n15229 ;
  assign n15231 = ( ~n2109 & n8298 ) | ( ~n2109 & n15230 ) | ( n8298 & n15230 ) ;
  assign n15232 = x139 & ~n15231 ;
  assign n15233 = n12242 & ~n14331 ;
  assign n15234 = x39 | n15233 ;
  assign n15235 = n7627 & ~n15173 ;
  assign n15236 = n10112 | n14356 ;
  assign n15237 = ~n15235 & n15236 ;
  assign n15238 = ~n5099 & n7628 ;
  assign n15239 = n10115 | n15238 ;
  assign n15240 = x232 & ~n15239 ;
  assign n15241 = n15237 & n15240 ;
  assign n15242 = ( x39 & n15180 ) | ( x39 & ~n15241 ) | ( n15180 & ~n15241 ) ;
  assign n15243 = ~n15180 & n15242 ;
  assign n15244 = ( n9901 & n15234 ) | ( n9901 & ~n15243 ) | ( n15234 & ~n15243 ) ;
  assign n15245 = ~n9901 & n15244 ;
  assign n15246 = ~x139 & n15245 ;
  assign n15247 = ( n15186 & n15232 ) | ( n15186 & ~n15246 ) | ( n15232 & ~n15246 ) ;
  assign n15248 = ~n15232 & n15247 ;
  assign n15249 = ~x139 & n8259 ;
  assign n15250 = n15245 & ~n15249 ;
  assign n15251 = n15186 | n15250 ;
  assign n15252 = ~n15231 & n15249 ;
  assign n15253 = ( ~n15248 & n15251 ) | ( ~n15248 & n15252 ) | ( n15251 & n15252 ) ;
  assign n15254 = ~n15248 & n15253 ;
  assign n15334 = n5069 | n5362 ;
  assign n15335 = ~x120 & n15334 ;
  assign n15336 = ( n1292 & n15334 ) | ( n1292 & n15335 ) | ( n15334 & n15335 ) ;
  assign n15337 = n1611 & ~n15336 ;
  assign n15510 = x621 & x1091 ;
  assign n15531 = n15337 & n15510 ;
  assign n15532 = ~n5075 & n15531 ;
  assign n15340 = ~n1292 & n1611 ;
  assign n15341 = x120 & ~n15340 ;
  assign n15339 = n5072 & n12778 ;
  assign n15342 = ( x120 & n15339 ) | ( x120 & n15341 ) | ( n15339 & n15341 ) ;
  assign n15343 = x1091 & ~n15342 ;
  assign n15549 = ( n15337 & n15341 ) | ( n15337 & n15343 ) | ( n15341 & n15343 ) ;
  assign n15557 = x621 & n15549 ;
  assign n15558 = n5075 & n15557 ;
  assign n15559 = ( x603 & n15532 ) | ( x603 & ~n15558 ) | ( n15532 & ~n15558 ) ;
  assign n15560 = ~n15532 & n15559 ;
  assign n15355 = n5075 | n15337 ;
  assign n15344 = x1091 | n15341 ;
  assign n15345 = x120 & x824 ;
  assign n15346 = n5072 & n15345 ;
  assign n15347 = ( ~n15343 & n15344 ) | ( ~n15343 & n15346 ) | ( n15344 & n15346 ) ;
  assign n15348 = ~n15343 & n15347 ;
  assign n15349 = n1611 & ~n15334 ;
  assign n15350 = ( x120 & ~n15348 ) | ( x120 & n15349 ) | ( ~n15348 & n15349 ) ;
  assign n15351 = ~n15348 & n15350 ;
  assign n15356 = n5075 & ~n15351 ;
  assign n15357 = n15355 & ~n15356 ;
  assign n15561 = n5078 & n15357 ;
  assign n15562 = ~n15560 & n15561 ;
  assign n15443 = n15337 ^ x603 ^ 1'b0 ;
  assign n15689 = x665 & x1091 ;
  assign n15697 = n15337 & ~n15689 ;
  assign n15698 = x603 & ~x665 ;
  assign n15699 = ( n15443 & n15697 ) | ( n15443 & n15698 ) | ( n15697 & n15698 ) ;
  assign n15750 = n15562 & n15699 ;
  assign n15382 = x661 | x681 ;
  assign n15383 = x662 | n15382 ;
  assign n15693 = x680 & n15383 ;
  assign n15524 = x603 & ~n15510 ;
  assign n15525 = n15337 & ~n15524 ;
  assign n15694 = n15525 & ~n15689 ;
  assign n15695 = x616 & ~n15694 ;
  assign n15696 = n15693 & ~n15695 ;
  assign n15526 = x614 | x642 ;
  assign n15527 = x616 | n15526 ;
  assign n15528 = n15525 & n15527 ;
  assign n15529 = x603 | n15337 ;
  assign n15530 = ~n15527 & n15529 ;
  assign n15563 = n15530 & ~n15560 ;
  assign n15564 = n15528 | n15563 ;
  assign n15751 = n15564 & ~n15689 ;
  assign n15752 = x616 | n15751 ;
  assign n15753 = n15696 & n15752 ;
  assign n15754 = n15750 | n15753 ;
  assign n15755 = ~n5061 & n15754 ;
  assign n15338 = n5075 & n15337 ;
  assign n15352 = ~n5075 & n15351 ;
  assign n15353 = n15338 | n15352 ;
  assign n15547 = n1611 & ~n15524 ;
  assign n15548 = n15353 & n15547 ;
  assign n15756 = n15548 & n15699 ;
  assign n15757 = x616 & ~n15756 ;
  assign n15758 = ~n15560 & n15699 ;
  assign n15759 = x642 | n15758 ;
  assign n15760 = n15756 & n15759 ;
  assign n15761 = n5080 | n15760 ;
  assign n15762 = x614 & ~x616 ;
  assign n15763 = ~n15756 & n15762 ;
  assign n15764 = n15761 & ~n15763 ;
  assign n15765 = ~n15757 & n15764 ;
  assign n15766 = n15383 & ~n15765 ;
  assign n15690 = n15524 | n15689 ;
  assign n15691 = x680 & ~n15690 ;
  assign n15767 = n15351 & n15691 ;
  assign n15768 = n15693 | n15767 ;
  assign n15769 = ~n15766 & n15768 ;
  assign n15770 = n5061 & n15769 ;
  assign n15771 = ( x215 & n15755 ) | ( x215 & ~n15770 ) | ( n15755 & ~n15770 ) ;
  assign n15772 = ~n15755 & n15771 ;
  assign n15436 = ~n2263 & n15337 ;
  assign n15692 = n15436 & n15691 ;
  assign n15415 = n1614 & n15349 ;
  assign n15409 = n5362 | n8852 ;
  assign n15410 = x1092 & ~n15409 ;
  assign n15416 = x829 & ~n15410 ;
  assign n15408 = ~x824 & n15334 ;
  assign n15411 = n9656 | n15410 ;
  assign n15412 = ~n15408 & n15411 ;
  assign n15417 = x829 | n15412 ;
  assign n15418 = ( n6422 & n15416 ) | ( n6422 & n15417 ) | ( n15416 & n15417 ) ;
  assign n15419 = ~n15416 & n15418 ;
  assign n15420 = ( x1091 & n15415 ) | ( x1091 & n15419 ) | ( n15415 & n15419 ) ;
  assign n15421 = n15419 ^ n15415 ^ 1'b0 ;
  assign n15422 = ( x1091 & n15420 ) | ( x1091 & n15421 ) | ( n15420 & n15421 ) ;
  assign n15423 = x120 | n15422 ;
  assign n15424 = ~n15341 & n15423 ;
  assign n15512 = n15424 & n15510 ;
  assign n15533 = n5075 & n15512 ;
  assign n15534 = ( x603 & n15532 ) | ( x603 & ~n15533 ) | ( n15532 & ~n15533 ) ;
  assign n15535 = ~n15532 & n15534 ;
  assign n15700 = ~n15535 & n15699 ;
  assign n15701 = ~n15526 & n15700 ;
  assign n15702 = n15526 & n15694 ;
  assign n15703 = ( x616 & ~n15701 ) | ( x616 & n15702 ) | ( ~n15701 & n15702 ) ;
  assign n15704 = n15701 | n15703 ;
  assign n15705 = n15696 & n15704 ;
  assign n15413 = ( x120 & n12552 ) | ( x120 & n15412 ) | ( n12552 & n15412 ) ;
  assign n15414 = ~n15344 & n15413 ;
  assign n15425 = n15414 | n15424 ;
  assign n15444 = n5075 | n15425 ;
  assign n15445 = n15444 ^ n15425 ^ n15355 ;
  assign n15706 = n15510 & n15698 ;
  assign n15707 = x603 & ~n15445 ;
  assign n15708 = n15706 | n15707 ;
  assign n15713 = n15337 & n15689 ;
  assign n15709 = n15338 & n15689 ;
  assign n15710 = n15424 & n15689 ;
  assign n15711 = ~n5075 & n15710 ;
  assign n15712 = n15709 | n15711 ;
  assign n15714 = n15713 ^ n15712 ^ n15710 ;
  assign n15715 = ( x603 & ~n15708 ) | ( x603 & n15714 ) | ( ~n15708 & n15714 ) ;
  assign n15716 = ~n15708 & n15715 ;
  assign n15717 = ( x681 & n5077 ) | ( x681 & ~n15716 ) | ( n5077 & ~n15716 ) ;
  assign n15718 = ~x681 & n15717 ;
  assign n15719 = n15445 & n15718 ;
  assign n15720 = n15705 | n15719 ;
  assign n15721 = ( n2263 & n5061 ) | ( n2263 & n15720 ) | ( n5061 & n15720 ) ;
  assign n15722 = n2263 & n15721 ;
  assign n15723 = x665 & ~n15414 ;
  assign n15724 = n15425 & ~n15723 ;
  assign n15725 = n5078 & n15724 ;
  assign n15726 = ~x665 & n15512 ;
  assign n15727 = x603 & ~n15726 ;
  assign n15728 = n15725 & ~n15727 ;
  assign n15729 = n15693 | n15728 ;
  assign n15730 = ~x662 & n15382 ;
  assign n15426 = ~n5075 & n15425 ;
  assign n15427 = n15338 | n15426 ;
  assign n15511 = n15338 & n15510 ;
  assign n15513 = ~n5075 & n15512 ;
  assign n15514 = ( x603 & n15511 ) | ( x603 & ~n15513 ) | ( n15511 & ~n15513 ) ;
  assign n15515 = ~n15511 & n15514 ;
  assign n15516 = n15427 & ~n15515 ;
  assign n15731 = n15697 | n15724 ;
  assign n15732 = n15516 & n15731 ;
  assign n15733 = x616 & ~n15732 ;
  assign n15734 = n15726 ^ x603 ^ 1'b0 ;
  assign n15735 = n15427 & n15731 ;
  assign n15736 = ( n15726 & ~n15734 ) | ( n15726 & n15735 ) | ( ~n15734 & n15735 ) ;
  assign n15737 = ~n15526 & n15736 ;
  assign n15738 = n15527 | n15736 ;
  assign n15739 = n15732 & n15738 ;
  assign n15740 = ( x616 & ~n15737 ) | ( x616 & n15739 ) | ( ~n15737 & n15739 ) ;
  assign n15741 = n15737 | n15740 ;
  assign n15742 = ~n15733 & n15741 ;
  assign n15743 = ( x662 & n15730 ) | ( x662 & ~n15742 ) | ( n15730 & ~n15742 ) ;
  assign n15744 = n15729 & ~n15743 ;
  assign n15745 = n15744 ^ n15722 ^ 1'b0 ;
  assign n15746 = ( ~n5061 & n15744 ) | ( ~n5061 & n15745 ) | ( n15744 & n15745 ) ;
  assign n15747 = ( n15722 & ~n15745 ) | ( n15722 & n15746 ) | ( ~n15745 & n15746 ) ;
  assign n15748 = ( x215 & ~n15692 ) | ( x215 & n15747 ) | ( ~n15692 & n15747 ) ;
  assign n15749 = n15692 | n15748 ;
  assign n15773 = n15772 ^ n15749 ^ 1'b0 ;
  assign n15774 = ( x299 & ~n15749 ) | ( x299 & n15772 ) | ( ~n15749 & n15772 ) ;
  assign n15775 = ( x299 & ~n15773 ) | ( x299 & n15774 ) | ( ~n15773 & n15774 ) ;
  assign n15478 = ~n1359 & n15337 ;
  assign n15626 = n15478 & n15524 ;
  assign n15776 = x223 | n15626 ;
  assign n15591 = n1611 & n15524 ;
  assign n15777 = x680 & ~n15689 ;
  assign n15778 = n1611 & n15777 ;
  assign n15779 = ( n1611 & n15591 ) | ( n1611 & n15778 ) | ( n15591 & n15778 ) ;
  assign n15780 = n15337 & n15779 ;
  assign n15781 = n1359 | n15780 ;
  assign n15782 = n5114 & n15744 ;
  assign n15783 = ~n5114 & n15720 ;
  assign n15784 = ( n1359 & n15782 ) | ( n1359 & ~n15783 ) | ( n15782 & ~n15783 ) ;
  assign n15785 = ~n15782 & n15784 ;
  assign n15786 = ( n15776 & n15781 ) | ( n15776 & ~n15785 ) | ( n15781 & ~n15785 ) ;
  assign n15787 = ~n15776 & n15786 ;
  assign n15788 = n5114 & ~n15769 ;
  assign n15789 = n5114 | n15754 ;
  assign n15790 = x223 & n15789 ;
  assign n15791 = n15790 ^ n15788 ^ 1'b0 ;
  assign n15792 = ( n15788 & n15790 ) | ( n15788 & n15791 ) | ( n15790 & n15791 ) ;
  assign n15793 = ( x299 & ~n15788 ) | ( x299 & n15792 ) | ( ~n15788 & n15792 ) ;
  assign n15794 = ( ~n15775 & n15787 ) | ( ~n15775 & n15793 ) | ( n15787 & n15793 ) ;
  assign n15795 = ~n15775 & n15794 ;
  assign n15796 = x140 & n15795 ;
  assign n15797 = x761 & ~n15796 ;
  assign n15595 = n15337 & n15524 ;
  assign n15608 = n15351 & n15595 ;
  assign n15798 = x665 & n15549 ;
  assign n15799 = n15608 | n15798 ;
  assign n15800 = ~x603 & n15709 ;
  assign n15801 = n15799 | n15800 ;
  assign n15609 = n15353 & n15595 ;
  assign n15802 = n15709 | n15798 ;
  assign n15803 = n15609 | n15802 ;
  assign n15804 = n15801 ^ n15527 ^ 1'b0 ;
  assign n15805 = ( n15801 & n15803 ) | ( n15801 & n15804 ) | ( n15803 & n15804 ) ;
  assign n15806 = n15693 & ~n15805 ;
  assign n15354 = n15337 ^ n5079 ^ 1'b0 ;
  assign n15358 = ( n15337 & n15354 ) | ( n15337 & n15357 ) | ( n15354 & n15357 ) ;
  assign n15359 = x614 | n15358 ;
  assign n15360 = n15353 & n15359 ;
  assign n15361 = ( x616 & n15353 ) | ( x616 & n15360 ) | ( n15353 & n15360 ) ;
  assign n15807 = x680 | n15361 ;
  assign n15808 = n5078 & ~n15799 ;
  assign n15809 = ( n15806 & n15807 ) | ( n15806 & ~n15808 ) | ( n15807 & ~n15808 ) ;
  assign n15810 = ~n15806 & n15809 ;
  assign n15811 = n5061 & ~n15810 ;
  assign n15607 = ~n15356 & n15595 ;
  assign n15812 = n5075 | n15713 ;
  assign n15813 = n5075 & ~n15798 ;
  assign n15814 = n15812 & ~n15813 ;
  assign n15815 = n5078 & ~n15814 ;
  assign n15816 = ~n15607 & n15815 ;
  assign n15367 = x616 & ~n15337 ;
  assign n15368 = ~x614 & n15351 ;
  assign n15369 = ( n15337 & n15359 ) | ( n15337 & n15368 ) | ( n15359 & n15368 ) ;
  assign n15370 = x616 | n15369 ;
  assign n15371 = ~n15367 & n15370 ;
  assign n15817 = x680 | n15371 ;
  assign n15818 = n15337 & n15690 ;
  assign n15819 = x616 & ~n15818 ;
  assign n15820 = x614 & ~n15818 ;
  assign n15821 = x642 & ~n15818 ;
  assign n15822 = x642 | n15814 ;
  assign n15823 = n15607 | n15822 ;
  assign n15824 = n15801 | n15823 ;
  assign n15825 = ~n15821 & n15824 ;
  assign n15826 = x614 | n15825 ;
  assign n15827 = ~n15820 & n15826 ;
  assign n15828 = x616 | n15827 ;
  assign n15829 = ~n15819 & n15828 ;
  assign n15830 = n15693 & ~n15829 ;
  assign n15831 = ( n15816 & n15817 ) | ( n15816 & ~n15830 ) | ( n15817 & ~n15830 ) ;
  assign n15832 = ~n15816 & n15831 ;
  assign n15833 = n5061 | n15832 ;
  assign n15834 = ( x215 & n15811 ) | ( x215 & n15833 ) | ( n15811 & n15833 ) ;
  assign n15835 = ~n15811 & n15834 ;
  assign n15446 = ( n15337 & n15443 ) | ( n15337 & n15445 ) | ( n15443 & n15445 ) ;
  assign n15447 = ( n15337 & n15354 ) | ( n15337 & n15446 ) | ( n15354 & n15446 ) ;
  assign n15463 = n15337 ^ x614 ^ 1'b0 ;
  assign n15464 = ( n15337 & n15447 ) | ( n15337 & ~n15463 ) | ( n15447 & ~n15463 ) ;
  assign n15465 = x616 | n15464 ;
  assign n15836 = ( x616 & n15465 ) | ( x616 & n15690 ) | ( n15465 & n15690 ) ;
  assign n15837 = ~n15819 & n15836 ;
  assign n15838 = n15693 & ~n15837 ;
  assign n15466 = ~n15367 & n15465 ;
  assign n15839 = x680 | n15466 ;
  assign n15840 = ( ~n15718 & n15838 ) | ( ~n15718 & n15839 ) | ( n15838 & n15839 ) ;
  assign n15841 = ~n15838 & n15840 ;
  assign n15428 = n15425 ^ n5081 ^ 1'b0 ;
  assign n15429 = ( n15425 & n15427 ) | ( n15425 & ~n15428 ) | ( n15427 & ~n15428 ) ;
  assign n15842 = n15429 & n15690 ;
  assign n15843 = n15693 & ~n15842 ;
  assign n15844 = x680 | n15429 ;
  assign n15517 = x621 & ~n15414 ;
  assign n15518 = n15425 & ~n15517 ;
  assign n15845 = x603 & n15518 ;
  assign n15846 = x603 & ~x621 ;
  assign n15847 = n15710 & ~n15846 ;
  assign n15848 = n5078 & ~n15847 ;
  assign n15849 = ~n15845 & n15848 ;
  assign n15850 = ( n15843 & n15844 ) | ( n15843 & ~n15849 ) | ( n15844 & ~n15849 ) ;
  assign n15851 = ~n15843 & n15850 ;
  assign n15852 = n15841 ^ n5061 ^ 1'b0 ;
  assign n15853 = ( n15841 & n15851 ) | ( n15841 & n15852 ) | ( n15851 & n15852 ) ;
  assign n15854 = ( x216 & x221 ) | ( x216 & ~n15853 ) | ( x221 & ~n15853 ) ;
  assign n15855 = ~n15853 & n15854 ;
  assign n15856 = n15337 & ~n15691 ;
  assign n15857 = n2263 | n15856 ;
  assign n15858 = ( x215 & ~n15855 ) | ( x215 & n15857 ) | ( ~n15855 & n15857 ) ;
  assign n15859 = ~x215 & n15858 ;
  assign n15860 = ( x299 & n15835 ) | ( x299 & ~n15859 ) | ( n15835 & ~n15859 ) ;
  assign n15861 = ~n15835 & n15860 ;
  assign n15862 = n5114 & ~n15810 ;
  assign n15863 = n5114 | n15832 ;
  assign n15864 = ( x223 & n15862 ) | ( x223 & n15863 ) | ( n15862 & n15863 ) ;
  assign n15865 = ~n15862 & n15864 ;
  assign n15866 = ~n5114 & n15841 ;
  assign n15867 = n5114 & n15851 ;
  assign n15868 = ( n1359 & n15866 ) | ( n1359 & ~n15867 ) | ( n15866 & ~n15867 ) ;
  assign n15869 = ~n15866 & n15868 ;
  assign n15870 = n1359 | n15856 ;
  assign n15871 = ~x223 & n15870 ;
  assign n15872 = n15871 ^ n15869 ^ 1'b0 ;
  assign n15873 = ( n15869 & n15871 ) | ( n15869 & n15872 ) | ( n15871 & n15872 ) ;
  assign n15874 = ( n15865 & ~n15869 ) | ( n15865 & n15873 ) | ( ~n15869 & n15873 ) ;
  assign n15875 = ( x299 & ~n15861 ) | ( x299 & n15874 ) | ( ~n15861 & n15874 ) ;
  assign n15876 = ~n15861 & n15875 ;
  assign n15877 = x140 | n15876 ;
  assign n15878 = n15797 & n15877 ;
  assign n15610 = ( n15527 & n15608 ) | ( n15527 & n15609 ) | ( n15608 & n15609 ) ;
  assign n15611 = ~n5078 & n15610 ;
  assign n15879 = n15608 | n15611 ;
  assign n15880 = n15353 & n15697 ;
  assign n15881 = ~n15356 & n15697 ;
  assign n15882 = n15383 | n15881 ;
  assign n15883 = x680 & n15882 ;
  assign n15884 = n15697 ^ n5081 ^ 1'b0 ;
  assign n15885 = ( n15697 & n15881 ) | ( n15697 & n15884 ) | ( n15881 & n15884 ) ;
  assign n15886 = n15883 & n15885 ;
  assign n15887 = n15880 & n15886 ;
  assign n15888 = n15879 | n15887 ;
  assign n15889 = n5061 & n15888 ;
  assign n15890 = n15689 & ~n15846 ;
  assign n15891 = n15337 & ~n15890 ;
  assign n15892 = n15527 & n15891 ;
  assign n15893 = n15693 & ~n15892 ;
  assign n15894 = n15607 | n15885 ;
  assign n15895 = ~n15527 & n15894 ;
  assign n15896 = n15893 & ~n15895 ;
  assign n15612 = n15607 | n15611 ;
  assign n15897 = ( n15612 & n15883 ) | ( n15612 & ~n15896 ) | ( n15883 & ~n15896 ) ;
  assign n15898 = ~n15896 & n15897 ;
  assign n15899 = ~n5061 & n15898 ;
  assign n15900 = ( x215 & n15889 ) | ( x215 & ~n15899 ) | ( n15889 & ~n15899 ) ;
  assign n15901 = ~n15889 & n15900 ;
  assign n15902 = n15736 | n15845 ;
  assign n15903 = ~n15527 & n15902 ;
  assign n15904 = n15427 & n15524 ;
  assign n15905 = n15735 | n15904 ;
  assign n15906 = n15527 & n15905 ;
  assign n15907 = ( n15693 & n15903 ) | ( n15693 & ~n15906 ) | ( n15903 & ~n15906 ) ;
  assign n15908 = ~n15903 & n15907 ;
  assign n15430 = n5078 & n15425 ;
  assign n15431 = ~n5078 & n15427 ;
  assign n15432 = n15430 | n15431 ;
  assign n15433 = ( n15425 & n15429 ) | ( n15425 & n15432 ) | ( n15429 & n15432 ) ;
  assign n15601 = n15433 & n15524 ;
  assign n15909 = n15693 | n15725 ;
  assign n15910 = ( n15601 & ~n15908 ) | ( n15601 & n15909 ) | ( ~n15908 & n15909 ) ;
  assign n15911 = ~n15908 & n15910 ;
  assign n15594 = n15445 & n15524 ;
  assign n15912 = n15445 & n15731 ;
  assign n15913 = n5078 & ~n15912 ;
  assign n15914 = ~n15594 & n15913 ;
  assign n15596 = n15594 ^ n15527 ^ 1'b0 ;
  assign n15597 = ( n15594 & n15595 ) | ( n15594 & n15596 ) | ( n15595 & n15596 ) ;
  assign n15915 = ( x680 & n15597 ) | ( x680 & ~n15914 ) | ( n15597 & ~n15914 ) ;
  assign n15916 = ~n15914 & n15915 ;
  assign n15917 = n15594 | n15700 ;
  assign n15918 = ~n15527 & n15917 ;
  assign n15919 = n15918 ^ n15916 ^ 1'b0 ;
  assign n15920 = ( ~n15893 & n15918 ) | ( ~n15893 & n15919 ) | ( n15918 & n15919 ) ;
  assign n15921 = ( n15916 & ~n15919 ) | ( n15916 & n15920 ) | ( ~n15919 & n15920 ) ;
  assign n15922 = n15911 ^ n5061 ^ 1'b0 ;
  assign n15923 = ( n15911 & n15921 ) | ( n15911 & ~n15922 ) | ( n15921 & ~n15922 ) ;
  assign n15924 = n2263 & n15923 ;
  assign n15925 = ~n2263 & n15780 ;
  assign n15926 = ( x215 & ~n15924 ) | ( x215 & n15925 ) | ( ~n15924 & n15925 ) ;
  assign n15927 = n15924 | n15926 ;
  assign n15928 = x299 & ~n15927 ;
  assign n15929 = ( x299 & n15901 ) | ( x299 & n15928 ) | ( n15901 & n15928 ) ;
  assign n15930 = n5114 | n15898 ;
  assign n15931 = n15930 ^ x299 ^ 1'b0 ;
  assign n15932 = n5114 & ~n15888 ;
  assign n15933 = x223 & ~n15932 ;
  assign n15934 = ( n15930 & ~n15931 ) | ( n15930 & n15933 ) | ( ~n15931 & n15933 ) ;
  assign n15935 = ( x299 & n15931 ) | ( x299 & n15934 ) | ( n15931 & n15934 ) ;
  assign n15936 = ~n5114 & n15921 ;
  assign n15937 = n5114 & n15911 ;
  assign n15938 = ( n1359 & n15936 ) | ( n1359 & ~n15937 ) | ( n15936 & ~n15937 ) ;
  assign n15939 = ~n15936 & n15938 ;
  assign n15940 = ( x223 & n15781 ) | ( x223 & ~n15939 ) | ( n15781 & ~n15939 ) ;
  assign n15941 = ~x223 & n15940 ;
  assign n15942 = ( ~n15929 & n15935 ) | ( ~n15929 & n15941 ) | ( n15935 & n15941 ) ;
  assign n15943 = ~n15929 & n15942 ;
  assign n15944 = x140 & n15943 ;
  assign n15945 = n15429 & ~n15524 ;
  assign n15946 = x680 | n15945 ;
  assign n15947 = ~n5081 & n15709 ;
  assign n15948 = ~n5490 & n15710 ;
  assign n15949 = n15947 | n15948 ;
  assign n15950 = n15890 & n15949 ;
  assign n15951 = n15693 & ~n15950 ;
  assign n15952 = ( n15848 & n15946 ) | ( n15848 & ~n15951 ) | ( n15946 & ~n15951 ) ;
  assign n15953 = ~n15848 & n15952 ;
  assign n15954 = n15713 & ~n15846 ;
  assign n15955 = n15527 & n15954 ;
  assign n15536 = n15530 & ~n15535 ;
  assign n15956 = n15536 & n15689 ;
  assign n15957 = ( n15693 & n15955 ) | ( n15693 & ~n15956 ) | ( n15955 & ~n15956 ) ;
  assign n15958 = ~n15955 & n15957 ;
  assign n15959 = n15714 & n15890 ;
  assign n15960 = n5078 & ~n15959 ;
  assign n15537 = n15528 | n15536 ;
  assign n15961 = x680 | n15537 ;
  assign n15962 = ( n15958 & ~n15960 ) | ( n15958 & n15961 ) | ( ~n15960 & n15961 ) ;
  assign n15963 = ~n15958 & n15962 ;
  assign n15964 = n15953 ^ n5114 ^ 1'b0 ;
  assign n15965 = ( n15953 & n15963 ) | ( n15953 & ~n15964 ) | ( n15963 & ~n15964 ) ;
  assign n15966 = n1359 & n15965 ;
  assign n15967 = n15524 | n15777 ;
  assign n15968 = n15340 & ~n15967 ;
  assign n15969 = ~n15335 & n15968 ;
  assign n15970 = ~n1359 & n15969 ;
  assign n15971 = ( x223 & ~n15966 ) | ( x223 & n15970 ) | ( ~n15966 & n15970 ) ;
  assign n15972 = n15966 | n15971 ;
  assign n15973 = x680 & ~n15798 ;
  assign n15974 = n15846 | n15973 ;
  assign n15975 = n5078 & n15974 ;
  assign n15550 = n5081 & ~n15549 ;
  assign n15551 = n15548 & ~n15550 ;
  assign n15976 = ( x680 & n15551 ) | ( x680 & ~n15975 ) | ( n15551 & ~n15975 ) ;
  assign n15977 = ~n15975 & n15976 ;
  assign n15978 = n15564 & n15802 ;
  assign n15979 = n15978 ^ n15977 ^ 1'b0 ;
  assign n15980 = ( ~n15693 & n15978 ) | ( ~n15693 & n15979 ) | ( n15978 & n15979 ) ;
  assign n15981 = ( n15977 & ~n15979 ) | ( n15977 & n15980 ) | ( ~n15979 & n15980 ) ;
  assign n15982 = n5114 & n15981 ;
  assign n15983 = n5078 & ~n15846 ;
  assign n15984 = n15814 & n15983 ;
  assign n15565 = ~n5078 & n15564 ;
  assign n15985 = n15565 & ~n15777 ;
  assign n15986 = n15984 | n15985 ;
  assign n15987 = ~n5114 & n15986 ;
  assign n15988 = x223 & ~n15987 ;
  assign n15989 = n15972 & ~n15988 ;
  assign n15990 = ( n15972 & n15982 ) | ( n15972 & n15989 ) | ( n15982 & n15989 ) ;
  assign n15991 = n15953 ^ n5061 ^ 1'b0 ;
  assign n15992 = ( n15953 & n15963 ) | ( n15953 & ~n15991 ) | ( n15963 & ~n15991 ) ;
  assign n15993 = n2263 & n15992 ;
  assign n15994 = ~n2263 & n15969 ;
  assign n15995 = ( x215 & ~n15993 ) | ( x215 & n15994 ) | ( ~n15993 & n15994 ) ;
  assign n15996 = n15993 | n15995 ;
  assign n15997 = n5061 & n15981 ;
  assign n15998 = ~n5061 & n15986 ;
  assign n15999 = x215 & ~n15998 ;
  assign n16000 = n15996 & ~n15999 ;
  assign n16001 = ( n15996 & n15997 ) | ( n15996 & n16000 ) | ( n15997 & n16000 ) ;
  assign n16002 = n15990 ^ x299 ^ 1'b0 ;
  assign n16003 = ( n15990 & n16001 ) | ( n15990 & n16002 ) | ( n16001 & n16002 ) ;
  assign n16004 = x140 | n16003 ;
  assign n16005 = ( x761 & ~n15944 ) | ( x761 & n16004 ) | ( ~n15944 & n16004 ) ;
  assign n16006 = ~x761 & n16005 ;
  assign n16007 = ( x39 & n15878 ) | ( x39 & n16006 ) | ( n15878 & n16006 ) ;
  assign n16008 = n16006 ^ n15878 ^ 1'b0 ;
  assign n16009 = ( x39 & n16007 ) | ( x39 & n16008 ) | ( n16007 & n16008 ) ;
  assign n16010 = x603 & x665 ;
  assign n15256 = x40 | n8835 ;
  assign n15257 = n1412 | n1450 ;
  assign n15258 = x98 | n1475 ;
  assign n15259 = x102 | n9932 ;
  assign n15260 = ~n15258 & n15259 ;
  assign n15261 = n6379 | n10855 ;
  assign n15262 = n15260 & ~n15261 ;
  assign n15263 = ~n7471 & n15262 ;
  assign n15264 = x47 | n15263 ;
  assign n15265 = x314 & n8820 ;
  assign n15266 = n15264 | n15265 ;
  assign n15267 = ~n15257 & n15266 ;
  assign n15268 = ( x35 & ~n15256 ) | ( x35 & n15267 ) | ( ~n15256 & n15267 ) ;
  assign n15269 = ~n15256 & n15268 ;
  assign n15270 = ( x252 & n1586 ) | ( x252 & ~n15269 ) | ( n1586 & ~n15269 ) ;
  assign n15271 = ~n1586 & n15270 ;
  assign n15272 = n7472 | n7786 ;
  assign n15273 = n15262 & ~n15272 ;
  assign n15274 = x40 | n15273 ;
  assign n15275 = ~n8890 & n15274 ;
  assign n15276 = ( x252 & ~n15271 ) | ( x252 & n15275 ) | ( ~n15271 & n15275 ) ;
  assign n15277 = ~n15271 & n15276 ;
  assign n15278 = ~n1289 & n15277 ;
  assign n15279 = x1092 & n8670 ;
  assign n15280 = n1614 & n15279 ;
  assign n15281 = n15278 & n15280 ;
  assign n15282 = n1615 | n15281 ;
  assign n15283 = x1092 & ~n10860 ;
  assign n15284 = n15278 & n15283 ;
  assign n15285 = ~x95 & n5020 ;
  assign n15286 = x32 & n5283 ;
  assign n15287 = n15285 & ~n15286 ;
  assign n15288 = x88 | n15260 ;
  assign n15289 = ~n9629 & n15288 ;
  assign n15290 = x252 | n7908 ;
  assign n15291 = n15289 & ~n15290 ;
  assign n15292 = x252 & ~n8835 ;
  assign n15293 = ~n1264 & n15289 ;
  assign n15294 = x47 | n15265 ;
  assign n15295 = n15293 | n15294 ;
  assign n15296 = n15295 ^ n15257 ^ 1'b0 ;
  assign n15297 = ( n15257 & n15295 ) | ( n15257 & n15296 ) | ( n15295 & n15296 ) ;
  assign n15298 = ( x35 & ~n15257 ) | ( x35 & n15297 ) | ( ~n15257 & n15297 ) ;
  assign n15299 = n15292 & n15298 ;
  assign n15300 = ( x40 & ~n15291 ) | ( x40 & n15299 ) | ( ~n15291 & n15299 ) ;
  assign n15301 = n15291 | n15300 ;
  assign n15302 = ~n2218 & n15301 ;
  assign n15303 = x32 | n15302 ;
  assign n15304 = n15287 & n15303 ;
  assign n15305 = x824 & n15304 ;
  assign n15306 = n15284 | n15305 ;
  assign n15307 = x32 | n15277 ;
  assign n15308 = n15287 & n15307 ;
  assign n15309 = ~x824 & x829 ;
  assign n15310 = n15308 & n15309 ;
  assign n15311 = ( x1093 & n15306 ) | ( x1093 & n15310 ) | ( n15306 & n15310 ) ;
  assign n15312 = n15310 ^ n15306 ^ 1'b0 ;
  assign n15313 = ( x1093 & n15311 ) | ( x1093 & n15312 ) | ( n15311 & n15312 ) ;
  assign n15314 = ( n1614 & n15282 ) | ( n1614 & n15313 ) | ( n15282 & n15313 ) ;
  assign n15315 = n15282 & n15314 ;
  assign n15490 = x621 & n15315 ;
  assign n15505 = x198 & n15490 ;
  assign n15319 = n6425 & ~n8890 ;
  assign n15320 = n15301 & n15319 ;
  assign n15321 = n15284 | n15320 ;
  assign n15322 = x1093 & n15321 ;
  assign n15324 = ( n15281 & n15282 ) | ( n15281 & n15322 ) | ( n15282 & n15322 ) ;
  assign n15491 = x621 & n15324 ;
  assign n15504 = x198 | n15491 ;
  assign n15506 = n15505 ^ n15504 ^ x198 ;
  assign n16011 = x603 & ~n15506 ;
  assign n16012 = n16010 | n16011 ;
  assign n15323 = ~x1091 & n15322 ;
  assign n16013 = ~x665 & n15324 ;
  assign n16014 = n15323 | n16013 ;
  assign n15316 = n6489 & n15306 ;
  assign n16015 = ~x665 & n15315 ;
  assign n16016 = n15316 | n16015 ;
  assign n16017 = n16014 ^ x198 ^ 1'b0 ;
  assign n16018 = ( n16014 & n16016 ) | ( n16014 & n16017 ) | ( n16016 & n16017 ) ;
  assign n16019 = x603 | n16018 ;
  assign n16020 = ~n16012 & n16019 ;
  assign n16021 = x680 & n16020 ;
  assign n15325 = n15323 | n15324 ;
  assign n15492 = n15325 ^ x210 ^ 1'b0 ;
  assign n15493 = ( n15490 & n15491 ) | ( n15490 & n15492 ) | ( n15491 & n15492 ) ;
  assign n15494 = x603 & ~n15493 ;
  assign n16022 = n15494 | n16010 ;
  assign n16023 = n16014 ^ x210 ^ 1'b0 ;
  assign n16024 = ( n16014 & n16016 ) | ( n16014 & n16023 ) | ( n16016 & n16023 ) ;
  assign n16025 = x603 | n16024 ;
  assign n16026 = ~n16022 & n16025 ;
  assign n16027 = x680 & n16026 ;
  assign n16028 = n16021 ^ x299 ^ 1'b0 ;
  assign n16029 = ( n16021 & n16027 ) | ( n16021 & n16028 ) | ( n16027 & n16028 ) ;
  assign n16030 = x140 & ~n16029 ;
  assign n15317 = n15315 | n15316 ;
  assign n15328 = x210 & ~n15317 ;
  assign n15329 = x210 | n15325 ;
  assign n15330 = ~n15328 & n15329 ;
  assign n16031 = x665 & n15315 ;
  assign n16032 = x665 & n15324 ;
  assign n16033 = ( n15492 & n16031 ) | ( n15492 & n16032 ) | ( n16031 & n16032 ) ;
  assign n16034 = x680 & ~n16033 ;
  assign n16035 = n15330 & ~n16034 ;
  assign n15318 = x198 & ~n15317 ;
  assign n15326 = x198 | n15325 ;
  assign n15327 = ~n15318 & n15326 ;
  assign n16036 = x198 & ~n16031 ;
  assign n16037 = x198 | n16032 ;
  assign n16038 = ~n16036 & n16037 ;
  assign n16039 = ( ~x680 & n15327 ) | ( ~x680 & n16038 ) | ( n15327 & n16038 ) ;
  assign n16040 = n16039 ^ x299 ^ 1'b0 ;
  assign n16041 = ( n16035 & n16039 ) | ( n16035 & n16040 ) | ( n16039 & n16040 ) ;
  assign n16042 = n16041 ^ x680 ^ 1'b0 ;
  assign n15496 = x621 & ~n15316 ;
  assign n15497 = n15317 & ~n15496 ;
  assign n15498 = x198 & ~n15497 ;
  assign n15499 = x621 & ~n15323 ;
  assign n15500 = n15325 & ~n15499 ;
  assign n15501 = x198 | n15500 ;
  assign n15502 = ~n15498 & n15501 ;
  assign n15633 = x603 & n15502 ;
  assign n15634 = n15500 ^ x210 ^ 1'b0 ;
  assign n15635 = ( n15497 & n15500 ) | ( n15497 & n15634 ) | ( n15500 & n15634 ) ;
  assign n15636 = x603 & n15635 ;
  assign n15637 = n15633 ^ x299 ^ 1'b0 ;
  assign n15638 = ( n15633 & n15636 ) | ( n15633 & n15637 ) | ( n15636 & n15637 ) ;
  assign n16043 = ( x680 & n15638 ) | ( x680 & ~n16042 ) | ( n15638 & ~n16042 ) ;
  assign n16044 = ( n16041 & n16042 ) | ( n16041 & n16043 ) | ( n16042 & n16043 ) ;
  assign n16045 = ~x140 & n16044 ;
  assign n16046 = ( x761 & n16030 ) | ( x761 & ~n16045 ) | ( n16030 & ~n16045 ) ;
  assign n16047 = ~n16030 & n16046 ;
  assign n15495 = n15330 & ~n15494 ;
  assign n15503 = ~x603 & n15502 ;
  assign n15507 = n15503 | n15506 ;
  assign n15508 = n15495 ^ x299 ^ 1'b0 ;
  assign n15509 = ( n15495 & n15507 ) | ( n15495 & ~n15508 ) | ( n15507 & ~n15508 ) ;
  assign n16048 = n15509 & n16041 ;
  assign n16049 = ~x140 & n16048 ;
  assign n16050 = x680 & n16018 ;
  assign n16051 = x680 & n16024 ;
  assign n16052 = n16050 ^ x299 ^ 1'b0 ;
  assign n16053 = ( n16050 & n16051 ) | ( n16050 & n16052 ) | ( n16051 & n16052 ) ;
  assign n16054 = n15638 | n16053 ;
  assign n16055 = x140 & ~n16054 ;
  assign n16056 = ( x761 & ~n16049 ) | ( x761 & n16055 ) | ( ~n16049 & n16055 ) ;
  assign n16057 = n16049 | n16056 ;
  assign n16058 = ( x39 & ~n16047 ) | ( x39 & n16057 ) | ( ~n16047 & n16057 ) ;
  assign n16059 = ~x39 & n16058 ;
  assign n16060 = ( x38 & ~n16009 ) | ( x38 & n16059 ) | ( ~n16009 & n16059 ) ;
  assign n16061 = n16009 | n16060 ;
  assign n16062 = x39 & x140 ;
  assign n16063 = x140 | n15968 ;
  assign n16064 = x140 & n15779 ;
  assign n16065 = ~n1292 & n16064 ;
  assign n16066 = ( x761 & n16063 ) | ( x761 & ~n16065 ) | ( n16063 & ~n16065 ) ;
  assign n16067 = ~x761 & n16066 ;
  assign n16068 = n15340 & n15691 ;
  assign n16069 = x140 | n15340 ;
  assign n16070 = x761 & n16069 ;
  assign n16071 = ~n16068 & n16070 ;
  assign n16072 = ( ~x39 & n16067 ) | ( ~x39 & n16071 ) | ( n16067 & n16071 ) ;
  assign n16073 = ~x39 & n16072 ;
  assign n16074 = ( x38 & n16062 ) | ( x38 & ~n16073 ) | ( n16062 & ~n16073 ) ;
  assign n16075 = ~n16062 & n16074 ;
  assign n16076 = ( x738 & n16061 ) | ( x738 & ~n16075 ) | ( n16061 & ~n16075 ) ;
  assign n16077 = n16076 ^ n16061 ^ 1'b0 ;
  assign n16078 = ( x738 & n16076 ) | ( x738 & ~n16077 ) | ( n16076 & ~n16077 ) ;
  assign n15331 = n15327 ^ x299 ^ 1'b0 ;
  assign n15332 = ( n15327 & n15330 ) | ( n15327 & n15331 ) | ( n15330 & n15331 ) ;
  assign n15333 = x39 | n15332 ;
  assign n15362 = x681 & ~n15361 ;
  assign n15363 = x661 & n15361 ;
  assign n15364 = n5076 & ~n15351 ;
  assign n15365 = n5075 & ~n15364 ;
  assign n15366 = n15365 ^ n15352 ^ 1'b0 ;
  assign n15372 = n5076 | n15371 ;
  assign n15373 = ( n15365 & ~n15366 ) | ( n15365 & n15372 ) | ( ~n15366 & n15372 ) ;
  assign n15374 = ( n15352 & n15366 ) | ( n15352 & n15373 ) | ( n15366 & n15373 ) ;
  assign n15375 = ~x661 & n15374 ;
  assign n15376 = ( x681 & ~n15363 ) | ( x681 & n15375 ) | ( ~n15363 & n15375 ) ;
  assign n15377 = n15363 | n15376 ;
  assign n15378 = ~n15362 & n15377 ;
  assign n15379 = n5055 & n15378 ;
  assign n15380 = n5060 & ~n15378 ;
  assign n15381 = x680 & ~n15357 ;
  assign n15384 = x616 | n15383 ;
  assign n15385 = n15381 | n15384 ;
  assign n15386 = x680 | n15370 ;
  assign n15387 = ~n15385 & n15386 ;
  assign n15388 = ~x616 & n15383 ;
  assign n15389 = n15387 ^ n15369 ^ 1'b0 ;
  assign n15390 = ( ~n15369 & n15388 ) | ( ~n15369 & n15389 ) | ( n15388 & n15389 ) ;
  assign n15391 = ( n15369 & n15387 ) | ( n15369 & n15390 ) | ( n15387 & n15390 ) ;
  assign n15392 = x616 & n15337 ;
  assign n15393 = n15383 & n15392 ;
  assign n15394 = x680 | n15337 ;
  assign n15395 = x616 & ~n15383 ;
  assign n15396 = n15394 & n15395 ;
  assign n15397 = ~n15381 & n15396 ;
  assign n15398 = n15393 | n15397 ;
  assign n15399 = x681 | n15398 ;
  assign n15400 = n15391 | n15399 ;
  assign n15401 = x681 & ~n15371 ;
  assign n15402 = n15400 & ~n15401 ;
  assign n15403 = n5060 | n15402 ;
  assign n15404 = ( n5055 & ~n15380 ) | ( n5055 & n15403 ) | ( ~n15380 & n15403 ) ;
  assign n15405 = ~n5055 & n15404 ;
  assign n15406 = n15379 | n15405 ;
  assign n15407 = x215 & ~n15406 ;
  assign n15434 = n5055 & n15433 ;
  assign n15435 = n2263 & n15434 ;
  assign n15437 = x215 | n15436 ;
  assign n15438 = n15435 | n15437 ;
  assign n15439 = n5060 & ~n15433 ;
  assign n15440 = n5055 | n15439 ;
  assign n15441 = x614 | n5078 ;
  assign n15442 = n15367 | n15441 ;
  assign n15448 = x616 | n15447 ;
  assign n15449 = ~n15442 & n15448 ;
  assign n15450 = n15449 ^ n15445 ^ 1'b0 ;
  assign n15451 = ~x614 & n5078 ;
  assign n15452 = ( n15445 & ~n15450 ) | ( n15445 & n15451 ) | ( ~n15450 & n15451 ) ;
  assign n15453 = ( n15449 & n15450 ) | ( n15449 & n15452 ) | ( n15450 & n15452 ) ;
  assign n15454 = x680 & ~n15445 ;
  assign n15455 = x614 & ~n15383 ;
  assign n15456 = n15394 & n15455 ;
  assign n15457 = ~n15454 & n15456 ;
  assign n15458 = x614 & n15337 ;
  assign n15459 = n15383 & n15458 ;
  assign n15460 = n15457 | n15459 ;
  assign n15461 = x681 | n15460 ;
  assign n15462 = n15453 | n15461 ;
  assign n15467 = x681 & ~n15466 ;
  assign n15468 = n15462 & ~n15467 ;
  assign n15469 = ( n5060 & ~n15440 ) | ( n5060 & n15468 ) | ( ~n15440 & n15468 ) ;
  assign n15470 = ~n15440 & n15469 ;
  assign n15471 = n2263 & n15470 ;
  assign n15472 = n15438 | n15471 ;
  assign n15473 = x299 & ~n15472 ;
  assign n15474 = ( x299 & n15407 ) | ( x299 & n15473 ) | ( n15407 & n15473 ) ;
  assign n15475 = n15468 ^ n5114 ^ 1'b0 ;
  assign n15476 = ( n15433 & n15468 ) | ( n15433 & n15475 ) | ( n15468 & n15475 ) ;
  assign n15477 = n1359 & n15476 ;
  assign n15479 = x223 | n15478 ;
  assign n15480 = n15477 | n15479 ;
  assign n15481 = n15378 ^ n5114 ^ 1'b0 ;
  assign n15482 = ( n15378 & n15402 ) | ( n15378 & ~n15481 ) | ( n15402 & ~n15481 ) ;
  assign n15483 = x223 & ~n15482 ;
  assign n15484 = n15480 & ~n15483 ;
  assign n15485 = x299 | n15484 ;
  assign n15486 = ~n15474 & n15485 ;
  assign n15487 = ~x39 & n15332 ;
  assign n15488 = ( n15333 & n15486 ) | ( n15333 & n15487 ) | ( n15486 & n15487 ) ;
  assign n15489 = x761 & n15488 ;
  assign n15519 = ~x603 & n15518 ;
  assign n15520 = n15512 | n15519 ;
  assign n15521 = ( n15433 & n15516 ) | ( n15433 & n15520 ) | ( n15516 & n15520 ) ;
  assign n15522 = n15433 & n15521 ;
  assign n15523 = n5061 & ~n15522 ;
  assign n15538 = n15445 & ~n15535 ;
  assign n15539 = n15537 ^ n5078 ^ 1'b0 ;
  assign n15540 = ( n15537 & n15538 ) | ( n15537 & n15539 ) | ( n15538 & n15539 ) ;
  assign n15541 = n5061 | n15540 ;
  assign n15542 = ( n2263 & n15523 ) | ( n2263 & n15541 ) | ( n15523 & n15541 ) ;
  assign n15543 = ~n15523 & n15542 ;
  assign n15544 = ~n2263 & n15525 ;
  assign n15545 = ( ~x215 & n15543 ) | ( ~x215 & n15544 ) | ( n15543 & n15544 ) ;
  assign n15546 = ~x215 & n15545 ;
  assign n15552 = n15351 & n15547 ;
  assign n15553 = n15551 ^ n5078 ^ 1'b0 ;
  assign n15554 = ( n15551 & n15552 ) | ( n15551 & n15553 ) | ( n15552 & n15553 ) ;
  assign n15555 = n5061 & ~n15554 ;
  assign n15556 = x215 & ~n15555 ;
  assign n15566 = n15562 | n15565 ;
  assign n15567 = n5061 | n15566 ;
  assign n15568 = n15556 & n15567 ;
  assign n15569 = ( x299 & n15546 ) | ( x299 & ~n15568 ) | ( n15546 & ~n15568 ) ;
  assign n15570 = ~n15546 & n15569 ;
  assign n15571 = n5114 & ~n15522 ;
  assign n15572 = n5114 | n15540 ;
  assign n15573 = ( n1359 & n15571 ) | ( n1359 & n15572 ) | ( n15571 & n15572 ) ;
  assign n15574 = ~n15571 & n15573 ;
  assign n15575 = ~n1359 & n15525 ;
  assign n15576 = ( ~x223 & n15574 ) | ( ~x223 & n15575 ) | ( n15574 & n15575 ) ;
  assign n15577 = ~x223 & n15576 ;
  assign n15578 = n5114 & ~n15554 ;
  assign n15579 = x223 & ~n15578 ;
  assign n15580 = n15579 ^ n15577 ^ 1'b0 ;
  assign n15581 = n5114 | n15566 ;
  assign n15582 = ( n15579 & ~n15580 ) | ( n15579 & n15581 ) | ( ~n15580 & n15581 ) ;
  assign n15583 = ( n15577 & n15580 ) | ( n15577 & n15582 ) | ( n15580 & n15582 ) ;
  assign n15584 = ( x299 & ~n15570 ) | ( x299 & n15583 ) | ( ~n15570 & n15583 ) ;
  assign n15585 = ~n15570 & n15584 ;
  assign n15586 = n15509 ^ x39 ^ 1'b0 ;
  assign n15587 = ( n15509 & n15585 ) | ( n15509 & n15586 ) | ( n15585 & n15586 ) ;
  assign n15588 = ~x761 & n15587 ;
  assign n15589 = ( x140 & ~n15489 ) | ( x140 & n15588 ) | ( ~n15489 & n15588 ) ;
  assign n15590 = n15489 | n15589 ;
  assign n15592 = n2263 | n15336 ;
  assign n15593 = n15591 & ~n15592 ;
  assign n15598 = n15594 ^ n5078 ^ 1'b0 ;
  assign n15599 = ( n15594 & n15597 ) | ( n15594 & ~n15598 ) | ( n15597 & ~n15598 ) ;
  assign n15600 = n5061 | n15599 ;
  assign n15602 = n5061 & ~n15601 ;
  assign n15603 = n2263 & ~n15602 ;
  assign n15604 = n15600 & n15603 ;
  assign n15605 = ( x215 & ~n15593 ) | ( x215 & n15604 ) | ( ~n15593 & n15604 ) ;
  assign n15606 = n15593 | n15605 ;
  assign n15613 = n5061 & ~n15353 ;
  assign n15614 = n15612 & ~n15613 ;
  assign n15615 = x215 & ~n15614 ;
  assign n15616 = x299 & ~n15615 ;
  assign n15617 = n15606 & n15616 ;
  assign n15618 = n5114 & ~n15353 ;
  assign n15619 = n15612 & ~n15618 ;
  assign n15620 = x223 & ~n15619 ;
  assign n15621 = x299 | n15620 ;
  assign n15622 = n5114 | n15599 ;
  assign n15623 = n5114 & ~n15601 ;
  assign n15624 = n1359 & ~n15623 ;
  assign n15625 = n15622 & n15624 ;
  assign n15627 = ( x223 & ~n15625 ) | ( x223 & n15626 ) | ( ~n15625 & n15626 ) ;
  assign n15628 = n15625 | n15627 ;
  assign n15629 = n15628 ^ n15621 ^ 1'b0 ;
  assign n15630 = ( n15621 & n15628 ) | ( n15621 & n15629 ) | ( n15628 & n15629 ) ;
  assign n15631 = ( n15617 & ~n15621 ) | ( n15617 & n15630 ) | ( ~n15621 & n15630 ) ;
  assign n15632 = x39 & ~n15631 ;
  assign n15639 = x39 | n15638 ;
  assign n15640 = ~n15632 & n15639 ;
  assign n15641 = x140 & ~x761 ;
  assign n15642 = n15590 & ~n15641 ;
  assign n15643 = ( n15590 & ~n15640 ) | ( n15590 & n15642 ) | ( ~n15640 & n15642 ) ;
  assign n15644 = n1611 & ~n5017 ;
  assign n15645 = x140 | n15644 ;
  assign n15646 = ~n5017 & n15591 ;
  assign n15647 = ~x761 & n15646 ;
  assign n15648 = n15645 & ~n15647 ;
  assign n15649 = n15643 ^ x38 ^ 1'b0 ;
  assign n15650 = ( n15643 & n15648 ) | ( n15643 & n15649 ) | ( n15648 & n15649 ) ;
  assign n16079 = x738 & ~n15650 ;
  assign n16080 = ( n2069 & n16078 ) | ( n2069 & ~n16079 ) | ( n16078 & ~n16079 ) ;
  assign n16081 = ~n2069 & n16080 ;
  assign n16082 = n16081 ^ x140 ^ 1'b0 ;
  assign n16083 = ( ~x140 & n2069 ) | ( ~x140 & n16082 ) | ( n2069 & n16082 ) ;
  assign n16084 = ( x140 & n16081 ) | ( x140 & n16083 ) | ( n16081 & n16083 ) ;
  assign n16085 = x625 & ~n16084 ;
  assign n15255 = x140 & n2069 ;
  assign n15651 = ~n2069 & n15650 ;
  assign n15652 = n15255 | n15651 ;
  assign n16086 = x625 | n15652 ;
  assign n16087 = ( x1153 & n16085 ) | ( x1153 & n16086 ) | ( n16085 & n16086 ) ;
  assign n16088 = ~n16085 & n16087 ;
  assign n15653 = n1611 & ~n5052 ;
  assign n15654 = n15488 ^ x38 ^ 1'b0 ;
  assign n15655 = ( n15488 & n15653 ) | ( n15488 & n15654 ) | ( n15653 & n15654 ) ;
  assign n15656 = ~n2069 & n15655 ;
  assign n15657 = x140 | n15656 ;
  assign n16089 = x625 & ~n15657 ;
  assign n16090 = x1153 | n16089 ;
  assign n16091 = x140 & n16053 ;
  assign n16092 = x39 | n16091 ;
  assign n16093 = ( x140 & n16041 ) | ( x140 & ~n16092 ) | ( n16041 & ~n16092 ) ;
  assign n16094 = ~n16092 & n16093 ;
  assign n16095 = ~n5081 & n15713 ;
  assign n16096 = x680 & ~n16095 ;
  assign n16097 = ~n15814 & n16096 ;
  assign n16098 = n15815 | n16097 ;
  assign n16099 = ~n15947 & n15973 ;
  assign n16100 = n15807 & ~n16099 ;
  assign n16101 = ~n16098 & n16100 ;
  assign n16102 = n5114 & n16101 ;
  assign n16103 = n15817 & ~n16098 ;
  assign n16104 = ~n5114 & n16103 ;
  assign n16105 = ( x223 & n16102 ) | ( x223 & ~n16104 ) | ( n16102 & ~n16104 ) ;
  assign n16106 = ~n16102 & n16105 ;
  assign n16107 = n15383 & n15949 ;
  assign n16108 = ~n15383 & n15710 ;
  assign n16109 = x680 & ~n16108 ;
  assign n16110 = n15844 & ~n16109 ;
  assign n16111 = ( n15844 & n16107 ) | ( n15844 & n16110 ) | ( n16107 & n16110 ) ;
  assign n16112 = n5114 & ~n16111 ;
  assign n16113 = n1359 & ~n16112 ;
  assign n16114 = x680 & ~n15714 ;
  assign n16115 = ( n15383 & n15839 ) | ( n15383 & ~n16114 ) | ( n15839 & ~n16114 ) ;
  assign n16116 = ~n15383 & n16115 ;
  assign n16117 = n5081 & n15714 ;
  assign n16118 = n16096 & ~n16117 ;
  assign n16119 = n15839 & ~n16118 ;
  assign n16120 = ( ~n15383 & n16115 ) | ( ~n15383 & n16119 ) | ( n16115 & n16119 ) ;
  assign n16121 = ( n15383 & n16116 ) | ( n15383 & n16120 ) | ( n16116 & n16120 ) ;
  assign n16122 = n5114 | n16121 ;
  assign n16123 = n16113 & n16122 ;
  assign n16124 = n1611 & ~n15777 ;
  assign n16125 = ( x223 & n15479 ) | ( x223 & n16124 ) | ( n15479 & n16124 ) ;
  assign n16126 = ( ~n16106 & n16123 ) | ( ~n16106 & n16125 ) | ( n16123 & n16125 ) ;
  assign n16127 = ~n16106 & n16126 ;
  assign n16128 = n5061 & n16101 ;
  assign n16129 = ~n5061 & n16103 ;
  assign n16130 = ( x215 & n16128 ) | ( x215 & ~n16129 ) | ( n16128 & ~n16129 ) ;
  assign n16131 = ~n16128 & n16130 ;
  assign n16132 = n5061 & ~n16111 ;
  assign n16133 = n2263 & ~n16132 ;
  assign n16134 = n5061 | n16121 ;
  assign n16135 = n16133 & n16134 ;
  assign n16136 = ~n15592 & n16124 ;
  assign n16137 = x215 | n16136 ;
  assign n16138 = ( ~n16131 & n16135 ) | ( ~n16131 & n16137 ) | ( n16135 & n16137 ) ;
  assign n16139 = ~n16131 & n16138 ;
  assign n16140 = n16127 ^ x299 ^ 1'b0 ;
  assign n16141 = ( n16127 & n16139 ) | ( n16127 & n16140 ) | ( n16139 & n16140 ) ;
  assign n16142 = x140 | n16141 ;
  assign n16143 = x680 & n15885 ;
  assign n16144 = ~n15618 & n16143 ;
  assign n16145 = n15478 & n15777 ;
  assign n16146 = ( n15697 & n15884 ) | ( n15697 & n15912 ) | ( n15884 & n15912 ) ;
  assign n16147 = n15383 & ~n16146 ;
  assign n16148 = n15383 | n15912 ;
  assign n16149 = ( x680 & n16147 ) | ( x680 & n16148 ) | ( n16147 & n16148 ) ;
  assign n16150 = ~n16147 & n16149 ;
  assign n16151 = n5114 | n16150 ;
  assign n16152 = n15429 & n15777 ;
  assign n16153 = n15383 & n16152 ;
  assign n16154 = n15725 | n16153 ;
  assign n16155 = n5114 & ~n16154 ;
  assign n16156 = n1359 & ~n16155 ;
  assign n16157 = n16151 & n16156 ;
  assign n16158 = ( ~x223 & n16145 ) | ( ~x223 & n16157 ) | ( n16145 & n16157 ) ;
  assign n16159 = ~x223 & n16158 ;
  assign n16160 = x223 & n15882 ;
  assign n16161 = n16159 ^ n16144 ^ 1'b0 ;
  assign n16162 = ( ~n16144 & n16160 ) | ( ~n16144 & n16161 ) | ( n16160 & n16161 ) ;
  assign n16163 = ( n16144 & n16159 ) | ( n16144 & n16162 ) | ( n16159 & n16162 ) ;
  assign n16164 = n15337 & n15777 ;
  assign n16165 = ~n2263 & n16164 ;
  assign n16166 = n5061 & ~n16154 ;
  assign n16167 = n5061 | n16150 ;
  assign n16168 = ( n2263 & n16166 ) | ( n2263 & n16167 ) | ( n16166 & n16167 ) ;
  assign n16169 = ~n16166 & n16168 ;
  assign n16170 = ( ~x215 & n16165 ) | ( ~x215 & n16169 ) | ( n16165 & n16169 ) ;
  assign n16171 = ~x215 & n16170 ;
  assign n16172 = ~n15613 & n16143 ;
  assign n16173 = n16172 ^ n16171 ^ 1'b0 ;
  assign n16174 = x215 & n15882 ;
  assign n16175 = ( n16172 & ~n16173 ) | ( n16172 & n16174 ) | ( ~n16173 & n16174 ) ;
  assign n16176 = ( n16171 & n16173 ) | ( n16171 & n16175 ) | ( n16173 & n16175 ) ;
  assign n16177 = n16163 ^ x299 ^ 1'b0 ;
  assign n16178 = ( n16163 & n16176 ) | ( n16163 & n16177 ) | ( n16176 & n16177 ) ;
  assign n16179 = x140 & n16178 ;
  assign n16180 = x39 & ~n16179 ;
  assign n16181 = n16142 & n16180 ;
  assign n16182 = ( ~x38 & n16094 ) | ( ~x38 & n16181 ) | ( n16094 & n16181 ) ;
  assign n16183 = ~x38 & n16182 ;
  assign n16184 = ~n5017 & n15778 ;
  assign n16185 = x38 & ~n16184 ;
  assign n16186 = n15645 & n16185 ;
  assign n16187 = ( x738 & ~n16183 ) | ( x738 & n16186 ) | ( ~n16183 & n16186 ) ;
  assign n16188 = n16183 | n16187 ;
  assign n16189 = ~x140 & x738 ;
  assign n16190 = ~n15655 & n16189 ;
  assign n16191 = n2069 | n16190 ;
  assign n16192 = ( n15255 & n16188 ) | ( n15255 & ~n16191 ) | ( n16188 & ~n16191 ) ;
  assign n16193 = n16192 ^ n16188 ^ 1'b0 ;
  assign n16194 = ( n15255 & n16192 ) | ( n15255 & ~n16193 ) | ( n16192 & ~n16193 ) ;
  assign n16195 = ( x625 & ~n16090 ) | ( x625 & n16194 ) | ( ~n16090 & n16194 ) ;
  assign n16196 = ~n16090 & n16195 ;
  assign n16197 = ( x608 & n16088 ) | ( x608 & ~n16196 ) | ( n16088 & ~n16196 ) ;
  assign n16198 = ~n16088 & n16197 ;
  assign n16199 = x625 & ~n16194 ;
  assign n16200 = x625 | n15657 ;
  assign n16201 = ( x1153 & n16199 ) | ( x1153 & n16200 ) | ( n16199 & n16200 ) ;
  assign n16202 = ~n16199 & n16201 ;
  assign n16203 = x608 | n16202 ;
  assign n16204 = x625 & ~n15652 ;
  assign n16205 = x1153 | n16204 ;
  assign n16206 = ( n16084 & n16085 ) | ( n16084 & ~n16205 ) | ( n16085 & ~n16205 ) ;
  assign n16207 = ( ~n16198 & n16203 ) | ( ~n16198 & n16206 ) | ( n16203 & n16206 ) ;
  assign n16208 = ~n16198 & n16207 ;
  assign n16209 = n16084 ^ x778 ^ 1'b0 ;
  assign n16210 = ( n16084 & n16208 ) | ( n16084 & n16209 ) | ( n16208 & n16209 ) ;
  assign n16211 = x609 & ~n16210 ;
  assign n16212 = n16196 | n16202 ;
  assign n16213 = n16194 ^ x778 ^ 1'b0 ;
  assign n16214 = ( n16194 & n16212 ) | ( n16194 & n16213 ) | ( n16212 & n16213 ) ;
  assign n16215 = x609 | n16214 ;
  assign n16216 = ( x1155 & n16211 ) | ( x1155 & n16215 ) | ( n16211 & n16215 ) ;
  assign n16217 = ~n16211 & n16216 ;
  assign n15658 = x1153 ^ x608 ^ 1'b0 ;
  assign n15659 = x778 & n15658 ;
  assign n15662 = x609 | n15659 ;
  assign n15663 = n15657 & n15662 ;
  assign n15664 = n15652 & ~n15659 ;
  assign n15665 = ~x609 & n15664 ;
  assign n15666 = n15663 | n15665 ;
  assign n16218 = ~x1155 & n15666 ;
  assign n16219 = ( x660 & n16217 ) | ( x660 & ~n16218 ) | ( n16217 & ~n16218 ) ;
  assign n16220 = ~n16217 & n16219 ;
  assign n15667 = x609 & n15664 ;
  assign n15668 = x609 & ~n15659 ;
  assign n15669 = n15657 & ~n15668 ;
  assign n15670 = n15667 | n15669 ;
  assign n16221 = x1155 & n15670 ;
  assign n16222 = x660 | n16221 ;
  assign n16223 = x609 & ~n16214 ;
  assign n16224 = x1155 | n16223 ;
  assign n16225 = ( n16210 & n16211 ) | ( n16210 & ~n16224 ) | ( n16211 & ~n16224 ) ;
  assign n16226 = ( ~n16220 & n16222 ) | ( ~n16220 & n16225 ) | ( n16222 & n16225 ) ;
  assign n16227 = ~n16220 & n16226 ;
  assign n16228 = n16210 ^ x785 ^ 1'b0 ;
  assign n16229 = ( n16210 & n16227 ) | ( n16210 & n16228 ) | ( n16227 & n16228 ) ;
  assign n16230 = x618 & ~n16229 ;
  assign n16231 = x660 | x1155 ;
  assign n16232 = x660 & x1155 ;
  assign n16233 = x785 & ~n16232 ;
  assign n16234 = n16231 & n16233 ;
  assign n16235 = n16234 ^ n15657 ^ 1'b0 ;
  assign n16236 = ( n15657 & n16214 ) | ( n15657 & ~n16235 ) | ( n16214 & ~n16235 ) ;
  assign n16237 = x618 | n16236 ;
  assign n16238 = ( x1154 & n16230 ) | ( x1154 & n16237 ) | ( n16230 & n16237 ) ;
  assign n16239 = ~n16230 & n16238 ;
  assign n15660 = n15659 ^ n15657 ^ 1'b0 ;
  assign n15661 = ( n15652 & n15657 ) | ( n15652 & ~n15660 ) | ( n15657 & ~n15660 ) ;
  assign n15671 = n15670 ^ x1155 ^ 1'b0 ;
  assign n15672 = ( n15666 & n15670 ) | ( n15666 & ~n15671 ) | ( n15670 & ~n15671 ) ;
  assign n15673 = n15661 ^ x785 ^ 1'b0 ;
  assign n15674 = ( n15661 & n15672 ) | ( n15661 & n15673 ) | ( n15672 & n15673 ) ;
  assign n15675 = x618 & ~n15674 ;
  assign n15679 = x618 & ~n15657 ;
  assign n15680 = x1154 | n15679 ;
  assign n15681 = ( n15674 & n15675 ) | ( n15674 & ~n15680 ) | ( n15675 & ~n15680 ) ;
  assign n16240 = ( x627 & ~n15681 ) | ( x627 & n16239 ) | ( ~n15681 & n16239 ) ;
  assign n16241 = ~n16239 & n16240 ;
  assign n15676 = x618 | n15657 ;
  assign n15677 = ( x1154 & n15675 ) | ( x1154 & n15676 ) | ( n15675 & n15676 ) ;
  assign n15678 = ~n15675 & n15677 ;
  assign n16242 = x627 | n15678 ;
  assign n16243 = x618 & ~n16236 ;
  assign n16244 = x1154 | n16243 ;
  assign n16245 = ( n16229 & n16230 ) | ( n16229 & ~n16244 ) | ( n16230 & ~n16244 ) ;
  assign n16246 = ( ~n16241 & n16242 ) | ( ~n16241 & n16245 ) | ( n16242 & n16245 ) ;
  assign n16247 = ~n16241 & n16246 ;
  assign n16248 = n16229 ^ x781 ^ 1'b0 ;
  assign n16249 = ( n16229 & n16247 ) | ( n16229 & n16248 ) | ( n16247 & n16248 ) ;
  assign n16250 = x619 & ~n16249 ;
  assign n16251 = x627 | x1154 ;
  assign n16252 = x627 & x1154 ;
  assign n16253 = x781 & ~n16252 ;
  assign n16254 = n16251 & n16253 ;
  assign n16255 = n16254 ^ n15657 ^ 1'b0 ;
  assign n16256 = ( n15657 & n16236 ) | ( n15657 & ~n16255 ) | ( n16236 & ~n16255 ) ;
  assign n16262 = x619 | n16256 ;
  assign n16263 = ( x1159 & n16250 ) | ( x1159 & n16262 ) | ( n16250 & n16262 ) ;
  assign n16264 = ~n16250 & n16263 ;
  assign n15682 = n15678 | n15681 ;
  assign n15683 = n15674 ^ x781 ^ 1'b0 ;
  assign n15684 = ( n15674 & n15682 ) | ( n15674 & n15683 ) | ( n15682 & n15683 ) ;
  assign n15685 = x619 & ~n15684 ;
  assign n16265 = x619 & ~n15657 ;
  assign n16266 = x1159 | n16265 ;
  assign n16267 = ( n15684 & n15685 ) | ( n15684 & ~n16266 ) | ( n15685 & ~n16266 ) ;
  assign n16268 = ( x648 & n16264 ) | ( x648 & ~n16267 ) | ( n16264 & ~n16267 ) ;
  assign n16269 = ~n16264 & n16268 ;
  assign n15686 = x619 | n15657 ;
  assign n15687 = ( x1159 & n15685 ) | ( x1159 & n15686 ) | ( n15685 & n15686 ) ;
  assign n15688 = ~n15685 & n15687 ;
  assign n16257 = x619 & ~n16256 ;
  assign n16258 = x1159 | n16257 ;
  assign n16259 = ( n16249 & n16250 ) | ( n16249 & ~n16258 ) | ( n16250 & ~n16258 ) ;
  assign n16260 = ( x648 & ~n15688 ) | ( x648 & n16259 ) | ( ~n15688 & n16259 ) ;
  assign n16261 = n15688 | n16260 ;
  assign n16270 = n16269 ^ n16261 ^ 1'b0 ;
  assign n16271 = ( x789 & ~n16261 ) | ( x789 & n16269 ) | ( ~n16261 & n16269 ) ;
  assign n16272 = ( x789 & ~n16270 ) | ( x789 & n16271 ) | ( ~n16270 & n16271 ) ;
  assign n16273 = ( x789 & n16249 ) | ( x789 & ~n16272 ) | ( n16249 & ~n16272 ) ;
  assign n16274 = ~n16272 & n16273 ;
  assign n16275 = ~x626 & n16274 ;
  assign n16276 = ~x648 & x1159 ;
  assign n16277 = x648 & ~x1159 ;
  assign n16278 = n16276 | n16277 ;
  assign n16279 = x789 & n16278 ;
  assign n16280 = n16279 ^ n15657 ^ 1'b0 ;
  assign n16281 = ( n15657 & n16256 ) | ( n15657 & ~n16280 ) | ( n16256 & ~n16280 ) ;
  assign n16282 = x626 & n16281 ;
  assign n16283 = ( x641 & ~n16275 ) | ( x641 & n16282 ) | ( ~n16275 & n16282 ) ;
  assign n16284 = n16275 | n16283 ;
  assign n16285 = ~x626 & n16281 ;
  assign n16286 = x626 & n16274 ;
  assign n16287 = ( x641 & n16285 ) | ( x641 & ~n16286 ) | ( n16285 & ~n16286 ) ;
  assign n16288 = ~n16285 & n16287 ;
  assign n16289 = x641 & x1158 ;
  assign n16290 = n15688 | n16267 ;
  assign n16291 = n15684 ^ x789 ^ 1'b0 ;
  assign n16292 = ( n15684 & n16290 ) | ( n15684 & n16291 ) | ( n16290 & n16291 ) ;
  assign n16293 = x626 & ~n16292 ;
  assign n16294 = x626 | n15657 ;
  assign n16295 = ( x1158 & n16293 ) | ( x1158 & n16294 ) | ( n16293 & n16294 ) ;
  assign n16296 = ~n16293 & n16295 ;
  assign n16297 = ( ~n16288 & n16289 ) | ( ~n16288 & n16296 ) | ( n16289 & n16296 ) ;
  assign n16298 = ~n16288 & n16297 ;
  assign n16299 = x641 | x1158 ;
  assign n16300 = x626 & ~n15657 ;
  assign n16301 = x1158 | n16300 ;
  assign n16302 = ( n16292 & n16293 ) | ( n16292 & ~n16301 ) | ( n16293 & ~n16301 ) ;
  assign n16303 = n16299 & ~n16302 ;
  assign n16304 = ~n16298 & n16303 ;
  assign n16305 = ( n16284 & n16298 ) | ( n16284 & ~n16304 ) | ( n16298 & ~n16304 ) ;
  assign n16306 = n16274 ^ x788 ^ 1'b0 ;
  assign n16307 = ( n16274 & n16305 ) | ( n16274 & n16306 ) | ( n16305 & n16306 ) ;
  assign n16308 = x628 & ~n16307 ;
  assign n16309 = n16296 | n16302 ;
  assign n16310 = n16292 ^ x788 ^ 1'b0 ;
  assign n16311 = ( n16292 & n16309 ) | ( n16292 & n16310 ) | ( n16309 & n16310 ) ;
  assign n16312 = x628 | n16311 ;
  assign n16313 = ( x1156 & n16308 ) | ( x1156 & n16312 ) | ( n16308 & n16312 ) ;
  assign n16314 = ~n16308 & n16313 ;
  assign n16315 = x628 & ~n15657 ;
  assign n16316 = x1156 | n16315 ;
  assign n16317 = x1158 ^ x641 ^ 1'b0 ;
  assign n16318 = x788 & n16317 ;
  assign n16319 = n16318 ^ n15657 ^ 1'b0 ;
  assign n16320 = ( n15657 & n16281 ) | ( n15657 & ~n16319 ) | ( n16281 & ~n16319 ) ;
  assign n16321 = x628 & ~n16320 ;
  assign n16322 = ( ~n16316 & n16320 ) | ( ~n16316 & n16321 ) | ( n16320 & n16321 ) ;
  assign n16323 = ( x629 & n16314 ) | ( x629 & ~n16322 ) | ( n16314 & ~n16322 ) ;
  assign n16324 = ~n16314 & n16323 ;
  assign n16325 = x628 | n15657 ;
  assign n16326 = ( x1156 & n16321 ) | ( x1156 & n16325 ) | ( n16321 & n16325 ) ;
  assign n16327 = ~n16321 & n16326 ;
  assign n16328 = x629 | n16327 ;
  assign n16329 = x628 & ~n16311 ;
  assign n16330 = x1156 | n16329 ;
  assign n16331 = ( n16307 & n16308 ) | ( n16307 & ~n16330 ) | ( n16308 & ~n16330 ) ;
  assign n16332 = ( ~n16324 & n16328 ) | ( ~n16324 & n16331 ) | ( n16328 & n16331 ) ;
  assign n16333 = ~n16324 & n16332 ;
  assign n16334 = n16307 ^ x792 ^ 1'b0 ;
  assign n16335 = ( n16307 & n16333 ) | ( n16307 & n16334 ) | ( n16333 & n16334 ) ;
  assign n16336 = x647 & ~n16335 ;
  assign n16337 = ~x629 & x1156 ;
  assign n16338 = x629 & ~x1156 ;
  assign n16339 = ( x792 & n16337 ) | ( x792 & n16338 ) | ( n16337 & n16338 ) ;
  assign n16340 = n16339 ^ n15657 ^ 1'b0 ;
  assign n16341 = ( n15657 & n16311 ) | ( n15657 & ~n16340 ) | ( n16311 & ~n16340 ) ;
  assign n16342 = x647 | n16341 ;
  assign n16343 = ( x1157 & n16336 ) | ( x1157 & n16342 ) | ( n16336 & n16342 ) ;
  assign n16344 = ~n16336 & n16343 ;
  assign n16345 = x647 & ~n15657 ;
  assign n16346 = x1157 | n16345 ;
  assign n16347 = n16322 | n16327 ;
  assign n16348 = n16320 ^ x792 ^ 1'b0 ;
  assign n16349 = ( n16320 & n16347 ) | ( n16320 & n16348 ) | ( n16347 & n16348 ) ;
  assign n16350 = x647 & ~n16349 ;
  assign n16351 = ( ~n16346 & n16349 ) | ( ~n16346 & n16350 ) | ( n16349 & n16350 ) ;
  assign n16352 = ( x630 & n16344 ) | ( x630 & ~n16351 ) | ( n16344 & ~n16351 ) ;
  assign n16353 = ~n16344 & n16352 ;
  assign n16354 = x647 | n15657 ;
  assign n16355 = ( x1157 & n16350 ) | ( x1157 & n16354 ) | ( n16350 & n16354 ) ;
  assign n16356 = ~n16350 & n16355 ;
  assign n16357 = x630 | n16356 ;
  assign n16358 = x647 & ~n16341 ;
  assign n16359 = x1157 | n16358 ;
  assign n16360 = ( n16335 & n16336 ) | ( n16335 & ~n16359 ) | ( n16336 & ~n16359 ) ;
  assign n16361 = ( ~n16353 & n16357 ) | ( ~n16353 & n16360 ) | ( n16357 & n16360 ) ;
  assign n16362 = ~n16353 & n16361 ;
  assign n16363 = n16335 ^ x787 ^ 1'b0 ;
  assign n16364 = ( n16335 & n16362 ) | ( n16335 & n16363 ) | ( n16362 & n16363 ) ;
  assign n16365 = x644 & ~n16364 ;
  assign n16366 = n16351 | n16356 ;
  assign n16367 = n16349 ^ x787 ^ 1'b0 ;
  assign n16368 = ( n16349 & n16366 ) | ( n16349 & n16367 ) | ( n16366 & n16367 ) ;
  assign n16369 = x644 | n16368 ;
  assign n16370 = ( x715 & n16365 ) | ( x715 & n16369 ) | ( n16365 & n16369 ) ;
  assign n16371 = ~n16365 & n16370 ;
  assign n16372 = x644 | n15657 ;
  assign n16373 = ~x630 & x1157 ;
  assign n16374 = x630 & ~x1157 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = x787 & n16375 ;
  assign n16377 = n16376 ^ n15657 ^ 1'b0 ;
  assign n16378 = ( n15657 & n16341 ) | ( n15657 & ~n16377 ) | ( n16341 & ~n16377 ) ;
  assign n16379 = x644 & ~n16378 ;
  assign n16380 = ( x715 & n16372 ) | ( x715 & ~n16379 ) | ( n16372 & ~n16379 ) ;
  assign n16381 = ~x715 & n16380 ;
  assign n16382 = ( x1160 & n16371 ) | ( x1160 & ~n16381 ) | ( n16371 & ~n16381 ) ;
  assign n16383 = ~n16371 & n16382 ;
  assign n16384 = x644 & ~n15657 ;
  assign n16385 = x715 & ~n16384 ;
  assign n16386 = ( n16378 & n16379 ) | ( n16378 & n16385 ) | ( n16379 & n16385 ) ;
  assign n16387 = x644 & ~n16368 ;
  assign n16388 = x715 | n16387 ;
  assign n16389 = ( n16364 & n16365 ) | ( n16364 & ~n16388 ) | ( n16365 & ~n16388 ) ;
  assign n16390 = ( x1160 & ~n16386 ) | ( x1160 & n16389 ) | ( ~n16386 & n16389 ) ;
  assign n16391 = n16386 | n16390 ;
  assign n16392 = ( x790 & n16383 ) | ( x790 & n16391 ) | ( n16383 & n16391 ) ;
  assign n16393 = ~n16383 & n16392 ;
  assign n16394 = ~x790 & n16364 ;
  assign n16395 = ( n7318 & ~n16393 ) | ( n7318 & n16394 ) | ( ~n16393 & n16394 ) ;
  assign n16396 = n16393 | n16395 ;
  assign n16397 = n1611 & n15659 ;
  assign n16398 = x140 | n1611 ;
  assign n16399 = ~x761 & n15591 ;
  assign n16400 = n16398 & ~n16399 ;
  assign n16401 = n16397 | n16400 ;
  assign n16402 = n1611 & ~n15668 ;
  assign n16403 = n16400 | n16402 ;
  assign n16404 = x1155 & n16403 ;
  assign n16405 = x609 & n1611 ;
  assign n16406 = n16401 | n16405 ;
  assign n16407 = ~x1155 & n16406 ;
  assign n16408 = n16404 | n16407 ;
  assign n16409 = n16401 ^ x785 ^ 1'b0 ;
  assign n16410 = ( n16401 & n16408 ) | ( n16401 & n16409 ) | ( n16408 & n16409 ) ;
  assign n16411 = ~x618 & n1611 ;
  assign n16412 = n16410 | n16411 ;
  assign n16413 = x1154 & n16412 ;
  assign n16414 = x618 & n1611 ;
  assign n16415 = n16410 | n16414 ;
  assign n16416 = ~x1154 & n16415 ;
  assign n16417 = n16413 | n16416 ;
  assign n16418 = n16410 ^ x781 ^ 1'b0 ;
  assign n16419 = ( n16410 & n16417 ) | ( n16410 & n16418 ) | ( n16417 & n16418 ) ;
  assign n16420 = x619 & ~n16419 ;
  assign n16421 = x619 | n16398 ;
  assign n16422 = ( x1159 & n16420 ) | ( x1159 & n16421 ) | ( n16420 & n16421 ) ;
  assign n16423 = ~n16420 & n16422 ;
  assign n16424 = x619 & ~n16398 ;
  assign n16425 = x1159 | n16424 ;
  assign n16426 = ( n16419 & n16420 ) | ( n16419 & ~n16425 ) | ( n16420 & ~n16425 ) ;
  assign n16427 = n16423 | n16426 ;
  assign n16428 = n16419 ^ x789 ^ 1'b0 ;
  assign n16429 = ( n16419 & n16427 ) | ( n16419 & n16428 ) | ( n16427 & n16428 ) ;
  assign n16430 = x626 & ~n16429 ;
  assign n16431 = x626 & ~n16398 ;
  assign n16432 = x1158 | n16431 ;
  assign n16433 = ( n16429 & n16430 ) | ( n16429 & ~n16432 ) | ( n16430 & ~n16432 ) ;
  assign n16434 = n16430 & ~n16433 ;
  assign n16435 = ( x1158 & n16398 ) | ( x1158 & n16431 ) | ( n16398 & n16431 ) ;
  assign n16436 = ( n16433 & ~n16434 ) | ( n16433 & n16435 ) | ( ~n16434 & n16435 ) ;
  assign n16437 = n16317 & ~n16436 ;
  assign n16438 = ~x738 & n15778 ;
  assign n16439 = n16398 & ~n16438 ;
  assign n16440 = ~x625 & n16438 ;
  assign n16441 = ~x1153 & n16398 ;
  assign n16442 = ~n16440 & n16441 ;
  assign n16443 = ( x1153 & n16439 ) | ( x1153 & n16440 ) | ( n16439 & n16440 ) ;
  assign n16444 = n16442 | n16443 ;
  assign n16445 = n16439 ^ x778 ^ 1'b0 ;
  assign n16446 = ( n16439 & n16444 ) | ( n16439 & n16445 ) | ( n16444 & n16445 ) ;
  assign n16447 = n1611 & n16234 ;
  assign n16448 = n16446 | n16447 ;
  assign n16449 = n1611 & n16254 ;
  assign n16450 = n16448 | n16449 ;
  assign n16451 = n1611 & n16279 ;
  assign n16452 = n16450 | n16451 ;
  assign n16453 = ~x626 & x1158 ;
  assign n16454 = x626 & ~x1158 ;
  assign n16455 = n16453 | n16454 ;
  assign n16456 = ~x626 & x641 ;
  assign n16457 = x626 & ~x641 ;
  assign n16458 = n16456 | n16457 ;
  assign n16459 = n16455 & n16458 ;
  assign n16460 = ~n16452 & n16459 ;
  assign n16461 = ( x788 & n16437 ) | ( x788 & n16460 ) | ( n16437 & n16460 ) ;
  assign n16462 = n16460 ^ n16437 ^ 1'b0 ;
  assign n16463 = ( x788 & n16461 ) | ( x788 & n16462 ) | ( n16461 & n16462 ) ;
  assign n16464 = x619 & ~n16450 ;
  assign n16465 = x1159 | n16464 ;
  assign n16466 = n15524 | n16439 ;
  assign n16467 = n16400 & n16466 ;
  assign n16468 = x625 & ~n16466 ;
  assign n16469 = x1153 & n16400 ;
  assign n16470 = ~n16468 & n16469 ;
  assign n16471 = ( x608 & n16442 ) | ( x608 & ~n16470 ) | ( n16442 & ~n16470 ) ;
  assign n16472 = ~n16442 & n16471 ;
  assign n16473 = x608 | n16443 ;
  assign n16474 = ( n16441 & n16467 ) | ( n16441 & n16468 ) | ( n16467 & n16468 ) ;
  assign n16475 = ( ~n16472 & n16473 ) | ( ~n16472 & n16474 ) | ( n16473 & n16474 ) ;
  assign n16476 = ~n16472 & n16475 ;
  assign n16477 = n16467 ^ x778 ^ 1'b0 ;
  assign n16478 = ( n16467 & n16476 ) | ( n16467 & n16477 ) | ( n16476 & n16477 ) ;
  assign n16479 = x609 & ~n16478 ;
  assign n16480 = x609 | n16446 ;
  assign n16481 = ( x1155 & n16479 ) | ( x1155 & n16480 ) | ( n16479 & n16480 ) ;
  assign n16482 = ~n16479 & n16481 ;
  assign n16483 = ( x660 & n16407 ) | ( x660 & ~n16482 ) | ( n16407 & ~n16482 ) ;
  assign n16484 = ~n16407 & n16483 ;
  assign n16485 = x660 | n16404 ;
  assign n16486 = x609 & ~n16446 ;
  assign n16487 = x1155 | n16486 ;
  assign n16488 = ( n16478 & n16479 ) | ( n16478 & ~n16487 ) | ( n16479 & ~n16487 ) ;
  assign n16489 = ( ~n16484 & n16485 ) | ( ~n16484 & n16488 ) | ( n16485 & n16488 ) ;
  assign n16490 = ~n16484 & n16489 ;
  assign n16491 = n16478 ^ x785 ^ 1'b0 ;
  assign n16492 = ( n16478 & n16490 ) | ( n16478 & n16491 ) | ( n16490 & n16491 ) ;
  assign n16493 = x618 & ~n16492 ;
  assign n16494 = x618 | n16448 ;
  assign n16495 = ( x1154 & n16493 ) | ( x1154 & n16494 ) | ( n16493 & n16494 ) ;
  assign n16496 = ~n16493 & n16495 ;
  assign n16497 = ( x627 & n16416 ) | ( x627 & ~n16496 ) | ( n16416 & ~n16496 ) ;
  assign n16498 = ~n16416 & n16497 ;
  assign n16499 = x627 | n16413 ;
  assign n16500 = x618 & ~n16448 ;
  assign n16501 = x1154 | n16500 ;
  assign n16502 = ( n16492 & n16493 ) | ( n16492 & ~n16501 ) | ( n16493 & ~n16501 ) ;
  assign n16503 = ( ~n16498 & n16499 ) | ( ~n16498 & n16502 ) | ( n16499 & n16502 ) ;
  assign n16504 = ~n16498 & n16503 ;
  assign n16505 = n16492 ^ x781 ^ 1'b0 ;
  assign n16506 = ( n16492 & n16504 ) | ( n16492 & n16505 ) | ( n16504 & n16505 ) ;
  assign n16507 = x619 & ~n16506 ;
  assign n16508 = ( ~n16465 & n16506 ) | ( ~n16465 & n16507 ) | ( n16506 & n16507 ) ;
  assign n16509 = ( x648 & n16423 ) | ( x648 & ~n16508 ) | ( n16423 & ~n16508 ) ;
  assign n16510 = n16508 | n16509 ;
  assign n16511 = x619 | n16450 ;
  assign n16512 = ( x1159 & n16507 ) | ( x1159 & n16511 ) | ( n16507 & n16511 ) ;
  assign n16513 = ~n16507 & n16512 ;
  assign n16514 = ( x648 & n16426 ) | ( x648 & ~n16513 ) | ( n16426 & ~n16513 ) ;
  assign n16515 = ~n16426 & n16514 ;
  assign n16516 = x789 & ~n16515 ;
  assign n16517 = n16510 & n16516 ;
  assign n16518 = x788 & n16455 ;
  assign n16519 = n16318 | n16518 ;
  assign n16520 = ~x789 & n16506 ;
  assign n16521 = n16519 | n16520 ;
  assign n16522 = ( ~n16463 & n16517 ) | ( ~n16463 & n16521 ) | ( n16517 & n16521 ) ;
  assign n16523 = ~n16463 & n16522 ;
  assign n16524 = x628 & ~n16523 ;
  assign n16525 = n16429 ^ x788 ^ 1'b0 ;
  assign n16526 = ( n16429 & n16436 ) | ( n16429 & n16525 ) | ( n16436 & n16525 ) ;
  assign n16527 = x628 | n16526 ;
  assign n16528 = ( x1156 & n16524 ) | ( x1156 & n16527 ) | ( n16524 & n16527 ) ;
  assign n16529 = ~n16524 & n16528 ;
  assign n16530 = n1611 & n16318 ;
  assign n16531 = n16452 | n16530 ;
  assign n16532 = x628 & n1611 ;
  assign n16533 = n16531 | n16532 ;
  assign n16534 = ~x1156 & n16533 ;
  assign n16535 = ( x629 & n16529 ) | ( x629 & ~n16534 ) | ( n16529 & ~n16534 ) ;
  assign n16536 = ~n16529 & n16535 ;
  assign n16537 = ~x628 & n1611 ;
  assign n16538 = n16531 | n16537 ;
  assign n16539 = x1156 & n16538 ;
  assign n16540 = x629 | n16539 ;
  assign n16541 = x628 & ~n16526 ;
  assign n16542 = x1156 | n16541 ;
  assign n16543 = ( n16523 & n16524 ) | ( n16523 & ~n16542 ) | ( n16524 & ~n16542 ) ;
  assign n16544 = ( ~n16536 & n16540 ) | ( ~n16536 & n16543 ) | ( n16540 & n16543 ) ;
  assign n16545 = ~n16536 & n16544 ;
  assign n16546 = n16523 ^ x792 ^ 1'b0 ;
  assign n16547 = ( n16523 & n16545 ) | ( n16523 & n16546 ) | ( n16545 & n16546 ) ;
  assign n16548 = x647 & ~n16547 ;
  assign n16549 = n16398 ^ n16339 ^ 1'b0 ;
  assign n16550 = ( n16398 & n16526 ) | ( n16398 & ~n16549 ) | ( n16526 & ~n16549 ) ;
  assign n16551 = x647 | n16550 ;
  assign n16552 = ( x1157 & n16548 ) | ( x1157 & n16551 ) | ( n16548 & n16551 ) ;
  assign n16553 = ~n16548 & n16552 ;
  assign n16554 = x647 & ~n16398 ;
  assign n16555 = x1157 | n16554 ;
  assign n16556 = ~x628 & x1156 ;
  assign n16557 = x628 & ~x1156 ;
  assign n16558 = n16556 | n16557 ;
  assign n16559 = x792 & n16558 ;
  assign n16560 = n1611 & n16559 ;
  assign n16561 = n16531 | n16560 ;
  assign n16562 = x647 & ~n16561 ;
  assign n16563 = ( ~n16555 & n16561 ) | ( ~n16555 & n16562 ) | ( n16561 & n16562 ) ;
  assign n16564 = ( x630 & n16553 ) | ( x630 & ~n16563 ) | ( n16553 & ~n16563 ) ;
  assign n16565 = ~n16553 & n16564 ;
  assign n16566 = x647 | n16398 ;
  assign n16567 = ( x1157 & n16562 ) | ( x1157 & n16566 ) | ( n16562 & n16566 ) ;
  assign n16568 = ~n16562 & n16567 ;
  assign n16569 = x630 | n16568 ;
  assign n16570 = x647 & ~n16550 ;
  assign n16571 = x1157 | n16570 ;
  assign n16572 = ( n16547 & n16548 ) | ( n16547 & ~n16571 ) | ( n16548 & ~n16571 ) ;
  assign n16573 = ( ~n16565 & n16569 ) | ( ~n16565 & n16572 ) | ( n16569 & n16572 ) ;
  assign n16574 = ~n16565 & n16573 ;
  assign n16575 = n16547 ^ x787 ^ 1'b0 ;
  assign n16576 = ( n16547 & n16574 ) | ( n16547 & n16575 ) | ( n16574 & n16575 ) ;
  assign n16577 = x644 & ~n16576 ;
  assign n16578 = n16563 | n16568 ;
  assign n16579 = n16561 ^ x787 ^ 1'b0 ;
  assign n16580 = ( n16561 & n16578 ) | ( n16561 & n16579 ) | ( n16578 & n16579 ) ;
  assign n16581 = x644 | n16580 ;
  assign n16582 = ( x715 & n16577 ) | ( x715 & n16581 ) | ( n16577 & n16581 ) ;
  assign n16583 = ~n16577 & n16582 ;
  assign n16584 = n16398 ^ n16376 ^ 1'b0 ;
  assign n16585 = ( n16398 & n16550 ) | ( n16398 & ~n16584 ) | ( n16550 & ~n16584 ) ;
  assign n16586 = x644 & ~n16585 ;
  assign n16587 = x644 | n16398 ;
  assign n16588 = ( x715 & ~n16586 ) | ( x715 & n16587 ) | ( ~n16586 & n16587 ) ;
  assign n16589 = ~x715 & n16588 ;
  assign n16590 = ( x1160 & n16583 ) | ( x1160 & ~n16589 ) | ( n16583 & ~n16589 ) ;
  assign n16591 = ~n16583 & n16590 ;
  assign n16592 = x644 & ~n16398 ;
  assign n16593 = x644 | n16585 ;
  assign n16594 = ( x715 & n16592 ) | ( x715 & n16593 ) | ( n16592 & n16593 ) ;
  assign n16595 = ~n16592 & n16594 ;
  assign n16596 = x644 & ~n16580 ;
  assign n16597 = x715 | n16596 ;
  assign n16598 = ( n16576 & n16577 ) | ( n16576 & ~n16597 ) | ( n16577 & ~n16597 ) ;
  assign n16599 = ( x1160 & ~n16595 ) | ( x1160 & n16598 ) | ( ~n16595 & n16598 ) ;
  assign n16600 = n16595 | n16599 ;
  assign n16601 = x790 & ~n16600 ;
  assign n16602 = ( x790 & n16591 ) | ( x790 & n16601 ) | ( n16591 & n16601 ) ;
  assign n16603 = x790 | n16576 ;
  assign n16604 = ( x832 & n16602 ) | ( x832 & n16603 ) | ( n16602 & n16603 ) ;
  assign n16605 = ~n16602 & n16604 ;
  assign n16606 = ~x140 & n7318 ;
  assign n16607 = x832 | n16606 ;
  assign n16608 = ~n16605 & n16607 ;
  assign n16609 = ( n16396 & n16605 ) | ( n16396 & ~n16608 ) | ( n16605 & ~n16608 ) ;
  assign n16611 = x141 | n15644 ;
  assign n16612 = x749 & n15646 ;
  assign n16613 = n16611 & ~n16612 ;
  assign n16658 = ~x39 & n16068 ;
  assign n16659 = x38 & ~n16658 ;
  assign n16660 = n16613 & n16659 ;
  assign n16624 = x141 | x749 ;
  assign n16661 = ( x749 & n15795 ) | ( x749 & n16624 ) | ( n15795 & n16624 ) ;
  assign n16662 = ( x141 & n15876 ) | ( x141 & ~n16661 ) | ( n15876 & ~n16661 ) ;
  assign n16663 = ~n16661 & n16662 ;
  assign n16664 = x141 | n16003 ;
  assign n16665 = x141 & n15943 ;
  assign n16666 = x749 & ~n16665 ;
  assign n16667 = n16664 & n16666 ;
  assign n16668 = ( x39 & n16663 ) | ( x39 & ~n16667 ) | ( n16663 & ~n16667 ) ;
  assign n16669 = ~n16663 & n16668 ;
  assign n16670 = x141 & n16054 ;
  assign n16671 = x141 | n16048 ;
  assign n16672 = ( x749 & n16670 ) | ( x749 & n16671 ) | ( n16670 & n16671 ) ;
  assign n16673 = ~n16670 & n16672 ;
  assign n16674 = x141 | n16044 ;
  assign n16675 = x141 & n16029 ;
  assign n16676 = ( x749 & n16674 ) | ( x749 & ~n16675 ) | ( n16674 & ~n16675 ) ;
  assign n16677 = ~x749 & n16676 ;
  assign n16678 = ( x39 & ~n16673 ) | ( x39 & n16677 ) | ( ~n16673 & n16677 ) ;
  assign n16679 = n16673 | n16678 ;
  assign n16680 = ( x38 & ~n16669 ) | ( x38 & n16679 ) | ( ~n16669 & n16679 ) ;
  assign n16681 = ~x38 & n16680 ;
  assign n16682 = ( x706 & n16660 ) | ( x706 & ~n16681 ) | ( n16660 & ~n16681 ) ;
  assign n16683 = ~n16660 & n16682 ;
  assign n16614 = x38 & ~n16613 ;
  assign n16615 = x141 & ~n15631 ;
  assign n16616 = ~x749 & n15486 ;
  assign n16617 = ( x39 & n16615 ) | ( x39 & n16616 ) | ( n16615 & n16616 ) ;
  assign n16618 = n16616 ^ n16615 ^ 1'b0 ;
  assign n16619 = ( x39 & n16617 ) | ( x39 & n16618 ) | ( n16617 & n16618 ) ;
  assign n16620 = x141 & ~n15639 ;
  assign n16621 = ~x141 & n15587 ;
  assign n16622 = ( x749 & n16620 ) | ( x749 & ~n16621 ) | ( n16620 & ~n16621 ) ;
  assign n16623 = ~n16620 & n16622 ;
  assign n16625 = n15487 | n16624 ;
  assign n16626 = n16625 ^ n16623 ^ 1'b0 ;
  assign n16627 = ( n16623 & n16625 ) | ( n16623 & n16626 ) | ( n16625 & n16626 ) ;
  assign n16628 = ( x38 & ~n16623 ) | ( x38 & n16627 ) | ( ~n16623 & n16627 ) ;
  assign n16629 = ( ~n16614 & n16619 ) | ( ~n16614 & n16628 ) | ( n16619 & n16628 ) ;
  assign n16630 = ~n16614 & n16629 ;
  assign n16684 = x706 | n16630 ;
  assign n16685 = ( n2069 & ~n16683 ) | ( n2069 & n16684 ) | ( ~n16683 & n16684 ) ;
  assign n16686 = ~n2069 & n16685 ;
  assign n16687 = n16686 ^ x141 ^ 1'b0 ;
  assign n16688 = ( ~x141 & n2069 ) | ( ~x141 & n16687 ) | ( n2069 & n16687 ) ;
  assign n16689 = ( x141 & n16686 ) | ( x141 & n16688 ) | ( n16686 & n16688 ) ;
  assign n16690 = x625 & ~n16689 ;
  assign n16610 = x141 & n2069 ;
  assign n16631 = ~n2069 & n16630 ;
  assign n16632 = n16610 | n16631 ;
  assign n16691 = x625 | n16632 ;
  assign n16692 = ( x1153 & n16690 ) | ( x1153 & n16691 ) | ( n16690 & n16691 ) ;
  assign n16693 = ~n16690 & n16692 ;
  assign n16633 = x141 | n15656 ;
  assign n16694 = x625 & ~n16633 ;
  assign n16695 = x1153 | n16694 ;
  assign n16698 = n16053 ^ x39 ^ 1'b0 ;
  assign n16699 = ( n16053 & n16178 ) | ( n16053 & n16698 ) | ( n16178 & n16698 ) ;
  assign n16700 = x38 | n16699 ;
  assign n16701 = ( x38 & x141 ) | ( x38 & n16700 ) | ( x141 & n16700 ) ;
  assign n16696 = n16041 ^ x39 ^ 1'b0 ;
  assign n16697 = ( n16041 & n16141 ) | ( n16041 & n16696 ) | ( n16141 & n16696 ) ;
  assign n16702 = ( x141 & n16697 ) | ( x141 & ~n16701 ) | ( n16697 & ~n16701 ) ;
  assign n16703 = ~n16701 & n16702 ;
  assign n16704 = n16185 & n16611 ;
  assign n16705 = ( x706 & n16703 ) | ( x706 & ~n16704 ) | ( n16703 & ~n16704 ) ;
  assign n16706 = ~n16703 & n16705 ;
  assign n16707 = x141 | x706 ;
  assign n16708 = ( ~n2069 & n15656 ) | ( ~n2069 & n16707 ) | ( n15656 & n16707 ) ;
  assign n16709 = n16708 ^ n16706 ^ 1'b0 ;
  assign n16710 = ( n16706 & n16708 ) | ( n16706 & n16709 ) | ( n16708 & n16709 ) ;
  assign n16711 = ( n16610 & ~n16706 ) | ( n16610 & n16710 ) | ( ~n16706 & n16710 ) ;
  assign n16712 = ( x625 & ~n16695 ) | ( x625 & n16711 ) | ( ~n16695 & n16711 ) ;
  assign n16713 = ~n16695 & n16712 ;
  assign n16714 = ( x608 & n16693 ) | ( x608 & ~n16713 ) | ( n16693 & ~n16713 ) ;
  assign n16715 = ~n16693 & n16714 ;
  assign n16716 = x625 & ~n16711 ;
  assign n16717 = x625 | n16633 ;
  assign n16718 = ( x1153 & n16716 ) | ( x1153 & n16717 ) | ( n16716 & n16717 ) ;
  assign n16719 = ~n16716 & n16718 ;
  assign n16720 = x608 | n16719 ;
  assign n16721 = x625 & ~n16632 ;
  assign n16722 = x1153 | n16721 ;
  assign n16723 = ( n16689 & n16690 ) | ( n16689 & ~n16722 ) | ( n16690 & ~n16722 ) ;
  assign n16724 = ( ~n16715 & n16720 ) | ( ~n16715 & n16723 ) | ( n16720 & n16723 ) ;
  assign n16725 = ~n16715 & n16724 ;
  assign n16726 = n16689 ^ x778 ^ 1'b0 ;
  assign n16727 = ( n16689 & n16725 ) | ( n16689 & n16726 ) | ( n16725 & n16726 ) ;
  assign n16728 = x609 & ~n16727 ;
  assign n16729 = n16713 | n16719 ;
  assign n16730 = n16711 ^ x778 ^ 1'b0 ;
  assign n16731 = ( n16711 & n16729 ) | ( n16711 & n16730 ) | ( n16729 & n16730 ) ;
  assign n16732 = x609 | n16731 ;
  assign n16733 = ( x1155 & n16728 ) | ( x1155 & n16732 ) | ( n16728 & n16732 ) ;
  assign n16734 = ~n16728 & n16733 ;
  assign n16636 = ~n15668 & n16633 ;
  assign n16637 = ( n15668 & n16610 ) | ( n15668 & n16631 ) | ( n16610 & n16631 ) ;
  assign n16638 = n16636 | n16637 ;
  assign n16634 = n16632 ^ n15659 ^ 1'b0 ;
  assign n16635 = ( n16632 & n16633 ) | ( n16632 & n16634 ) | ( n16633 & n16634 ) ;
  assign n16640 = n16638 ^ n16635 ^ n16633 ;
  assign n16735 = ~x1155 & n16640 ;
  assign n16736 = ( x660 & n16734 ) | ( x660 & ~n16735 ) | ( n16734 & ~n16735 ) ;
  assign n16737 = ~n16734 & n16736 ;
  assign n16738 = x1155 & n16638 ;
  assign n16739 = x660 | n16738 ;
  assign n16740 = x609 & ~n16731 ;
  assign n16741 = x1155 | n16740 ;
  assign n16742 = ( n16727 & n16728 ) | ( n16727 & ~n16741 ) | ( n16728 & ~n16741 ) ;
  assign n16743 = ( ~n16737 & n16739 ) | ( ~n16737 & n16742 ) | ( n16739 & n16742 ) ;
  assign n16744 = ~n16737 & n16743 ;
  assign n16745 = n16727 ^ x785 ^ 1'b0 ;
  assign n16746 = ( n16727 & n16744 ) | ( n16727 & n16745 ) | ( n16744 & n16745 ) ;
  assign n16747 = x618 & ~n16746 ;
  assign n16748 = n16633 ^ n16234 ^ 1'b0 ;
  assign n16749 = ( n16633 & n16731 ) | ( n16633 & ~n16748 ) | ( n16731 & ~n16748 ) ;
  assign n16750 = x618 | n16749 ;
  assign n16751 = ( x1154 & n16747 ) | ( x1154 & n16750 ) | ( n16747 & n16750 ) ;
  assign n16752 = ~n16747 & n16751 ;
  assign n16639 = n16638 ^ x1155 ^ 1'b0 ;
  assign n16641 = ( n16638 & ~n16639 ) | ( n16638 & n16640 ) | ( ~n16639 & n16640 ) ;
  assign n16642 = n16635 ^ x785 ^ 1'b0 ;
  assign n16643 = ( n16635 & n16641 ) | ( n16635 & n16642 ) | ( n16641 & n16642 ) ;
  assign n16644 = x618 & ~n16643 ;
  assign n16648 = x618 & ~n16633 ;
  assign n16649 = x1154 | n16648 ;
  assign n16650 = ( n16643 & n16644 ) | ( n16643 & ~n16649 ) | ( n16644 & ~n16649 ) ;
  assign n16753 = ( x627 & ~n16650 ) | ( x627 & n16752 ) | ( ~n16650 & n16752 ) ;
  assign n16754 = ~n16752 & n16753 ;
  assign n16645 = x618 | n16633 ;
  assign n16646 = ( x1154 & n16644 ) | ( x1154 & n16645 ) | ( n16644 & n16645 ) ;
  assign n16647 = ~n16644 & n16646 ;
  assign n16755 = x627 | n16647 ;
  assign n16756 = x618 & ~n16749 ;
  assign n16757 = x1154 | n16756 ;
  assign n16758 = ( n16746 & n16747 ) | ( n16746 & ~n16757 ) | ( n16747 & ~n16757 ) ;
  assign n16759 = ( ~n16754 & n16755 ) | ( ~n16754 & n16758 ) | ( n16755 & n16758 ) ;
  assign n16760 = ~n16754 & n16759 ;
  assign n16761 = n16746 ^ x781 ^ 1'b0 ;
  assign n16762 = ( n16746 & n16760 ) | ( n16746 & n16761 ) | ( n16760 & n16761 ) ;
  assign n16763 = x619 & ~n16762 ;
  assign n16764 = n16633 ^ n16254 ^ 1'b0 ;
  assign n16765 = ( n16633 & n16749 ) | ( n16633 & ~n16764 ) | ( n16749 & ~n16764 ) ;
  assign n16771 = x619 | n16765 ;
  assign n16772 = ( x1159 & n16763 ) | ( x1159 & n16771 ) | ( n16763 & n16771 ) ;
  assign n16773 = ~n16763 & n16772 ;
  assign n16651 = n16647 | n16650 ;
  assign n16652 = n16643 ^ x781 ^ 1'b0 ;
  assign n16653 = ( n16643 & n16651 ) | ( n16643 & n16652 ) | ( n16651 & n16652 ) ;
  assign n16654 = x619 & ~n16653 ;
  assign n16774 = x619 & ~n16633 ;
  assign n16775 = x1159 | n16774 ;
  assign n16776 = ( n16653 & n16654 ) | ( n16653 & ~n16775 ) | ( n16654 & ~n16775 ) ;
  assign n16777 = ( x648 & n16773 ) | ( x648 & ~n16776 ) | ( n16773 & ~n16776 ) ;
  assign n16778 = ~n16773 & n16777 ;
  assign n16655 = x619 | n16633 ;
  assign n16656 = ( x1159 & n16654 ) | ( x1159 & n16655 ) | ( n16654 & n16655 ) ;
  assign n16657 = ~n16654 & n16656 ;
  assign n16766 = x619 & ~n16765 ;
  assign n16767 = x1159 | n16766 ;
  assign n16768 = ( n16762 & n16763 ) | ( n16762 & ~n16767 ) | ( n16763 & ~n16767 ) ;
  assign n16769 = ( x648 & ~n16657 ) | ( x648 & n16768 ) | ( ~n16657 & n16768 ) ;
  assign n16770 = n16657 | n16769 ;
  assign n16779 = n16778 ^ n16770 ^ 1'b0 ;
  assign n16780 = ( x789 & ~n16770 ) | ( x789 & n16778 ) | ( ~n16770 & n16778 ) ;
  assign n16781 = ( x789 & ~n16779 ) | ( x789 & n16780 ) | ( ~n16779 & n16780 ) ;
  assign n16782 = ( x789 & n16762 ) | ( x789 & ~n16781 ) | ( n16762 & ~n16781 ) ;
  assign n16783 = ~n16781 & n16782 ;
  assign n16784 = ~x626 & n16783 ;
  assign n16785 = n16633 ^ n16279 ^ 1'b0 ;
  assign n16786 = ( n16633 & n16765 ) | ( n16633 & ~n16785 ) | ( n16765 & ~n16785 ) ;
  assign n16787 = x626 & n16786 ;
  assign n16788 = ( x641 & ~n16784 ) | ( x641 & n16787 ) | ( ~n16784 & n16787 ) ;
  assign n16789 = n16784 | n16788 ;
  assign n16790 = ~x626 & n16786 ;
  assign n16791 = x626 & n16783 ;
  assign n16792 = ( x641 & n16790 ) | ( x641 & ~n16791 ) | ( n16790 & ~n16791 ) ;
  assign n16793 = ~n16790 & n16792 ;
  assign n16794 = n16657 | n16776 ;
  assign n16795 = n16653 ^ x789 ^ 1'b0 ;
  assign n16796 = ( n16653 & n16794 ) | ( n16653 & n16795 ) | ( n16794 & n16795 ) ;
  assign n16797 = x626 & ~n16796 ;
  assign n16798 = x626 | n16633 ;
  assign n16799 = ( x1158 & n16797 ) | ( x1158 & n16798 ) | ( n16797 & n16798 ) ;
  assign n16800 = ~n16797 & n16799 ;
  assign n16801 = n16289 | n16800 ;
  assign n16802 = ~n16793 & n16801 ;
  assign n16803 = x626 & ~n16633 ;
  assign n16804 = x1158 | n16803 ;
  assign n16805 = ( n16796 & n16797 ) | ( n16796 & ~n16804 ) | ( n16797 & ~n16804 ) ;
  assign n16806 = n16299 & ~n16805 ;
  assign n16807 = ~n16802 & n16806 ;
  assign n16808 = ( n16789 & n16802 ) | ( n16789 & ~n16807 ) | ( n16802 & ~n16807 ) ;
  assign n16809 = n16783 ^ x788 ^ 1'b0 ;
  assign n16810 = ( n16783 & n16808 ) | ( n16783 & n16809 ) | ( n16808 & n16809 ) ;
  assign n16811 = x628 & ~n16810 ;
  assign n16812 = n16800 | n16805 ;
  assign n16813 = n16796 ^ x788 ^ 1'b0 ;
  assign n16814 = ( n16796 & n16812 ) | ( n16796 & n16813 ) | ( n16812 & n16813 ) ;
  assign n16815 = x628 | n16814 ;
  assign n16816 = ( x1156 & n16811 ) | ( x1156 & n16815 ) | ( n16811 & n16815 ) ;
  assign n16817 = ~n16811 & n16816 ;
  assign n16818 = x628 & ~n16633 ;
  assign n16819 = x1156 | n16818 ;
  assign n16820 = n16633 ^ n16318 ^ 1'b0 ;
  assign n16821 = ( n16633 & n16786 ) | ( n16633 & ~n16820 ) | ( n16786 & ~n16820 ) ;
  assign n16822 = x628 & ~n16821 ;
  assign n16823 = ( ~n16819 & n16821 ) | ( ~n16819 & n16822 ) | ( n16821 & n16822 ) ;
  assign n16824 = ( x629 & n16817 ) | ( x629 & ~n16823 ) | ( n16817 & ~n16823 ) ;
  assign n16825 = ~n16817 & n16824 ;
  assign n16826 = x628 | n16633 ;
  assign n16827 = ( x1156 & n16822 ) | ( x1156 & n16826 ) | ( n16822 & n16826 ) ;
  assign n16828 = ~n16822 & n16827 ;
  assign n16829 = x629 | n16828 ;
  assign n16830 = x628 & ~n16814 ;
  assign n16831 = x1156 | n16830 ;
  assign n16832 = ( n16810 & n16811 ) | ( n16810 & ~n16831 ) | ( n16811 & ~n16831 ) ;
  assign n16833 = ( ~n16825 & n16829 ) | ( ~n16825 & n16832 ) | ( n16829 & n16832 ) ;
  assign n16834 = ~n16825 & n16833 ;
  assign n16835 = n16810 ^ x792 ^ 1'b0 ;
  assign n16836 = ( n16810 & n16834 ) | ( n16810 & n16835 ) | ( n16834 & n16835 ) ;
  assign n16837 = x647 & ~n16836 ;
  assign n16838 = n16633 ^ n16339 ^ 1'b0 ;
  assign n16839 = ( n16633 & n16814 ) | ( n16633 & ~n16838 ) | ( n16814 & ~n16838 ) ;
  assign n16840 = x647 | n16839 ;
  assign n16841 = ( x1157 & n16837 ) | ( x1157 & n16840 ) | ( n16837 & n16840 ) ;
  assign n16842 = ~n16837 & n16841 ;
  assign n16843 = x647 & ~n16633 ;
  assign n16844 = x1157 | n16843 ;
  assign n16845 = n16823 | n16828 ;
  assign n16846 = n16821 ^ x792 ^ 1'b0 ;
  assign n16847 = ( n16821 & n16845 ) | ( n16821 & n16846 ) | ( n16845 & n16846 ) ;
  assign n16848 = x647 & ~n16847 ;
  assign n16849 = ( ~n16844 & n16847 ) | ( ~n16844 & n16848 ) | ( n16847 & n16848 ) ;
  assign n16850 = ( x630 & n16842 ) | ( x630 & ~n16849 ) | ( n16842 & ~n16849 ) ;
  assign n16851 = ~n16842 & n16850 ;
  assign n16852 = x647 | n16633 ;
  assign n16853 = ( x1157 & n16848 ) | ( x1157 & n16852 ) | ( n16848 & n16852 ) ;
  assign n16854 = ~n16848 & n16853 ;
  assign n16855 = x630 | n16854 ;
  assign n16856 = x647 & ~n16839 ;
  assign n16857 = x1157 | n16856 ;
  assign n16858 = ( n16836 & n16837 ) | ( n16836 & ~n16857 ) | ( n16837 & ~n16857 ) ;
  assign n16859 = ( ~n16851 & n16855 ) | ( ~n16851 & n16858 ) | ( n16855 & n16858 ) ;
  assign n16860 = ~n16851 & n16859 ;
  assign n16861 = n16836 ^ x787 ^ 1'b0 ;
  assign n16862 = ( n16836 & n16860 ) | ( n16836 & n16861 ) | ( n16860 & n16861 ) ;
  assign n16863 = x644 & ~n16862 ;
  assign n16864 = n16849 | n16854 ;
  assign n16865 = n16847 ^ x787 ^ 1'b0 ;
  assign n16866 = ( n16847 & n16864 ) | ( n16847 & n16865 ) | ( n16864 & n16865 ) ;
  assign n16867 = x644 | n16866 ;
  assign n16868 = ( x715 & n16863 ) | ( x715 & n16867 ) | ( n16863 & n16867 ) ;
  assign n16869 = ~n16863 & n16868 ;
  assign n16870 = x644 | n16633 ;
  assign n16871 = n16633 ^ n16376 ^ 1'b0 ;
  assign n16872 = ( n16633 & n16839 ) | ( n16633 & ~n16871 ) | ( n16839 & ~n16871 ) ;
  assign n16873 = x644 & ~n16872 ;
  assign n16874 = ( x715 & n16870 ) | ( x715 & ~n16873 ) | ( n16870 & ~n16873 ) ;
  assign n16875 = ~x715 & n16874 ;
  assign n16876 = ( x1160 & n16869 ) | ( x1160 & ~n16875 ) | ( n16869 & ~n16875 ) ;
  assign n16877 = ~n16869 & n16876 ;
  assign n16878 = x644 & ~n16633 ;
  assign n16879 = x715 & ~n16878 ;
  assign n16880 = ( n16872 & n16873 ) | ( n16872 & n16879 ) | ( n16873 & n16879 ) ;
  assign n16881 = x644 & ~n16866 ;
  assign n16882 = x715 | n16881 ;
  assign n16883 = ( n16862 & n16863 ) | ( n16862 & ~n16882 ) | ( n16863 & ~n16882 ) ;
  assign n16884 = ( x1160 & ~n16880 ) | ( x1160 & n16883 ) | ( ~n16880 & n16883 ) ;
  assign n16885 = n16880 | n16884 ;
  assign n16886 = ( x790 & n16877 ) | ( x790 & n16885 ) | ( n16877 & n16885 ) ;
  assign n16887 = ~n16877 & n16886 ;
  assign n16888 = ~x790 & n16862 ;
  assign n16889 = ( n7318 & ~n16887 ) | ( n7318 & n16888 ) | ( ~n16887 & n16888 ) ;
  assign n16890 = n16887 | n16889 ;
  assign n16891 = x141 | n1611 ;
  assign n16892 = x749 & n15591 ;
  assign n16893 = n16891 & ~n16892 ;
  assign n16894 = n16397 | n16893 ;
  assign n16895 = n16402 | n16893 ;
  assign n16896 = x1155 & n16895 ;
  assign n16897 = n16405 | n16894 ;
  assign n16898 = ~x1155 & n16897 ;
  assign n16899 = n16896 | n16898 ;
  assign n16900 = n16894 ^ x785 ^ 1'b0 ;
  assign n16901 = ( n16894 & n16899 ) | ( n16894 & n16900 ) | ( n16899 & n16900 ) ;
  assign n16902 = n16411 | n16901 ;
  assign n16903 = x1154 & n16902 ;
  assign n16904 = n16414 | n16901 ;
  assign n16905 = ~x1154 & n16904 ;
  assign n16906 = n16903 | n16905 ;
  assign n16907 = n16901 ^ x781 ^ 1'b0 ;
  assign n16908 = ( n16901 & n16906 ) | ( n16901 & n16907 ) | ( n16906 & n16907 ) ;
  assign n16909 = x619 & ~n16908 ;
  assign n16910 = x619 | n16891 ;
  assign n16911 = ( x1159 & n16909 ) | ( x1159 & n16910 ) | ( n16909 & n16910 ) ;
  assign n16912 = ~n16909 & n16911 ;
  assign n16913 = x619 & ~n16891 ;
  assign n16914 = x1159 | n16913 ;
  assign n16915 = ( n16908 & n16909 ) | ( n16908 & ~n16914 ) | ( n16909 & ~n16914 ) ;
  assign n16916 = n16912 | n16915 ;
  assign n16917 = n16908 ^ x789 ^ 1'b0 ;
  assign n16918 = ( n16908 & n16916 ) | ( n16908 & n16917 ) | ( n16916 & n16917 ) ;
  assign n16919 = x626 & ~n16918 ;
  assign n16920 = x626 & ~n16891 ;
  assign n16921 = x1158 | n16920 ;
  assign n16922 = ( n16918 & n16919 ) | ( n16918 & ~n16921 ) | ( n16919 & ~n16921 ) ;
  assign n16923 = n16919 & ~n16922 ;
  assign n16924 = ( x1158 & n16891 ) | ( x1158 & n16920 ) | ( n16891 & n16920 ) ;
  assign n16925 = ( n16922 & ~n16923 ) | ( n16922 & n16924 ) | ( ~n16923 & n16924 ) ;
  assign n16926 = n16317 & ~n16925 ;
  assign n16927 = x706 & n15778 ;
  assign n16928 = n16891 & ~n16927 ;
  assign n16929 = ~x625 & n16927 ;
  assign n16930 = ~x1153 & n16891 ;
  assign n16931 = ~n16929 & n16930 ;
  assign n16932 = ( x1153 & n16928 ) | ( x1153 & n16929 ) | ( n16928 & n16929 ) ;
  assign n16933 = n16931 | n16932 ;
  assign n16934 = n16928 ^ x778 ^ 1'b0 ;
  assign n16935 = ( n16928 & n16933 ) | ( n16928 & n16934 ) | ( n16933 & n16934 ) ;
  assign n16936 = n16447 | n16935 ;
  assign n16937 = n16449 | n16936 ;
  assign n16938 = n16451 | n16937 ;
  assign n16939 = n16459 & ~n16938 ;
  assign n16940 = ( x788 & n16926 ) | ( x788 & n16939 ) | ( n16926 & n16939 ) ;
  assign n16941 = n16939 ^ n16926 ^ 1'b0 ;
  assign n16942 = ( x788 & n16940 ) | ( x788 & n16941 ) | ( n16940 & n16941 ) ;
  assign n16943 = x619 & ~n16937 ;
  assign n16944 = x1159 | n16943 ;
  assign n16945 = n15524 | n16928 ;
  assign n16946 = n16893 & n16945 ;
  assign n16947 = x625 & ~n16945 ;
  assign n16948 = x1153 & n16893 ;
  assign n16949 = ~n16947 & n16948 ;
  assign n16950 = ( x608 & n16931 ) | ( x608 & ~n16949 ) | ( n16931 & ~n16949 ) ;
  assign n16951 = ~n16931 & n16950 ;
  assign n16952 = x608 | n16932 ;
  assign n16953 = ( n16930 & n16946 ) | ( n16930 & n16947 ) | ( n16946 & n16947 ) ;
  assign n16954 = ( ~n16951 & n16952 ) | ( ~n16951 & n16953 ) | ( n16952 & n16953 ) ;
  assign n16955 = ~n16951 & n16954 ;
  assign n16956 = n16946 ^ x778 ^ 1'b0 ;
  assign n16957 = ( n16946 & n16955 ) | ( n16946 & n16956 ) | ( n16955 & n16956 ) ;
  assign n16958 = x609 & ~n16957 ;
  assign n16959 = x609 | n16935 ;
  assign n16960 = ( x1155 & n16958 ) | ( x1155 & n16959 ) | ( n16958 & n16959 ) ;
  assign n16961 = ~n16958 & n16960 ;
  assign n16962 = ( x660 & n16898 ) | ( x660 & ~n16961 ) | ( n16898 & ~n16961 ) ;
  assign n16963 = ~n16898 & n16962 ;
  assign n16964 = x660 | n16896 ;
  assign n16965 = x609 & ~n16935 ;
  assign n16966 = x1155 | n16965 ;
  assign n16967 = ( n16957 & n16958 ) | ( n16957 & ~n16966 ) | ( n16958 & ~n16966 ) ;
  assign n16968 = ( ~n16963 & n16964 ) | ( ~n16963 & n16967 ) | ( n16964 & n16967 ) ;
  assign n16969 = ~n16963 & n16968 ;
  assign n16970 = n16957 ^ x785 ^ 1'b0 ;
  assign n16971 = ( n16957 & n16969 ) | ( n16957 & n16970 ) | ( n16969 & n16970 ) ;
  assign n16972 = x618 & ~n16971 ;
  assign n16973 = x618 | n16936 ;
  assign n16974 = ( x1154 & n16972 ) | ( x1154 & n16973 ) | ( n16972 & n16973 ) ;
  assign n16975 = ~n16972 & n16974 ;
  assign n16976 = ( x627 & n16905 ) | ( x627 & ~n16975 ) | ( n16905 & ~n16975 ) ;
  assign n16977 = ~n16905 & n16976 ;
  assign n16978 = x627 | n16903 ;
  assign n16979 = x618 & ~n16936 ;
  assign n16980 = x1154 | n16979 ;
  assign n16981 = ( n16971 & n16972 ) | ( n16971 & ~n16980 ) | ( n16972 & ~n16980 ) ;
  assign n16982 = ( ~n16977 & n16978 ) | ( ~n16977 & n16981 ) | ( n16978 & n16981 ) ;
  assign n16983 = ~n16977 & n16982 ;
  assign n16984 = n16971 ^ x781 ^ 1'b0 ;
  assign n16985 = ( n16971 & n16983 ) | ( n16971 & n16984 ) | ( n16983 & n16984 ) ;
  assign n16986 = x619 & ~n16985 ;
  assign n16987 = ( ~n16944 & n16985 ) | ( ~n16944 & n16986 ) | ( n16985 & n16986 ) ;
  assign n16988 = ( x648 & n16912 ) | ( x648 & ~n16987 ) | ( n16912 & ~n16987 ) ;
  assign n16989 = n16987 | n16988 ;
  assign n16990 = x619 | n16937 ;
  assign n16991 = ( x1159 & n16986 ) | ( x1159 & n16990 ) | ( n16986 & n16990 ) ;
  assign n16992 = ~n16986 & n16991 ;
  assign n16993 = ( x648 & n16915 ) | ( x648 & ~n16992 ) | ( n16915 & ~n16992 ) ;
  assign n16994 = ~n16915 & n16993 ;
  assign n16995 = x789 & ~n16994 ;
  assign n16996 = n16989 & n16995 ;
  assign n16997 = ~x789 & n16985 ;
  assign n16998 = n16519 | n16997 ;
  assign n16999 = ( ~n16942 & n16996 ) | ( ~n16942 & n16998 ) | ( n16996 & n16998 ) ;
  assign n17000 = ~n16942 & n16999 ;
  assign n17001 = x628 & ~n17000 ;
  assign n17002 = n16918 ^ x788 ^ 1'b0 ;
  assign n17003 = ( n16918 & n16925 ) | ( n16918 & n17002 ) | ( n16925 & n17002 ) ;
  assign n17004 = x628 | n17003 ;
  assign n17005 = ( x1156 & n17001 ) | ( x1156 & n17004 ) | ( n17001 & n17004 ) ;
  assign n17006 = ~n17001 & n17005 ;
  assign n17007 = n16530 | n16938 ;
  assign n17008 = n16532 | n17007 ;
  assign n17009 = ~x1156 & n17008 ;
  assign n17010 = ( x629 & n17006 ) | ( x629 & ~n17009 ) | ( n17006 & ~n17009 ) ;
  assign n17011 = ~n17006 & n17010 ;
  assign n17012 = n16537 | n17007 ;
  assign n17013 = x1156 & n17012 ;
  assign n17014 = x629 | n17013 ;
  assign n17015 = x628 & ~n17003 ;
  assign n17016 = x1156 | n17015 ;
  assign n17017 = ( n17000 & n17001 ) | ( n17000 & ~n17016 ) | ( n17001 & ~n17016 ) ;
  assign n17018 = ( ~n17011 & n17014 ) | ( ~n17011 & n17017 ) | ( n17014 & n17017 ) ;
  assign n17019 = ~n17011 & n17018 ;
  assign n17020 = n17000 ^ x792 ^ 1'b0 ;
  assign n17021 = ( n17000 & n17019 ) | ( n17000 & n17020 ) | ( n17019 & n17020 ) ;
  assign n17022 = x647 & ~n17021 ;
  assign n17023 = n16891 ^ n16339 ^ 1'b0 ;
  assign n17024 = ( n16891 & n17003 ) | ( n16891 & ~n17023 ) | ( n17003 & ~n17023 ) ;
  assign n17025 = x647 | n17024 ;
  assign n17026 = ( x1157 & n17022 ) | ( x1157 & n17025 ) | ( n17022 & n17025 ) ;
  assign n17027 = ~n17022 & n17026 ;
  assign n17028 = x647 & ~n16891 ;
  assign n17029 = x1157 | n17028 ;
  assign n17030 = n16560 | n17007 ;
  assign n17031 = x647 & ~n17030 ;
  assign n17032 = ( ~n17029 & n17030 ) | ( ~n17029 & n17031 ) | ( n17030 & n17031 ) ;
  assign n17033 = ( x630 & n17027 ) | ( x630 & ~n17032 ) | ( n17027 & ~n17032 ) ;
  assign n17034 = ~n17027 & n17033 ;
  assign n17035 = x647 | n16891 ;
  assign n17036 = ( x1157 & n17031 ) | ( x1157 & n17035 ) | ( n17031 & n17035 ) ;
  assign n17037 = ~n17031 & n17036 ;
  assign n17038 = x630 | n17037 ;
  assign n17039 = x647 & ~n17024 ;
  assign n17040 = x1157 | n17039 ;
  assign n17041 = ( n17021 & n17022 ) | ( n17021 & ~n17040 ) | ( n17022 & ~n17040 ) ;
  assign n17042 = ( ~n17034 & n17038 ) | ( ~n17034 & n17041 ) | ( n17038 & n17041 ) ;
  assign n17043 = ~n17034 & n17042 ;
  assign n17044 = n17021 ^ x787 ^ 1'b0 ;
  assign n17045 = ( n17021 & n17043 ) | ( n17021 & n17044 ) | ( n17043 & n17044 ) ;
  assign n17046 = x644 & ~n17045 ;
  assign n17047 = n17032 | n17037 ;
  assign n17048 = n17030 ^ x787 ^ 1'b0 ;
  assign n17049 = ( n17030 & n17047 ) | ( n17030 & n17048 ) | ( n17047 & n17048 ) ;
  assign n17050 = x644 | n17049 ;
  assign n17051 = ( x715 & n17046 ) | ( x715 & n17050 ) | ( n17046 & n17050 ) ;
  assign n17052 = ~n17046 & n17051 ;
  assign n17053 = n16891 ^ n16376 ^ 1'b0 ;
  assign n17054 = ( n16891 & n17024 ) | ( n16891 & ~n17053 ) | ( n17024 & ~n17053 ) ;
  assign n17055 = x644 & ~n17054 ;
  assign n17056 = x644 | n16891 ;
  assign n17057 = ( x715 & ~n17055 ) | ( x715 & n17056 ) | ( ~n17055 & n17056 ) ;
  assign n17058 = ~x715 & n17057 ;
  assign n17059 = ( x1160 & n17052 ) | ( x1160 & ~n17058 ) | ( n17052 & ~n17058 ) ;
  assign n17060 = ~n17052 & n17059 ;
  assign n17061 = x644 & ~n16891 ;
  assign n17062 = x644 | n17054 ;
  assign n17063 = ( x715 & n17061 ) | ( x715 & n17062 ) | ( n17061 & n17062 ) ;
  assign n17064 = ~n17061 & n17063 ;
  assign n17065 = x644 & ~n17049 ;
  assign n17066 = x715 | n17065 ;
  assign n17067 = ( n17045 & n17046 ) | ( n17045 & ~n17066 ) | ( n17046 & ~n17066 ) ;
  assign n17068 = ( x1160 & ~n17064 ) | ( x1160 & n17067 ) | ( ~n17064 & n17067 ) ;
  assign n17069 = n17064 | n17068 ;
  assign n17070 = x790 & ~n17069 ;
  assign n17071 = ( x790 & n17060 ) | ( x790 & n17070 ) | ( n17060 & n17070 ) ;
  assign n17072 = x790 | n17045 ;
  assign n17073 = ( x832 & n17071 ) | ( x832 & n17072 ) | ( n17071 & n17072 ) ;
  assign n17074 = ~n17071 & n17073 ;
  assign n17075 = ~x141 & n7318 ;
  assign n17076 = x832 | n17075 ;
  assign n17077 = ~n17074 & n17076 ;
  assign n17078 = ( n16890 & n17074 ) | ( n16890 & ~n17077 ) | ( n17074 & ~n17077 ) ;
  assign n17079 = x142 & ~n1611 ;
  assign n17080 = x1157 | n17079 ;
  assign n17081 = x735 & n15778 ;
  assign n17082 = x1153 ^ x625 ^ 1'b0 ;
  assign n17083 = x778 & n17082 ;
  assign n17084 = n17081 & ~n17083 ;
  assign n17085 = n17079 | n17084 ;
  assign n17086 = n16279 | n16318 ;
  assign n17087 = n16234 | n16254 ;
  assign n17088 = n17086 | n17087 ;
  assign n17089 = n17085 & ~n17088 ;
  assign n17090 = x628 | x1156 ;
  assign n17091 = x628 & x1156 ;
  assign n17092 = x792 & ~n17091 ;
  assign n17093 = n17090 & n17092 ;
  assign n17094 = n17089 & ~n17093 ;
  assign n17095 = ~x647 & n17094 ;
  assign n17096 = n17080 | n17095 ;
  assign n17097 = x1155 & ~n17079 ;
  assign n17098 = x743 & n15591 ;
  assign n17099 = ~n15659 & n17098 ;
  assign n17100 = x609 & n17099 ;
  assign n17101 = n17097 & ~n17100 ;
  assign n17102 = x1155 | n17079 ;
  assign n17103 = ~x609 & n17099 ;
  assign n17104 = n17102 | n17103 ;
  assign n17105 = ~n17101 & n17104 ;
  assign n17106 = x785 & ~n17105 ;
  assign n17107 = x785 | n17079 ;
  assign n17108 = n17099 | n17107 ;
  assign n17109 = ~n17106 & n17108 ;
  assign n17110 = ~x618 & n17079 ;
  assign n17111 = x618 & n17109 ;
  assign n17112 = ( x1154 & n17110 ) | ( x1154 & ~n17111 ) | ( n17110 & ~n17111 ) ;
  assign n17113 = ~n17110 & n17112 ;
  assign n17114 = ~x618 & n17109 ;
  assign n17115 = x618 & n17079 ;
  assign n17116 = ( x1154 & ~n17114 ) | ( x1154 & n17115 ) | ( ~n17114 & n17115 ) ;
  assign n17117 = n17114 | n17116 ;
  assign n17118 = ~n17113 & n17117 ;
  assign n17119 = n17109 ^ x781 ^ 1'b0 ;
  assign n17120 = ( n17109 & n17118 ) | ( n17109 & n17119 ) | ( n17118 & n17119 ) ;
  assign n17121 = ~x619 & n17079 ;
  assign n17122 = x619 & n17120 ;
  assign n17123 = ( x1159 & n17121 ) | ( x1159 & ~n17122 ) | ( n17121 & ~n17122 ) ;
  assign n17124 = ~n17121 & n17123 ;
  assign n17125 = ~x619 & n17120 ;
  assign n17126 = x619 & n17079 ;
  assign n17127 = ( x1159 & ~n17125 ) | ( x1159 & n17126 ) | ( ~n17125 & n17126 ) ;
  assign n17128 = n17125 | n17127 ;
  assign n17129 = ~n17124 & n17128 ;
  assign n17130 = n17120 ^ x789 ^ 1'b0 ;
  assign n17131 = ( n17120 & n17129 ) | ( n17120 & n17130 ) | ( n17129 & n17130 ) ;
  assign n17132 = ~x626 & n17079 ;
  assign n17133 = x626 & n17131 ;
  assign n17134 = ( x1158 & n17132 ) | ( x1158 & ~n17133 ) | ( n17132 & ~n17133 ) ;
  assign n17135 = ~n17132 & n17134 ;
  assign n17136 = x626 & n17079 ;
  assign n17137 = x1158 | n17136 ;
  assign n17138 = ~x626 & n17131 ;
  assign n17139 = ( ~n17135 & n17137 ) | ( ~n17135 & n17138 ) | ( n17137 & n17138 ) ;
  assign n17140 = ~n17135 & n17139 ;
  assign n17141 = n17131 ^ x788 ^ 1'b0 ;
  assign n17142 = ( n17131 & n17140 ) | ( n17131 & n17141 ) | ( n17140 & n17141 ) ;
  assign n17143 = n17079 ^ n16339 ^ 1'b0 ;
  assign n17144 = ( n17079 & n17142 ) | ( n17079 & ~n17143 ) | ( n17142 & ~n17143 ) ;
  assign n17145 = ~x647 & n17144 ;
  assign n17146 = ~n16234 & n17085 ;
  assign n17147 = ~n16254 & n17146 ;
  assign n17148 = n17079 | n17147 ;
  assign n17149 = ~x619 & n17148 ;
  assign n17150 = n17079 | n17146 ;
  assign n17151 = ~x618 & n17150 ;
  assign n17152 = ~x609 & n17085 ;
  assign n17153 = x625 | x1153 ;
  assign n17154 = n17081 & ~n17153 ;
  assign n17155 = n17079 | n17154 ;
  assign n17156 = ~n15524 & n15778 ;
  assign n17157 = x735 & n17156 ;
  assign n17158 = x625 & n17157 ;
  assign n17159 = ( x1153 & n17098 ) | ( x1153 & n17158 ) | ( n17098 & n17158 ) ;
  assign n17160 = ( x608 & n17155 ) | ( x608 & n17159 ) | ( n17155 & n17159 ) ;
  assign n17161 = n17159 ^ n17155 ^ 1'b0 ;
  assign n17162 = ( x608 & n17160 ) | ( x608 & n17161 ) | ( n17160 & n17161 ) ;
  assign n17163 = x1153 & ~n17079 ;
  assign n17164 = x625 & n17081 ;
  assign n17165 = ( x608 & n17163 ) | ( x608 & ~n17164 ) | ( n17163 & ~n17164 ) ;
  assign n17166 = n17165 ^ n17163 ^ 1'b0 ;
  assign n17167 = ( x608 & n17165 ) | ( x608 & ~n17166 ) | ( n17165 & ~n17166 ) ;
  assign n17168 = n17157 ^ n17098 ^ n17079 ;
  assign n17169 = ~n17158 & n17168 ;
  assign n17170 = ( x1153 & ~n17167 ) | ( x1153 & n17169 ) | ( ~n17167 & n17169 ) ;
  assign n17171 = ~n17167 & n17170 ;
  assign n17172 = ( x778 & n17162 ) | ( x778 & ~n17171 ) | ( n17162 & ~n17171 ) ;
  assign n17173 = ~n17162 & n17172 ;
  assign n17174 = ( x778 & n17168 ) | ( x778 & ~n17173 ) | ( n17168 & ~n17173 ) ;
  assign n17175 = ~n17173 & n17174 ;
  assign n17176 = x609 & n17175 ;
  assign n17177 = ( x1155 & n17152 ) | ( x1155 & ~n17176 ) | ( n17152 & ~n17176 ) ;
  assign n17178 = ~n17152 & n17177 ;
  assign n17179 = ( x660 & n17104 ) | ( x660 & n17178 ) | ( n17104 & n17178 ) ;
  assign n17180 = ~n17178 & n17179 ;
  assign n17181 = ~x609 & n17175 ;
  assign n17182 = x609 & n17085 ;
  assign n17183 = ( x1155 & ~n17181 ) | ( x1155 & n17182 ) | ( ~n17181 & n17182 ) ;
  assign n17184 = n17181 | n17183 ;
  assign n17185 = ( x660 & ~n17101 ) | ( x660 & n17184 ) | ( ~n17101 & n17184 ) ;
  assign n17186 = ~x660 & n17185 ;
  assign n17187 = ( x785 & n17180 ) | ( x785 & ~n17186 ) | ( n17180 & ~n17186 ) ;
  assign n17188 = ~n17180 & n17187 ;
  assign n17189 = ( x785 & n17175 ) | ( x785 & ~n17188 ) | ( n17175 & ~n17188 ) ;
  assign n17190 = ~n17188 & n17189 ;
  assign n17191 = x618 & n17190 ;
  assign n17192 = ( x1154 & n17151 ) | ( x1154 & ~n17191 ) | ( n17151 & ~n17191 ) ;
  assign n17193 = ~n17151 & n17192 ;
  assign n17194 = ( x627 & n17117 ) | ( x627 & n17193 ) | ( n17117 & n17193 ) ;
  assign n17195 = ~n17193 & n17194 ;
  assign n17196 = ~x618 & n17190 ;
  assign n17197 = x618 & n17150 ;
  assign n17198 = ( x1154 & ~n17196 ) | ( x1154 & n17197 ) | ( ~n17196 & n17197 ) ;
  assign n17199 = n17196 | n17198 ;
  assign n17200 = ( x627 & ~n17113 ) | ( x627 & n17199 ) | ( ~n17113 & n17199 ) ;
  assign n17201 = ~x627 & n17200 ;
  assign n17202 = ( x781 & n17195 ) | ( x781 & ~n17201 ) | ( n17195 & ~n17201 ) ;
  assign n17203 = ~n17195 & n17202 ;
  assign n17204 = ( x781 & n17190 ) | ( x781 & ~n17203 ) | ( n17190 & ~n17203 ) ;
  assign n17205 = ~n17203 & n17204 ;
  assign n17206 = x619 & n17205 ;
  assign n17207 = ( x1159 & n17149 ) | ( x1159 & ~n17206 ) | ( n17149 & ~n17206 ) ;
  assign n17208 = ~n17149 & n17207 ;
  assign n17209 = ( x648 & n17128 ) | ( x648 & n17208 ) | ( n17128 & n17208 ) ;
  assign n17210 = ~n17208 & n17209 ;
  assign n17211 = ~x619 & n17205 ;
  assign n17212 = x619 & n17148 ;
  assign n17213 = ( x1159 & ~n17211 ) | ( x1159 & n17212 ) | ( ~n17211 & n17212 ) ;
  assign n17214 = n17211 | n17213 ;
  assign n17215 = ( x648 & ~n17124 ) | ( x648 & n17214 ) | ( ~n17124 & n17214 ) ;
  assign n17216 = ~x648 & n17215 ;
  assign n17217 = ( x789 & n17210 ) | ( x789 & ~n17216 ) | ( n17210 & ~n17216 ) ;
  assign n17218 = ~n17210 & n17217 ;
  assign n17219 = x789 | n17205 ;
  assign n17220 = ( n16519 & ~n17218 ) | ( n16519 & n17219 ) | ( ~n17218 & n17219 ) ;
  assign n17221 = ~n16519 & n17220 ;
  assign n17222 = n16279 & ~n17079 ;
  assign n17223 = n16459 & ~n17222 ;
  assign n17224 = n17148 & n17223 ;
  assign n17225 = n17224 ^ n16317 ^ 1'b0 ;
  assign n17226 = ( ~n16317 & n17140 ) | ( ~n16317 & n17225 ) | ( n17140 & n17225 ) ;
  assign n17227 = ( n16317 & n17224 ) | ( n16317 & n17226 ) | ( n17224 & n17226 ) ;
  assign n17228 = n17221 ^ x788 ^ 1'b0 ;
  assign n17229 = ( ~x788 & n17227 ) | ( ~x788 & n17228 ) | ( n17227 & n17228 ) ;
  assign n17230 = ( x788 & n17221 ) | ( x788 & n17229 ) | ( n17221 & n17229 ) ;
  assign n17231 = x628 & ~n17230 ;
  assign n17232 = x628 | n17142 ;
  assign n17233 = ( x1156 & n17231 ) | ( x1156 & n17232 ) | ( n17231 & n17232 ) ;
  assign n17234 = ~n17231 & n17233 ;
  assign n17235 = ~x628 & n17089 ;
  assign n17236 = ( ~x1156 & n17079 ) | ( ~x1156 & n17235 ) | ( n17079 & n17235 ) ;
  assign n17237 = ~x1156 & n17236 ;
  assign n17238 = ( x629 & n17234 ) | ( x629 & ~n17237 ) | ( n17234 & ~n17237 ) ;
  assign n17239 = ~n17234 & n17238 ;
  assign n17240 = x1156 ^ x629 ^ 1'b0 ;
  assign n17241 = x628 & n17089 ;
  assign n17242 = n17079 | n17241 ;
  assign n17243 = ( x1156 & ~n17240 ) | ( x1156 & n17242 ) | ( ~n17240 & n17242 ) ;
  assign n17244 = ( x629 & n17240 ) | ( x629 & n17243 ) | ( n17240 & n17243 ) ;
  assign n17245 = x628 & ~n17142 ;
  assign n17246 = x1156 | n17245 ;
  assign n17247 = ( n17230 & n17231 ) | ( n17230 & ~n17246 ) | ( n17231 & ~n17246 ) ;
  assign n17248 = ( ~n17239 & n17244 ) | ( ~n17239 & n17247 ) | ( n17244 & n17247 ) ;
  assign n17249 = ~n17239 & n17248 ;
  assign n17250 = n17230 ^ x792 ^ 1'b0 ;
  assign n17251 = ( n17230 & n17249 ) | ( n17230 & n17250 ) | ( n17249 & n17250 ) ;
  assign n17252 = x647 & n17251 ;
  assign n17253 = ( x1157 & n17145 ) | ( x1157 & ~n17252 ) | ( n17145 & ~n17252 ) ;
  assign n17254 = ~n17145 & n17253 ;
  assign n17255 = x630 & ~n17254 ;
  assign n17256 = n17096 & n17255 ;
  assign n17257 = ~x647 & n17251 ;
  assign n17258 = x647 & n17144 ;
  assign n17259 = ( x1157 & ~n17257 ) | ( x1157 & n17258 ) | ( ~n17257 & n17258 ) ;
  assign n17260 = n17257 | n17259 ;
  assign n17261 = x1157 & ~n17079 ;
  assign n17262 = x647 & n17094 ;
  assign n17263 = n17261 & ~n17262 ;
  assign n17264 = ( x630 & n17260 ) | ( x630 & ~n17263 ) | ( n17260 & ~n17263 ) ;
  assign n17265 = ~x630 & n17264 ;
  assign n17266 = ( x787 & n17256 ) | ( x787 & ~n17265 ) | ( n17256 & ~n17265 ) ;
  assign n17267 = ~n17256 & n17266 ;
  assign n17268 = ( x787 & n17251 ) | ( x787 & ~n17267 ) | ( n17251 & ~n17267 ) ;
  assign n17269 = ~n17267 & n17268 ;
  assign n17270 = ~x790 & n17269 ;
  assign n17271 = ~x644 & n17269 ;
  assign n17272 = x1157 ^ x647 ^ 1'b0 ;
  assign n17273 = x787 & n17272 ;
  assign n17274 = n17094 & ~n17273 ;
  assign n17275 = n17079 | n17274 ;
  assign n17276 = x644 & n17275 ;
  assign n17277 = ( x715 & ~n17271 ) | ( x715 & n17276 ) | ( ~n17271 & n17276 ) ;
  assign n17278 = n17271 | n17277 ;
  assign n17279 = x644 & n17079 ;
  assign n17280 = n17079 ^ n16376 ^ 1'b0 ;
  assign n17281 = ( n17079 & n17144 ) | ( n17079 & ~n17280 ) | ( n17144 & ~n17280 ) ;
  assign n17282 = ~x644 & n17281 ;
  assign n17283 = ( x715 & n17279 ) | ( x715 & ~n17282 ) | ( n17279 & ~n17282 ) ;
  assign n17284 = ~n17279 & n17283 ;
  assign n17285 = ( x1160 & n17278 ) | ( x1160 & ~n17284 ) | ( n17278 & ~n17284 ) ;
  assign n17286 = ~x1160 & n17285 ;
  assign n17287 = x644 & n17281 ;
  assign n17288 = ~x644 & n17079 ;
  assign n17289 = ( x715 & ~n17287 ) | ( x715 & n17288 ) | ( ~n17287 & n17288 ) ;
  assign n17290 = n17287 | n17289 ;
  assign n17291 = ~x644 & n17275 ;
  assign n17292 = x644 & n17269 ;
  assign n17293 = ( x715 & n17291 ) | ( x715 & ~n17292 ) | ( n17291 & ~n17292 ) ;
  assign n17294 = ~n17291 & n17293 ;
  assign n17295 = x1160 & ~n17294 ;
  assign n17296 = n17290 & n17295 ;
  assign n17297 = ( x790 & n17286 ) | ( x790 & n17296 ) | ( n17286 & n17296 ) ;
  assign n17298 = n17296 ^ n17286 ^ 1'b0 ;
  assign n17299 = ( x790 & n17297 ) | ( x790 & n17298 ) | ( n17297 & n17298 ) ;
  assign n17300 = ( x832 & n17270 ) | ( x832 & ~n17299 ) | ( n17270 & ~n17299 ) ;
  assign n17301 = ~n17270 & n17300 ;
  assign n17302 = ~x142 & n5193 ;
  assign n17303 = x142 & ~n15402 ;
  assign n17304 = n5061 | n17303 ;
  assign n17305 = x215 & n17304 ;
  assign n17306 = x142 & ~n15337 ;
  assign n17307 = n2263 | n17306 ;
  assign n17308 = x142 & ~n15468 ;
  assign n17309 = x142 & ~n15433 ;
  assign n17310 = n17308 ^ n5061 ^ 1'b0 ;
  assign n17311 = ( n17308 & n17309 ) | ( n17308 & n17310 ) | ( n17309 & n17310 ) ;
  assign n17312 = ( x216 & x221 ) | ( x216 & ~n17311 ) | ( x221 & ~n17311 ) ;
  assign n17313 = ~n17311 & n17312 ;
  assign n17314 = ( x215 & n17307 ) | ( x215 & ~n17313 ) | ( n17307 & ~n17313 ) ;
  assign n17315 = ~x215 & n17314 ;
  assign n17316 = x142 & ~n15378 ;
  assign n17317 = n5061 & ~n17316 ;
  assign n17318 = ~n17315 & n17317 ;
  assign n17319 = ( n17305 & n17315 ) | ( n17305 & ~n17318 ) | ( n17315 & ~n17318 ) ;
  assign n17320 = ( ~x39 & x299 ) | ( ~x39 & n17319 ) | ( x299 & n17319 ) ;
  assign n17321 = x39 & n17320 ;
  assign n17322 = x39 & n15485 ;
  assign n17323 = x142 & ~n15487 ;
  assign n17324 = ~n17322 & n17323 ;
  assign n17325 = ( ~n15102 & n17321 ) | ( ~n15102 & n17324 ) | ( n17321 & n17324 ) ;
  assign n17326 = ~n15102 & n17325 ;
  assign n17327 = x38 & ~n15653 ;
  assign n17328 = n2069 | n17327 ;
  assign n17329 = n17326 ^ x142 ^ 1'b0 ;
  assign n17330 = ( ~x142 & n17328 ) | ( ~x142 & n17329 ) | ( n17328 & n17329 ) ;
  assign n17331 = ( x142 & n17326 ) | ( x142 & n17330 ) | ( n17326 & n17330 ) ;
  assign n17332 = ~x142 & n15886 ;
  assign n17333 = x735 & ~n17332 ;
  assign n17334 = x142 & ~n16103 ;
  assign n17335 = n17333 & ~n17334 ;
  assign n17336 = ( x735 & n17303 ) | ( x735 & ~n17335 ) | ( n17303 & ~n17335 ) ;
  assign n17337 = ~n17335 & n17336 ;
  assign n17338 = n5061 | n17337 ;
  assign n17339 = x142 & ~n16101 ;
  assign n17340 = n15880 & n17332 ;
  assign n17341 = ( x735 & n17339 ) | ( x735 & ~n17340 ) | ( n17339 & ~n17340 ) ;
  assign n17342 = ~n17339 & n17341 ;
  assign n17343 = ( x735 & n17316 ) | ( x735 & ~n17342 ) | ( n17316 & ~n17342 ) ;
  assign n17344 = ~n17342 & n17343 ;
  assign n17345 = n5061 & ~n17344 ;
  assign n17346 = x215 & ~n17345 ;
  assign n17347 = n17338 & n17346 ;
  assign n17348 = n16154 ^ x142 ^ 1'b0 ;
  assign n17349 = ( ~n16111 & n16154 ) | ( ~n16111 & n17348 ) | ( n16154 & n17348 ) ;
  assign n17350 = n17309 ^ x735 ^ 1'b0 ;
  assign n17351 = ( n17309 & n17349 ) | ( n17309 & n17350 ) | ( n17349 & n17350 ) ;
  assign n17352 = n5061 & n17351 ;
  assign n17353 = n16150 ^ x142 ^ 1'b0 ;
  assign n17354 = ( ~n16121 & n16150 ) | ( ~n16121 & n17353 ) | ( n16150 & n17353 ) ;
  assign n17355 = n17308 ^ x735 ^ 1'b0 ;
  assign n17356 = ( n17308 & n17354 ) | ( n17308 & n17355 ) | ( n17354 & n17355 ) ;
  assign n17357 = ~n5061 & n17356 ;
  assign n17358 = ( n2263 & n17352 ) | ( n2263 & ~n17357 ) | ( n17352 & ~n17357 ) ;
  assign n17359 = ~n17352 & n17358 ;
  assign n17360 = ~n15336 & n17081 ;
  assign n17361 = n17306 | n17360 ;
  assign n17362 = n2263 | n17361 ;
  assign n17363 = ( x215 & ~n17359 ) | ( x215 & n17362 ) | ( ~n17359 & n17362 ) ;
  assign n17364 = ~x215 & n17363 ;
  assign n17365 = ( x299 & n17347 ) | ( x299 & ~n17364 ) | ( n17347 & ~n17364 ) ;
  assign n17366 = ~n17347 & n17365 ;
  assign n17367 = n5114 & n17351 ;
  assign n17368 = ~n5114 & n17356 ;
  assign n17369 = ( n1359 & n17367 ) | ( n1359 & ~n17368 ) | ( n17367 & ~n17368 ) ;
  assign n17370 = ~n17367 & n17369 ;
  assign n17371 = n1359 | n17361 ;
  assign n17372 = ( x223 & ~n17370 ) | ( x223 & n17371 ) | ( ~n17370 & n17371 ) ;
  assign n17373 = ~x223 & n17372 ;
  assign n17374 = n5114 | n17337 ;
  assign n17375 = n5114 & ~n17344 ;
  assign n17376 = x223 & ~n17375 ;
  assign n17377 = n17374 & n17376 ;
  assign n17378 = ( x299 & ~n17373 ) | ( x299 & n17377 ) | ( ~n17373 & n17377 ) ;
  assign n17379 = n17373 | n17378 ;
  assign n17380 = ( x39 & n17366 ) | ( x39 & n17379 ) | ( n17366 & n17379 ) ;
  assign n17381 = ~n17366 & n17380 ;
  assign n17382 = x142 & ~x735 ;
  assign n17383 = ~n15332 & n17382 ;
  assign n17384 = x142 | n16053 ;
  assign n17385 = x142 & n16041 ;
  assign n17386 = x735 & ~n17385 ;
  assign n17387 = n17384 & n17386 ;
  assign n17388 = ( ~x39 & n17383 ) | ( ~x39 & n17387 ) | ( n17383 & n17387 ) ;
  assign n17389 = ~x39 & n17388 ;
  assign n17390 = ( x38 & ~n17381 ) | ( x38 & n17389 ) | ( ~n17381 & n17389 ) ;
  assign n17391 = n17381 | n17390 ;
  assign n17392 = x39 & x142 ;
  assign n17393 = x142 & ~n15340 ;
  assign n17394 = ~n1292 & n17081 ;
  assign n17395 = ( ~x39 & n17393 ) | ( ~x39 & n17394 ) | ( n17393 & n17394 ) ;
  assign n17396 = ~x39 & n17395 ;
  assign n17397 = ( x38 & n17392 ) | ( x38 & ~n17396 ) | ( n17392 & ~n17396 ) ;
  assign n17398 = ~n17392 & n17397 ;
  assign n17399 = ( n2069 & n17391 ) | ( n2069 & ~n17398 ) | ( n17391 & ~n17398 ) ;
  assign n17400 = ~n2069 & n17399 ;
  assign n17401 = n17400 ^ x142 ^ 1'b0 ;
  assign n17402 = ( ~x142 & n2069 ) | ( ~x142 & n17401 ) | ( n2069 & n17401 ) ;
  assign n17403 = ( x142 & n17400 ) | ( x142 & n17402 ) | ( n17400 & n17402 ) ;
  assign n17404 = x625 & ~n17331 ;
  assign n17405 = x1153 | n17404 ;
  assign n17406 = ( x625 & n17403 ) | ( x625 & ~n17405 ) | ( n17403 & ~n17405 ) ;
  assign n17407 = ~n17405 & n17406 ;
  assign n17408 = x625 & ~n17403 ;
  assign n17409 = x625 | n17331 ;
  assign n17410 = ( x1153 & n17408 ) | ( x1153 & n17409 ) | ( n17408 & n17409 ) ;
  assign n17411 = ~n17408 & n17410 ;
  assign n17412 = n17407 | n17411 ;
  assign n17413 = n17403 ^ x778 ^ 1'b0 ;
  assign n17414 = ( n17403 & n17412 ) | ( n17403 & n17413 ) | ( n17412 & n17413 ) ;
  assign n17415 = n17331 ^ n16234 ^ 1'b0 ;
  assign n17416 = ( n17331 & n17414 ) | ( n17331 & ~n17415 ) | ( n17414 & ~n17415 ) ;
  assign n17417 = n17331 ^ n16254 ^ 1'b0 ;
  assign n17418 = ( n17331 & n17416 ) | ( n17331 & ~n17417 ) | ( n17416 & ~n17417 ) ;
  assign n17419 = n17331 ^ n16279 ^ 1'b0 ;
  assign n17420 = ( n17331 & n17418 ) | ( n17331 & ~n17419 ) | ( n17418 & ~n17419 ) ;
  assign n17437 = ~x626 & n17420 ;
  assign n17442 = x142 & n15495 ;
  assign n17438 = x142 | n15636 ;
  assign n17439 = x142 & ~n15330 ;
  assign n17440 = ( x743 & n17438 ) | ( x743 & n17439 ) | ( n17438 & n17439 ) ;
  assign n17441 = n17438 & n17440 ;
  assign n17443 = n17442 ^ n17441 ^ 1'b0 ;
  assign n17444 = ( x299 & ~n17441 ) | ( x299 & n17442 ) | ( ~n17441 & n17442 ) ;
  assign n17445 = ( x299 & ~n17443 ) | ( x299 & n17444 ) | ( ~n17443 & n17444 ) ;
  assign n17446 = x142 & ~x743 ;
  assign n17447 = ~n15327 & n17446 ;
  assign n17448 = x299 | n17447 ;
  assign n17449 = x142 & n15507 ;
  assign n17450 = x142 | n15633 ;
  assign n17451 = x743 & n17450 ;
  assign n17452 = ~n17449 & n17451 ;
  assign n17453 = ( ~n17445 & n17448 ) | ( ~n17445 & n17452 ) | ( n17448 & n17452 ) ;
  assign n17454 = ~n17445 & n17453 ;
  assign n17544 = ~x735 & n17454 ;
  assign n17546 = ~n16034 & n17442 ;
  assign n17545 = n16051 | n17438 ;
  assign n17547 = n17546 ^ n17545 ^ 1'b0 ;
  assign n17548 = ( x743 & ~n17545 ) | ( x743 & n17546 ) | ( ~n17545 & n17546 ) ;
  assign n17549 = ( x743 & ~n17547 ) | ( x743 & n17548 ) | ( ~n17547 & n17548 ) ;
  assign n17550 = ~x142 & n16027 ;
  assign n17551 = x142 & ~n16035 ;
  assign n17552 = ~n15636 & n17551 ;
  assign n17553 = ( x743 & ~n17550 ) | ( x743 & n17552 ) | ( ~n17550 & n17552 ) ;
  assign n17554 = n17550 | n17553 ;
  assign n17555 = ( x299 & n17549 ) | ( x299 & n17554 ) | ( n17549 & n17554 ) ;
  assign n17556 = ~n17549 & n17555 ;
  assign n17557 = n16039 & n17449 ;
  assign n17558 = n16050 | n17450 ;
  assign n17559 = x743 & ~n17558 ;
  assign n17560 = ( x743 & n17557 ) | ( x743 & n17559 ) | ( n17557 & n17559 ) ;
  assign n17561 = ~x142 & n16021 ;
  assign n17562 = x142 & ~n16039 ;
  assign n17563 = ~n15633 & n17562 ;
  assign n17564 = ( x743 & ~n17561 ) | ( x743 & n17563 ) | ( ~n17561 & n17563 ) ;
  assign n17565 = n17561 | n17564 ;
  assign n17566 = ( x299 & ~n17560 ) | ( x299 & n17565 ) | ( ~n17560 & n17565 ) ;
  assign n17567 = ~x299 & n17566 ;
  assign n17568 = ( x735 & n17556 ) | ( x735 & n17567 ) | ( n17556 & n17567 ) ;
  assign n17569 = n17567 ^ n17556 ^ 1'b0 ;
  assign n17570 = ( x735 & n17568 ) | ( x735 & n17569 ) | ( n17568 & n17569 ) ;
  assign n17571 = ( x39 & ~n17544 ) | ( x39 & n17570 ) | ( ~n17544 & n17570 ) ;
  assign n17572 = n17544 | n17571 ;
  assign n17573 = x142 | n15888 ;
  assign n17574 = x142 & n15981 ;
  assign n17575 = x743 & ~n17574 ;
  assign n17576 = n17573 & n17575 ;
  assign n17577 = x142 & n15810 ;
  assign n17578 = x743 | n17577 ;
  assign n17579 = ( x142 & n15769 ) | ( x142 & ~n17578 ) | ( n15769 & ~n17578 ) ;
  assign n17580 = ~n17578 & n17579 ;
  assign n17581 = ( x735 & n17576 ) | ( x735 & n17580 ) | ( n17576 & n17580 ) ;
  assign n17582 = n17580 ^ n17576 ^ 1'b0 ;
  assign n17583 = ( x735 & n17581 ) | ( x735 & n17582 ) | ( n17581 & n17582 ) ;
  assign n17480 = x743 & ~n15879 ;
  assign n17481 = x142 & ~n15554 ;
  assign n17482 = n17480 & ~n17481 ;
  assign n17483 = ( x743 & n17316 ) | ( x743 & ~n17482 ) | ( n17316 & ~n17482 ) ;
  assign n17484 = ~n17482 & n17483 ;
  assign n17584 = x735 | n17484 ;
  assign n17585 = ( ~x735 & n17583 ) | ( ~x735 & n17584 ) | ( n17583 & n17584 ) ;
  assign n17586 = n5114 & ~n17585 ;
  assign n17474 = x743 & ~n15612 ;
  assign n17475 = x142 & ~n15566 ;
  assign n17476 = n17474 & ~n17475 ;
  assign n17477 = ( x743 & n17303 ) | ( x743 & ~n17476 ) | ( n17303 & ~n17476 ) ;
  assign n17478 = ~n17476 & n17477 ;
  assign n17587 = x142 | n15898 ;
  assign n17588 = x743 & n17587 ;
  assign n17589 = x142 | n15754 ;
  assign n17590 = x142 & n15832 ;
  assign n17591 = ( x743 & n17589 ) | ( x743 & ~n17590 ) | ( n17589 & ~n17590 ) ;
  assign n17592 = ~x743 & n17591 ;
  assign n17593 = x142 & n15986 ;
  assign n17594 = ~n17592 & n17593 ;
  assign n17595 = ( n17588 & n17592 ) | ( n17588 & ~n17594 ) | ( n17592 & ~n17594 ) ;
  assign n17596 = n17595 ^ x735 ^ 1'b0 ;
  assign n17597 = ( n17478 & n17595 ) | ( n17478 & ~n17596 ) | ( n17595 & ~n17596 ) ;
  assign n17598 = n5114 | n17597 ;
  assign n17599 = ( x223 & n17586 ) | ( x223 & n17598 ) | ( n17586 & n17598 ) ;
  assign n17600 = ~n17586 & n17599 ;
  assign n17456 = x142 & ~n15522 ;
  assign n17457 = x743 & ~n15601 ;
  assign n17458 = ~n17456 & n17457 ;
  assign n17459 = ( x743 & n17309 ) | ( x743 & ~n17458 ) | ( n17309 & ~n17458 ) ;
  assign n17460 = ~n17458 & n17459 ;
  assign n17601 = x142 & n15953 ;
  assign n17602 = x743 & ~n17601 ;
  assign n17603 = x142 | n15744 ;
  assign n17604 = x142 & n15851 ;
  assign n17605 = ( x743 & n17603 ) | ( x743 & ~n17604 ) | ( n17603 & ~n17604 ) ;
  assign n17606 = ~x743 & n17605 ;
  assign n17607 = x142 | n15911 ;
  assign n17608 = n17606 ^ n17602 ^ 1'b0 ;
  assign n17609 = ( ~n17602 & n17607 ) | ( ~n17602 & n17608 ) | ( n17607 & n17608 ) ;
  assign n17610 = ( n17602 & n17606 ) | ( n17602 & n17609 ) | ( n17606 & n17609 ) ;
  assign n17611 = n17610 ^ x735 ^ 1'b0 ;
  assign n17612 = ( n17460 & n17610 ) | ( n17460 & ~n17611 ) | ( n17610 & ~n17611 ) ;
  assign n17613 = n5114 & n17612 ;
  assign n17614 = x142 & n15963 ;
  assign n17615 = x743 & ~n17614 ;
  assign n17616 = x142 | n15921 ;
  assign n17617 = n17615 & n17616 ;
  assign n17618 = x142 | n15720 ;
  assign n17619 = x142 & n15841 ;
  assign n17620 = ( x743 & n17618 ) | ( x743 & ~n17619 ) | ( n17618 & ~n17619 ) ;
  assign n17621 = ~x743 & n17620 ;
  assign n17622 = ( x735 & n17617 ) | ( x735 & ~n17621 ) | ( n17617 & ~n17621 ) ;
  assign n17623 = ~n17617 & n17622 ;
  assign n17462 = n15599 ^ x142 ^ 1'b0 ;
  assign n17463 = ( ~n15540 & n15599 ) | ( ~n15540 & n17462 ) | ( n15599 & n17462 ) ;
  assign n17464 = n17463 ^ x743 ^ 1'b0 ;
  assign n17465 = ( n17308 & n17463 ) | ( n17308 & ~n17464 ) | ( n17463 & ~n17464 ) ;
  assign n17624 = ( x735 & n17465 ) | ( x735 & ~n17623 ) | ( n17465 & ~n17623 ) ;
  assign n17625 = ~n17623 & n17624 ;
  assign n17626 = ~n5114 & n17625 ;
  assign n17627 = ( n1359 & n17613 ) | ( n1359 & ~n17626 ) | ( n17613 & ~n17626 ) ;
  assign n17628 = ~n17613 & n17627 ;
  assign n17507 = ~n1292 & n17098 ;
  assign n17508 = n17393 | n17507 ;
  assign n17629 = n16068 | n17508 ;
  assign n17630 = ~n15335 & n17629 ;
  assign n17631 = ( x735 & n17306 ) | ( x735 & ~n17630 ) | ( n17306 & ~n17630 ) ;
  assign n17632 = ~n17306 & n17631 ;
  assign n17469 = x743 & n15595 ;
  assign n17470 = n17306 | n17469 ;
  assign n17633 = ( x735 & n17470 ) | ( x735 & ~n17632 ) | ( n17470 & ~n17632 ) ;
  assign n17634 = ~n17632 & n17633 ;
  assign n17635 = n1359 | n17634 ;
  assign n17636 = ( x223 & ~n17628 ) | ( x223 & n17635 ) | ( ~n17628 & n17635 ) ;
  assign n17637 = ~x223 & n17636 ;
  assign n17638 = ( ~x299 & n17600 ) | ( ~x299 & n17637 ) | ( n17600 & n17637 ) ;
  assign n17639 = ~x299 & n17638 ;
  assign n17640 = ~n5061 & n17625 ;
  assign n17641 = n5061 & n17612 ;
  assign n17642 = ( n2263 & n17640 ) | ( n2263 & ~n17641 ) | ( n17640 & ~n17641 ) ;
  assign n17643 = ~n17640 & n17642 ;
  assign n17644 = n2263 | n17634 ;
  assign n17645 = ( x215 & ~n17643 ) | ( x215 & n17644 ) | ( ~n17643 & n17644 ) ;
  assign n17646 = ~x215 & n17645 ;
  assign n17647 = n5061 | n17597 ;
  assign n17648 = n5061 & ~n17585 ;
  assign n17649 = x215 & ~n17648 ;
  assign n17650 = n17647 & n17649 ;
  assign n17651 = ( x299 & n17646 ) | ( x299 & n17650 ) | ( n17646 & n17650 ) ;
  assign n17652 = n17650 ^ n17646 ^ 1'b0 ;
  assign n17653 = ( x299 & n17651 ) | ( x299 & n17652 ) | ( n17651 & n17652 ) ;
  assign n17654 = ( x39 & n17639 ) | ( x39 & ~n17653 ) | ( n17639 & ~n17653 ) ;
  assign n17655 = ~n17639 & n17654 ;
  assign n17656 = ( x38 & n17572 ) | ( x38 & ~n17655 ) | ( n17572 & ~n17655 ) ;
  assign n17657 = n17656 ^ n17572 ^ 1'b0 ;
  assign n17658 = ( x38 & n17656 ) | ( x38 & ~n17657 ) | ( n17656 & ~n17657 ) ;
  assign n17659 = x735 & n16068 ;
  assign n17660 = ( ~x39 & n17508 ) | ( ~x39 & n17659 ) | ( n17508 & n17659 ) ;
  assign n17661 = ~x39 & n17660 ;
  assign n17662 = ( x38 & n17392 ) | ( x38 & ~n17661 ) | ( n17392 & ~n17661 ) ;
  assign n17663 = ~n17392 & n17662 ;
  assign n17664 = ( n2069 & n17658 ) | ( n2069 & ~n17663 ) | ( n17658 & ~n17663 ) ;
  assign n17665 = ~n2069 & n17664 ;
  assign n17666 = n17665 ^ x142 ^ 1'b0 ;
  assign n17667 = ( ~x142 & n2069 ) | ( ~x142 & n17666 ) | ( n2069 & n17666 ) ;
  assign n17668 = ( x142 & n17665 ) | ( x142 & n17667 ) | ( n17665 & n17667 ) ;
  assign n17669 = x625 & ~n17668 ;
  assign n17455 = ~x39 & n17454 ;
  assign n17461 = n5114 & n17460 ;
  assign n17466 = ~n5114 & n17465 ;
  assign n17467 = ( n1359 & n17461 ) | ( n1359 & ~n17466 ) | ( n17461 & ~n17466 ) ;
  assign n17468 = ~n17461 & n17467 ;
  assign n17471 = n1359 | n17470 ;
  assign n17472 = ( x223 & ~n17468 ) | ( x223 & n17471 ) | ( ~n17468 & n17471 ) ;
  assign n17473 = ~x223 & n17472 ;
  assign n17479 = n5114 | n17478 ;
  assign n17485 = n5114 & ~n17484 ;
  assign n17486 = x223 & ~n17485 ;
  assign n17487 = n17479 & n17486 ;
  assign n17488 = ( x299 & ~n17473 ) | ( x299 & n17487 ) | ( ~n17473 & n17487 ) ;
  assign n17489 = n17473 | n17488 ;
  assign n17490 = ~n5061 & n17478 ;
  assign n17491 = n5061 & n17484 ;
  assign n17492 = ( x215 & n17490 ) | ( x215 & ~n17491 ) | ( n17490 & ~n17491 ) ;
  assign n17493 = ~n17490 & n17492 ;
  assign n17494 = n17465 ^ n5061 ^ 1'b0 ;
  assign n17495 = ( n17460 & n17465 ) | ( n17460 & n17494 ) | ( n17465 & n17494 ) ;
  assign n17496 = n2263 & n17495 ;
  assign n17497 = ~n2263 & n17470 ;
  assign n17498 = ( x215 & ~n17496 ) | ( x215 & n17497 ) | ( ~n17496 & n17497 ) ;
  assign n17499 = n17496 | n17498 ;
  assign n17500 = x299 & ~n17499 ;
  assign n17501 = ( x299 & n17493 ) | ( x299 & n17500 ) | ( n17493 & n17500 ) ;
  assign n17502 = x39 & ~n17501 ;
  assign n17503 = n17489 & n17502 ;
  assign n17504 = ( x38 & ~n17455 ) | ( x38 & n17503 ) | ( ~n17455 & n17503 ) ;
  assign n17505 = n17455 | n17504 ;
  assign n17506 = x38 & ~n17392 ;
  assign n17509 = ~x39 & n17508 ;
  assign n17510 = n17506 & ~n17509 ;
  assign n17511 = ( n2069 & n17505 ) | ( n2069 & ~n17510 ) | ( n17505 & ~n17510 ) ;
  assign n17512 = ~n2069 & n17511 ;
  assign n17513 = n17512 ^ x142 ^ 1'b0 ;
  assign n17514 = ( ~x142 & n2069 ) | ( ~x142 & n17513 ) | ( n2069 & n17513 ) ;
  assign n17515 = ( x142 & n17512 ) | ( x142 & n17514 ) | ( n17512 & n17514 ) ;
  assign n17670 = x625 | n17515 ;
  assign n17671 = ( x1153 & n17669 ) | ( x1153 & n17670 ) | ( n17669 & n17670 ) ;
  assign n17672 = ~n17669 & n17671 ;
  assign n17673 = ( x608 & ~n17407 ) | ( x608 & n17672 ) | ( ~n17407 & n17672 ) ;
  assign n17674 = ~n17672 & n17673 ;
  assign n17675 = x625 & ~n17515 ;
  assign n17676 = x1153 | n17675 ;
  assign n17677 = ( n17668 & n17669 ) | ( n17668 & ~n17676 ) | ( n17669 & ~n17676 ) ;
  assign n17678 = ( x608 & ~n17411 ) | ( x608 & n17677 ) | ( ~n17411 & n17677 ) ;
  assign n17679 = n17411 | n17678 ;
  assign n17680 = x778 & ~n17679 ;
  assign n17681 = ( x778 & n17674 ) | ( x778 & n17680 ) | ( n17674 & n17680 ) ;
  assign n17682 = ( x778 & n17668 ) | ( x778 & ~n17681 ) | ( n17668 & ~n17681 ) ;
  assign n17683 = ~n17681 & n17682 ;
  assign n17684 = x609 & ~n17683 ;
  assign n17690 = x609 | n17414 ;
  assign n17691 = ( x1155 & n17684 ) | ( x1155 & n17690 ) | ( n17684 & n17690 ) ;
  assign n17692 = ~n17684 & n17691 ;
  assign n17518 = ~n15659 & n17515 ;
  assign n17519 = ~x609 & n17518 ;
  assign n17520 = n15662 & n17331 ;
  assign n17521 = n17519 | n17520 ;
  assign n17693 = ~x1155 & n17521 ;
  assign n17694 = ( x660 & n17692 ) | ( x660 & ~n17693 ) | ( n17692 & ~n17693 ) ;
  assign n17695 = ~n17692 & n17694 ;
  assign n17522 = x609 & n17518 ;
  assign n17523 = ~n15668 & n17331 ;
  assign n17524 = n17522 | n17523 ;
  assign n17543 = x1155 & n17524 ;
  assign n17685 = x609 & ~n17414 ;
  assign n17686 = x1155 | n17685 ;
  assign n17687 = ( n17683 & n17684 ) | ( n17683 & ~n17686 ) | ( n17684 & ~n17686 ) ;
  assign n17688 = ( x660 & ~n17543 ) | ( x660 & n17687 ) | ( ~n17543 & n17687 ) ;
  assign n17689 = n17543 | n17688 ;
  assign n17696 = n17695 ^ n17689 ^ 1'b0 ;
  assign n17697 = ( x785 & ~n17689 ) | ( x785 & n17695 ) | ( ~n17689 & n17695 ) ;
  assign n17698 = ( x785 & ~n17696 ) | ( x785 & n17697 ) | ( ~n17696 & n17697 ) ;
  assign n17699 = ( x785 & n17683 ) | ( x785 & ~n17698 ) | ( n17683 & ~n17698 ) ;
  assign n17700 = ~n17698 & n17699 ;
  assign n17701 = x618 & ~n17700 ;
  assign n17707 = x618 | n17416 ;
  assign n17708 = ( x1154 & n17701 ) | ( x1154 & n17707 ) | ( n17701 & n17707 ) ;
  assign n17709 = ~n17701 & n17708 ;
  assign n17516 = n17515 ^ n15659 ^ 1'b0 ;
  assign n17517 = ( n17331 & n17515 ) | ( n17331 & n17516 ) | ( n17515 & n17516 ) ;
  assign n17525 = n17524 ^ x1155 ^ 1'b0 ;
  assign n17526 = ( n17521 & n17524 ) | ( n17521 & ~n17525 ) | ( n17524 & ~n17525 ) ;
  assign n17527 = n17517 ^ x785 ^ 1'b0 ;
  assign n17528 = ( n17517 & n17526 ) | ( n17517 & n17527 ) | ( n17526 & n17527 ) ;
  assign n17529 = x618 & ~n17528 ;
  assign n17533 = x618 & ~n17331 ;
  assign n17534 = x1154 | n17533 ;
  assign n17535 = ( n17528 & n17529 ) | ( n17528 & ~n17534 ) | ( n17529 & ~n17534 ) ;
  assign n17710 = ( x627 & ~n17535 ) | ( x627 & n17709 ) | ( ~n17535 & n17709 ) ;
  assign n17711 = ~n17709 & n17710 ;
  assign n17530 = x618 | n17331 ;
  assign n17531 = ( x1154 & n17529 ) | ( x1154 & n17530 ) | ( n17529 & n17530 ) ;
  assign n17532 = ~n17529 & n17531 ;
  assign n17702 = x618 & ~n17416 ;
  assign n17703 = x1154 | n17702 ;
  assign n17704 = ( n17700 & n17701 ) | ( n17700 & ~n17703 ) | ( n17701 & ~n17703 ) ;
  assign n17705 = ( x627 & ~n17532 ) | ( x627 & n17704 ) | ( ~n17532 & n17704 ) ;
  assign n17706 = n17532 | n17705 ;
  assign n17712 = n17711 ^ n17706 ^ 1'b0 ;
  assign n17713 = ( x781 & ~n17706 ) | ( x781 & n17711 ) | ( ~n17706 & n17711 ) ;
  assign n17714 = ( x781 & ~n17712 ) | ( x781 & n17713 ) | ( ~n17712 & n17713 ) ;
  assign n17715 = ( x781 & n17700 ) | ( x781 & ~n17714 ) | ( n17700 & ~n17714 ) ;
  assign n17716 = ~n17714 & n17715 ;
  assign n17717 = x619 & ~n17716 ;
  assign n17723 = x619 | n17418 ;
  assign n17724 = ( x1159 & n17717 ) | ( x1159 & n17723 ) | ( n17717 & n17723 ) ;
  assign n17725 = ~n17717 & n17724 ;
  assign n17536 = n17532 | n17535 ;
  assign n17537 = n17528 ^ x781 ^ 1'b0 ;
  assign n17538 = ( n17528 & n17536 ) | ( n17528 & n17537 ) | ( n17536 & n17537 ) ;
  assign n17539 = x619 & ~n17538 ;
  assign n17726 = x619 & ~n17331 ;
  assign n17727 = x1159 | n17726 ;
  assign n17728 = ( n17538 & n17539 ) | ( n17538 & ~n17727 ) | ( n17539 & ~n17727 ) ;
  assign n17729 = ( x648 & n17725 ) | ( x648 & ~n17728 ) | ( n17725 & ~n17728 ) ;
  assign n17730 = ~n17725 & n17729 ;
  assign n17540 = x619 | n17331 ;
  assign n17541 = ( x1159 & n17539 ) | ( x1159 & n17540 ) | ( n17539 & n17540 ) ;
  assign n17542 = ~n17539 & n17541 ;
  assign n17718 = x619 & ~n17418 ;
  assign n17719 = x1159 | n17718 ;
  assign n17720 = ( n17716 & n17717 ) | ( n17716 & ~n17719 ) | ( n17717 & ~n17719 ) ;
  assign n17721 = ( x648 & ~n17542 ) | ( x648 & n17720 ) | ( ~n17542 & n17720 ) ;
  assign n17722 = n17542 | n17721 ;
  assign n17731 = n17730 ^ n17722 ^ 1'b0 ;
  assign n17732 = ( x789 & ~n17722 ) | ( x789 & n17730 ) | ( ~n17722 & n17730 ) ;
  assign n17733 = ( x789 & ~n17731 ) | ( x789 & n17732 ) | ( ~n17731 & n17732 ) ;
  assign n17734 = ( x789 & n17716 ) | ( x789 & ~n17733 ) | ( n17716 & ~n17733 ) ;
  assign n17735 = ~n17733 & n17734 ;
  assign n17736 = x626 & n17735 ;
  assign n17737 = ( x641 & n17437 ) | ( x641 & ~n17736 ) | ( n17437 & ~n17736 ) ;
  assign n17738 = ~n17437 & n17737 ;
  assign n17739 = n17542 | n17728 ;
  assign n17740 = n17538 ^ x789 ^ 1'b0 ;
  assign n17741 = ( n17538 & n17739 ) | ( n17538 & n17740 ) | ( n17739 & n17740 ) ;
  assign n17742 = x626 & ~n17741 ;
  assign n17743 = x626 | n17331 ;
  assign n17744 = ( x1158 & n17742 ) | ( x1158 & n17743 ) | ( n17742 & n17743 ) ;
  assign n17745 = ~n17742 & n17744 ;
  assign n17746 = n16289 | n17745 ;
  assign n17747 = ~n17738 & n17746 ;
  assign n17748 = ~x626 & n17735 ;
  assign n17749 = x626 & n17420 ;
  assign n17750 = ( x641 & ~n17748 ) | ( x641 & n17749 ) | ( ~n17748 & n17749 ) ;
  assign n17751 = n17748 | n17750 ;
  assign n17752 = x626 & ~n17331 ;
  assign n17753 = x1158 | n17752 ;
  assign n17754 = ( n17741 & n17742 ) | ( n17741 & ~n17753 ) | ( n17742 & ~n17753 ) ;
  assign n17755 = ( ~n16299 & n17751 ) | ( ~n16299 & n17754 ) | ( n17751 & n17754 ) ;
  assign n17756 = n17751 ^ n16299 ^ 1'b0 ;
  assign n17757 = ( n17751 & n17755 ) | ( n17751 & n17756 ) | ( n17755 & n17756 ) ;
  assign n17758 = ( x788 & n17747 ) | ( x788 & ~n17757 ) | ( n17747 & ~n17757 ) ;
  assign n17759 = ~n17747 & n17758 ;
  assign n17760 = ( x788 & n17735 ) | ( x788 & ~n17759 ) | ( n17735 & ~n17759 ) ;
  assign n17761 = ~n17759 & n17760 ;
  assign n17762 = x628 & ~n17761 ;
  assign n17763 = n17745 | n17754 ;
  assign n17764 = n17741 ^ x788 ^ 1'b0 ;
  assign n17765 = ( n17741 & n17763 ) | ( n17741 & n17764 ) | ( n17763 & n17764 ) ;
  assign n17771 = x628 | n17765 ;
  assign n17772 = ( x1156 & n17762 ) | ( x1156 & n17771 ) | ( n17762 & n17771 ) ;
  assign n17773 = ~n17762 & n17772 ;
  assign n17421 = n17331 ^ n16318 ^ 1'b0 ;
  assign n17422 = ( n17331 & n17420 ) | ( n17331 & ~n17421 ) | ( n17420 & ~n17421 ) ;
  assign n17423 = x628 & ~n17422 ;
  assign n17427 = x628 & ~n17331 ;
  assign n17428 = x1156 | n17427 ;
  assign n17429 = ( n17422 & n17423 ) | ( n17422 & ~n17428 ) | ( n17423 & ~n17428 ) ;
  assign n17774 = ( x629 & ~n17429 ) | ( x629 & n17773 ) | ( ~n17429 & n17773 ) ;
  assign n17775 = ~n17773 & n17774 ;
  assign n17424 = x628 | n17331 ;
  assign n17425 = ( x1156 & n17423 ) | ( x1156 & n17424 ) | ( n17423 & n17424 ) ;
  assign n17426 = ~n17423 & n17425 ;
  assign n17766 = x628 & ~n17765 ;
  assign n17767 = x1156 | n17766 ;
  assign n17768 = ( n17761 & n17762 ) | ( n17761 & ~n17767 ) | ( n17762 & ~n17767 ) ;
  assign n17769 = ( x629 & ~n17426 ) | ( x629 & n17768 ) | ( ~n17426 & n17768 ) ;
  assign n17770 = n17426 | n17769 ;
  assign n17776 = n17775 ^ n17770 ^ 1'b0 ;
  assign n17777 = ( x792 & ~n17770 ) | ( x792 & n17775 ) | ( ~n17770 & n17775 ) ;
  assign n17778 = ( x792 & ~n17776 ) | ( x792 & n17777 ) | ( ~n17776 & n17777 ) ;
  assign n17779 = ( x792 & n17761 ) | ( x792 & ~n17778 ) | ( n17761 & ~n17778 ) ;
  assign n17780 = ~n17778 & n17779 ;
  assign n17781 = x647 & ~n17780 ;
  assign n17782 = n17331 ^ n16339 ^ 1'b0 ;
  assign n17783 = ( n17331 & n17765 ) | ( n17331 & ~n17782 ) | ( n17765 & ~n17782 ) ;
  assign n17789 = x647 | n17783 ;
  assign n17790 = ( x1157 & n17781 ) | ( x1157 & n17789 ) | ( n17781 & n17789 ) ;
  assign n17791 = ~n17781 & n17790 ;
  assign n17430 = n17426 | n17429 ;
  assign n17431 = n17422 ^ x792 ^ 1'b0 ;
  assign n17432 = ( n17422 & n17430 ) | ( n17422 & n17431 ) | ( n17430 & n17431 ) ;
  assign n17433 = x647 & ~n17432 ;
  assign n17792 = x647 & ~n17331 ;
  assign n17793 = x1157 | n17792 ;
  assign n17794 = ( n17432 & n17433 ) | ( n17432 & ~n17793 ) | ( n17433 & ~n17793 ) ;
  assign n17795 = ( x630 & n17791 ) | ( x630 & ~n17794 ) | ( n17791 & ~n17794 ) ;
  assign n17796 = ~n17791 & n17795 ;
  assign n17434 = x647 | n17331 ;
  assign n17435 = ( x1157 & n17433 ) | ( x1157 & n17434 ) | ( n17433 & n17434 ) ;
  assign n17436 = ~n17433 & n17435 ;
  assign n17784 = x647 & ~n17783 ;
  assign n17785 = x1157 | n17784 ;
  assign n17786 = ( n17780 & n17781 ) | ( n17780 & ~n17785 ) | ( n17781 & ~n17785 ) ;
  assign n17787 = ( x630 & ~n17436 ) | ( x630 & n17786 ) | ( ~n17436 & n17786 ) ;
  assign n17788 = n17436 | n17787 ;
  assign n17797 = n17796 ^ n17788 ^ 1'b0 ;
  assign n17798 = ( x787 & ~n17788 ) | ( x787 & n17796 ) | ( ~n17788 & n17796 ) ;
  assign n17799 = ( x787 & ~n17797 ) | ( x787 & n17798 ) | ( ~n17797 & n17798 ) ;
  assign n17800 = ( x787 & n17780 ) | ( x787 & ~n17799 ) | ( n17780 & ~n17799 ) ;
  assign n17801 = ~n17799 & n17800 ;
  assign n17802 = ~x790 & n17801 ;
  assign n17810 = x644 & ~n17331 ;
  assign n17811 = x715 & ~n17810 ;
  assign n17812 = n17331 ^ n16376 ^ 1'b0 ;
  assign n17813 = ( n17331 & n17783 ) | ( n17331 & ~n17812 ) | ( n17783 & ~n17812 ) ;
  assign n17814 = x644 & ~n17813 ;
  assign n17815 = ( n17811 & n17813 ) | ( n17811 & n17814 ) | ( n17813 & n17814 ) ;
  assign n17803 = x644 | n17801 ;
  assign n17804 = n17436 | n17794 ;
  assign n17805 = n17432 ^ x787 ^ 1'b0 ;
  assign n17806 = ( n17432 & n17804 ) | ( n17432 & n17805 ) | ( n17804 & n17805 ) ;
  assign n17807 = x644 & ~n17806 ;
  assign n17808 = ( x715 & n17803 ) | ( x715 & ~n17807 ) | ( n17803 & ~n17807 ) ;
  assign n17809 = ~x715 & n17808 ;
  assign n17816 = ( x1160 & n17809 ) | ( x1160 & ~n17815 ) | ( n17809 & ~n17815 ) ;
  assign n17817 = n17815 | n17816 ;
  assign n17818 = x644 & ~n17801 ;
  assign n17819 = x644 | n17806 ;
  assign n17820 = ( x715 & n17818 ) | ( x715 & n17819 ) | ( n17818 & n17819 ) ;
  assign n17821 = ~n17818 & n17820 ;
  assign n17822 = x644 | n17331 ;
  assign n17823 = ( x715 & ~n17814 ) | ( x715 & n17822 ) | ( ~n17814 & n17822 ) ;
  assign n17824 = ~x715 & n17823 ;
  assign n17825 = ( x1160 & n17821 ) | ( x1160 & ~n17824 ) | ( n17821 & ~n17824 ) ;
  assign n17826 = ~n17821 & n17825 ;
  assign n17827 = x790 & ~n17826 ;
  assign n17828 = n17817 & n17827 ;
  assign n17829 = ( n5193 & ~n17802 ) | ( n5193 & n17828 ) | ( ~n17802 & n17828 ) ;
  assign n17830 = n17802 | n17829 ;
  assign n17831 = ( x57 & ~n17302 ) | ( x57 & n17830 ) | ( ~n17302 & n17830 ) ;
  assign n17832 = ~x57 & n17831 ;
  assign n17833 = x57 & x142 ;
  assign n17834 = x832 | n17833 ;
  assign n17835 = ( ~n17301 & n17832 ) | ( ~n17301 & n17834 ) | ( n17832 & n17834 ) ;
  assign n17836 = ~n17301 & n17835 ;
  assign n17838 = ~n5052 & n15591 ;
  assign n17839 = x38 & n17838 ;
  assign n17840 = ~n5017 & n15547 ;
  assign n17841 = x38 & ~n17840 ;
  assign n17842 = x38 | n15587 ;
  assign n17843 = ~n17841 & n17842 ;
  assign n17844 = x143 | x774 ;
  assign n17845 = n17843 & ~n17844 ;
  assign n17846 = ~x38 & n15640 ;
  assign n17847 = x143 & ~n17846 ;
  assign n17848 = ( ~n17839 & n17845 ) | ( ~n17839 & n17847 ) | ( n17845 & n17847 ) ;
  assign n17849 = ~n17839 & n17848 ;
  assign n17850 = x143 | n15655 ;
  assign n17851 = n17849 ^ x774 ^ 1'b0 ;
  assign n17852 = ( ~x774 & n17850 ) | ( ~x774 & n17851 ) | ( n17850 & n17851 ) ;
  assign n17853 = ( x774 & n17849 ) | ( x774 & n17852 ) | ( n17849 & n17852 ) ;
  assign n17881 = x687 | n17853 ;
  assign n17882 = x38 & n16658 ;
  assign n17883 = x774 & ~n17882 ;
  assign n17884 = n15795 ^ x39 ^ 1'b0 ;
  assign n17885 = ( n15795 & n16029 ) | ( n15795 & ~n17884 ) | ( n16029 & ~n17884 ) ;
  assign n17886 = ~x38 & n17885 ;
  assign n17887 = x143 & n17886 ;
  assign n17888 = n17883 & ~n17887 ;
  assign n17889 = n15644 & ~n15691 ;
  assign n17890 = n15876 ^ x39 ^ 1'b0 ;
  assign n17891 = ( n15876 & n16044 ) | ( n15876 & ~n17890 ) | ( n16044 & ~n17890 ) ;
  assign n17892 = n17889 ^ x38 ^ 1'b0 ;
  assign n17893 = ( n17889 & n17891 ) | ( n17889 & ~n17892 ) | ( n17891 & ~n17892 ) ;
  assign n17894 = x143 | n17893 ;
  assign n17895 = n17888 & n17894 ;
  assign n17896 = x39 | n16048 ;
  assign n17897 = ~x39 & n15968 ;
  assign n17898 = n17896 ^ x38 ^ 1'b0 ;
  assign n17899 = ( n17896 & n17897 ) | ( n17896 & n17898 ) | ( n17897 & n17898 ) ;
  assign n17900 = n17899 ^ n16003 ^ 1'b0 ;
  assign n17901 = ( ~x39 & n16003 ) | ( ~x39 & n17900 ) | ( n16003 & n17900 ) ;
  assign n17902 = ( n17899 & ~n17900 ) | ( n17899 & n17901 ) | ( ~n17900 & n17901 ) ;
  assign n17903 = x143 | n17902 ;
  assign n17904 = ~n5017 & n15779 ;
  assign n17905 = x38 & ~n17904 ;
  assign n17906 = x39 & ~n15943 ;
  assign n17907 = n15639 | n16053 ;
  assign n17908 = ~n17906 & n17907 ;
  assign n17909 = x38 | n17908 ;
  assign n17910 = ~n17905 & n17909 ;
  assign n17911 = x143 & n17910 ;
  assign n17912 = ( x774 & n17903 ) | ( x774 & ~n17911 ) | ( n17903 & ~n17911 ) ;
  assign n17913 = ~x774 & n17912 ;
  assign n17914 = ( x687 & n17895 ) | ( x687 & ~n17913 ) | ( n17895 & ~n17913 ) ;
  assign n17915 = ~n17895 & n17914 ;
  assign n17916 = ( n2069 & n17881 ) | ( n2069 & ~n17915 ) | ( n17881 & ~n17915 ) ;
  assign n17917 = ~n2069 & n17916 ;
  assign n17918 = n17917 ^ x143 ^ 1'b0 ;
  assign n17919 = ( ~x143 & n2069 ) | ( ~x143 & n17918 ) | ( n2069 & n17918 ) ;
  assign n17920 = ( x143 & n17917 ) | ( x143 & n17919 ) | ( n17917 & n17919 ) ;
  assign n17921 = x625 & ~n17920 ;
  assign n17837 = x143 & n2069 ;
  assign n17854 = ~n2069 & n17853 ;
  assign n17855 = n17837 | n17854 ;
  assign n17922 = x625 | n17855 ;
  assign n17923 = ( x1153 & n17921 ) | ( x1153 & n17922 ) | ( n17921 & n17922 ) ;
  assign n17924 = ~n17921 & n17923 ;
  assign n17856 = x143 | n15656 ;
  assign n17925 = x625 & ~n17856 ;
  assign n17926 = x1153 | n17925 ;
  assign n17927 = ( x38 & x143 ) | ( x38 & n16700 ) | ( x143 & n16700 ) ;
  assign n17928 = ( x143 & n16697 ) | ( x143 & ~n17927 ) | ( n16697 & ~n17927 ) ;
  assign n17929 = ~n17927 & n17928 ;
  assign n17930 = x143 | n15644 ;
  assign n17931 = n16185 & n17930 ;
  assign n17932 = ( x687 & n17929 ) | ( x687 & ~n17931 ) | ( n17929 & ~n17931 ) ;
  assign n17933 = ~n17929 & n17932 ;
  assign n17934 = x687 | n17850 ;
  assign n17935 = ~n2069 & n17934 ;
  assign n17936 = n17935 ^ n17933 ^ 1'b0 ;
  assign n17937 = ( n17933 & n17935 ) | ( n17933 & n17936 ) | ( n17935 & n17936 ) ;
  assign n17938 = ( n17837 & ~n17933 ) | ( n17837 & n17937 ) | ( ~n17933 & n17937 ) ;
  assign n17939 = ( x625 & ~n17926 ) | ( x625 & n17938 ) | ( ~n17926 & n17938 ) ;
  assign n17940 = ~n17926 & n17939 ;
  assign n17941 = ( x608 & n17924 ) | ( x608 & ~n17940 ) | ( n17924 & ~n17940 ) ;
  assign n17942 = ~n17924 & n17941 ;
  assign n17943 = x625 & ~n17938 ;
  assign n17944 = x625 | n17856 ;
  assign n17945 = ( x1153 & n17943 ) | ( x1153 & n17944 ) | ( n17943 & n17944 ) ;
  assign n17946 = ~n17943 & n17945 ;
  assign n17947 = x608 | n17946 ;
  assign n17948 = x625 & ~n17855 ;
  assign n17949 = x1153 | n17948 ;
  assign n17950 = ( n17920 & n17921 ) | ( n17920 & ~n17949 ) | ( n17921 & ~n17949 ) ;
  assign n17951 = ( ~n17942 & n17947 ) | ( ~n17942 & n17950 ) | ( n17947 & n17950 ) ;
  assign n17952 = ~n17942 & n17951 ;
  assign n17953 = n17920 ^ x778 ^ 1'b0 ;
  assign n17954 = ( n17920 & n17952 ) | ( n17920 & n17953 ) | ( n17952 & n17953 ) ;
  assign n17955 = x609 & ~n17954 ;
  assign n17956 = n17940 | n17946 ;
  assign n17957 = n17938 ^ x778 ^ 1'b0 ;
  assign n17958 = ( n17938 & n17956 ) | ( n17938 & n17957 ) | ( n17956 & n17957 ) ;
  assign n17959 = x609 | n17958 ;
  assign n17960 = ( x1155 & n17955 ) | ( x1155 & n17959 ) | ( n17955 & n17959 ) ;
  assign n17961 = ~n17955 & n17960 ;
  assign n17859 = ~n15668 & n17856 ;
  assign n17860 = ( n15668 & n17837 ) | ( n15668 & n17854 ) | ( n17837 & n17854 ) ;
  assign n17861 = n17859 | n17860 ;
  assign n17857 = n17855 ^ n15659 ^ 1'b0 ;
  assign n17858 = ( n17855 & n17856 ) | ( n17855 & n17857 ) | ( n17856 & n17857 ) ;
  assign n17863 = n17861 ^ n17858 ^ n17856 ;
  assign n17962 = ~x1155 & n17863 ;
  assign n17963 = ( x660 & n17961 ) | ( x660 & ~n17962 ) | ( n17961 & ~n17962 ) ;
  assign n17964 = ~n17961 & n17963 ;
  assign n17965 = x1155 & n17861 ;
  assign n17966 = x660 | n17965 ;
  assign n17967 = x609 & ~n17958 ;
  assign n17968 = x1155 | n17967 ;
  assign n17969 = ( n17954 & n17955 ) | ( n17954 & ~n17968 ) | ( n17955 & ~n17968 ) ;
  assign n17970 = ( ~n17964 & n17966 ) | ( ~n17964 & n17969 ) | ( n17966 & n17969 ) ;
  assign n17971 = ~n17964 & n17970 ;
  assign n17972 = n17954 ^ x785 ^ 1'b0 ;
  assign n17973 = ( n17954 & n17971 ) | ( n17954 & n17972 ) | ( n17971 & n17972 ) ;
  assign n17974 = x618 & ~n17973 ;
  assign n17975 = n17856 ^ n16234 ^ 1'b0 ;
  assign n17976 = ( n17856 & n17958 ) | ( n17856 & ~n17975 ) | ( n17958 & ~n17975 ) ;
  assign n17977 = x618 | n17976 ;
  assign n17978 = ( x1154 & n17974 ) | ( x1154 & n17977 ) | ( n17974 & n17977 ) ;
  assign n17979 = ~n17974 & n17978 ;
  assign n17862 = n17861 ^ x1155 ^ 1'b0 ;
  assign n17864 = ( n17861 & ~n17862 ) | ( n17861 & n17863 ) | ( ~n17862 & n17863 ) ;
  assign n17865 = n17858 ^ x785 ^ 1'b0 ;
  assign n17866 = ( n17858 & n17864 ) | ( n17858 & n17865 ) | ( n17864 & n17865 ) ;
  assign n17867 = x618 & ~n17866 ;
  assign n17871 = x618 & ~n17856 ;
  assign n17872 = x1154 | n17871 ;
  assign n17873 = ( n17866 & n17867 ) | ( n17866 & ~n17872 ) | ( n17867 & ~n17872 ) ;
  assign n17980 = ( x627 & ~n17873 ) | ( x627 & n17979 ) | ( ~n17873 & n17979 ) ;
  assign n17981 = ~n17979 & n17980 ;
  assign n17868 = x618 | n17856 ;
  assign n17869 = ( x1154 & n17867 ) | ( x1154 & n17868 ) | ( n17867 & n17868 ) ;
  assign n17870 = ~n17867 & n17869 ;
  assign n17982 = x627 | n17870 ;
  assign n17983 = x618 & ~n17976 ;
  assign n17984 = x1154 | n17983 ;
  assign n17985 = ( n17973 & n17974 ) | ( n17973 & ~n17984 ) | ( n17974 & ~n17984 ) ;
  assign n17986 = ( ~n17981 & n17982 ) | ( ~n17981 & n17985 ) | ( n17982 & n17985 ) ;
  assign n17987 = ~n17981 & n17986 ;
  assign n17988 = n17973 ^ x781 ^ 1'b0 ;
  assign n17989 = ( n17973 & n17987 ) | ( n17973 & n17988 ) | ( n17987 & n17988 ) ;
  assign n17990 = x619 & ~n17989 ;
  assign n17991 = n17856 ^ n16254 ^ 1'b0 ;
  assign n17992 = ( n17856 & n17976 ) | ( n17856 & ~n17991 ) | ( n17976 & ~n17991 ) ;
  assign n17998 = x619 | n17992 ;
  assign n17999 = ( x1159 & n17990 ) | ( x1159 & n17998 ) | ( n17990 & n17998 ) ;
  assign n18000 = ~n17990 & n17999 ;
  assign n17874 = n17870 | n17873 ;
  assign n17875 = n17866 ^ x781 ^ 1'b0 ;
  assign n17876 = ( n17866 & n17874 ) | ( n17866 & n17875 ) | ( n17874 & n17875 ) ;
  assign n17877 = x619 & ~n17876 ;
  assign n18001 = x619 & ~n17856 ;
  assign n18002 = x1159 | n18001 ;
  assign n18003 = ( n17876 & n17877 ) | ( n17876 & ~n18002 ) | ( n17877 & ~n18002 ) ;
  assign n18004 = ( x648 & n18000 ) | ( x648 & ~n18003 ) | ( n18000 & ~n18003 ) ;
  assign n18005 = ~n18000 & n18004 ;
  assign n17878 = x619 | n17856 ;
  assign n17879 = ( x1159 & n17877 ) | ( x1159 & n17878 ) | ( n17877 & n17878 ) ;
  assign n17880 = ~n17877 & n17879 ;
  assign n17993 = x619 & ~n17992 ;
  assign n17994 = x1159 | n17993 ;
  assign n17995 = ( n17989 & n17990 ) | ( n17989 & ~n17994 ) | ( n17990 & ~n17994 ) ;
  assign n17996 = ( x648 & ~n17880 ) | ( x648 & n17995 ) | ( ~n17880 & n17995 ) ;
  assign n17997 = n17880 | n17996 ;
  assign n18006 = n18005 ^ n17997 ^ 1'b0 ;
  assign n18007 = ( x789 & ~n17997 ) | ( x789 & n18005 ) | ( ~n17997 & n18005 ) ;
  assign n18008 = ( x789 & ~n18006 ) | ( x789 & n18007 ) | ( ~n18006 & n18007 ) ;
  assign n18009 = ( x789 & n17989 ) | ( x789 & ~n18008 ) | ( n17989 & ~n18008 ) ;
  assign n18010 = ~n18008 & n18009 ;
  assign n18011 = ~x626 & n18010 ;
  assign n18012 = n17856 ^ n16279 ^ 1'b0 ;
  assign n18013 = ( n17856 & n17992 ) | ( n17856 & ~n18012 ) | ( n17992 & ~n18012 ) ;
  assign n18014 = x626 & n18013 ;
  assign n18015 = ( x641 & ~n18011 ) | ( x641 & n18014 ) | ( ~n18011 & n18014 ) ;
  assign n18016 = n18011 | n18015 ;
  assign n18017 = ~x626 & n18013 ;
  assign n18018 = x626 & n18010 ;
  assign n18019 = ( x641 & n18017 ) | ( x641 & ~n18018 ) | ( n18017 & ~n18018 ) ;
  assign n18020 = ~n18017 & n18019 ;
  assign n18021 = n17880 | n18003 ;
  assign n18022 = n17876 ^ x789 ^ 1'b0 ;
  assign n18023 = ( n17876 & n18021 ) | ( n17876 & n18022 ) | ( n18021 & n18022 ) ;
  assign n18024 = x626 & ~n18023 ;
  assign n18025 = x626 | n17856 ;
  assign n18026 = ( x1158 & n18024 ) | ( x1158 & n18025 ) | ( n18024 & n18025 ) ;
  assign n18027 = ~n18024 & n18026 ;
  assign n18028 = n16289 | n18027 ;
  assign n18029 = ~n18020 & n18028 ;
  assign n18030 = x626 & ~n17856 ;
  assign n18031 = x1158 | n18030 ;
  assign n18032 = ( n18023 & n18024 ) | ( n18023 & ~n18031 ) | ( n18024 & ~n18031 ) ;
  assign n18033 = n16299 & ~n18032 ;
  assign n18034 = ~n18029 & n18033 ;
  assign n18035 = ( n18016 & n18029 ) | ( n18016 & ~n18034 ) | ( n18029 & ~n18034 ) ;
  assign n18036 = n18010 ^ x788 ^ 1'b0 ;
  assign n18037 = ( n18010 & n18035 ) | ( n18010 & n18036 ) | ( n18035 & n18036 ) ;
  assign n18038 = x628 & ~n18037 ;
  assign n18039 = n18027 | n18032 ;
  assign n18040 = n18023 ^ x788 ^ 1'b0 ;
  assign n18041 = ( n18023 & n18039 ) | ( n18023 & n18040 ) | ( n18039 & n18040 ) ;
  assign n18042 = x628 | n18041 ;
  assign n18043 = ( x1156 & n18038 ) | ( x1156 & n18042 ) | ( n18038 & n18042 ) ;
  assign n18044 = ~n18038 & n18043 ;
  assign n18045 = x628 & ~n17856 ;
  assign n18046 = x1156 | n18045 ;
  assign n18047 = n17856 ^ n16318 ^ 1'b0 ;
  assign n18048 = ( n17856 & n18013 ) | ( n17856 & ~n18047 ) | ( n18013 & ~n18047 ) ;
  assign n18049 = x628 & ~n18048 ;
  assign n18050 = ( ~n18046 & n18048 ) | ( ~n18046 & n18049 ) | ( n18048 & n18049 ) ;
  assign n18051 = ( x629 & n18044 ) | ( x629 & ~n18050 ) | ( n18044 & ~n18050 ) ;
  assign n18052 = ~n18044 & n18051 ;
  assign n18053 = x628 | n17856 ;
  assign n18054 = ( x1156 & n18049 ) | ( x1156 & n18053 ) | ( n18049 & n18053 ) ;
  assign n18055 = ~n18049 & n18054 ;
  assign n18056 = x629 | n18055 ;
  assign n18057 = x628 & ~n18041 ;
  assign n18058 = x1156 | n18057 ;
  assign n18059 = ( n18037 & n18038 ) | ( n18037 & ~n18058 ) | ( n18038 & ~n18058 ) ;
  assign n18060 = ( ~n18052 & n18056 ) | ( ~n18052 & n18059 ) | ( n18056 & n18059 ) ;
  assign n18061 = ~n18052 & n18060 ;
  assign n18062 = n18037 ^ x792 ^ 1'b0 ;
  assign n18063 = ( n18037 & n18061 ) | ( n18037 & n18062 ) | ( n18061 & n18062 ) ;
  assign n18064 = x647 & ~n18063 ;
  assign n18065 = n17856 ^ n16339 ^ 1'b0 ;
  assign n18066 = ( n17856 & n18041 ) | ( n17856 & ~n18065 ) | ( n18041 & ~n18065 ) ;
  assign n18067 = x647 | n18066 ;
  assign n18068 = ( x1157 & n18064 ) | ( x1157 & n18067 ) | ( n18064 & n18067 ) ;
  assign n18069 = ~n18064 & n18068 ;
  assign n18070 = x647 & ~n17856 ;
  assign n18071 = x1157 | n18070 ;
  assign n18072 = n18050 | n18055 ;
  assign n18073 = n18048 ^ x792 ^ 1'b0 ;
  assign n18074 = ( n18048 & n18072 ) | ( n18048 & n18073 ) | ( n18072 & n18073 ) ;
  assign n18075 = x647 & ~n18074 ;
  assign n18076 = ( ~n18071 & n18074 ) | ( ~n18071 & n18075 ) | ( n18074 & n18075 ) ;
  assign n18077 = ( x630 & n18069 ) | ( x630 & ~n18076 ) | ( n18069 & ~n18076 ) ;
  assign n18078 = ~n18069 & n18077 ;
  assign n18079 = x647 | n17856 ;
  assign n18080 = ( x1157 & n18075 ) | ( x1157 & n18079 ) | ( n18075 & n18079 ) ;
  assign n18081 = ~n18075 & n18080 ;
  assign n18082 = x630 | n18081 ;
  assign n18083 = x647 & ~n18066 ;
  assign n18084 = x1157 | n18083 ;
  assign n18085 = ( n18063 & n18064 ) | ( n18063 & ~n18084 ) | ( n18064 & ~n18084 ) ;
  assign n18086 = ( ~n18078 & n18082 ) | ( ~n18078 & n18085 ) | ( n18082 & n18085 ) ;
  assign n18087 = ~n18078 & n18086 ;
  assign n18088 = n18063 ^ x787 ^ 1'b0 ;
  assign n18089 = ( n18063 & n18087 ) | ( n18063 & n18088 ) | ( n18087 & n18088 ) ;
  assign n18090 = x644 & ~n18089 ;
  assign n18091 = n18076 | n18081 ;
  assign n18092 = n18074 ^ x787 ^ 1'b0 ;
  assign n18093 = ( n18074 & n18091 ) | ( n18074 & n18092 ) | ( n18091 & n18092 ) ;
  assign n18094 = x644 | n18093 ;
  assign n18095 = ( x715 & n18090 ) | ( x715 & n18094 ) | ( n18090 & n18094 ) ;
  assign n18096 = ~n18090 & n18095 ;
  assign n18097 = x644 | n17856 ;
  assign n18098 = n17856 ^ n16376 ^ 1'b0 ;
  assign n18099 = ( n17856 & n18066 ) | ( n17856 & ~n18098 ) | ( n18066 & ~n18098 ) ;
  assign n18100 = x644 & ~n18099 ;
  assign n18101 = ( x715 & n18097 ) | ( x715 & ~n18100 ) | ( n18097 & ~n18100 ) ;
  assign n18102 = ~x715 & n18101 ;
  assign n18103 = ( x1160 & n18096 ) | ( x1160 & ~n18102 ) | ( n18096 & ~n18102 ) ;
  assign n18104 = ~n18096 & n18103 ;
  assign n18105 = x644 & ~n17856 ;
  assign n18106 = x715 & ~n18105 ;
  assign n18107 = ( n18099 & n18100 ) | ( n18099 & n18106 ) | ( n18100 & n18106 ) ;
  assign n18108 = x644 & ~n18093 ;
  assign n18109 = x715 | n18108 ;
  assign n18110 = ( n18089 & n18090 ) | ( n18089 & ~n18109 ) | ( n18090 & ~n18109 ) ;
  assign n18111 = ( x1160 & ~n18107 ) | ( x1160 & n18110 ) | ( ~n18107 & n18110 ) ;
  assign n18112 = n18107 | n18111 ;
  assign n18113 = ( x790 & n18104 ) | ( x790 & n18112 ) | ( n18104 & n18112 ) ;
  assign n18114 = ~n18104 & n18113 ;
  assign n18115 = ~x790 & n18089 ;
  assign n18116 = ( n7318 & ~n18114 ) | ( n7318 & n18115 ) | ( ~n18114 & n18115 ) ;
  assign n18117 = n18114 | n18116 ;
  assign n18118 = x143 | n1611 ;
  assign n18119 = ~x774 & n15591 ;
  assign n18120 = n18118 & ~n18119 ;
  assign n18121 = n16397 | n18120 ;
  assign n18122 = n16402 | n18120 ;
  assign n18123 = x1155 & n18122 ;
  assign n18124 = n16405 | n18121 ;
  assign n18125 = ~x1155 & n18124 ;
  assign n18126 = n18123 | n18125 ;
  assign n18127 = n18121 ^ x785 ^ 1'b0 ;
  assign n18128 = ( n18121 & n18126 ) | ( n18121 & n18127 ) | ( n18126 & n18127 ) ;
  assign n18129 = n16411 | n18128 ;
  assign n18130 = x1154 & n18129 ;
  assign n18131 = n16414 | n18128 ;
  assign n18132 = ~x1154 & n18131 ;
  assign n18133 = n18130 | n18132 ;
  assign n18134 = n18128 ^ x781 ^ 1'b0 ;
  assign n18135 = ( n18128 & n18133 ) | ( n18128 & n18134 ) | ( n18133 & n18134 ) ;
  assign n18136 = x619 & ~n18135 ;
  assign n18137 = x619 | n18118 ;
  assign n18138 = ( x1159 & n18136 ) | ( x1159 & n18137 ) | ( n18136 & n18137 ) ;
  assign n18139 = ~n18136 & n18138 ;
  assign n18140 = x619 & ~n18118 ;
  assign n18141 = x1159 | n18140 ;
  assign n18142 = ( n18135 & n18136 ) | ( n18135 & ~n18141 ) | ( n18136 & ~n18141 ) ;
  assign n18143 = n18139 | n18142 ;
  assign n18144 = n18135 ^ x789 ^ 1'b0 ;
  assign n18145 = ( n18135 & n18143 ) | ( n18135 & n18144 ) | ( n18143 & n18144 ) ;
  assign n18146 = x626 & ~n18145 ;
  assign n18147 = x626 & ~n18118 ;
  assign n18148 = x1158 | n18147 ;
  assign n18149 = ( n18145 & n18146 ) | ( n18145 & ~n18148 ) | ( n18146 & ~n18148 ) ;
  assign n18150 = n18146 & ~n18149 ;
  assign n18151 = ( x1158 & n18118 ) | ( x1158 & n18147 ) | ( n18118 & n18147 ) ;
  assign n18152 = ( n18149 & ~n18150 ) | ( n18149 & n18151 ) | ( ~n18150 & n18151 ) ;
  assign n18153 = n16317 & ~n18152 ;
  assign n18154 = x687 & n15778 ;
  assign n18155 = n18118 & ~n18154 ;
  assign n18156 = ~x625 & n18154 ;
  assign n18157 = ~x1153 & n18118 ;
  assign n18158 = ~n18156 & n18157 ;
  assign n18159 = ( x1153 & n18155 ) | ( x1153 & n18156 ) | ( n18155 & n18156 ) ;
  assign n18160 = n18158 | n18159 ;
  assign n18161 = n18155 ^ x778 ^ 1'b0 ;
  assign n18162 = ( n18155 & n18160 ) | ( n18155 & n18161 ) | ( n18160 & n18161 ) ;
  assign n18163 = n16447 | n18162 ;
  assign n18164 = n16449 | n18163 ;
  assign n18165 = n16451 | n18164 ;
  assign n18166 = n16459 & ~n18165 ;
  assign n18167 = ( x788 & n18153 ) | ( x788 & n18166 ) | ( n18153 & n18166 ) ;
  assign n18168 = n18166 ^ n18153 ^ 1'b0 ;
  assign n18169 = ( x788 & n18167 ) | ( x788 & n18168 ) | ( n18167 & n18168 ) ;
  assign n18170 = x619 & ~n18164 ;
  assign n18171 = x1159 | n18170 ;
  assign n18172 = n15524 | n18155 ;
  assign n18173 = n18120 & n18172 ;
  assign n18174 = x625 & ~n18172 ;
  assign n18175 = x1153 & n18120 ;
  assign n18176 = ~n18174 & n18175 ;
  assign n18177 = ( x608 & n18158 ) | ( x608 & ~n18176 ) | ( n18158 & ~n18176 ) ;
  assign n18178 = ~n18158 & n18177 ;
  assign n18179 = x608 | n18159 ;
  assign n18180 = ( n18157 & n18173 ) | ( n18157 & n18174 ) | ( n18173 & n18174 ) ;
  assign n18181 = ( ~n18178 & n18179 ) | ( ~n18178 & n18180 ) | ( n18179 & n18180 ) ;
  assign n18182 = ~n18178 & n18181 ;
  assign n18183 = n18173 ^ x778 ^ 1'b0 ;
  assign n18184 = ( n18173 & n18182 ) | ( n18173 & n18183 ) | ( n18182 & n18183 ) ;
  assign n18185 = x609 & ~n18184 ;
  assign n18186 = x609 | n18162 ;
  assign n18187 = ( x1155 & n18185 ) | ( x1155 & n18186 ) | ( n18185 & n18186 ) ;
  assign n18188 = ~n18185 & n18187 ;
  assign n18189 = ( x660 & n18125 ) | ( x660 & ~n18188 ) | ( n18125 & ~n18188 ) ;
  assign n18190 = ~n18125 & n18189 ;
  assign n18191 = x660 | n18123 ;
  assign n18192 = x609 & ~n18162 ;
  assign n18193 = x1155 | n18192 ;
  assign n18194 = ( n18184 & n18185 ) | ( n18184 & ~n18193 ) | ( n18185 & ~n18193 ) ;
  assign n18195 = ( ~n18190 & n18191 ) | ( ~n18190 & n18194 ) | ( n18191 & n18194 ) ;
  assign n18196 = ~n18190 & n18195 ;
  assign n18197 = n18184 ^ x785 ^ 1'b0 ;
  assign n18198 = ( n18184 & n18196 ) | ( n18184 & n18197 ) | ( n18196 & n18197 ) ;
  assign n18199 = x618 & ~n18198 ;
  assign n18200 = x618 | n18163 ;
  assign n18201 = ( x1154 & n18199 ) | ( x1154 & n18200 ) | ( n18199 & n18200 ) ;
  assign n18202 = ~n18199 & n18201 ;
  assign n18203 = ( x627 & n18132 ) | ( x627 & ~n18202 ) | ( n18132 & ~n18202 ) ;
  assign n18204 = ~n18132 & n18203 ;
  assign n18205 = x627 | n18130 ;
  assign n18206 = x618 & ~n18163 ;
  assign n18207 = x1154 | n18206 ;
  assign n18208 = ( n18198 & n18199 ) | ( n18198 & ~n18207 ) | ( n18199 & ~n18207 ) ;
  assign n18209 = ( ~n18204 & n18205 ) | ( ~n18204 & n18208 ) | ( n18205 & n18208 ) ;
  assign n18210 = ~n18204 & n18209 ;
  assign n18211 = n18198 ^ x781 ^ 1'b0 ;
  assign n18212 = ( n18198 & n18210 ) | ( n18198 & n18211 ) | ( n18210 & n18211 ) ;
  assign n18213 = x619 & ~n18212 ;
  assign n18214 = ( ~n18171 & n18212 ) | ( ~n18171 & n18213 ) | ( n18212 & n18213 ) ;
  assign n18215 = ( x648 & n18139 ) | ( x648 & ~n18214 ) | ( n18139 & ~n18214 ) ;
  assign n18216 = n18214 | n18215 ;
  assign n18217 = x619 | n18164 ;
  assign n18218 = ( x1159 & n18213 ) | ( x1159 & n18217 ) | ( n18213 & n18217 ) ;
  assign n18219 = ~n18213 & n18218 ;
  assign n18220 = ( x648 & n18142 ) | ( x648 & ~n18219 ) | ( n18142 & ~n18219 ) ;
  assign n18221 = ~n18142 & n18220 ;
  assign n18222 = x789 & ~n18221 ;
  assign n18223 = n18216 & n18222 ;
  assign n18224 = ~x789 & n18212 ;
  assign n18225 = n16519 | n18224 ;
  assign n18226 = ( ~n18169 & n18223 ) | ( ~n18169 & n18225 ) | ( n18223 & n18225 ) ;
  assign n18227 = ~n18169 & n18226 ;
  assign n18228 = x628 & ~n18227 ;
  assign n18229 = n18145 ^ x788 ^ 1'b0 ;
  assign n18230 = ( n18145 & n18152 ) | ( n18145 & n18229 ) | ( n18152 & n18229 ) ;
  assign n18231 = x628 | n18230 ;
  assign n18232 = ( x1156 & n18228 ) | ( x1156 & n18231 ) | ( n18228 & n18231 ) ;
  assign n18233 = ~n18228 & n18232 ;
  assign n18234 = n16530 | n18165 ;
  assign n18235 = n16532 | n18234 ;
  assign n18236 = ~x1156 & n18235 ;
  assign n18237 = ( x629 & n18233 ) | ( x629 & ~n18236 ) | ( n18233 & ~n18236 ) ;
  assign n18238 = ~n18233 & n18237 ;
  assign n18239 = n16537 | n18234 ;
  assign n18240 = ( x1156 & ~n17240 ) | ( x1156 & n18239 ) | ( ~n17240 & n18239 ) ;
  assign n18241 = ( x629 & n17240 ) | ( x629 & n18240 ) | ( n17240 & n18240 ) ;
  assign n18242 = x628 & ~n18230 ;
  assign n18243 = x1156 | n18242 ;
  assign n18244 = ( n18227 & n18228 ) | ( n18227 & ~n18243 ) | ( n18228 & ~n18243 ) ;
  assign n18245 = ( ~n18238 & n18241 ) | ( ~n18238 & n18244 ) | ( n18241 & n18244 ) ;
  assign n18246 = ~n18238 & n18245 ;
  assign n18247 = n18227 ^ x792 ^ 1'b0 ;
  assign n18248 = ( n18227 & n18246 ) | ( n18227 & n18247 ) | ( n18246 & n18247 ) ;
  assign n18249 = x647 & ~n18248 ;
  assign n18250 = n18118 ^ n16339 ^ 1'b0 ;
  assign n18251 = ( n18118 & n18230 ) | ( n18118 & ~n18250 ) | ( n18230 & ~n18250 ) ;
  assign n18252 = x647 | n18251 ;
  assign n18253 = ( x1157 & n18249 ) | ( x1157 & n18252 ) | ( n18249 & n18252 ) ;
  assign n18254 = ~n18249 & n18253 ;
  assign n18255 = x647 & ~n18118 ;
  assign n18256 = x1157 | n18255 ;
  assign n18257 = n16560 | n18234 ;
  assign n18258 = x647 & ~n18257 ;
  assign n18259 = ( ~n18256 & n18257 ) | ( ~n18256 & n18258 ) | ( n18257 & n18258 ) ;
  assign n18260 = ( x630 & n18254 ) | ( x630 & ~n18259 ) | ( n18254 & ~n18259 ) ;
  assign n18261 = ~n18254 & n18260 ;
  assign n18262 = x647 | n18118 ;
  assign n18263 = ( x1157 & n18258 ) | ( x1157 & n18262 ) | ( n18258 & n18262 ) ;
  assign n18264 = ~n18258 & n18263 ;
  assign n18265 = x630 | n18264 ;
  assign n18266 = x647 & ~n18251 ;
  assign n18267 = x1157 | n18266 ;
  assign n18268 = ( n18248 & n18249 ) | ( n18248 & ~n18267 ) | ( n18249 & ~n18267 ) ;
  assign n18269 = ( ~n18261 & n18265 ) | ( ~n18261 & n18268 ) | ( n18265 & n18268 ) ;
  assign n18270 = ~n18261 & n18269 ;
  assign n18271 = n18248 ^ x787 ^ 1'b0 ;
  assign n18272 = ( n18248 & n18270 ) | ( n18248 & n18271 ) | ( n18270 & n18271 ) ;
  assign n18273 = x644 & ~n18272 ;
  assign n18274 = n18259 | n18264 ;
  assign n18275 = n18257 ^ x787 ^ 1'b0 ;
  assign n18276 = ( n18257 & n18274 ) | ( n18257 & n18275 ) | ( n18274 & n18275 ) ;
  assign n18277 = x644 | n18276 ;
  assign n18278 = ( x715 & n18273 ) | ( x715 & n18277 ) | ( n18273 & n18277 ) ;
  assign n18279 = ~n18273 & n18278 ;
  assign n18280 = n18118 ^ n16376 ^ 1'b0 ;
  assign n18281 = ( n18118 & n18251 ) | ( n18118 & ~n18280 ) | ( n18251 & ~n18280 ) ;
  assign n18282 = x644 & ~n18281 ;
  assign n18283 = x644 | n18118 ;
  assign n18284 = ( x715 & ~n18282 ) | ( x715 & n18283 ) | ( ~n18282 & n18283 ) ;
  assign n18285 = ~x715 & n18284 ;
  assign n18286 = ( x1160 & n18279 ) | ( x1160 & ~n18285 ) | ( n18279 & ~n18285 ) ;
  assign n18287 = ~n18279 & n18286 ;
  assign n18288 = x644 & ~n18118 ;
  assign n18289 = x644 | n18281 ;
  assign n18290 = ( x715 & n18288 ) | ( x715 & n18289 ) | ( n18288 & n18289 ) ;
  assign n18291 = ~n18288 & n18290 ;
  assign n18292 = x644 & ~n18276 ;
  assign n18293 = x715 | n18292 ;
  assign n18294 = ( n18272 & n18273 ) | ( n18272 & ~n18293 ) | ( n18273 & ~n18293 ) ;
  assign n18295 = ( x1160 & ~n18291 ) | ( x1160 & n18294 ) | ( ~n18291 & n18294 ) ;
  assign n18296 = n18291 | n18295 ;
  assign n18297 = x790 & ~n18296 ;
  assign n18298 = ( x790 & n18287 ) | ( x790 & n18297 ) | ( n18287 & n18297 ) ;
  assign n18299 = x790 | n18272 ;
  assign n18300 = ( x832 & n18298 ) | ( x832 & n18299 ) | ( n18298 & n18299 ) ;
  assign n18301 = ~n18298 & n18300 ;
  assign n18302 = ~x143 & n7318 ;
  assign n18303 = x832 | n18302 ;
  assign n18304 = ~n18301 & n18303 ;
  assign n18305 = ( n18117 & n18301 ) | ( n18117 & ~n18304 ) | ( n18301 & ~n18304 ) ;
  assign n18326 = x144 & ~n1611 ;
  assign n18327 = x736 & n15778 ;
  assign n18328 = n18326 | n18327 ;
  assign n18329 = x625 & n18327 ;
  assign n18330 = n18329 ^ n18327 ^ n18326 ;
  assign n18331 = x1153 | n18330 ;
  assign n18332 = x1153 & ~n18326 ;
  assign n18333 = ~n18329 & n18332 ;
  assign n18334 = n18331 & ~n18333 ;
  assign n18335 = n18328 ^ x778 ^ 1'b0 ;
  assign n18336 = ( n18328 & n18334 ) | ( n18328 & n18335 ) | ( n18334 & n18335 ) ;
  assign n18337 = ~n17088 & n18336 ;
  assign n18338 = ~n17093 & n18337 ;
  assign n18339 = x630 & ~n18338 ;
  assign n18340 = ( x647 & n18338 ) | ( x647 & n18339 ) | ( n18338 & n18339 ) ;
  assign n18306 = x609 & x1155 ;
  assign n18307 = x609 | x1155 ;
  assign n18308 = x785 & n18307 ;
  assign n18309 = ~n18306 & n18308 ;
  assign n18310 = x758 & n15591 ;
  assign n18311 = ~n18309 & n18310 ;
  assign n18312 = x618 & x1154 ;
  assign n18313 = x618 | x1154 ;
  assign n18314 = x781 & n18313 ;
  assign n18315 = ~n18312 & n18314 ;
  assign n18316 = ~x619 & x1159 ;
  assign n18317 = x619 & ~x1159 ;
  assign n18318 = n18316 | n18317 ;
  assign n18319 = x789 & n18318 ;
  assign n18320 = n15659 | n18319 ;
  assign n18321 = n18315 | n18320 ;
  assign n18322 = n18311 & ~n18321 ;
  assign n18323 = ~n16518 & n18322 ;
  assign n18324 = ~n16339 & n18323 ;
  assign n18325 = x630 & n18324 ;
  assign n18341 = ( x1157 & ~n18325 ) | ( x1157 & n18340 ) | ( ~n18325 & n18340 ) ;
  assign n18342 = ~n18340 & n18341 ;
  assign n18343 = ~x630 & n18324 ;
  assign n18344 = ~n18339 & n18343 ;
  assign n18345 = ( x647 & n18339 ) | ( x647 & ~n18344 ) | ( n18339 & ~n18344 ) ;
  assign n18346 = ( ~x1157 & n18342 ) | ( ~x1157 & n18345 ) | ( n18342 & n18345 ) ;
  assign n18347 = n18342 ^ x1157 ^ 1'b0 ;
  assign n18348 = ( n18342 & n18346 ) | ( n18342 & ~n18347 ) | ( n18346 & ~n18347 ) ;
  assign n18349 = x787 & ~n18326 ;
  assign n18350 = n18348 & n18349 ;
  assign n18351 = ~x626 & n18322 ;
  assign n18352 = n18326 | n18351 ;
  assign n18353 = ( x641 & x1158 ) | ( x641 & ~n18352 ) | ( x1158 & ~n18352 ) ;
  assign n18354 = ( x641 & ~n16317 ) | ( x641 & n18353 ) | ( ~n16317 & n18353 ) ;
  assign n18355 = n16279 & ~n18326 ;
  assign n18356 = ~n16234 & n18336 ;
  assign n18357 = ~n16254 & n18356 ;
  assign n18358 = n18326 | n18357 ;
  assign n18359 = ~n18355 & n18358 ;
  assign n18360 = ( n16453 & ~n18354 ) | ( n16453 & n18359 ) | ( ~n18354 & n18359 ) ;
  assign n18361 = n18360 ^ n18354 ^ 1'b0 ;
  assign n18362 = ( n18354 & ~n18360 ) | ( n18354 & n18361 ) | ( ~n18360 & n18361 ) ;
  assign n18363 = x626 & n18322 ;
  assign n18364 = n18326 | n18363 ;
  assign n18365 = ( x1158 & ~n16317 ) | ( x1158 & n18364 ) | ( ~n16317 & n18364 ) ;
  assign n18366 = ( x641 & n16317 ) | ( x641 & n18365 ) | ( n16317 & n18365 ) ;
  assign n18367 = n18366 ^ n16454 ^ 1'b0 ;
  assign n18368 = ( ~n16454 & n18359 ) | ( ~n16454 & n18367 ) | ( n18359 & n18367 ) ;
  assign n18369 = ( n16454 & n18366 ) | ( n16454 & n18368 ) | ( n18366 & n18368 ) ;
  assign n18370 = ( x788 & n18362 ) | ( x788 & n18369 ) | ( n18362 & n18369 ) ;
  assign n18371 = ~n18362 & n18370 ;
  assign n18372 = x1159 | n18326 ;
  assign n18373 = n18311 & ~n18315 ;
  assign n18374 = x619 | n15659 ;
  assign n18375 = n18373 & ~n18374 ;
  assign n18376 = n18372 | n18375 ;
  assign n18377 = x1154 | n18326 ;
  assign n18378 = x618 | n15659 ;
  assign n18379 = n18311 & ~n18378 ;
  assign n18380 = n18377 | n18379 ;
  assign n18381 = n18326 | n18356 ;
  assign n18382 = ~x618 & n18381 ;
  assign n18383 = x608 | n18333 ;
  assign n18384 = n18310 | n18326 ;
  assign n18385 = x736 & n17156 ;
  assign n18386 = n18384 | n18385 ;
  assign n18387 = x625 & n18385 ;
  assign n18388 = n18386 & ~n18387 ;
  assign n18389 = ( x1153 & ~n18383 ) | ( x1153 & n18388 ) | ( ~n18383 & n18388 ) ;
  assign n18390 = ~n18383 & n18389 ;
  assign n18391 = x1153 & ~n18384 ;
  assign n18392 = ~n18387 & n18391 ;
  assign n18393 = ( x608 & n18331 ) | ( x608 & n18392 ) | ( n18331 & n18392 ) ;
  assign n18394 = ~n18392 & n18393 ;
  assign n18395 = ( x778 & n18390 ) | ( x778 & ~n18394 ) | ( n18390 & ~n18394 ) ;
  assign n18396 = ~n18390 & n18395 ;
  assign n18397 = ( x778 & n18386 ) | ( x778 & ~n18396 ) | ( n18386 & ~n18396 ) ;
  assign n18398 = ~n18396 & n18397 ;
  assign n18399 = ~x609 & n18398 ;
  assign n18400 = x609 & n18336 ;
  assign n18401 = ( x1155 & ~n18399 ) | ( x1155 & n18400 ) | ( ~n18399 & n18400 ) ;
  assign n18402 = n18399 | n18401 ;
  assign n18403 = x1155 | n18326 ;
  assign n18404 = ~n15662 & n18310 ;
  assign n18405 = n18403 | n18404 ;
  assign n18406 = ~x609 & n18336 ;
  assign n18407 = x609 & n18398 ;
  assign n18408 = ( x1155 & n18406 ) | ( x1155 & ~n18407 ) | ( n18406 & ~n18407 ) ;
  assign n18409 = ~n18406 & n18408 ;
  assign n18410 = x660 & ~n18409 ;
  assign n18411 = n18405 & n18410 ;
  assign n18412 = x1155 & ~n18326 ;
  assign n18413 = n15668 & n18310 ;
  assign n18414 = ( x660 & n18412 ) | ( x660 & ~n18413 ) | ( n18412 & ~n18413 ) ;
  assign n18415 = n18414 ^ n18412 ^ 1'b0 ;
  assign n18416 = ( x660 & n18414 ) | ( x660 & ~n18415 ) | ( n18414 & ~n18415 ) ;
  assign n18417 = ~n18411 & n18416 ;
  assign n18418 = ( n18402 & n18411 ) | ( n18402 & ~n18417 ) | ( n18411 & ~n18417 ) ;
  assign n18419 = n18398 ^ x785 ^ 1'b0 ;
  assign n18420 = ( n18398 & n18418 ) | ( n18398 & n18419 ) | ( n18418 & n18419 ) ;
  assign n18421 = x618 & n18420 ;
  assign n18422 = ( x1154 & n18382 ) | ( x1154 & ~n18421 ) | ( n18382 & ~n18421 ) ;
  assign n18423 = ~n18382 & n18422 ;
  assign n18424 = x627 & ~n18423 ;
  assign n18425 = n18380 & n18424 ;
  assign n18426 = ~x618 & n18420 ;
  assign n18427 = x618 & n18381 ;
  assign n18428 = ( x1154 & ~n18426 ) | ( x1154 & n18427 ) | ( ~n18426 & n18427 ) ;
  assign n18429 = n18426 | n18428 ;
  assign n18430 = x1154 & ~n18326 ;
  assign n18431 = x618 & ~n15659 ;
  assign n18432 = n18311 & n18431 ;
  assign n18433 = n18430 & ~n18432 ;
  assign n18434 = ( x627 & n18429 ) | ( x627 & ~n18433 ) | ( n18429 & ~n18433 ) ;
  assign n18435 = ~x627 & n18434 ;
  assign n18436 = ( x781 & n18425 ) | ( x781 & ~n18435 ) | ( n18425 & ~n18435 ) ;
  assign n18437 = ~n18425 & n18436 ;
  assign n18438 = ( x781 & n18420 ) | ( x781 & ~n18437 ) | ( n18420 & ~n18437 ) ;
  assign n18439 = ~n18437 & n18438 ;
  assign n18440 = x619 & n18439 ;
  assign n18441 = ~x619 & n18358 ;
  assign n18442 = ( x1159 & n18440 ) | ( x1159 & ~n18441 ) | ( n18440 & ~n18441 ) ;
  assign n18443 = ~n18440 & n18442 ;
  assign n18444 = x648 & ~n18443 ;
  assign n18445 = n18376 & n18444 ;
  assign n18446 = ~x619 & n18439 ;
  assign n18447 = x619 & n18358 ;
  assign n18448 = ( x1159 & ~n18446 ) | ( x1159 & n18447 ) | ( ~n18446 & n18447 ) ;
  assign n18449 = n18446 | n18448 ;
  assign n18450 = x1159 & ~n18326 ;
  assign n18451 = x619 & ~n15659 ;
  assign n18452 = n18373 & n18451 ;
  assign n18453 = n18450 & ~n18452 ;
  assign n18454 = ( x648 & n18449 ) | ( x648 & ~n18453 ) | ( n18449 & ~n18453 ) ;
  assign n18455 = ~x648 & n18454 ;
  assign n18456 = ( x789 & n18445 ) | ( x789 & ~n18455 ) | ( n18445 & ~n18455 ) ;
  assign n18457 = ~n18445 & n18456 ;
  assign n18458 = x789 | n18439 ;
  assign n18459 = ~n16519 & n18458 ;
  assign n18460 = n18459 ^ n18457 ^ 1'b0 ;
  assign n18461 = ( n18457 & n18459 ) | ( n18457 & n18460 ) | ( n18459 & n18460 ) ;
  assign n18462 = ( n18371 & ~n18457 ) | ( n18371 & n18461 ) | ( ~n18457 & n18461 ) ;
  assign n18463 = ~x628 & n18337 ;
  assign n18464 = x629 & ~n18463 ;
  assign n18465 = x628 & ~n18323 ;
  assign n18466 = ( ~x1156 & n18464 ) | ( ~x1156 & n18465 ) | ( n18464 & n18465 ) ;
  assign n18467 = ~x1156 & n18466 ;
  assign n18468 = x628 | n18323 ;
  assign n18469 = ( x629 & ~x1156 ) | ( x629 & n18468 ) | ( ~x1156 & n18468 ) ;
  assign n18470 = ( x1156 & n17240 ) | ( x1156 & ~n18469 ) | ( n17240 & ~n18469 ) ;
  assign n18471 = ( x628 & n18337 ) | ( x628 & ~n18470 ) | ( n18337 & ~n18470 ) ;
  assign n18472 = n18471 ^ n18470 ^ 1'b0 ;
  assign n18473 = ( n18470 & ~n18471 ) | ( n18470 & n18472 ) | ( ~n18471 & n18472 ) ;
  assign n18474 = ( ~n18326 & n18467 ) | ( ~n18326 & n18473 ) | ( n18467 & n18473 ) ;
  assign n18475 = ~n18326 & n18474 ;
  assign n18476 = ( x792 & ~n18462 ) | ( x792 & n18475 ) | ( ~n18462 & n18475 ) ;
  assign n18477 = n18476 ^ n18462 ^ 1'b0 ;
  assign n18478 = ( n18462 & ~n18476 ) | ( n18462 & n18477 ) | ( ~n18476 & n18477 ) ;
  assign n18479 = x629 & n17091 ;
  assign n18480 = x792 & ~n18479 ;
  assign n18481 = x629 | n17090 ;
  assign n18482 = n18480 & n18481 ;
  assign n18483 = ~n18475 & n18482 ;
  assign n18484 = ( x787 & n16376 ) | ( x787 & n17273 ) | ( n16376 & n17273 ) ;
  assign n18485 = n18483 | n18484 ;
  assign n18486 = ( ~n18350 & n18478 ) | ( ~n18350 & n18485 ) | ( n18478 & n18485 ) ;
  assign n18487 = ~n18350 & n18486 ;
  assign n18488 = ~x790 & n18487 ;
  assign n18489 = ~x644 & n18487 ;
  assign n18490 = ~n17273 & n18338 ;
  assign n18491 = n18326 | n18490 ;
  assign n18492 = x644 & n18491 ;
  assign n18493 = ( x715 & ~n18489 ) | ( x715 & n18492 ) | ( ~n18489 & n18492 ) ;
  assign n18494 = n18489 | n18493 ;
  assign n18495 = x715 & ~n18326 ;
  assign n18496 = ~n16376 & n18324 ;
  assign n18497 = ~x644 & n18496 ;
  assign n18498 = n18495 & ~n18497 ;
  assign n18499 = ( x1160 & n18494 ) | ( x1160 & ~n18498 ) | ( n18494 & ~n18498 ) ;
  assign n18500 = ~x1160 & n18499 ;
  assign n18501 = x715 | n18326 ;
  assign n18502 = x644 & n18496 ;
  assign n18503 = n18501 | n18502 ;
  assign n18504 = ~x644 & n18491 ;
  assign n18505 = x644 & n18487 ;
  assign n18506 = ( x715 & n18504 ) | ( x715 & ~n18505 ) | ( n18504 & ~n18505 ) ;
  assign n18507 = ~n18504 & n18506 ;
  assign n18508 = x1160 & ~n18507 ;
  assign n18509 = n18503 & n18508 ;
  assign n18510 = ( x790 & n18500 ) | ( x790 & n18509 ) | ( n18500 & n18509 ) ;
  assign n18511 = n18509 ^ n18500 ^ 1'b0 ;
  assign n18512 = ( x790 & n18510 ) | ( x790 & n18511 ) | ( n18510 & n18511 ) ;
  assign n18513 = ( x832 & n18488 ) | ( x832 & ~n18512 ) | ( n18488 & ~n18512 ) ;
  assign n18514 = ~n18488 & n18513 ;
  assign n18515 = ~x144 & n5193 ;
  assign n18516 = x144 & ~n15656 ;
  assign n18517 = x144 | n16699 ;
  assign n18518 = x144 & n16697 ;
  assign n18519 = ( x38 & n18517 ) | ( x38 & ~n18518 ) | ( n18517 & ~n18518 ) ;
  assign n18520 = ~x38 & n18519 ;
  assign n18521 = x736 & ~n2069 ;
  assign n18522 = x144 | n15644 ;
  assign n18523 = n15644 & ~n15777 ;
  assign n18524 = x38 & ~n18523 ;
  assign n18525 = n18522 & n18524 ;
  assign n18526 = ( n18520 & n18521 ) | ( n18520 & ~n18525 ) | ( n18521 & ~n18525 ) ;
  assign n18527 = ~n18520 & n18526 ;
  assign n18528 = ( n18516 & n18521 ) | ( n18516 & ~n18527 ) | ( n18521 & ~n18527 ) ;
  assign n18529 = ~n18527 & n18528 ;
  assign n18530 = x625 & ~n18529 ;
  assign n18531 = x625 | n18516 ;
  assign n18532 = ( x1153 & n18530 ) | ( x1153 & n18531 ) | ( n18530 & n18531 ) ;
  assign n18533 = ~n18530 & n18532 ;
  assign n18534 = x625 & ~n18516 ;
  assign n18535 = x1153 | n18534 ;
  assign n18536 = ( x625 & n18529 ) | ( x625 & ~n18535 ) | ( n18529 & ~n18535 ) ;
  assign n18537 = ~n18535 & n18536 ;
  assign n18538 = n18533 | n18537 ;
  assign n18539 = n18529 ^ x778 ^ 1'b0 ;
  assign n18540 = ( n18529 & n18538 ) | ( n18529 & n18539 ) | ( n18538 & n18539 ) ;
  assign n18541 = n18516 ^ n16234 ^ 1'b0 ;
  assign n18542 = ( n18516 & n18540 ) | ( n18516 & ~n18541 ) | ( n18540 & ~n18541 ) ;
  assign n18543 = n18516 ^ n16254 ^ 1'b0 ;
  assign n18544 = ( n18516 & n18542 ) | ( n18516 & ~n18543 ) | ( n18542 & ~n18543 ) ;
  assign n18545 = n18516 ^ n16279 ^ 1'b0 ;
  assign n18546 = ( n18516 & n18544 ) | ( n18516 & ~n18545 ) | ( n18544 & ~n18545 ) ;
  assign n18563 = ~x626 & n18546 ;
  assign n18565 = x758 & n15524 ;
  assign n18566 = n15644 & ~n18565 ;
  assign n18567 = x38 & ~n18566 ;
  assign n18568 = n18522 & n18567 ;
  assign n18614 = x144 & n16048 ;
  assign n18615 = x144 | n16054 ;
  assign n18616 = ( x758 & n18614 ) | ( x758 & n18615 ) | ( n18614 & n18615 ) ;
  assign n18617 = ~n18614 & n18616 ;
  assign n18618 = x144 | n16029 ;
  assign n18619 = x144 & n16044 ;
  assign n18620 = ( x758 & n18618 ) | ( x758 & ~n18619 ) | ( n18618 & ~n18619 ) ;
  assign n18621 = ~x758 & n18620 ;
  assign n18622 = ( x39 & ~n18617 ) | ( x39 & n18621 ) | ( ~n18617 & n18621 ) ;
  assign n18623 = n18617 | n18622 ;
  assign n18624 = x144 | n15795 ;
  assign n18625 = x144 & n15876 ;
  assign n18626 = ( x758 & n18624 ) | ( x758 & ~n18625 ) | ( n18624 & ~n18625 ) ;
  assign n18627 = ~x758 & n18626 ;
  assign n18628 = x144 & n16003 ;
  assign n18629 = x144 | n15943 ;
  assign n18630 = ( x758 & n18628 ) | ( x758 & n18629 ) | ( n18628 & n18629 ) ;
  assign n18631 = ~n18628 & n18630 ;
  assign n18632 = ( x39 & n18627 ) | ( x39 & ~n18631 ) | ( n18627 & ~n18631 ) ;
  assign n18633 = ~n18627 & n18632 ;
  assign n18634 = ( x38 & n18623 ) | ( x38 & ~n18633 ) | ( n18623 & ~n18633 ) ;
  assign n18635 = ~x38 & n18634 ;
  assign n18636 = x736 & ~n17882 ;
  assign n18637 = ( n18568 & ~n18635 ) | ( n18568 & n18636 ) | ( ~n18635 & n18636 ) ;
  assign n18638 = ~n18568 & n18637 ;
  assign n18639 = ( n2051 & n2068 ) | ( n2051 & ~n18638 ) | ( n2068 & ~n18638 ) ;
  assign n18640 = n18638 | n18639 ;
  assign n18569 = ~x144 & x758 ;
  assign n18570 = n15640 & n18569 ;
  assign n18571 = ~x758 & n15332 ;
  assign n18572 = x758 & n15509 ;
  assign n18573 = ( x39 & ~n18571 ) | ( x39 & n18572 ) | ( ~n18571 & n18572 ) ;
  assign n18574 = n18571 | n18573 ;
  assign n18575 = x758 & ~n15585 ;
  assign n18576 = x758 | n15486 ;
  assign n18577 = ~n18575 & n18576 ;
  assign n18578 = n18577 ^ n18574 ^ 1'b0 ;
  assign n18579 = ( ~x39 & n18577 ) | ( ~x39 & n18578 ) | ( n18577 & n18578 ) ;
  assign n18580 = ( n18574 & ~n18578 ) | ( n18574 & n18579 ) | ( ~n18578 & n18579 ) ;
  assign n18581 = ~n18570 & n18580 ;
  assign n18582 = ( x144 & n18570 ) | ( x144 & ~n18581 ) | ( n18570 & ~n18581 ) ;
  assign n18583 = ( ~x38 & n18568 ) | ( ~x38 & n18582 ) | ( n18568 & n18582 ) ;
  assign n18584 = n18568 ^ x38 ^ 1'b0 ;
  assign n18585 = ( n18568 & n18583 ) | ( n18568 & ~n18584 ) | ( n18583 & ~n18584 ) ;
  assign n18641 = ( x736 & n18585 ) | ( x736 & ~n18640 ) | ( n18585 & ~n18640 ) ;
  assign n18642 = ~n18640 & n18641 ;
  assign n18643 = n18642 ^ x144 ^ 1'b0 ;
  assign n18644 = ( ~x144 & n2069 ) | ( ~x144 & n18643 ) | ( n2069 & n18643 ) ;
  assign n18645 = ( x144 & n18642 ) | ( x144 & n18644 ) | ( n18642 & n18644 ) ;
  assign n18646 = x625 & ~n18645 ;
  assign n18564 = x144 & n2069 ;
  assign n18586 = ~n2069 & n18585 ;
  assign n18587 = n18564 | n18586 ;
  assign n18652 = x625 | n18587 ;
  assign n18653 = ( x1153 & n18646 ) | ( x1153 & n18652 ) | ( n18646 & n18652 ) ;
  assign n18654 = ~n18646 & n18653 ;
  assign n18655 = ( x608 & ~n18537 ) | ( x608 & n18654 ) | ( ~n18537 & n18654 ) ;
  assign n18656 = ~n18654 & n18655 ;
  assign n18647 = x625 & ~n18587 ;
  assign n18648 = x1153 | n18647 ;
  assign n18649 = ( n18645 & n18646 ) | ( n18645 & ~n18648 ) | ( n18646 & ~n18648 ) ;
  assign n18650 = ( x608 & ~n18533 ) | ( x608 & n18649 ) | ( ~n18533 & n18649 ) ;
  assign n18651 = n18533 | n18650 ;
  assign n18657 = n18656 ^ n18651 ^ 1'b0 ;
  assign n18658 = ( x778 & ~n18651 ) | ( x778 & n18656 ) | ( ~n18651 & n18656 ) ;
  assign n18659 = ( x778 & ~n18657 ) | ( x778 & n18658 ) | ( ~n18657 & n18658 ) ;
  assign n18660 = ( x778 & n18645 ) | ( x778 & ~n18659 ) | ( n18645 & ~n18659 ) ;
  assign n18661 = ~n18659 & n18660 ;
  assign n18662 = x609 & ~n18661 ;
  assign n18668 = x609 | n18540 ;
  assign n18669 = ( x1155 & n18662 ) | ( x1155 & n18668 ) | ( n18662 & n18668 ) ;
  assign n18670 = ~n18662 & n18669 ;
  assign n18588 = n18587 ^ n15659 ^ 1'b0 ;
  assign n18589 = ( n18516 & n18587 ) | ( n18516 & n18588 ) | ( n18587 & n18588 ) ;
  assign n18590 = x609 & ~n18589 ;
  assign n18594 = x609 & ~n18516 ;
  assign n18595 = x1155 | n18594 ;
  assign n18596 = ( n18589 & n18590 ) | ( n18589 & ~n18595 ) | ( n18590 & ~n18595 ) ;
  assign n18671 = ( x660 & ~n18596 ) | ( x660 & n18670 ) | ( ~n18596 & n18670 ) ;
  assign n18672 = ~n18670 & n18671 ;
  assign n18591 = x609 | n18516 ;
  assign n18592 = ( x1155 & n18590 ) | ( x1155 & n18591 ) | ( n18590 & n18591 ) ;
  assign n18593 = ~n18590 & n18592 ;
  assign n18663 = x609 & ~n18540 ;
  assign n18664 = x1155 | n18663 ;
  assign n18665 = ( n18661 & n18662 ) | ( n18661 & ~n18664 ) | ( n18662 & ~n18664 ) ;
  assign n18666 = ( x660 & ~n18593 ) | ( x660 & n18665 ) | ( ~n18593 & n18665 ) ;
  assign n18667 = n18593 | n18666 ;
  assign n18673 = n18672 ^ n18667 ^ 1'b0 ;
  assign n18674 = ( x785 & ~n18667 ) | ( x785 & n18672 ) | ( ~n18667 & n18672 ) ;
  assign n18675 = ( x785 & ~n18673 ) | ( x785 & n18674 ) | ( ~n18673 & n18674 ) ;
  assign n18676 = ( x785 & n18661 ) | ( x785 & ~n18675 ) | ( n18661 & ~n18675 ) ;
  assign n18677 = ~n18675 & n18676 ;
  assign n18678 = x618 & ~n18677 ;
  assign n18684 = x618 | n18542 ;
  assign n18685 = ( x1154 & n18678 ) | ( x1154 & n18684 ) | ( n18678 & n18684 ) ;
  assign n18686 = ~n18678 & n18685 ;
  assign n18597 = n18593 | n18596 ;
  assign n18598 = n18589 ^ x785 ^ 1'b0 ;
  assign n18599 = ( n18589 & n18597 ) | ( n18589 & n18598 ) | ( n18597 & n18598 ) ;
  assign n18600 = x618 & ~n18599 ;
  assign n18604 = x618 & ~n18516 ;
  assign n18605 = x1154 | n18604 ;
  assign n18606 = ( n18599 & n18600 ) | ( n18599 & ~n18605 ) | ( n18600 & ~n18605 ) ;
  assign n18687 = ( x627 & ~n18606 ) | ( x627 & n18686 ) | ( ~n18606 & n18686 ) ;
  assign n18688 = ~n18686 & n18687 ;
  assign n18601 = x618 | n18516 ;
  assign n18602 = ( x1154 & n18600 ) | ( x1154 & n18601 ) | ( n18600 & n18601 ) ;
  assign n18603 = ~n18600 & n18602 ;
  assign n18679 = x618 & ~n18542 ;
  assign n18680 = x1154 | n18679 ;
  assign n18681 = ( n18677 & n18678 ) | ( n18677 & ~n18680 ) | ( n18678 & ~n18680 ) ;
  assign n18682 = ( x627 & ~n18603 ) | ( x627 & n18681 ) | ( ~n18603 & n18681 ) ;
  assign n18683 = n18603 | n18682 ;
  assign n18689 = n18688 ^ n18683 ^ 1'b0 ;
  assign n18690 = ( x781 & ~n18683 ) | ( x781 & n18688 ) | ( ~n18683 & n18688 ) ;
  assign n18691 = ( x781 & ~n18689 ) | ( x781 & n18690 ) | ( ~n18689 & n18690 ) ;
  assign n18692 = ( x781 & n18677 ) | ( x781 & ~n18691 ) | ( n18677 & ~n18691 ) ;
  assign n18693 = ~n18691 & n18692 ;
  assign n18694 = x619 & ~n18693 ;
  assign n18700 = x619 | n18544 ;
  assign n18701 = ( x1159 & n18694 ) | ( x1159 & n18700 ) | ( n18694 & n18700 ) ;
  assign n18702 = ~n18694 & n18701 ;
  assign n18607 = n18603 | n18606 ;
  assign n18608 = n18599 ^ x781 ^ 1'b0 ;
  assign n18609 = ( n18599 & n18607 ) | ( n18599 & n18608 ) | ( n18607 & n18608 ) ;
  assign n18610 = x619 & ~n18609 ;
  assign n18703 = x619 & ~n18516 ;
  assign n18704 = x1159 | n18703 ;
  assign n18705 = ( n18609 & n18610 ) | ( n18609 & ~n18704 ) | ( n18610 & ~n18704 ) ;
  assign n18706 = ( x648 & n18702 ) | ( x648 & ~n18705 ) | ( n18702 & ~n18705 ) ;
  assign n18707 = ~n18702 & n18706 ;
  assign n18611 = x619 | n18516 ;
  assign n18612 = ( x1159 & n18610 ) | ( x1159 & n18611 ) | ( n18610 & n18611 ) ;
  assign n18613 = ~n18610 & n18612 ;
  assign n18695 = x619 & ~n18544 ;
  assign n18696 = x1159 | n18695 ;
  assign n18697 = ( n18693 & n18694 ) | ( n18693 & ~n18696 ) | ( n18694 & ~n18696 ) ;
  assign n18698 = ( x648 & ~n18613 ) | ( x648 & n18697 ) | ( ~n18613 & n18697 ) ;
  assign n18699 = n18613 | n18698 ;
  assign n18708 = n18707 ^ n18699 ^ 1'b0 ;
  assign n18709 = ( x789 & ~n18699 ) | ( x789 & n18707 ) | ( ~n18699 & n18707 ) ;
  assign n18710 = ( x789 & ~n18708 ) | ( x789 & n18709 ) | ( ~n18708 & n18709 ) ;
  assign n18711 = ( x789 & n18693 ) | ( x789 & ~n18710 ) | ( n18693 & ~n18710 ) ;
  assign n18712 = ~n18710 & n18711 ;
  assign n18713 = x626 & n18712 ;
  assign n18714 = ( x641 & n18563 ) | ( x641 & ~n18713 ) | ( n18563 & ~n18713 ) ;
  assign n18715 = ~n18563 & n18714 ;
  assign n18716 = n18613 | n18705 ;
  assign n18717 = n18609 ^ x789 ^ 1'b0 ;
  assign n18718 = ( n18609 & n18716 ) | ( n18609 & n18717 ) | ( n18716 & n18717 ) ;
  assign n18719 = x626 & ~n18718 ;
  assign n18720 = x626 | n18516 ;
  assign n18721 = ( x1158 & n18719 ) | ( x1158 & n18720 ) | ( n18719 & n18720 ) ;
  assign n18722 = ~n18719 & n18721 ;
  assign n18723 = n16289 | n18722 ;
  assign n18724 = ~n18715 & n18723 ;
  assign n18725 = ~x626 & n18712 ;
  assign n18726 = x626 & n18546 ;
  assign n18727 = ( x641 & ~n18725 ) | ( x641 & n18726 ) | ( ~n18725 & n18726 ) ;
  assign n18728 = n18725 | n18727 ;
  assign n18729 = x626 & ~n18516 ;
  assign n18730 = x1158 | n18729 ;
  assign n18731 = ( n18718 & n18719 ) | ( n18718 & ~n18730 ) | ( n18719 & ~n18730 ) ;
  assign n18732 = ( ~n16299 & n18728 ) | ( ~n16299 & n18731 ) | ( n18728 & n18731 ) ;
  assign n18733 = n18728 ^ n16299 ^ 1'b0 ;
  assign n18734 = ( n18728 & n18732 ) | ( n18728 & n18733 ) | ( n18732 & n18733 ) ;
  assign n18735 = ( x788 & n18724 ) | ( x788 & ~n18734 ) | ( n18724 & ~n18734 ) ;
  assign n18736 = ~n18724 & n18735 ;
  assign n18737 = ( x788 & n18712 ) | ( x788 & ~n18736 ) | ( n18712 & ~n18736 ) ;
  assign n18738 = ~n18736 & n18737 ;
  assign n18739 = x628 & ~n18738 ;
  assign n18740 = n18722 | n18731 ;
  assign n18741 = n18718 ^ x788 ^ 1'b0 ;
  assign n18742 = ( n18718 & n18740 ) | ( n18718 & n18741 ) | ( n18740 & n18741 ) ;
  assign n18748 = x628 | n18742 ;
  assign n18749 = ( x1156 & n18739 ) | ( x1156 & n18748 ) | ( n18739 & n18748 ) ;
  assign n18750 = ~n18739 & n18749 ;
  assign n18547 = n18516 ^ n16318 ^ 1'b0 ;
  assign n18548 = ( n18516 & n18546 ) | ( n18516 & ~n18547 ) | ( n18546 & ~n18547 ) ;
  assign n18549 = x628 & ~n18548 ;
  assign n18553 = x628 & ~n18516 ;
  assign n18554 = x1156 | n18553 ;
  assign n18555 = ( n18548 & n18549 ) | ( n18548 & ~n18554 ) | ( n18549 & ~n18554 ) ;
  assign n18751 = ( x629 & ~n18555 ) | ( x629 & n18750 ) | ( ~n18555 & n18750 ) ;
  assign n18752 = ~n18750 & n18751 ;
  assign n18550 = x628 | n18516 ;
  assign n18551 = ( x1156 & n18549 ) | ( x1156 & n18550 ) | ( n18549 & n18550 ) ;
  assign n18552 = ~n18549 & n18551 ;
  assign n18743 = x628 & ~n18742 ;
  assign n18744 = x1156 | n18743 ;
  assign n18745 = ( n18738 & n18739 ) | ( n18738 & ~n18744 ) | ( n18739 & ~n18744 ) ;
  assign n18746 = ( x629 & ~n18552 ) | ( x629 & n18745 ) | ( ~n18552 & n18745 ) ;
  assign n18747 = n18552 | n18746 ;
  assign n18753 = n18752 ^ n18747 ^ 1'b0 ;
  assign n18754 = ( x792 & ~n18747 ) | ( x792 & n18752 ) | ( ~n18747 & n18752 ) ;
  assign n18755 = ( x792 & ~n18753 ) | ( x792 & n18754 ) | ( ~n18753 & n18754 ) ;
  assign n18756 = ( x792 & n18738 ) | ( x792 & ~n18755 ) | ( n18738 & ~n18755 ) ;
  assign n18757 = ~n18755 & n18756 ;
  assign n18758 = x647 & ~n18757 ;
  assign n18759 = n18516 ^ n16339 ^ 1'b0 ;
  assign n18760 = ( n18516 & n18742 ) | ( n18516 & ~n18759 ) | ( n18742 & ~n18759 ) ;
  assign n18766 = x647 | n18760 ;
  assign n18767 = ( x1157 & n18758 ) | ( x1157 & n18766 ) | ( n18758 & n18766 ) ;
  assign n18768 = ~n18758 & n18767 ;
  assign n18556 = n18552 | n18555 ;
  assign n18557 = n18548 ^ x792 ^ 1'b0 ;
  assign n18558 = ( n18548 & n18556 ) | ( n18548 & n18557 ) | ( n18556 & n18557 ) ;
  assign n18559 = x647 & ~n18558 ;
  assign n18769 = x647 & ~n18516 ;
  assign n18770 = x1157 | n18769 ;
  assign n18771 = ( n18558 & n18559 ) | ( n18558 & ~n18770 ) | ( n18559 & ~n18770 ) ;
  assign n18772 = ( x630 & n18768 ) | ( x630 & ~n18771 ) | ( n18768 & ~n18771 ) ;
  assign n18773 = ~n18768 & n18772 ;
  assign n18560 = x647 | n18516 ;
  assign n18561 = ( x1157 & n18559 ) | ( x1157 & n18560 ) | ( n18559 & n18560 ) ;
  assign n18562 = ~n18559 & n18561 ;
  assign n18761 = x647 & ~n18760 ;
  assign n18762 = x1157 | n18761 ;
  assign n18763 = ( n18757 & n18758 ) | ( n18757 & ~n18762 ) | ( n18758 & ~n18762 ) ;
  assign n18764 = ( x630 & ~n18562 ) | ( x630 & n18763 ) | ( ~n18562 & n18763 ) ;
  assign n18765 = n18562 | n18764 ;
  assign n18774 = n18773 ^ n18765 ^ 1'b0 ;
  assign n18775 = ( x787 & ~n18765 ) | ( x787 & n18773 ) | ( ~n18765 & n18773 ) ;
  assign n18776 = ( x787 & ~n18774 ) | ( x787 & n18775 ) | ( ~n18774 & n18775 ) ;
  assign n18777 = ( x787 & n18757 ) | ( x787 & ~n18776 ) | ( n18757 & ~n18776 ) ;
  assign n18778 = ~n18776 & n18777 ;
  assign n18779 = ~x790 & n18778 ;
  assign n18787 = x644 & ~n18516 ;
  assign n18788 = x715 & ~n18787 ;
  assign n18789 = n18516 ^ n16376 ^ 1'b0 ;
  assign n18790 = ( n18516 & n18760 ) | ( n18516 & ~n18789 ) | ( n18760 & ~n18789 ) ;
  assign n18791 = x644 & ~n18790 ;
  assign n18792 = ( n18788 & n18790 ) | ( n18788 & n18791 ) | ( n18790 & n18791 ) ;
  assign n18780 = x644 | n18778 ;
  assign n18781 = n18562 | n18771 ;
  assign n18782 = n18558 ^ x787 ^ 1'b0 ;
  assign n18783 = ( n18558 & n18781 ) | ( n18558 & n18782 ) | ( n18781 & n18782 ) ;
  assign n18784 = x644 & ~n18783 ;
  assign n18785 = ( x715 & n18780 ) | ( x715 & ~n18784 ) | ( n18780 & ~n18784 ) ;
  assign n18786 = ~x715 & n18785 ;
  assign n18793 = ( x1160 & n18786 ) | ( x1160 & ~n18792 ) | ( n18786 & ~n18792 ) ;
  assign n18794 = n18792 | n18793 ;
  assign n18795 = x644 & ~n18778 ;
  assign n18796 = x644 | n18783 ;
  assign n18797 = ( x715 & n18795 ) | ( x715 & n18796 ) | ( n18795 & n18796 ) ;
  assign n18798 = ~n18795 & n18797 ;
  assign n18799 = x644 | n18516 ;
  assign n18800 = ( x715 & ~n18791 ) | ( x715 & n18799 ) | ( ~n18791 & n18799 ) ;
  assign n18801 = ~x715 & n18800 ;
  assign n18802 = ( x1160 & n18798 ) | ( x1160 & ~n18801 ) | ( n18798 & ~n18801 ) ;
  assign n18803 = ~n18798 & n18802 ;
  assign n18804 = x790 & ~n18803 ;
  assign n18805 = n18794 & n18804 ;
  assign n18806 = ( n5193 & ~n18779 ) | ( n5193 & n18805 ) | ( ~n18779 & n18805 ) ;
  assign n18807 = n18779 | n18806 ;
  assign n18808 = ( x57 & ~n18515 ) | ( x57 & n18807 ) | ( ~n18515 & n18807 ) ;
  assign n18809 = ~x57 & n18808 ;
  assign n18810 = x57 & x144 ;
  assign n18811 = x832 | n18810 ;
  assign n18812 = ( ~n18514 & n18809 ) | ( ~n18514 & n18811 ) | ( n18809 & n18811 ) ;
  assign n18813 = ~n18514 & n18812 ;
  assign n18814 = ~x145 & n7318 ;
  assign n18815 = x832 | n18814 ;
  assign n18816 = x145 | n15656 ;
  assign n18817 = x145 | n15644 ;
  assign n18818 = x38 & n18817 ;
  assign n18819 = x145 | x767 ;
  assign n18820 = n15587 & ~n18819 ;
  assign n18821 = n15640 & ~n18820 ;
  assign n18822 = ( x145 & n18820 ) | ( x145 & ~n18821 ) | ( n18820 & ~n18821 ) ;
  assign n18823 = x145 | n15488 ;
  assign n18824 = x767 & n18823 ;
  assign n18825 = ( ~x38 & n18822 ) | ( ~x38 & n18824 ) | ( n18822 & n18824 ) ;
  assign n18826 = ~x38 & n18825 ;
  assign n18827 = ~x767 & n15646 ;
  assign n18828 = ~n18826 & n18827 ;
  assign n18829 = ( n18818 & n18826 ) | ( n18818 & ~n18828 ) | ( n18826 & ~n18828 ) ;
  assign n18830 = ~n2069 & n18829 ;
  assign n18831 = x145 & n2069 ;
  assign n18832 = n18830 | n18831 ;
  assign n18833 = n18816 ^ n15659 ^ 1'b0 ;
  assign n18834 = ( n18816 & n18832 ) | ( n18816 & ~n18833 ) | ( n18832 & ~n18833 ) ;
  assign n18835 = ~n15659 & n18832 ;
  assign n18836 = x609 & n18835 ;
  assign n18837 = ~n15668 & n18816 ;
  assign n18838 = n18836 | n18837 ;
  assign n18839 = ~x609 & n18835 ;
  assign n18840 = n15662 & n18816 ;
  assign n18841 = n18839 | n18840 ;
  assign n18842 = n18838 ^ x1155 ^ 1'b0 ;
  assign n18843 = ( n18838 & n18841 ) | ( n18838 & ~n18842 ) | ( n18841 & ~n18842 ) ;
  assign n18844 = n18834 ^ x785 ^ 1'b0 ;
  assign n18845 = ( n18834 & n18843 ) | ( n18834 & n18844 ) | ( n18843 & n18844 ) ;
  assign n18846 = x618 & ~n18845 ;
  assign n18847 = x618 | n18816 ;
  assign n18848 = ( x1154 & n18846 ) | ( x1154 & n18847 ) | ( n18846 & n18847 ) ;
  assign n18849 = ~n18846 & n18848 ;
  assign n18850 = x618 & ~n18816 ;
  assign n18851 = x1154 | n18850 ;
  assign n18852 = ( n18845 & n18846 ) | ( n18845 & ~n18851 ) | ( n18846 & ~n18851 ) ;
  assign n18853 = n18849 | n18852 ;
  assign n18854 = n18845 ^ x781 ^ 1'b0 ;
  assign n18855 = ( n18845 & n18853 ) | ( n18845 & n18854 ) | ( n18853 & n18854 ) ;
  assign n18856 = x619 & ~n18855 ;
  assign n18857 = x619 | n18816 ;
  assign n18858 = ( x1159 & n18856 ) | ( x1159 & n18857 ) | ( n18856 & n18857 ) ;
  assign n18859 = ~n18856 & n18858 ;
  assign n18860 = x619 & ~n18816 ;
  assign n18861 = x1159 | n18860 ;
  assign n18862 = ( n18855 & n18856 ) | ( n18855 & ~n18861 ) | ( n18856 & ~n18861 ) ;
  assign n18863 = n18859 | n18862 ;
  assign n18864 = n18855 ^ x789 ^ 1'b0 ;
  assign n18865 = ( n18855 & n18863 ) | ( n18855 & n18864 ) | ( n18863 & n18864 ) ;
  assign n18866 = x626 & ~n18865 ;
  assign n18867 = x626 & ~n18816 ;
  assign n18868 = x1158 | n18867 ;
  assign n18869 = ( n18865 & n18866 ) | ( n18865 & ~n18868 ) | ( n18866 & ~n18868 ) ;
  assign n18870 = n18866 & ~n18869 ;
  assign n18871 = ( x1158 & n18816 ) | ( x1158 & n18867 ) | ( n18816 & n18867 ) ;
  assign n18872 = ( n18869 & ~n18870 ) | ( n18869 & n18871 ) | ( ~n18870 & n18871 ) ;
  assign n18873 = n18865 ^ x788 ^ 1'b0 ;
  assign n18874 = ( n18865 & n18872 ) | ( n18865 & n18873 ) | ( n18872 & n18873 ) ;
  assign n18875 = n18816 ^ n16339 ^ 1'b0 ;
  assign n18876 = ( n18816 & n18874 ) | ( n18816 & ~n18875 ) | ( n18874 & ~n18875 ) ;
  assign n18877 = n18816 ^ n16376 ^ 1'b0 ;
  assign n18878 = ( n18816 & n18876 ) | ( n18816 & ~n18877 ) | ( n18876 & ~n18877 ) ;
  assign n18879 = x644 & ~n18878 ;
  assign n18880 = x644 & ~n18816 ;
  assign n18881 = ( ~x715 & n18816 ) | ( ~x715 & n18880 ) | ( n18816 & n18880 ) ;
  assign n18882 = x1160 & ~n18881 ;
  assign n18883 = ( x1160 & n18879 ) | ( x1160 & n18882 ) | ( n18879 & n18882 ) ;
  assign n18884 = n16185 & n18817 ;
  assign n18885 = ( x38 & x145 ) | ( x38 & n16700 ) | ( x145 & n16700 ) ;
  assign n18886 = ~n2069 & n18885 ;
  assign n18887 = ( x145 & n16697 ) | ( x145 & ~n18886 ) | ( n16697 & ~n18886 ) ;
  assign n18888 = ~n18886 & n18887 ;
  assign n18889 = ( x698 & ~n18884 ) | ( x698 & n18888 ) | ( ~n18884 & n18888 ) ;
  assign n18890 = n18884 | n18889 ;
  assign n18891 = n18890 ^ n18816 ^ 1'b0 ;
  assign n18892 = x698 | n2069 ;
  assign n18893 = ( n18816 & n18891 ) | ( n18816 & ~n18892 ) | ( n18891 & ~n18892 ) ;
  assign n18894 = ( n18890 & ~n18891 ) | ( n18890 & n18893 ) | ( ~n18891 & n18893 ) ;
  assign n18895 = x625 & ~n18894 ;
  assign n18896 = x625 | n18816 ;
  assign n18897 = ( x1153 & n18895 ) | ( x1153 & n18896 ) | ( n18895 & n18896 ) ;
  assign n18898 = ~n18895 & n18897 ;
  assign n18899 = x625 & ~n18816 ;
  assign n18900 = x1153 | n18899 ;
  assign n18901 = ( x625 & n18894 ) | ( x625 & ~n18900 ) | ( n18894 & ~n18900 ) ;
  assign n18902 = ~n18900 & n18901 ;
  assign n18903 = n18898 | n18902 ;
  assign n18904 = n18894 ^ x778 ^ 1'b0 ;
  assign n18905 = ( n18894 & n18903 ) | ( n18894 & n18904 ) | ( n18903 & n18904 ) ;
  assign n18906 = n18816 ^ n16234 ^ 1'b0 ;
  assign n18907 = ( n18816 & n18905 ) | ( n18816 & ~n18906 ) | ( n18905 & ~n18906 ) ;
  assign n18908 = n18816 ^ n16254 ^ 1'b0 ;
  assign n18909 = ( n18816 & n18907 ) | ( n18816 & ~n18908 ) | ( n18907 & ~n18908 ) ;
  assign n18910 = n18816 ^ n16279 ^ 1'b0 ;
  assign n18911 = ( n18816 & n18909 ) | ( n18816 & ~n18910 ) | ( n18909 & ~n18910 ) ;
  assign n18912 = n18816 ^ n16318 ^ 1'b0 ;
  assign n18913 = ( n18816 & n18911 ) | ( n18816 & ~n18912 ) | ( n18911 & ~n18912 ) ;
  assign n18914 = x628 & ~n18913 ;
  assign n18915 = x628 | n18816 ;
  assign n18916 = ( x1156 & n18914 ) | ( x1156 & n18915 ) | ( n18914 & n18915 ) ;
  assign n18917 = ~n18914 & n18916 ;
  assign n18918 = x628 & ~n18816 ;
  assign n18919 = x1156 | n18918 ;
  assign n18920 = ( n18913 & n18914 ) | ( n18913 & ~n18919 ) | ( n18914 & ~n18919 ) ;
  assign n18921 = n18917 | n18920 ;
  assign n18922 = n18913 ^ x792 ^ 1'b0 ;
  assign n18923 = ( n18913 & n18921 ) | ( n18913 & n18922 ) | ( n18921 & n18922 ) ;
  assign n18924 = n18816 ^ x647 ^ 1'b0 ;
  assign n18925 = ( n18816 & n18923 ) | ( n18816 & ~n18924 ) | ( n18923 & ~n18924 ) ;
  assign n18926 = ( n18816 & n18923 ) | ( n18816 & n18924 ) | ( n18923 & n18924 ) ;
  assign n18927 = n18925 ^ x1157 ^ 1'b0 ;
  assign n18928 = ( n18925 & n18926 ) | ( n18925 & n18927 ) | ( n18926 & n18927 ) ;
  assign n18929 = n18923 ^ x787 ^ 1'b0 ;
  assign n18930 = ( n18923 & n18928 ) | ( n18923 & n18929 ) | ( n18928 & n18929 ) ;
  assign n18931 = x644 & ~n18930 ;
  assign n18932 = ( x715 & n18930 ) | ( x715 & n18931 ) | ( n18930 & n18931 ) ;
  assign n18933 = n18883 & ~n18932 ;
  assign n19065 = x715 & ~n18880 ;
  assign n19066 = ( n18878 & n18879 ) | ( n18878 & n19065 ) | ( n18879 & n19065 ) ;
  assign n18934 = x715 | n18931 ;
  assign n18935 = x698 & ~n18829 ;
  assign n18936 = x145 & ~n16054 ;
  assign n18937 = ~x145 & n16048 ;
  assign n18938 = ( x767 & ~n18936 ) | ( x767 & n18937 ) | ( ~n18936 & n18937 ) ;
  assign n18939 = n18936 | n18938 ;
  assign n18940 = ~x145 & n16044 ;
  assign n18941 = x145 & ~n16029 ;
  assign n18942 = ( x767 & n18940 ) | ( x767 & ~n18941 ) | ( n18940 & ~n18941 ) ;
  assign n18943 = ~n18940 & n18942 ;
  assign n18944 = ( x39 & n18939 ) | ( x39 & ~n18943 ) | ( n18939 & ~n18943 ) ;
  assign n18945 = n18944 ^ n18939 ^ 1'b0 ;
  assign n18946 = ( x39 & n18944 ) | ( x39 & ~n18945 ) | ( n18944 & ~n18945 ) ;
  assign n18947 = x145 & n15795 ;
  assign n18948 = x767 & ~n18947 ;
  assign n18949 = x145 | n15876 ;
  assign n18950 = n18948 & n18949 ;
  assign n18951 = x145 & n15943 ;
  assign n18952 = x145 | n16003 ;
  assign n18953 = ( x767 & ~n18951 ) | ( x767 & n18952 ) | ( ~n18951 & n18952 ) ;
  assign n18954 = ~x767 & n18953 ;
  assign n18955 = ( x39 & n18950 ) | ( x39 & ~n18954 ) | ( n18950 & ~n18954 ) ;
  assign n18956 = ~n18950 & n18955 ;
  assign n18957 = ( x38 & n18946 ) | ( x38 & ~n18956 ) | ( n18946 & ~n18956 ) ;
  assign n18958 = ~x38 & n18957 ;
  assign n18959 = ~x767 & n15591 ;
  assign n18960 = n17156 | n18959 ;
  assign n18961 = x145 & ~n5017 ;
  assign n18962 = n18960 & n18961 ;
  assign n18963 = x38 & ~n18962 ;
  assign n18964 = n18963 ^ x698 ^ 1'b0 ;
  assign n18965 = x767 | n15968 ;
  assign n18966 = n17889 & n18965 ;
  assign n18967 = x145 | n18966 ;
  assign n18968 = ( n18963 & ~n18964 ) | ( n18963 & n18967 ) | ( ~n18964 & n18967 ) ;
  assign n18969 = ( x698 & n18964 ) | ( x698 & n18968 ) | ( n18964 & n18968 ) ;
  assign n18970 = ( ~n2069 & n18958 ) | ( ~n2069 & n18969 ) | ( n18958 & n18969 ) ;
  assign n18971 = ~n2069 & n18970 ;
  assign n18972 = n18971 ^ n18935 ^ 1'b0 ;
  assign n18973 = ( n18935 & n18971 ) | ( n18935 & n18972 ) | ( n18971 & n18972 ) ;
  assign n18974 = ( n18831 & ~n18935 ) | ( n18831 & n18973 ) | ( ~n18935 & n18973 ) ;
  assign n18975 = x625 & ~n18974 ;
  assign n18976 = x625 | n18832 ;
  assign n18977 = ( x1153 & n18975 ) | ( x1153 & n18976 ) | ( n18975 & n18976 ) ;
  assign n18978 = ~n18975 & n18977 ;
  assign n18979 = ( x608 & n18902 ) | ( x608 & ~n18978 ) | ( n18902 & ~n18978 ) ;
  assign n18980 = ~n18902 & n18979 ;
  assign n18981 = x608 | n18898 ;
  assign n18982 = x625 & ~n18832 ;
  assign n18983 = x1153 | n18982 ;
  assign n18984 = ( n18974 & n18975 ) | ( n18974 & ~n18983 ) | ( n18975 & ~n18983 ) ;
  assign n18985 = ( ~n18980 & n18981 ) | ( ~n18980 & n18984 ) | ( n18981 & n18984 ) ;
  assign n18986 = ~n18980 & n18985 ;
  assign n18987 = n18974 ^ x778 ^ 1'b0 ;
  assign n18988 = ( n18974 & n18986 ) | ( n18974 & n18987 ) | ( n18986 & n18987 ) ;
  assign n18989 = x609 & ~n18988 ;
  assign n18990 = x609 | n18905 ;
  assign n18991 = ( x1155 & n18989 ) | ( x1155 & n18990 ) | ( n18989 & n18990 ) ;
  assign n18992 = ~n18989 & n18991 ;
  assign n18993 = ~x1155 & n18841 ;
  assign n18994 = ( x660 & n18992 ) | ( x660 & ~n18993 ) | ( n18992 & ~n18993 ) ;
  assign n18995 = ~n18992 & n18994 ;
  assign n18996 = x1155 & n18838 ;
  assign n18997 = x660 | n18996 ;
  assign n18998 = x609 & ~n18905 ;
  assign n18999 = x1155 | n18998 ;
  assign n19000 = ( n18988 & n18989 ) | ( n18988 & ~n18999 ) | ( n18989 & ~n18999 ) ;
  assign n19001 = ( ~n18995 & n18997 ) | ( ~n18995 & n19000 ) | ( n18997 & n19000 ) ;
  assign n19002 = ~n18995 & n19001 ;
  assign n19003 = n18988 ^ x785 ^ 1'b0 ;
  assign n19004 = ( n18988 & n19002 ) | ( n18988 & n19003 ) | ( n19002 & n19003 ) ;
  assign n19005 = x618 & ~n19004 ;
  assign n19006 = x618 | n18907 ;
  assign n19007 = ( x1154 & n19005 ) | ( x1154 & n19006 ) | ( n19005 & n19006 ) ;
  assign n19008 = ~n19005 & n19007 ;
  assign n19009 = ( x627 & n18852 ) | ( x627 & ~n19008 ) | ( n18852 & ~n19008 ) ;
  assign n19010 = ~n18852 & n19009 ;
  assign n19011 = x627 | n18849 ;
  assign n19012 = x618 & ~n18907 ;
  assign n19013 = x1154 | n19012 ;
  assign n19014 = ( n19004 & n19005 ) | ( n19004 & ~n19013 ) | ( n19005 & ~n19013 ) ;
  assign n19015 = ( ~n19010 & n19011 ) | ( ~n19010 & n19014 ) | ( n19011 & n19014 ) ;
  assign n19016 = ~n19010 & n19015 ;
  assign n19017 = n19004 ^ x781 ^ 1'b0 ;
  assign n19018 = ( n19004 & n19016 ) | ( n19004 & n19017 ) | ( n19016 & n19017 ) ;
  assign n19019 = x619 | n19018 ;
  assign n19020 = x619 & ~n18909 ;
  assign n19021 = ( x1159 & n19019 ) | ( x1159 & ~n19020 ) | ( n19019 & ~n19020 ) ;
  assign n19022 = ~x1159 & n19021 ;
  assign n19023 = ( x648 & n18859 ) | ( x648 & ~n19022 ) | ( n18859 & ~n19022 ) ;
  assign n19024 = n19022 | n19023 ;
  assign n19025 = x619 & ~n19018 ;
  assign n19026 = x619 | n18909 ;
  assign n19027 = ( x1159 & n19025 ) | ( x1159 & n19026 ) | ( n19025 & n19026 ) ;
  assign n19028 = ~n19025 & n19027 ;
  assign n19029 = ( x648 & n18862 ) | ( x648 & ~n19028 ) | ( n18862 & ~n19028 ) ;
  assign n19030 = ~n18862 & n19029 ;
  assign n19031 = x789 & ~n19030 ;
  assign n19032 = n19024 & n19031 ;
  assign n19033 = ~x789 & n19018 ;
  assign n19034 = ( n16519 & ~n19032 ) | ( n16519 & n19033 ) | ( ~n19032 & n19033 ) ;
  assign n19035 = n19032 | n19034 ;
  assign n19036 = n16317 & ~n18872 ;
  assign n19037 = n16459 & ~n18911 ;
  assign n19038 = ( x788 & n19036 ) | ( x788 & n19037 ) | ( n19036 & n19037 ) ;
  assign n19039 = n19037 ^ n19036 ^ 1'b0 ;
  assign n19040 = ( x788 & n19038 ) | ( x788 & n19039 ) | ( n19038 & n19039 ) ;
  assign n19041 = ( n18482 & n19035 ) | ( n18482 & ~n19040 ) | ( n19035 & ~n19040 ) ;
  assign n19042 = ~n18482 & n19041 ;
  assign n19043 = n18917 ^ x629 ^ 1'b0 ;
  assign n19044 = ( n18917 & n18920 ) | ( n18917 & n19043 ) | ( n18920 & n19043 ) ;
  assign n19045 = ( x628 & x629 ) | ( x628 & ~x1156 ) | ( x629 & ~x1156 ) ;
  assign n19046 = n19045 ^ x629 ^ 1'b0 ;
  assign n19047 = n18874 & n19046 ;
  assign n19048 = ( x792 & n19044 ) | ( x792 & n19047 ) | ( n19044 & n19047 ) ;
  assign n19049 = n19047 ^ n19044 ^ 1'b0 ;
  assign n19050 = ( x792 & n19048 ) | ( x792 & n19049 ) | ( n19048 & n19049 ) ;
  assign n19051 = ( ~n18484 & n19042 ) | ( ~n18484 & n19050 ) | ( n19042 & n19050 ) ;
  assign n19052 = ~n18484 & n19051 ;
  assign n19053 = n16374 & n18925 ;
  assign n19054 = ( x630 & x647 ) | ( x630 & x1157 ) | ( x647 & x1157 ) ;
  assign n19055 = n19054 ^ x647 ^ 1'b0 ;
  assign n19056 = n18876 & n19055 ;
  assign n19057 = n16373 & n18926 ;
  assign n19058 = ( ~n19053 & n19056 ) | ( ~n19053 & n19057 ) | ( n19056 & n19057 ) ;
  assign n19059 = n19053 | n19058 ;
  assign n19060 = n19052 ^ x787 ^ 1'b0 ;
  assign n19061 = ( ~x787 & n19059 ) | ( ~x787 & n19060 ) | ( n19059 & n19060 ) ;
  assign n19062 = ( x787 & n19052 ) | ( x787 & n19061 ) | ( n19052 & n19061 ) ;
  assign n19063 = ( x644 & ~n18934 ) | ( x644 & n19062 ) | ( ~n18934 & n19062 ) ;
  assign n19064 = ~n18934 & n19063 ;
  assign n19067 = ( x1160 & n19064 ) | ( x1160 & ~n19066 ) | ( n19064 & ~n19066 ) ;
  assign n19068 = n19066 | n19067 ;
  assign n19069 = x790 & ~n19068 ;
  assign n19070 = ( x790 & n18933 ) | ( x790 & n19069 ) | ( n18933 & n19069 ) ;
  assign n19071 = x644 & n18883 ;
  assign n19072 = x790 & ~n19071 ;
  assign n19073 = ( n19062 & ~n19070 ) | ( n19062 & n19072 ) | ( ~n19070 & n19072 ) ;
  assign n19074 = ~n19070 & n19073 ;
  assign n19075 = ( n7318 & ~n18815 ) | ( n7318 & n19074 ) | ( ~n18815 & n19074 ) ;
  assign n19076 = ~n18815 & n19075 ;
  assign n19077 = x145 | n1611 ;
  assign n19078 = ~n18959 & n19077 ;
  assign n19079 = n16397 | n19078 ;
  assign n19080 = n16402 | n19078 ;
  assign n19081 = x1155 & n19080 ;
  assign n19082 = n16405 | n19079 ;
  assign n19083 = ~x1155 & n19082 ;
  assign n19084 = n19081 | n19083 ;
  assign n19085 = n19079 ^ x785 ^ 1'b0 ;
  assign n19086 = ( n19079 & n19084 ) | ( n19079 & n19085 ) | ( n19084 & n19085 ) ;
  assign n19087 = n16411 | n19086 ;
  assign n19088 = x1154 & n19087 ;
  assign n19089 = n16414 | n19086 ;
  assign n19090 = ~x1154 & n19089 ;
  assign n19091 = n19088 | n19090 ;
  assign n19092 = n19086 ^ x781 ^ 1'b0 ;
  assign n19093 = ( n19086 & n19091 ) | ( n19086 & n19092 ) | ( n19091 & n19092 ) ;
  assign n19094 = x619 & ~n19093 ;
  assign n19095 = x619 | n19077 ;
  assign n19096 = ( x1159 & n19094 ) | ( x1159 & n19095 ) | ( n19094 & n19095 ) ;
  assign n19097 = ~n19094 & n19096 ;
  assign n19098 = x619 & ~n19077 ;
  assign n19099 = x1159 | n19098 ;
  assign n19100 = ( n19093 & n19094 ) | ( n19093 & ~n19099 ) | ( n19094 & ~n19099 ) ;
  assign n19101 = n19097 | n19100 ;
  assign n19102 = n19093 ^ x789 ^ 1'b0 ;
  assign n19103 = ( n19093 & n19101 ) | ( n19093 & n19102 ) | ( n19101 & n19102 ) ;
  assign n19104 = x626 & ~n19103 ;
  assign n19105 = x626 & ~n19077 ;
  assign n19106 = x1158 | n19105 ;
  assign n19107 = ( n19103 & n19104 ) | ( n19103 & ~n19106 ) | ( n19104 & ~n19106 ) ;
  assign n19108 = n19104 & ~n19107 ;
  assign n19109 = ( x1158 & n19077 ) | ( x1158 & n19105 ) | ( n19077 & n19105 ) ;
  assign n19110 = ( n19107 & ~n19108 ) | ( n19107 & n19109 ) | ( ~n19108 & n19109 ) ;
  assign n19111 = n19103 ^ x788 ^ 1'b0 ;
  assign n19112 = ( n19103 & n19110 ) | ( n19103 & n19111 ) | ( n19110 & n19111 ) ;
  assign n19113 = n19077 ^ n16339 ^ 1'b0 ;
  assign n19114 = ( n19077 & n19112 ) | ( n19077 & ~n19113 ) | ( n19112 & ~n19113 ) ;
  assign n19115 = n19055 & n19114 ;
  assign n19116 = x647 & ~n19077 ;
  assign n19117 = x1157 | n19116 ;
  assign n19118 = ~x698 & n15778 ;
  assign n19119 = n19077 & ~n19118 ;
  assign n19120 = ~x625 & n19118 ;
  assign n19121 = ~x1153 & n19077 ;
  assign n19122 = ~n19120 & n19121 ;
  assign n19123 = ( x1153 & n19119 ) | ( x1153 & n19120 ) | ( n19119 & n19120 ) ;
  assign n19124 = n19122 | n19123 ;
  assign n19125 = n19119 ^ x778 ^ 1'b0 ;
  assign n19126 = ( n19119 & n19124 ) | ( n19119 & n19125 ) | ( n19124 & n19125 ) ;
  assign n19127 = n16447 | n19126 ;
  assign n19128 = n16449 | n19127 ;
  assign n19129 = n16451 | n19128 ;
  assign n19130 = n16530 | n19129 ;
  assign n19131 = n16560 | n19130 ;
  assign n19132 = ( x647 & ~n19117 ) | ( x647 & n19131 ) | ( ~n19117 & n19131 ) ;
  assign n19133 = ~n19117 & n19132 ;
  assign n19134 = n19077 ^ x647 ^ 1'b0 ;
  assign n19135 = ( n19077 & n19131 ) | ( n19077 & n19134 ) | ( n19131 & n19134 ) ;
  assign n19136 = x1157 & n19135 ;
  assign n19137 = ( n16375 & n19133 ) | ( n16375 & n19136 ) | ( n19133 & n19136 ) ;
  assign n19138 = ( x787 & n19115 ) | ( x787 & n19137 ) | ( n19115 & n19137 ) ;
  assign n19139 = n19137 ^ n19115 ^ 1'b0 ;
  assign n19140 = ( x787 & n19138 ) | ( x787 & n19139 ) | ( n19138 & n19139 ) ;
  assign n19141 = n16459 & ~n19129 ;
  assign n19142 = n16317 & ~n19110 ;
  assign n19143 = ( x788 & n19141 ) | ( x788 & n19142 ) | ( n19141 & n19142 ) ;
  assign n19144 = n19142 ^ n19141 ^ 1'b0 ;
  assign n19145 = ( x788 & n19143 ) | ( x788 & n19144 ) | ( n19143 & n19144 ) ;
  assign n19146 = n15524 | n19119 ;
  assign n19147 = n19078 & n19146 ;
  assign n19148 = x625 & ~n19146 ;
  assign n19149 = ( n19121 & n19147 ) | ( n19121 & n19148 ) | ( n19147 & n19148 ) ;
  assign n19150 = ( x608 & n19123 ) | ( x608 & ~n19149 ) | ( n19123 & ~n19149 ) ;
  assign n19151 = n19149 | n19150 ;
  assign n19152 = x1153 & n19078 ;
  assign n19153 = ~n19148 & n19152 ;
  assign n19154 = x608 & ~n19122 ;
  assign n19155 = n19151 & ~n19154 ;
  assign n19156 = ( n19151 & n19153 ) | ( n19151 & n19155 ) | ( n19153 & n19155 ) ;
  assign n19157 = n19147 ^ x778 ^ 1'b0 ;
  assign n19158 = ( n19147 & n19156 ) | ( n19147 & n19157 ) | ( n19156 & n19157 ) ;
  assign n19159 = x609 & ~n19158 ;
  assign n19160 = x609 | n19126 ;
  assign n19161 = ( x1155 & n19159 ) | ( x1155 & n19160 ) | ( n19159 & n19160 ) ;
  assign n19162 = ~n19159 & n19161 ;
  assign n19163 = ( x660 & n19083 ) | ( x660 & ~n19162 ) | ( n19083 & ~n19162 ) ;
  assign n19164 = ~n19083 & n19163 ;
  assign n19165 = x660 | n19081 ;
  assign n19166 = x609 & ~n19126 ;
  assign n19167 = x1155 | n19166 ;
  assign n19168 = ( n19158 & n19159 ) | ( n19158 & ~n19167 ) | ( n19159 & ~n19167 ) ;
  assign n19169 = ( ~n19164 & n19165 ) | ( ~n19164 & n19168 ) | ( n19165 & n19168 ) ;
  assign n19170 = ~n19164 & n19169 ;
  assign n19171 = n19158 ^ x785 ^ 1'b0 ;
  assign n19172 = ( n19158 & n19170 ) | ( n19158 & n19171 ) | ( n19170 & n19171 ) ;
  assign n19173 = x618 & ~n19172 ;
  assign n19174 = x618 | n19127 ;
  assign n19175 = ( x1154 & n19173 ) | ( x1154 & n19174 ) | ( n19173 & n19174 ) ;
  assign n19176 = ~n19173 & n19175 ;
  assign n19177 = ( x627 & n19090 ) | ( x627 & ~n19176 ) | ( n19090 & ~n19176 ) ;
  assign n19178 = ~n19090 & n19177 ;
  assign n19179 = x627 | n19088 ;
  assign n19180 = x618 & ~n19127 ;
  assign n19181 = x1154 | n19180 ;
  assign n19182 = ( n19172 & n19173 ) | ( n19172 & ~n19181 ) | ( n19173 & ~n19181 ) ;
  assign n19183 = ( ~n19178 & n19179 ) | ( ~n19178 & n19182 ) | ( n19179 & n19182 ) ;
  assign n19184 = ~n19178 & n19183 ;
  assign n19185 = n19172 ^ x781 ^ 1'b0 ;
  assign n19186 = ( n19172 & n19184 ) | ( n19172 & n19185 ) | ( n19184 & n19185 ) ;
  assign n19187 = ~x789 & n19186 ;
  assign n19188 = x619 & ~n19128 ;
  assign n19189 = x1159 | n19188 ;
  assign n19190 = x619 & ~n19186 ;
  assign n19191 = ( n19186 & ~n19189 ) | ( n19186 & n19190 ) | ( ~n19189 & n19190 ) ;
  assign n19192 = ( x648 & n19097 ) | ( x648 & ~n19191 ) | ( n19097 & ~n19191 ) ;
  assign n19193 = n19191 | n19192 ;
  assign n19194 = x619 | n19128 ;
  assign n19195 = x1159 & ~n19190 ;
  assign n19196 = n19194 & n19195 ;
  assign n19197 = ( x648 & n19100 ) | ( x648 & ~n19196 ) | ( n19100 & ~n19196 ) ;
  assign n19198 = ~n19100 & n19197 ;
  assign n19199 = x789 & ~n19198 ;
  assign n19200 = n19193 & n19199 ;
  assign n19201 = ( n16519 & ~n19187 ) | ( n16519 & n19200 ) | ( ~n19187 & n19200 ) ;
  assign n19202 = n19187 | n19201 ;
  assign n19203 = n19202 ^ n19145 ^ 1'b0 ;
  assign n19204 = ( n19145 & n19202 ) | ( n19145 & n19203 ) | ( n19202 & n19203 ) ;
  assign n19205 = ( n18482 & ~n19145 ) | ( n18482 & n19204 ) | ( ~n19145 & n19204 ) ;
  assign n19206 = n18484 ^ x792 ^ 1'b0 ;
  assign n19207 = n16556 & ~n19112 ;
  assign n19208 = x1156 | n16532 ;
  assign n19209 = n19130 | n19208 ;
  assign n19210 = ( x629 & n19207 ) | ( x629 & n19209 ) | ( n19207 & n19209 ) ;
  assign n19211 = ~n19207 & n19210 ;
  assign n19212 = x1156 & ~n16537 ;
  assign n19213 = ~n19130 & n19212 ;
  assign n19214 = n16557 & ~n19112 ;
  assign n19215 = n19213 | n19214 ;
  assign n19216 = ( x629 & ~n19211 ) | ( x629 & n19215 ) | ( ~n19211 & n19215 ) ;
  assign n19217 = ~n19211 & n19216 ;
  assign n19218 = ( x792 & ~n19206 ) | ( x792 & n19217 ) | ( ~n19206 & n19217 ) ;
  assign n19219 = ( n18484 & n19206 ) | ( n18484 & n19218 ) | ( n19206 & n19218 ) ;
  assign n19220 = ( n19140 & n19205 ) | ( n19140 & ~n19219 ) | ( n19205 & ~n19219 ) ;
  assign n19221 = n19220 ^ n19205 ^ 1'b0 ;
  assign n19222 = ( n19140 & n19220 ) | ( n19140 & ~n19221 ) | ( n19220 & ~n19221 ) ;
  assign n19223 = x790 | n19222 ;
  assign n19224 = x832 & n19223 ;
  assign n19225 = x644 & ~n19222 ;
  assign n19226 = ( x787 & n19133 ) | ( x787 & ~n19136 ) | ( n19133 & ~n19136 ) ;
  assign n19227 = ~n19133 & n19226 ;
  assign n19228 = ( x787 & n19131 ) | ( x787 & ~n19227 ) | ( n19131 & ~n19227 ) ;
  assign n19229 = ~n19227 & n19228 ;
  assign n19230 = x644 | n19229 ;
  assign n19231 = ( x715 & n19225 ) | ( x715 & n19230 ) | ( n19225 & n19230 ) ;
  assign n19232 = ~n19225 & n19231 ;
  assign n19233 = x644 | n19077 ;
  assign n19234 = n19077 ^ n16376 ^ 1'b0 ;
  assign n19235 = ( n19077 & n19114 ) | ( n19077 & ~n19234 ) | ( n19114 & ~n19234 ) ;
  assign n19236 = x644 & ~n19235 ;
  assign n19237 = ( x715 & n19233 ) | ( x715 & ~n19236 ) | ( n19233 & ~n19236 ) ;
  assign n19238 = ~x715 & n19237 ;
  assign n19239 = ( x1160 & n19232 ) | ( x1160 & ~n19238 ) | ( n19232 & ~n19238 ) ;
  assign n19240 = ~n19232 & n19239 ;
  assign n19241 = x644 & ~n19077 ;
  assign n19242 = x715 & ~n19241 ;
  assign n19243 = ( n19235 & n19236 ) | ( n19235 & n19242 ) | ( n19236 & n19242 ) ;
  assign n19244 = x644 & ~n19229 ;
  assign n19245 = x715 | n19244 ;
  assign n19246 = ( n19222 & n19225 ) | ( n19222 & ~n19245 ) | ( n19225 & ~n19245 ) ;
  assign n19247 = ( x1160 & ~n19243 ) | ( x1160 & n19246 ) | ( ~n19243 & n19246 ) ;
  assign n19248 = n19243 | n19247 ;
  assign n19249 = x790 & ~n19248 ;
  assign n19250 = ( x790 & n19240 ) | ( x790 & n19249 ) | ( n19240 & n19249 ) ;
  assign n19251 = ( n19076 & n19224 ) | ( n19076 & ~n19250 ) | ( n19224 & ~n19250 ) ;
  assign n19252 = n19251 ^ n19224 ^ 1'b0 ;
  assign n19253 = ( n19076 & n19251 ) | ( n19076 & ~n19252 ) | ( n19251 & ~n19252 ) ;
  assign n19256 = x907 & ~x947 ;
  assign n19257 = x735 & n19256 ;
  assign n19258 = x743 & x947 ;
  assign n19259 = n19257 | n19258 ;
  assign n19278 = n15378 & n19259 ;
  assign n19287 = x215 & ~n19278 ;
  assign n19288 = x146 & ~n15406 ;
  assign n19289 = n19287 & ~n19288 ;
  assign n19290 = x735 & x907 ;
  assign n19291 = n15433 & n19290 ;
  assign n19262 = x146 & ~n15468 ;
  assign n19292 = x907 | n5060 ;
  assign n19293 = n19262 & ~n19292 ;
  assign n19294 = ( x947 & ~n19291 ) | ( x947 & n19293 ) | ( ~n19291 & n19293 ) ;
  assign n19295 = n19291 | n19294 ;
  assign n19296 = x743 & n15433 ;
  assign n19254 = x146 & ~n15433 ;
  assign n19297 = x947 & ~n19254 ;
  assign n19298 = n19295 & ~n19297 ;
  assign n19299 = ( n19295 & n19296 ) | ( n19295 & n19298 ) | ( n19296 & n19298 ) ;
  assign n19300 = n19254 & n19292 ;
  assign n19301 = ( n2263 & n19299 ) | ( n2263 & n19300 ) | ( n19299 & n19300 ) ;
  assign n19302 = n19300 ^ n19299 ^ 1'b0 ;
  assign n19303 = ( n2263 & n19301 ) | ( n2263 & n19302 ) | ( n19301 & n19302 ) ;
  assign n19269 = n15337 ^ x146 ^ 1'b0 ;
  assign n19270 = ( x146 & n19259 ) | ( x146 & n19269 ) | ( n19259 & n19269 ) ;
  assign n19304 = ~n2263 & n19270 ;
  assign n19305 = ( x215 & ~n19303 ) | ( x215 & n19304 ) | ( ~n19303 & n19304 ) ;
  assign n19306 = n19303 | n19305 ;
  assign n19307 = x299 & ~n19306 ;
  assign n19308 = ( x299 & n19289 ) | ( x299 & n19307 ) | ( n19289 & n19307 ) ;
  assign n19255 = n5114 & ~n19254 ;
  assign n19260 = n15433 & n19259 ;
  assign n19261 = n19255 & ~n19260 ;
  assign n19263 = n5114 | n19262 ;
  assign n19264 = n15468 & n19259 ;
  assign n19265 = ( ~n19261 & n19263 ) | ( ~n19261 & n19264 ) | ( n19263 & n19264 ) ;
  assign n19266 = ~n19261 & n19265 ;
  assign n19267 = ( x222 & x224 ) | ( x222 & ~n19266 ) | ( x224 & ~n19266 ) ;
  assign n19268 = ~n19266 & n19267 ;
  assign n19271 = n1359 | n19270 ;
  assign n19272 = ( x223 & ~n19268 ) | ( x223 & n19271 ) | ( ~n19268 & n19271 ) ;
  assign n19273 = ~x223 & n19272 ;
  assign n19274 = n15402 & ~n19259 ;
  assign n19275 = x146 | n15402 ;
  assign n19276 = ( n5114 & ~n19274 ) | ( n5114 & n19275 ) | ( ~n19274 & n19275 ) ;
  assign n19277 = ~n5114 & n19276 ;
  assign n19279 = x146 & ~n15378 ;
  assign n19280 = n19278 | n19279 ;
  assign n19281 = n5114 & n19280 ;
  assign n19282 = ( x223 & n19277 ) | ( x223 & n19281 ) | ( n19277 & n19281 ) ;
  assign n19283 = n19281 ^ n19277 ^ 1'b0 ;
  assign n19284 = ( x223 & n19282 ) | ( x223 & n19283 ) | ( n19282 & n19283 ) ;
  assign n19285 = ( x299 & ~n19273 ) | ( x299 & n19284 ) | ( ~n19273 & n19284 ) ;
  assign n19286 = n19273 | n19285 ;
  assign n19309 = n19308 ^ n19286 ^ 1'b0 ;
  assign n19310 = ( x39 & ~n19286 ) | ( x39 & n19308 ) | ( ~n19286 & n19308 ) ;
  assign n19311 = ( x39 & ~n19309 ) | ( x39 & n19310 ) | ( ~n19309 & n19310 ) ;
  assign n19312 = x146 | n15330 ;
  assign n19313 = n15330 & ~n19259 ;
  assign n19314 = x299 & ~n19313 ;
  assign n19315 = n19312 & n19314 ;
  assign n19316 = x146 | n15327 ;
  assign n19317 = n15327 & ~n19259 ;
  assign n19318 = ( x299 & n19316 ) | ( x299 & ~n19317 ) | ( n19316 & ~n19317 ) ;
  assign n19319 = ~x299 & n19318 ;
  assign n19320 = ( x39 & ~n19315 ) | ( x39 & n19319 ) | ( ~n19315 & n19319 ) ;
  assign n19321 = n19315 | n19320 ;
  assign n19322 = ( x38 & ~n19311 ) | ( x38 & n19321 ) | ( ~n19311 & n19321 ) ;
  assign n19323 = ~x38 & n19322 ;
  assign n19324 = n1611 & ~n19259 ;
  assign n19325 = ~n5017 & n19324 ;
  assign n19326 = x146 | n15644 ;
  assign n19327 = ( x38 & n19325 ) | ( x38 & n19326 ) | ( n19325 & n19326 ) ;
  assign n19328 = ~n19325 & n19327 ;
  assign n19329 = ( n8793 & ~n19323 ) | ( n8793 & n19328 ) | ( ~n19323 & n19328 ) ;
  assign n19330 = n19323 | n19329 ;
  assign n19331 = x146 | n1611 ;
  assign n19332 = x832 & ~n19324 ;
  assign n19333 = n19331 & n19332 ;
  assign n19334 = ~x146 & n8793 ;
  assign n19335 = x832 | n19334 ;
  assign n19336 = ~n19333 & n19335 ;
  assign n19337 = ( n19330 & n19333 ) | ( n19330 & ~n19336 ) | ( n19333 & ~n19336 ) ;
  assign n19338 = x147 | n1611 ;
  assign n19339 = x832 & n19338 ;
  assign n19340 = ~x147 & n8793 ;
  assign n19341 = ~n5055 & n15653 ;
  assign n19342 = x147 | n19341 ;
  assign n19343 = n5055 & n15644 ;
  assign n19344 = x38 & ~n19343 ;
  assign n19345 = n19342 & n19344 ;
  assign n19346 = n5055 & n15332 ;
  assign n19347 = x215 & ~n15379 ;
  assign n19348 = ( x215 & n5055 ) | ( x215 & n15438 ) | ( n5055 & n15438 ) ;
  assign n19349 = ( x299 & n19347 ) | ( x299 & n19348 ) | ( n19347 & n19348 ) ;
  assign n19350 = ~n19347 & n19349 ;
  assign n19351 = n5055 & n15484 ;
  assign n19352 = ( ~x299 & n19350 ) | ( ~x299 & n19351 ) | ( n19350 & n19351 ) ;
  assign n19353 = n19350 ^ x299 ^ 1'b0 ;
  assign n19354 = ( n19350 & n19352 ) | ( n19350 & ~n19353 ) | ( n19352 & ~n19353 ) ;
  assign n19355 = n19346 ^ x39 ^ 1'b0 ;
  assign n19356 = ( n19346 & n19354 ) | ( n19346 & n19355 ) | ( n19354 & n19355 ) ;
  assign n19357 = x147 & n19356 ;
  assign n19358 = x38 | n19357 ;
  assign n19359 = ( ~n5055 & n15477 ) | ( ~n5055 & n15478 ) | ( n15477 & n15478 ) ;
  assign n19360 = x223 | n19359 ;
  assign n19361 = ~x947 & n15482 ;
  assign n19362 = x223 & ~n19361 ;
  assign n19363 = ( x223 & n15483 ) | ( x223 & n19256 ) | ( n15483 & n19256 ) ;
  assign n19364 = n19362 | n19363 ;
  assign n19365 = ( x299 & n19360 ) | ( x299 & ~n19364 ) | ( n19360 & ~n19364 ) ;
  assign n19366 = n19365 ^ n19360 ^ 1'b0 ;
  assign n19367 = ( x299 & n19365 ) | ( x299 & ~n19366 ) | ( n19365 & ~n19366 ) ;
  assign n19368 = x215 & ~n15405 ;
  assign n19369 = n15436 & ~n19256 ;
  assign n19370 = x947 & n15433 ;
  assign n19371 = n15470 | n19370 ;
  assign n19372 = n2263 & n19371 ;
  assign n19373 = x215 | n19372 ;
  assign n19374 = n19369 | n19373 ;
  assign n19375 = ~n19368 & n19374 ;
  assign n19376 = ~x947 & n19375 ;
  assign n19377 = x299 & ~n19376 ;
  assign n19378 = n19367 & ~n19377 ;
  assign n19379 = x39 & n19378 ;
  assign n19380 = x39 | n19346 ;
  assign n19381 = n15332 & ~n19380 ;
  assign n19382 = n19379 | n19381 ;
  assign n19383 = ( x147 & ~n19358 ) | ( x147 & n19382 ) | ( ~n19358 & n19382 ) ;
  assign n19384 = ~n19358 & n19383 ;
  assign n19385 = ( x770 & ~n19345 ) | ( x770 & n19384 ) | ( ~n19345 & n19384 ) ;
  assign n19386 = n19345 | n19385 ;
  assign n19397 = n15332 & n19256 ;
  assign n19398 = n15378 & n19256 ;
  assign n19399 = n15433 & n19256 ;
  assign n19400 = x907 & n15337 ;
  assign n19401 = ~x947 & n19400 ;
  assign n19402 = n19399 ^ n2263 ^ 1'b0 ;
  assign n19403 = ( n19399 & n19401 ) | ( n19399 & ~n19402 ) | ( n19401 & ~n19402 ) ;
  assign n19404 = n19398 ^ x215 ^ 1'b0 ;
  assign n19405 = ( n19398 & n19403 ) | ( n19398 & ~n19404 ) | ( n19403 & ~n19404 ) ;
  assign n19406 = x299 & n19405 ;
  assign n19391 = ~x299 & n15484 ;
  assign n19407 = n19391 | n19406 ;
  assign n19408 = n15484 & n19256 ;
  assign n19409 = x299 | n19408 ;
  assign n19410 = ( n19406 & n19407 ) | ( n19406 & n19409 ) | ( n19407 & n19409 ) ;
  assign n19411 = n19410 ^ x39 ^ 1'b0 ;
  assign n19412 = ( n19397 & n19410 ) | ( n19397 & ~n19411 ) | ( n19410 & ~n19411 ) ;
  assign n19413 = x38 | n19412 ;
  assign n19414 = ( x38 & x147 ) | ( x38 & n19413 ) | ( x147 & n19413 ) ;
  assign n19387 = x215 & x947 ;
  assign n19388 = n15378 & n19387 ;
  assign n19389 = n19375 | n19388 ;
  assign n19390 = x299 & n19389 ;
  assign n19392 = ~n19256 & n19391 ;
  assign n19393 = n19390 | n19392 ;
  assign n19394 = n15332 & ~n19256 ;
  assign n19395 = n19393 ^ x39 ^ 1'b0 ;
  assign n19396 = ( n19393 & n19394 ) | ( n19393 & ~n19395 ) | ( n19394 & ~n19395 ) ;
  assign n19415 = ( x147 & n19396 ) | ( x147 & ~n19414 ) | ( n19396 & ~n19414 ) ;
  assign n19416 = ~n19414 & n19415 ;
  assign n19417 = n15644 & n19256 ;
  assign n19418 = x38 & ~n19417 ;
  assign n19419 = n15644 & n19418 ;
  assign n19420 = ( x147 & n19418 ) | ( x147 & n19419 ) | ( n19418 & n19419 ) ;
  assign n19421 = ( x770 & n19416 ) | ( x770 & ~n19420 ) | ( n19416 & ~n19420 ) ;
  assign n19422 = ~n19416 & n19421 ;
  assign n19423 = x726 & ~n19422 ;
  assign n19424 = n19386 & n19423 ;
  assign n19425 = ( x38 & ~x947 ) | ( x38 & n17327 ) | ( ~x947 & n17327 ) ;
  assign n19426 = x947 & n15332 ;
  assign n19427 = x947 & n15484 ;
  assign n19428 = x299 | n19427 ;
  assign n19429 = x299 & ~n19388 ;
  assign n19430 = x947 & n15337 ;
  assign n19431 = n2263 | n19430 ;
  assign n19432 = ~x215 & n19431 ;
  assign n19433 = n2263 & ~n19370 ;
  assign n19434 = n19432 & ~n19433 ;
  assign n19435 = n19429 & ~n19434 ;
  assign n19436 = n19428 & ~n19435 ;
  assign n19437 = n19426 ^ x39 ^ 1'b0 ;
  assign n19438 = ( n19426 & n19436 ) | ( n19426 & n19437 ) | ( n19436 & n19437 ) ;
  assign n19439 = x38 | n19438 ;
  assign n19440 = ~n19425 & n19439 ;
  assign n19441 = x147 & ~x770 ;
  assign n19442 = n19440 & n19441 ;
  assign n19443 = ~x947 & n15332 ;
  assign n19444 = x947 & n19391 ;
  assign n19445 = n19368 & ~n19398 ;
  assign n19446 = ~x947 & n15436 ;
  assign n19447 = n15470 | n19399 ;
  assign n19448 = n2263 & n19447 ;
  assign n19449 = x215 | n19448 ;
  assign n19450 = n19446 | n19449 ;
  assign n19451 = ~n19445 & n19450 ;
  assign n19452 = ( n15485 & n19391 ) | ( n15485 & n19451 ) | ( n19391 & n19451 ) ;
  assign n19453 = ~n19444 & n19452 ;
  assign n19454 = n19443 ^ x39 ^ 1'b0 ;
  assign n19455 = ( n19443 & n19453 ) | ( n19443 & n19454 ) | ( n19453 & n19454 ) ;
  assign n19456 = ~x38 & n19455 ;
  assign n19457 = x38 & ~x947 ;
  assign n19458 = n15653 & n19457 ;
  assign n19459 = n19456 | n19458 ;
  assign n19460 = ~x770 & n19459 ;
  assign n19461 = x770 & n15655 ;
  assign n19462 = ( x147 & ~n19460 ) | ( x147 & n19461 ) | ( ~n19460 & n19461 ) ;
  assign n19463 = n19460 | n19462 ;
  assign n19464 = ( x726 & ~n19442 ) | ( x726 & n19463 ) | ( ~n19442 & n19463 ) ;
  assign n19465 = ~x726 & n19464 ;
  assign n19466 = ( n8793 & ~n19424 ) | ( n8793 & n19465 ) | ( ~n19424 & n19465 ) ;
  assign n19467 = n19424 | n19466 ;
  assign n19468 = ( x832 & ~n19340 ) | ( x832 & n19467 ) | ( ~n19340 & n19467 ) ;
  assign n19469 = ~x832 & n19468 ;
  assign n19470 = x726 & n19256 ;
  assign n19471 = ~x770 & x947 ;
  assign n19472 = ( n1611 & n19470 ) | ( n1611 & n19471 ) | ( n19470 & n19471 ) ;
  assign n19473 = n19471 ^ n19470 ^ 1'b0 ;
  assign n19474 = ( n1611 & n19472 ) | ( n1611 & n19473 ) | ( n19472 & n19473 ) ;
  assign n19475 = ~n19469 & n19474 ;
  assign n19476 = ( n19339 & n19469 ) | ( n19339 & ~n19475 ) | ( n19469 & ~n19475 ) ;
  assign n19477 = x749 & x947 ;
  assign n19478 = n1611 & ~n19477 ;
  assign n19479 = x706 & n19256 ;
  assign n19480 = n19478 & ~n19479 ;
  assign n19481 = x148 & ~n1611 ;
  assign n19482 = ( x832 & n19480 ) | ( x832 & ~n19481 ) | ( n19480 & ~n19481 ) ;
  assign n19483 = ~n19480 & n19482 ;
  assign n19484 = x57 & x148 ;
  assign n19485 = x832 | n19484 ;
  assign n19487 = ~x749 & x947 ;
  assign n19488 = n19343 & ~n19487 ;
  assign n19486 = x148 | n15644 ;
  assign n19489 = n19488 ^ n19486 ^ 1'b0 ;
  assign n19490 = ( x38 & ~n19486 ) | ( x38 & n19488 ) | ( ~n19486 & n19488 ) ;
  assign n19491 = ( x38 & ~n19489 ) | ( x38 & n19490 ) | ( ~n19489 & n19490 ) ;
  assign n19492 = x148 & ~n19407 ;
  assign n19493 = ~n8318 & n19393 ;
  assign n19494 = ( x749 & ~n19492 ) | ( x749 & n19493 ) | ( ~n19492 & n19493 ) ;
  assign n19495 = n19492 | n19494 ;
  assign n19496 = x148 & ~n19354 ;
  assign n19497 = ~x148 & n19378 ;
  assign n19498 = ( x749 & n19496 ) | ( x749 & ~n19497 ) | ( n19496 & ~n19497 ) ;
  assign n19499 = ~n19496 & n19498 ;
  assign n19500 = x39 & ~n19499 ;
  assign n19501 = n19495 & n19500 ;
  assign n19502 = n19346 & ~n19487 ;
  assign n19503 = ( ~x39 & x148 ) | ( ~x39 & n15487 ) | ( x148 & n15487 ) ;
  assign n19504 = ~n19502 & n19503 ;
  assign n19505 = ( x38 & ~n19501 ) | ( x38 & n19504 ) | ( ~n19501 & n19504 ) ;
  assign n19506 = n19501 | n19505 ;
  assign n19507 = ( x706 & n19491 ) | ( x706 & n19506 ) | ( n19491 & n19506 ) ;
  assign n19508 = ~n19491 & n19507 ;
  assign n19509 = n2069 | n5193 ;
  assign n19510 = x148 & ~n15653 ;
  assign n19511 = n15644 & ~n19477 ;
  assign n19512 = x38 & ~n19511 ;
  assign n19513 = n19512 ^ n19510 ^ 1'b0 ;
  assign n19514 = ( n19510 & n19512 ) | ( n19510 & n19513 ) | ( n19512 & n19513 ) ;
  assign n19515 = ( x706 & ~n19510 ) | ( x706 & n19514 ) | ( ~n19510 & n19514 ) ;
  assign n19516 = n19388 | n19434 ;
  assign n19517 = x148 & n19516 ;
  assign n19518 = x299 & ~n19517 ;
  assign n19519 = x148 | n19451 ;
  assign n19520 = n19518 & n19519 ;
  assign n19521 = x148 | n15484 ;
  assign n19522 = ~n19428 & n19521 ;
  assign n19523 = ( x749 & n19520 ) | ( x749 & ~n19522 ) | ( n19520 & ~n19522 ) ;
  assign n19524 = ~n19520 & n19523 ;
  assign n19525 = x148 | x749 ;
  assign n19526 = n15486 | n19525 ;
  assign n19527 = ( x39 & n19524 ) | ( x39 & n19526 ) | ( n19524 & n19526 ) ;
  assign n19528 = ~n19524 & n19527 ;
  assign n19529 = n15332 & n19477 ;
  assign n19530 = n19503 & ~n19529 ;
  assign n19531 = x38 | n19530 ;
  assign n19532 = ( ~n19515 & n19528 ) | ( ~n19515 & n19531 ) | ( n19528 & n19531 ) ;
  assign n19533 = ~n19515 & n19532 ;
  assign n19534 = ( ~n19508 & n19509 ) | ( ~n19508 & n19533 ) | ( n19509 & n19533 ) ;
  assign n19535 = n19508 | n19534 ;
  assign n19536 = ~x148 & n19509 ;
  assign n19537 = ( x57 & n19535 ) | ( x57 & ~n19536 ) | ( n19535 & ~n19536 ) ;
  assign n19538 = ~x57 & n19537 ;
  assign n19539 = ( ~n19483 & n19485 ) | ( ~n19483 & n19538 ) | ( n19485 & n19538 ) ;
  assign n19540 = ~n19483 & n19539 ;
  assign n19541 = x149 | n1611 ;
  assign n19542 = x832 & n19541 ;
  assign n19544 = ~x755 & x947 ;
  assign n19561 = n15644 & ~n19544 ;
  assign n19562 = x149 & ~n15653 ;
  assign n19563 = ( x38 & n19561 ) | ( x38 & ~n19562 ) | ( n19561 & ~n19562 ) ;
  assign n19564 = ~n19561 & n19563 ;
  assign n19543 = x149 | n15332 ;
  assign n19545 = n15332 & n19544 ;
  assign n19546 = ( x39 & n19543 ) | ( x39 & ~n19545 ) | ( n19543 & ~n19545 ) ;
  assign n19547 = ~x39 & n19546 ;
  assign n19548 = ~x149 & x755 ;
  assign n19549 = ~n15486 & n19548 ;
  assign n19550 = x39 & ~n19549 ;
  assign n19551 = x149 | n15484 ;
  assign n19552 = ~n19428 & n19551 ;
  assign n19553 = x149 | n19451 ;
  assign n19554 = ( x299 & n14736 ) | ( x299 & n19435 ) | ( n14736 & n19435 ) ;
  assign n19555 = n19553 & n19554 ;
  assign n19556 = ( x755 & ~n19552 ) | ( x755 & n19555 ) | ( ~n19552 & n19555 ) ;
  assign n19557 = n19552 | n19556 ;
  assign n19558 = n19550 & n19557 ;
  assign n19559 = ( x38 & ~n19547 ) | ( x38 & n19558 ) | ( ~n19547 & n19558 ) ;
  assign n19560 = n19547 | n19559 ;
  assign n19565 = n19564 ^ n19560 ^ 1'b0 ;
  assign n19566 = ( x725 & ~n19560 ) | ( x725 & n19564 ) | ( ~n19560 & n19564 ) ;
  assign n19567 = ( x725 & ~n19565 ) | ( x725 & n19566 ) | ( ~n19565 & n19566 ) ;
  assign n19568 = n5055 & n15340 ;
  assign n19569 = x755 & x947 ;
  assign n19570 = x39 | n19569 ;
  assign n19571 = n19568 & ~n19570 ;
  assign n19572 = x149 | n15644 ;
  assign n19573 = x38 & n19572 ;
  assign n19574 = n19573 ^ n19571 ^ 1'b0 ;
  assign n19575 = ( n19571 & n19573 ) | ( n19571 & n19574 ) | ( n19573 & n19574 ) ;
  assign n19576 = ( x725 & ~n19571 ) | ( x725 & n19575 ) | ( ~n19571 & n19575 ) ;
  assign n19577 = ~x149 & n19390 ;
  assign n19578 = x755 & ~n19392 ;
  assign n19579 = x149 & ~n19407 ;
  assign n19580 = ( n19577 & n19578 ) | ( n19577 & ~n19579 ) | ( n19578 & ~n19579 ) ;
  assign n19581 = ~n19577 & n19580 ;
  assign n19582 = ~x149 & n19378 ;
  assign n19583 = x149 & ~n19354 ;
  assign n19584 = ( x755 & ~n19582 ) | ( x755 & n19583 ) | ( ~n19582 & n19583 ) ;
  assign n19585 = n19582 | n19584 ;
  assign n19586 = ( x39 & n19581 ) | ( x39 & n19585 ) | ( n19581 & n19585 ) ;
  assign n19587 = ~n19581 & n19586 ;
  assign n19588 = ~n19397 & n19547 ;
  assign n19589 = ( ~x38 & n19587 ) | ( ~x38 & n19588 ) | ( n19587 & n19588 ) ;
  assign n19590 = ~x38 & n19589 ;
  assign n19591 = ( ~n19567 & n19576 ) | ( ~n19567 & n19590 ) | ( n19576 & n19590 ) ;
  assign n19592 = ~n19567 & n19591 ;
  assign n19593 = ( n2069 & n7318 ) | ( n2069 & ~n19592 ) | ( n7318 & ~n19592 ) ;
  assign n19594 = n19592 | n19593 ;
  assign n19595 = ~x149 & n8793 ;
  assign n19596 = ( x832 & n19594 ) | ( x832 & ~n19595 ) | ( n19594 & ~n19595 ) ;
  assign n19597 = ~x832 & n19596 ;
  assign n19598 = ~x725 & n19256 ;
  assign n19599 = n19544 | n19598 ;
  assign n19600 = n1611 & n19599 ;
  assign n19601 = ~n19597 & n19600 ;
  assign n19602 = ( n19542 & n19597 ) | ( n19542 & ~n19601 ) | ( n19597 & ~n19601 ) ;
  assign n19603 = ~x751 & x947 ;
  assign n19604 = n15644 & ~n19603 ;
  assign n19605 = x150 & ~n15653 ;
  assign n19606 = ( x38 & n19604 ) | ( x38 & n19605 ) | ( n19604 & n19605 ) ;
  assign n19607 = n19605 ^ n19604 ^ 1'b0 ;
  assign n19608 = ( x38 & n19606 ) | ( x38 & n19607 ) | ( n19606 & n19607 ) ;
  assign n19609 = ~x150 & x751 ;
  assign n19610 = ~n15486 & n19609 ;
  assign n19611 = ~x150 & n19453 ;
  assign n19612 = x150 & ~n19436 ;
  assign n19613 = ( x751 & ~n19611 ) | ( x751 & n19612 ) | ( ~n19611 & n19612 ) ;
  assign n19614 = n19611 | n19613 ;
  assign n19615 = x39 & ~n19614 ;
  assign n19616 = ( x39 & n19610 ) | ( x39 & n19615 ) | ( n19610 & n19615 ) ;
  assign n19617 = n15332 ^ x751 ^ 1'b0 ;
  assign n19618 = ( x150 & x751 ) | ( x150 & ~n19617 ) | ( x751 & ~n19617 ) ;
  assign n19619 = ( x39 & n19443 ) | ( x39 & ~n19618 ) | ( n19443 & ~n19618 ) ;
  assign n19620 = n19618 | n19619 ;
  assign n19621 = ( x38 & ~n19616 ) | ( x38 & n19620 ) | ( ~n19616 & n19620 ) ;
  assign n19622 = ~x38 & n19621 ;
  assign n19623 = ( x701 & n19608 ) | ( x701 & ~n19622 ) | ( n19608 & ~n19622 ) ;
  assign n19624 = ~n19608 & n19623 ;
  assign n19625 = x751 & x947 ;
  assign n19626 = ( x39 & n19568 ) | ( x39 & ~n19625 ) | ( n19568 & ~n19625 ) ;
  assign n19627 = ~x39 & n19626 ;
  assign n19628 = x150 | n15644 ;
  assign n19629 = x38 & n19628 ;
  assign n19630 = n19629 ^ n19627 ^ 1'b0 ;
  assign n19631 = ( n19627 & n19629 ) | ( n19627 & n19630 ) | ( n19629 & n19630 ) ;
  assign n19632 = ( x701 & ~n19627 ) | ( x701 & n19631 ) | ( ~n19627 & n19631 ) ;
  assign n19637 = x150 & ~n19410 ;
  assign n19638 = ~x150 & n19393 ;
  assign n19639 = ( x751 & n19637 ) | ( x751 & ~n19638 ) | ( n19637 & ~n19638 ) ;
  assign n19640 = ~n19637 & n19639 ;
  assign n19633 = ~x150 & n19378 ;
  assign n19634 = x150 & ~n19354 ;
  assign n19635 = ( x751 & ~n19633 ) | ( x751 & n19634 ) | ( ~n19633 & n19634 ) ;
  assign n19636 = n19633 | n19635 ;
  assign n19641 = n19640 ^ n19636 ^ 1'b0 ;
  assign n19642 = ( x39 & ~n19636 ) | ( x39 & n19640 ) | ( ~n19636 & n19640 ) ;
  assign n19643 = ( x39 & ~n19641 ) | ( x39 & n19642 ) | ( ~n19641 & n19642 ) ;
  assign n19644 = x150 & ~n15332 ;
  assign n19645 = n19394 & ~n19603 ;
  assign n19646 = ( x39 & ~n19644 ) | ( x39 & n19645 ) | ( ~n19644 & n19645 ) ;
  assign n19647 = n19644 | n19646 ;
  assign n19648 = ( x38 & ~n19643 ) | ( x38 & n19647 ) | ( ~n19643 & n19647 ) ;
  assign n19649 = ~x38 & n19648 ;
  assign n19650 = ( ~n19624 & n19632 ) | ( ~n19624 & n19649 ) | ( n19632 & n19649 ) ;
  assign n19651 = ~n19624 & n19650 ;
  assign n19652 = ( n2069 & n7318 ) | ( n2069 & ~n19651 ) | ( n7318 & ~n19651 ) ;
  assign n19653 = n19651 | n19652 ;
  assign n19654 = ~x701 & n19256 ;
  assign n19655 = n19603 | n19654 ;
  assign n19656 = n1611 & n19655 ;
  assign n19657 = x150 | n1611 ;
  assign n19658 = ( x832 & n19656 ) | ( x832 & n19657 ) | ( n19656 & n19657 ) ;
  assign n19659 = ~n19656 & n19658 ;
  assign n19660 = ~x150 & n8793 ;
  assign n19661 = x832 | n19660 ;
  assign n19662 = ~n19659 & n19661 ;
  assign n19663 = ( n19653 & n19659 ) | ( n19653 & ~n19662 ) | ( n19659 & ~n19662 ) ;
  assign n19664 = x151 | n1611 ;
  assign n19665 = x832 & n19664 ;
  assign n19666 = ~x745 & n19426 ;
  assign n19667 = x151 | n15332 ;
  assign n19668 = ~n19666 & n19667 ;
  assign n19669 = x39 | n19668 ;
  assign n19673 = n15405 | n19398 ;
  assign n19674 = x151 | n19673 ;
  assign n19675 = ~n15379 & n19674 ;
  assign n19676 = x215 & ~n19675 ;
  assign n19677 = ( n15405 & n19445 ) | ( n15405 & n19676 ) | ( n19445 & n19676 ) ;
  assign n19678 = x299 & ~n19677 ;
  assign n19679 = x151 | n15337 ;
  assign n19680 = ~n19431 & n19679 ;
  assign n19681 = x151 & n2263 ;
  assign n19682 = n15434 | n19681 ;
  assign n19683 = ( ~n15434 & n15471 ) | ( ~n15434 & n19682 ) | ( n15471 & n19682 ) ;
  assign n19684 = ( n19449 & ~n19680 ) | ( n19449 & n19683 ) | ( ~n19680 & n19683 ) ;
  assign n19685 = n19680 | n19684 ;
  assign n19686 = n19678 & n19685 ;
  assign n19687 = ( x745 & n19428 ) | ( x745 & ~n19686 ) | ( n19428 & ~n19686 ) ;
  assign n19688 = ~x745 & n19687 ;
  assign n19670 = ~x745 & n15485 ;
  assign n19671 = x151 | n15486 ;
  assign n19672 = n19670 | n19671 ;
  assign n19689 = n19688 ^ n19672 ^ 1'b0 ;
  assign n19690 = ( x39 & ~n19672 ) | ( x39 & n19688 ) | ( ~n19672 & n19688 ) ;
  assign n19691 = ( x39 & ~n19689 ) | ( x39 & n19690 ) | ( ~n19689 & n19690 ) ;
  assign n19692 = ( x38 & n19669 ) | ( x38 & ~n19691 ) | ( n19669 & ~n19691 ) ;
  assign n19693 = ~x38 & n19692 ;
  assign n19694 = ~x745 & x947 ;
  assign n19695 = n15644 & ~n19694 ;
  assign n19696 = x151 & ~n15653 ;
  assign n19697 = ( x38 & n19695 ) | ( x38 & n19696 ) | ( n19695 & n19696 ) ;
  assign n19698 = n19696 ^ n19695 ^ 1'b0 ;
  assign n19699 = ( x38 & n19697 ) | ( x38 & n19698 ) | ( n19697 & n19698 ) ;
  assign n19700 = ( x723 & n19693 ) | ( x723 & ~n19699 ) | ( n19693 & ~n19699 ) ;
  assign n19701 = ~n19693 & n19700 ;
  assign n19702 = x745 & x947 ;
  assign n19703 = ( x39 & n19568 ) | ( x39 & ~n19702 ) | ( n19568 & ~n19702 ) ;
  assign n19704 = ~x39 & n19703 ;
  assign n19705 = x151 | n15644 ;
  assign n19706 = x38 & n19705 ;
  assign n19707 = n19706 ^ n19704 ^ 1'b0 ;
  assign n19708 = ( n19704 & n19706 ) | ( n19704 & n19707 ) | ( n19706 & n19707 ) ;
  assign n19709 = ( x723 & ~n19704 ) | ( x723 & n19708 ) | ( ~n19704 & n19708 ) ;
  assign n19710 = n2263 | n19401 ;
  assign n19711 = n19679 & ~n19710 ;
  assign n19712 = n19683 | n19711 ;
  assign n19713 = n19373 | n19712 ;
  assign n19714 = ~n19676 & n19713 ;
  assign n19715 = ( x299 & n19388 ) | ( x299 & n19714 ) | ( n19388 & n19714 ) ;
  assign n19716 = n19714 ^ n19388 ^ 1'b0 ;
  assign n19717 = ( x299 & n19715 ) | ( x299 & n19716 ) | ( n19715 & n19716 ) ;
  assign n19718 = ( x151 & n19392 ) | ( x151 & ~n19409 ) | ( n19392 & ~n19409 ) ;
  assign n19719 = ( x745 & n19717 ) | ( x745 & ~n19718 ) | ( n19717 & ~n19718 ) ;
  assign n19720 = ~n19717 & n19719 ;
  assign n19721 = ( n2264 & ~n19432 ) | ( n2264 & n19711 ) | ( ~n19432 & n19711 ) ;
  assign n19722 = n19683 | n19721 ;
  assign n19723 = n19722 ^ n19676 ^ 1'b0 ;
  assign n19724 = ( x299 & n19676 ) | ( x299 & ~n19722 ) | ( n19676 & ~n19722 ) ;
  assign n19725 = ( x299 & ~n19723 ) | ( x299 & n19724 ) | ( ~n19723 & n19724 ) ;
  assign n19726 = x151 & ~n19351 ;
  assign n19727 = n19367 | n19726 ;
  assign n19728 = n19727 ^ n19725 ^ 1'b0 ;
  assign n19729 = ( n19725 & n19727 ) | ( n19725 & n19728 ) | ( n19727 & n19728 ) ;
  assign n19730 = ( x745 & ~n19725 ) | ( x745 & n19729 ) | ( ~n19725 & n19729 ) ;
  assign n19731 = ( x39 & n19720 ) | ( x39 & n19730 ) | ( n19720 & n19730 ) ;
  assign n19732 = ~n19720 & n19731 ;
  assign n19733 = x39 | n19397 ;
  assign n19734 = n19668 & ~n19733 ;
  assign n19735 = ( ~x38 & n19732 ) | ( ~x38 & n19734 ) | ( n19732 & n19734 ) ;
  assign n19736 = ~x38 & n19735 ;
  assign n19737 = ( ~n19701 & n19709 ) | ( ~n19701 & n19736 ) | ( n19709 & n19736 ) ;
  assign n19738 = ~n19701 & n19737 ;
  assign n19739 = ( n2069 & n7318 ) | ( n2069 & ~n19738 ) | ( n7318 & ~n19738 ) ;
  assign n19740 = n19738 | n19739 ;
  assign n19741 = ~x151 & n8793 ;
  assign n19742 = ( x832 & n19740 ) | ( x832 & ~n19741 ) | ( n19740 & ~n19741 ) ;
  assign n19743 = ~x832 & n19742 ;
  assign n19744 = ~x723 & n19256 ;
  assign n19745 = n19694 | n19744 ;
  assign n19746 = n1611 & n19745 ;
  assign n19747 = ~n19743 & n19746 ;
  assign n19748 = ( n19665 & n19743 ) | ( n19665 & ~n19747 ) | ( n19743 & ~n19747 ) ;
  assign n19749 = ~x152 & n8793 ;
  assign n19750 = x832 | n19749 ;
  assign n19751 = x759 & x947 ;
  assign n19752 = x39 | n19751 ;
  assign n19753 = n15333 & n19752 ;
  assign n19754 = x152 & ~n15332 ;
  assign n19755 = n19753 | n19754 ;
  assign n19756 = n19397 | n19755 ;
  assign n19757 = x152 | n15482 ;
  assign n19758 = n19362 & n19757 ;
  assign n19759 = x299 | n19758 ;
  assign n19760 = x152 | n15337 ;
  assign n19761 = ~n5055 & n15337 ;
  assign n19762 = n19760 & ~n19761 ;
  assign n19763 = n1359 | n19762 ;
  assign n19764 = x152 | n15476 ;
  assign n19765 = ~x947 & n15476 ;
  assign n19766 = n1359 & ~n19765 ;
  assign n19767 = n19764 & n19766 ;
  assign n19768 = n5055 & n15476 ;
  assign n19769 = n1359 & ~n19768 ;
  assign n19770 = ~n19767 & n19769 ;
  assign n19771 = ( x223 & n19763 ) | ( x223 & ~n19770 ) | ( n19763 & ~n19770 ) ;
  assign n19772 = ~x223 & n19771 ;
  assign n19773 = n19363 & n19757 ;
  assign n19774 = ( ~n19759 & n19772 ) | ( ~n19759 & n19773 ) | ( n19772 & n19773 ) ;
  assign n19775 = n19759 | n19774 ;
  assign n19776 = n2263 | n19762 ;
  assign n19777 = ~x215 & n19776 ;
  assign n19778 = n2263 & ~n19399 ;
  assign n19779 = x152 & ~n19371 ;
  assign n19780 = n19778 & ~n19779 ;
  assign n19781 = ~n15434 & n19780 ;
  assign n19782 = n19777 & ~n19781 ;
  assign n19783 = x152 | n15379 ;
  assign n19784 = n19368 & n19783 ;
  assign n19785 = ( x299 & n19782 ) | ( x299 & ~n19784 ) | ( n19782 & ~n19784 ) ;
  assign n19786 = ~n19782 & n19785 ;
  assign n19787 = x759 & ~n19786 ;
  assign n19788 = n19775 & n19787 ;
  assign n19789 = n15476 & ~n19256 ;
  assign n19790 = n1359 & ~n19789 ;
  assign n19791 = n19764 & n19790 ;
  assign n19792 = ~n1359 & n19430 ;
  assign n19793 = n19792 ^ n19763 ^ n1359 ;
  assign n19794 = ( ~x223 & n19791 ) | ( ~x223 & n19793 ) | ( n19791 & n19793 ) ;
  assign n19795 = ~x223 & n19794 ;
  assign n19796 = ( x299 & n19773 ) | ( x299 & ~n19795 ) | ( n19773 & ~n19795 ) ;
  assign n19797 = n19795 | n19796 ;
  assign n19798 = ~n19369 & n19777 ;
  assign n19799 = ~n19780 & n19798 ;
  assign n19800 = n19256 | n19347 ;
  assign n19801 = n19784 & n19800 ;
  assign n19802 = ( x299 & n19799 ) | ( x299 & ~n19801 ) | ( n19799 & ~n19801 ) ;
  assign n19803 = ~n19799 & n19802 ;
  assign n19804 = ( x759 & n19797 ) | ( x759 & ~n19803 ) | ( n19797 & ~n19803 ) ;
  assign n19805 = ~x759 & n19804 ;
  assign n19806 = ( x39 & n19788 ) | ( x39 & ~n19805 ) | ( n19788 & ~n19805 ) ;
  assign n19807 = ~n19788 & n19806 ;
  assign n19808 = ( x38 & n19756 ) | ( x38 & ~n19807 ) | ( n19756 & ~n19807 ) ;
  assign n19809 = ~x38 & n19808 ;
  assign n19810 = x152 | n15644 ;
  assign n19811 = n15340 & ~n19256 ;
  assign n19812 = ~n19752 & n19811 ;
  assign n19813 = x38 & ~n19812 ;
  assign n19814 = n19810 & n19813 ;
  assign n19815 = ( x696 & n19809 ) | ( x696 & ~n19814 ) | ( n19809 & ~n19814 ) ;
  assign n19816 = ~n19809 & n19815 ;
  assign n19817 = x152 | n15653 ;
  assign n19818 = n19817 ^ x696 ^ 1'b0 ;
  assign n19819 = n15644 & ~n19751 ;
  assign n19820 = x38 & ~n19819 ;
  assign n19821 = ( n19817 & ~n19818 ) | ( n19817 & n19820 ) | ( ~n19818 & n19820 ) ;
  assign n19822 = ( x696 & n19818 ) | ( x696 & n19821 ) | ( n19818 & n19821 ) ;
  assign n19823 = x759 | n15486 ;
  assign n19824 = x152 & ~n19823 ;
  assign n19825 = ~x947 & n15337 ;
  assign n19826 = n19760 & ~n19825 ;
  assign n19827 = ~n1359 & n19826 ;
  assign n19828 = n19767 | n19827 ;
  assign n19829 = x223 | n19828 ;
  assign n19830 = ( ~x223 & n19759 ) | ( ~x223 & n19829 ) | ( n19759 & n19829 ) ;
  assign n19831 = x152 & n19445 ;
  assign n19832 = n2263 | n19826 ;
  assign n19833 = ( n19399 & n19433 ) | ( n19399 & n19780 ) | ( n19433 & n19780 ) ;
  assign n19834 = ( x215 & n19832 ) | ( x215 & ~n19833 ) | ( n19832 & ~n19833 ) ;
  assign n19835 = ~x215 & n19834 ;
  assign n19836 = ( n19429 & n19831 ) | ( n19429 & ~n19835 ) | ( n19831 & ~n19835 ) ;
  assign n19837 = ~n19831 & n19836 ;
  assign n19838 = x759 & ~n19837 ;
  assign n19839 = n19830 & n19838 ;
  assign n19840 = ( x39 & n19824 ) | ( x39 & ~n19839 ) | ( n19824 & ~n19839 ) ;
  assign n19841 = ~n19824 & n19840 ;
  assign n19842 = ( x38 & n19755 ) | ( x38 & ~n19841 ) | ( n19755 & ~n19841 ) ;
  assign n19843 = ~x38 & n19842 ;
  assign n19844 = ( ~n19816 & n19822 ) | ( ~n19816 & n19843 ) | ( n19822 & n19843 ) ;
  assign n19845 = ~n19816 & n19844 ;
  assign n19846 = ( n8793 & ~n19750 ) | ( n8793 & n19845 ) | ( ~n19750 & n19845 ) ;
  assign n19847 = ~n19750 & n19846 ;
  assign n19848 = n1611 & ~n19751 ;
  assign n19849 = x696 & n19256 ;
  assign n19850 = n19848 & ~n19849 ;
  assign n19851 = x152 | n1611 ;
  assign n19852 = x832 & n19851 ;
  assign n19853 = n19852 ^ n19850 ^ 1'b0 ;
  assign n19854 = ( n19850 & n19852 ) | ( n19850 & n19853 ) | ( n19852 & n19853 ) ;
  assign n19855 = ( n19847 & ~n19850 ) | ( n19847 & n19854 ) | ( ~n19850 & n19854 ) ;
  assign n19856 = x766 & x947 ;
  assign n19857 = n1611 & ~n19856 ;
  assign n19858 = x700 & n19256 ;
  assign n19859 = n19857 & ~n19858 ;
  assign n19860 = x153 & ~n1611 ;
  assign n19861 = ( x832 & n19859 ) | ( x832 & ~n19860 ) | ( n19859 & ~n19860 ) ;
  assign n19862 = ~n19859 & n19861 ;
  assign n19863 = x57 & x153 ;
  assign n19864 = x832 | n19863 ;
  assign n19865 = ~x766 & x947 ;
  assign n19866 = ( x39 & n19568 ) | ( x39 & ~n19865 ) | ( n19568 & ~n19865 ) ;
  assign n19867 = ~x39 & n19866 ;
  assign n19868 = x153 | n15644 ;
  assign n19869 = ( x38 & n19867 ) | ( x38 & n19868 ) | ( n19867 & n19868 ) ;
  assign n19870 = ~n19867 & n19869 ;
  assign n19871 = x153 | n15484 ;
  assign n19872 = ~n19409 & n19871 ;
  assign n19873 = x153 & n2263 ;
  assign n19874 = n15434 | n19873 ;
  assign n19875 = ( ~n15434 & n15471 ) | ( ~n15434 & n19874 ) | ( n15471 & n19874 ) ;
  assign n19876 = x153 | n15337 ;
  assign n19877 = ~n19710 & n19876 ;
  assign n19878 = n19372 | n19877 ;
  assign n19879 = ( ~x215 & n19875 ) | ( ~x215 & n19878 ) | ( n19875 & n19878 ) ;
  assign n19880 = ~x215 & n19879 ;
  assign n19881 = x153 & ~n15379 ;
  assign n19882 = n19368 & ~n19881 ;
  assign n19883 = n19882 ^ n19388 ^ x215 ;
  assign n19884 = ( x299 & n19880 ) | ( x299 & n19883 ) | ( n19880 & n19883 ) ;
  assign n19885 = n19883 ^ n19880 ^ 1'b0 ;
  assign n19886 = ( x299 & n19884 ) | ( x299 & n19885 ) | ( n19884 & n19885 ) ;
  assign n19887 = ( x766 & ~n19872 ) | ( x766 & n19886 ) | ( ~n19872 & n19886 ) ;
  assign n19888 = n19872 | n19887 ;
  assign n19891 = ( n2264 & ~n19432 ) | ( n2264 & n19877 ) | ( ~n19432 & n19877 ) ;
  assign n19892 = n19875 | n19891 ;
  assign n19893 = n19892 ^ n19882 ^ 1'b0 ;
  assign n19894 = ( x299 & n19882 ) | ( x299 & ~n19892 ) | ( n19882 & ~n19892 ) ;
  assign n19895 = ( x299 & ~n19893 ) | ( x299 & n19894 ) | ( ~n19893 & n19894 ) ;
  assign n19889 = x153 & ~n19351 ;
  assign n19890 = n19367 | n19889 ;
  assign n19896 = n19895 ^ n19890 ^ 1'b0 ;
  assign n19897 = ( x766 & ~n19890 ) | ( x766 & n19895 ) | ( ~n19890 & n19895 ) ;
  assign n19898 = ( x766 & ~n19896 ) | ( x766 & n19897 ) | ( ~n19896 & n19897 ) ;
  assign n19899 = x39 & ~n19898 ;
  assign n19900 = n19888 & n19899 ;
  assign n19901 = x39 | n19426 ;
  assign n19902 = ~x766 & n15487 ;
  assign n19903 = n19901 & ~n19902 ;
  assign n19904 = x153 | n15332 ;
  assign n19905 = ~n19903 & n19904 ;
  assign n19906 = ~n19397 & n19905 ;
  assign n19907 = ( ~x38 & n19900 ) | ( ~x38 & n19906 ) | ( n19900 & n19906 ) ;
  assign n19908 = ~x38 & n19907 ;
  assign n19909 = ( x700 & n19870 ) | ( x700 & n19908 ) | ( n19870 & n19908 ) ;
  assign n19910 = n19908 ^ n19870 ^ 1'b0 ;
  assign n19911 = ( x700 & n19909 ) | ( x700 & n19910 ) | ( n19909 & n19910 ) ;
  assign n19912 = x153 & ~n15653 ;
  assign n19913 = ~n5017 & n19857 ;
  assign n19914 = x38 & ~n19913 ;
  assign n19915 = n19914 ^ n19912 ^ 1'b0 ;
  assign n19916 = ( n19912 & n19914 ) | ( n19912 & n19915 ) | ( n19914 & n19915 ) ;
  assign n19917 = ( x700 & ~n19912 ) | ( x700 & n19916 ) | ( ~n19912 & n19916 ) ;
  assign n19918 = ~n19428 & n19871 ;
  assign n19919 = n19445 & ~n19881 ;
  assign n19920 = ~n19431 & n19876 ;
  assign n19921 = n19875 | n19920 ;
  assign n19922 = n19449 | n19921 ;
  assign n19923 = ( x299 & n19919 ) | ( x299 & n19922 ) | ( n19919 & n19922 ) ;
  assign n19924 = ~n19919 & n19923 ;
  assign n19925 = ( x766 & n19918 ) | ( x766 & ~n19924 ) | ( n19918 & ~n19924 ) ;
  assign n19926 = ~n19918 & n19925 ;
  assign n19927 = x153 | x766 ;
  assign n19928 = n15486 | n19927 ;
  assign n19929 = ( x39 & n19926 ) | ( x39 & n19928 ) | ( n19926 & n19928 ) ;
  assign n19930 = ~n19926 & n19929 ;
  assign n19931 = x38 | n19905 ;
  assign n19932 = ( ~n19917 & n19930 ) | ( ~n19917 & n19931 ) | ( n19930 & n19931 ) ;
  assign n19933 = ~n19917 & n19932 ;
  assign n19934 = ( n19509 & ~n19911 ) | ( n19509 & n19933 ) | ( ~n19911 & n19933 ) ;
  assign n19935 = n19911 | n19934 ;
  assign n19936 = ~x153 & n19509 ;
  assign n19937 = ( x57 & n19935 ) | ( x57 & ~n19936 ) | ( n19935 & ~n19936 ) ;
  assign n19938 = ~x57 & n19937 ;
  assign n19939 = ( ~n19862 & n19864 ) | ( ~n19862 & n19938 ) | ( n19864 & n19938 ) ;
  assign n19940 = ~n19862 & n19939 ;
  assign n19941 = x154 | n1611 ;
  assign n19942 = x832 & n19941 ;
  assign n19943 = x154 & n19354 ;
  assign n19944 = x154 | n19378 ;
  assign n19945 = ( x39 & n19943 ) | ( x39 & n19944 ) | ( n19943 & n19944 ) ;
  assign n19946 = ~n19943 & n19945 ;
  assign n19947 = x154 | n15332 ;
  assign n19948 = ~n19733 & n19947 ;
  assign n19949 = ~n19346 & n19948 ;
  assign n19950 = ( ~x38 & n19946 ) | ( ~x38 & n19949 ) | ( n19946 & n19949 ) ;
  assign n19951 = ~x38 & n19950 ;
  assign n19952 = x154 | n15644 ;
  assign n19953 = n19344 & n19952 ;
  assign n19954 = ( x742 & ~n19951 ) | ( x742 & n19953 ) | ( ~n19951 & n19953 ) ;
  assign n19955 = n19951 | n19954 ;
  assign n19956 = x154 & n19410 ;
  assign n19957 = x39 & ~n19956 ;
  assign n19958 = x154 | n19393 ;
  assign n19959 = n19957 & n19958 ;
  assign n19960 = ( ~x38 & n19948 ) | ( ~x38 & n19959 ) | ( n19948 & n19959 ) ;
  assign n19961 = ~x38 & n19960 ;
  assign n19962 = n19418 & n19952 ;
  assign n19963 = ( x742 & n19961 ) | ( x742 & ~n19962 ) | ( n19961 & ~n19962 ) ;
  assign n19964 = ~n19961 & n19963 ;
  assign n19965 = ( x704 & n19955 ) | ( x704 & ~n19964 ) | ( n19955 & ~n19964 ) ;
  assign n19966 = ~x704 & n19965 ;
  assign n19967 = ~x154 & x742 ;
  assign n19968 = ~n15655 & n19967 ;
  assign n19969 = x154 & n19436 ;
  assign n19970 = x154 | n19453 ;
  assign n19971 = ( x39 & n19969 ) | ( x39 & n19970 ) | ( n19969 & n19970 ) ;
  assign n19972 = ~n19969 & n19971 ;
  assign n19973 = ~n19901 & n19947 ;
  assign n19974 = ( ~x38 & n19972 ) | ( ~x38 & n19973 ) | ( n19972 & n19973 ) ;
  assign n19975 = ~x38 & n19974 ;
  assign n19976 = x154 | n15653 ;
  assign n19977 = n19425 & n19976 ;
  assign n19978 = ( x742 & ~n19975 ) | ( x742 & n19977 ) | ( ~n19975 & n19977 ) ;
  assign n19979 = n19975 | n19978 ;
  assign n19980 = ( x704 & n19968 ) | ( x704 & n19979 ) | ( n19968 & n19979 ) ;
  assign n19981 = ~n19968 & n19980 ;
  assign n19982 = ( n8793 & ~n19966 ) | ( n8793 & n19981 ) | ( ~n19966 & n19981 ) ;
  assign n19983 = n19966 | n19982 ;
  assign n19984 = ~x154 & n8793 ;
  assign n19985 = ( x832 & n19983 ) | ( x832 & ~n19984 ) | ( n19983 & ~n19984 ) ;
  assign n19986 = ~x832 & n19985 ;
  assign n19987 = ~x704 & n19256 ;
  assign n19988 = ~x742 & x947 ;
  assign n19989 = ( n1611 & n19987 ) | ( n1611 & n19988 ) | ( n19987 & n19988 ) ;
  assign n19990 = n19988 ^ n19987 ^ 1'b0 ;
  assign n19991 = ( n1611 & n19989 ) | ( n1611 & n19990 ) | ( n19989 & n19990 ) ;
  assign n19992 = ~n19986 & n19991 ;
  assign n19993 = ( n19942 & n19986 ) | ( n19942 & ~n19992 ) | ( n19986 & ~n19992 ) ;
  assign n19994 = x155 | n1611 ;
  assign n19995 = x832 & n19994 ;
  assign n19996 = ~x757 & n19440 ;
  assign n19997 = x686 & ~n19996 ;
  assign n19998 = n8793 | n19997 ;
  assign n19999 = n19413 & ~n19418 ;
  assign n20000 = x757 & n19999 ;
  assign n20001 = n19356 ^ x38 ^ 1'b0 ;
  assign n20002 = ( n19343 & n19356 ) | ( n19343 & n20001 ) | ( n19356 & n20001 ) ;
  assign n20003 = ~x757 & n20002 ;
  assign n20004 = ( x686 & ~n20000 ) | ( x686 & n20003 ) | ( ~n20000 & n20003 ) ;
  assign n20005 = n20000 | n20004 ;
  assign n20006 = x155 & ~n20005 ;
  assign n20007 = ( x155 & n19998 ) | ( x155 & n20006 ) | ( n19998 & n20006 ) ;
  assign n20008 = x757 & ~n15655 ;
  assign n20009 = x686 & ~n20008 ;
  assign n20010 = ~x38 & n19396 ;
  assign n20011 = n19419 | n20010 ;
  assign n20012 = x757 & ~n20011 ;
  assign n20013 = n19382 ^ x38 ^ 1'b0 ;
  assign n20014 = ( n19341 & n19382 ) | ( n19341 & n20013 ) | ( n19382 & n20013 ) ;
  assign n20015 = x757 | n20014 ;
  assign n20016 = ( x686 & ~n20012 ) | ( x686 & n20015 ) | ( ~n20012 & n20015 ) ;
  assign n20017 = ~x686 & n20016 ;
  assign n20018 = x757 | n19459 ;
  assign n20019 = n20017 ^ n20009 ^ 1'b0 ;
  assign n20020 = ( ~n20009 & n20018 ) | ( ~n20009 & n20019 ) | ( n20018 & n20019 ) ;
  assign n20021 = ( n20009 & n20017 ) | ( n20009 & n20020 ) | ( n20017 & n20020 ) ;
  assign n20022 = ( x155 & ~n8793 ) | ( x155 & n20021 ) | ( ~n8793 & n20021 ) ;
  assign n20023 = ~x155 & n20022 ;
  assign n20024 = ( ~x832 & n20007 ) | ( ~x832 & n20023 ) | ( n20007 & n20023 ) ;
  assign n20025 = ~x832 & n20024 ;
  assign n20026 = ~x686 & n19256 ;
  assign n20027 = ~x757 & x947 ;
  assign n20028 = ( n1611 & n20026 ) | ( n1611 & n20027 ) | ( n20026 & n20027 ) ;
  assign n20029 = n20027 ^ n20026 ^ 1'b0 ;
  assign n20030 = ( n1611 & n20028 ) | ( n1611 & n20029 ) | ( n20028 & n20029 ) ;
  assign n20031 = ~n20025 & n20030 ;
  assign n20032 = ( n19995 & n20025 ) | ( n19995 & ~n20031 ) | ( n20025 & ~n20031 ) ;
  assign n20033 = x156 | n1611 ;
  assign n20034 = x832 & n20033 ;
  assign n20035 = ~x741 & n20014 ;
  assign n20036 = x741 & n20011 ;
  assign n20037 = ( x724 & ~n20035 ) | ( x724 & n20036 ) | ( ~n20035 & n20036 ) ;
  assign n20038 = n20035 | n20037 ;
  assign n20039 = ~x741 & n19459 ;
  assign n20040 = x741 & n15655 ;
  assign n20041 = x724 & ~n20040 ;
  assign n20042 = n20041 ^ n20039 ^ 1'b0 ;
  assign n20043 = ( n20039 & n20041 ) | ( n20039 & n20042 ) | ( n20041 & n20042 ) ;
  assign n20044 = ( n8793 & ~n20039 ) | ( n8793 & n20043 ) | ( ~n20039 & n20043 ) ;
  assign n20045 = ( x156 & n20038 ) | ( x156 & ~n20044 ) | ( n20038 & ~n20044 ) ;
  assign n20046 = n20045 ^ n20038 ^ 1'b0 ;
  assign n20047 = ( x156 & n20045 ) | ( x156 & ~n20046 ) | ( n20045 & ~n20046 ) ;
  assign n20048 = x741 & ~n19999 ;
  assign n20049 = x741 | n20002 ;
  assign n20050 = ( x724 & ~n20048 ) | ( x724 & n20049 ) | ( ~n20048 & n20049 ) ;
  assign n20051 = ~x724 & n20050 ;
  assign n20052 = x724 & ~x741 ;
  assign n20053 = n20051 ^ n19440 ^ 1'b0 ;
  assign n20054 = ( ~n19440 & n20052 ) | ( ~n19440 & n20053 ) | ( n20052 & n20053 ) ;
  assign n20055 = ( n19440 & n20051 ) | ( n19440 & n20054 ) | ( n20051 & n20054 ) ;
  assign n20056 = x156 & ~n8793 ;
  assign n20057 = n20055 & n20056 ;
  assign n20058 = ( x832 & n20047 ) | ( x832 & ~n20057 ) | ( n20047 & ~n20057 ) ;
  assign n20059 = ~x832 & n20058 ;
  assign n20060 = ~x724 & n19256 ;
  assign n20061 = ~x741 & x947 ;
  assign n20062 = ( n1611 & n20060 ) | ( n1611 & n20061 ) | ( n20060 & n20061 ) ;
  assign n20063 = n20061 ^ n20060 ^ 1'b0 ;
  assign n20064 = ( n1611 & n20062 ) | ( n1611 & n20063 ) | ( n20062 & n20063 ) ;
  assign n20065 = ~n20059 & n20064 ;
  assign n20066 = ( n20034 & n20059 ) | ( n20034 & ~n20065 ) | ( n20059 & ~n20065 ) ;
  assign n20067 = x157 | n1611 ;
  assign n20068 = x832 & n20067 ;
  assign n20070 = ~x760 & x947 ;
  assign n20087 = n15644 & ~n20070 ;
  assign n20088 = x157 & ~n15653 ;
  assign n20089 = ( x38 & n20087 ) | ( x38 & ~n20088 ) | ( n20087 & ~n20088 ) ;
  assign n20090 = ~n20087 & n20089 ;
  assign n20069 = x157 | n15332 ;
  assign n20071 = n15332 & n20070 ;
  assign n20072 = ( x39 & n20069 ) | ( x39 & ~n20071 ) | ( n20069 & ~n20071 ) ;
  assign n20073 = ~x39 & n20072 ;
  assign n20074 = ~x157 & x760 ;
  assign n20075 = ~n15486 & n20074 ;
  assign n20076 = x39 & ~n20075 ;
  assign n20077 = x157 | n15484 ;
  assign n20078 = ~n19428 & n20077 ;
  assign n20079 = n12320 | n19435 ;
  assign n20080 = x157 | n19451 ;
  assign n20081 = n20079 & n20080 ;
  assign n20082 = ( x760 & ~n20078 ) | ( x760 & n20081 ) | ( ~n20078 & n20081 ) ;
  assign n20083 = n20078 | n20082 ;
  assign n20084 = n20076 & n20083 ;
  assign n20085 = ( x38 & ~n20073 ) | ( x38 & n20084 ) | ( ~n20073 & n20084 ) ;
  assign n20086 = n20073 | n20085 ;
  assign n20091 = n20090 ^ n20086 ^ 1'b0 ;
  assign n20092 = ( x688 & ~n20086 ) | ( x688 & n20090 ) | ( ~n20086 & n20090 ) ;
  assign n20093 = ( x688 & ~n20091 ) | ( x688 & n20092 ) | ( ~n20091 & n20092 ) ;
  assign n20094 = x760 & x947 ;
  assign n20095 = ( x39 & n19568 ) | ( x39 & ~n20094 ) | ( n19568 & ~n20094 ) ;
  assign n20096 = ~x39 & n20095 ;
  assign n20097 = x157 | n15644 ;
  assign n20098 = x38 & n20097 ;
  assign n20099 = n20098 ^ n20096 ^ 1'b0 ;
  assign n20100 = ( n20096 & n20098 ) | ( n20096 & n20099 ) | ( n20098 & n20099 ) ;
  assign n20101 = ( x688 & ~n20096 ) | ( x688 & n20100 ) | ( ~n20096 & n20100 ) ;
  assign n20102 = x760 | n19354 ;
  assign n20103 = x760 & ~n19410 ;
  assign n20104 = x157 & ~n20103 ;
  assign n20105 = n20102 & n20104 ;
  assign n20106 = ~x760 & n19378 ;
  assign n20107 = x760 & n19393 ;
  assign n20108 = ( x157 & ~n20106 ) | ( x157 & n20107 ) | ( ~n20106 & n20107 ) ;
  assign n20109 = n20106 | n20108 ;
  assign n20110 = ( x39 & n20105 ) | ( x39 & n20109 ) | ( n20105 & n20109 ) ;
  assign n20111 = ~n20105 & n20110 ;
  assign n20112 = ~n19397 & n20073 ;
  assign n20113 = ( ~x38 & n20111 ) | ( ~x38 & n20112 ) | ( n20111 & n20112 ) ;
  assign n20114 = ~x38 & n20113 ;
  assign n20115 = ( ~n20093 & n20101 ) | ( ~n20093 & n20114 ) | ( n20101 & n20114 ) ;
  assign n20116 = ~n20093 & n20115 ;
  assign n20117 = ( n2069 & n7318 ) | ( n2069 & ~n20116 ) | ( n7318 & ~n20116 ) ;
  assign n20118 = n20116 | n20117 ;
  assign n20119 = ~x157 & n8793 ;
  assign n20120 = ( x832 & n20118 ) | ( x832 & ~n20119 ) | ( n20118 & ~n20119 ) ;
  assign n20121 = ~x832 & n20120 ;
  assign n20122 = ~x688 & n19256 ;
  assign n20123 = n20070 | n20122 ;
  assign n20124 = n1611 & n20123 ;
  assign n20125 = ~n20121 & n20124 ;
  assign n20126 = ( n20068 & n20121 ) | ( n20068 & ~n20125 ) | ( n20121 & ~n20125 ) ;
  assign n20127 = ~x753 & x947 ;
  assign n20128 = n15644 & ~n20127 ;
  assign n20129 = x158 & ~n15653 ;
  assign n20130 = ( x38 & n20128 ) | ( x38 & n20129 ) | ( n20128 & n20129 ) ;
  assign n20131 = n20129 ^ n20128 ^ 1'b0 ;
  assign n20132 = ( x38 & n20130 ) | ( x38 & n20131 ) | ( n20130 & n20131 ) ;
  assign n20133 = ~x158 & x753 ;
  assign n20134 = ~n15486 & n20133 ;
  assign n20135 = ~x158 & n19453 ;
  assign n20136 = x158 & ~n19436 ;
  assign n20137 = ( x753 & ~n20135 ) | ( x753 & n20136 ) | ( ~n20135 & n20136 ) ;
  assign n20138 = n20135 | n20137 ;
  assign n20139 = x39 & ~n20138 ;
  assign n20140 = ( x39 & n20134 ) | ( x39 & n20139 ) | ( n20134 & n20139 ) ;
  assign n20141 = n15332 ^ x753 ^ 1'b0 ;
  assign n20142 = ( x158 & x753 ) | ( x158 & ~n20141 ) | ( x753 & ~n20141 ) ;
  assign n20143 = ( x39 & n19443 ) | ( x39 & ~n20142 ) | ( n19443 & ~n20142 ) ;
  assign n20144 = n20142 | n20143 ;
  assign n20145 = ( x38 & ~n20140 ) | ( x38 & n20144 ) | ( ~n20140 & n20144 ) ;
  assign n20146 = ~x38 & n20145 ;
  assign n20147 = ( x702 & n20132 ) | ( x702 & ~n20146 ) | ( n20132 & ~n20146 ) ;
  assign n20148 = ~n20132 & n20147 ;
  assign n20149 = x753 & x947 ;
  assign n20150 = ( x39 & n19568 ) | ( x39 & ~n20149 ) | ( n19568 & ~n20149 ) ;
  assign n20151 = ~x39 & n20150 ;
  assign n20152 = x158 | n15644 ;
  assign n20153 = x38 & n20152 ;
  assign n20154 = n20153 ^ n20151 ^ 1'b0 ;
  assign n20155 = ( n20151 & n20153 ) | ( n20151 & n20154 ) | ( n20153 & n20154 ) ;
  assign n20156 = ( x702 & ~n20151 ) | ( x702 & n20155 ) | ( ~n20151 & n20155 ) ;
  assign n20161 = x158 & ~n19410 ;
  assign n20162 = ~x158 & n19393 ;
  assign n20163 = ( x753 & n20161 ) | ( x753 & ~n20162 ) | ( n20161 & ~n20162 ) ;
  assign n20164 = ~n20161 & n20163 ;
  assign n20157 = ~x158 & n19378 ;
  assign n20158 = x158 & ~n19354 ;
  assign n20159 = ( x753 & ~n20157 ) | ( x753 & n20158 ) | ( ~n20157 & n20158 ) ;
  assign n20160 = n20157 | n20159 ;
  assign n20165 = n20164 ^ n20160 ^ 1'b0 ;
  assign n20166 = ( x39 & ~n20160 ) | ( x39 & n20164 ) | ( ~n20160 & n20164 ) ;
  assign n20167 = ( x39 & ~n20165 ) | ( x39 & n20166 ) | ( ~n20165 & n20166 ) ;
  assign n20168 = x158 & ~n15332 ;
  assign n20169 = n19394 & ~n20127 ;
  assign n20170 = ( x39 & ~n20168 ) | ( x39 & n20169 ) | ( ~n20168 & n20169 ) ;
  assign n20171 = n20168 | n20170 ;
  assign n20172 = ( x38 & ~n20167 ) | ( x38 & n20171 ) | ( ~n20167 & n20171 ) ;
  assign n20173 = ~x38 & n20172 ;
  assign n20174 = ( ~n20148 & n20156 ) | ( ~n20148 & n20173 ) | ( n20156 & n20173 ) ;
  assign n20175 = ~n20148 & n20174 ;
  assign n20176 = ( n2069 & n7318 ) | ( n2069 & ~n20175 ) | ( n7318 & ~n20175 ) ;
  assign n20177 = n20175 | n20176 ;
  assign n20178 = ~x702 & n19256 ;
  assign n20179 = n20127 | n20178 ;
  assign n20180 = n1611 & n20179 ;
  assign n20181 = x158 | n1611 ;
  assign n20182 = ( x832 & n20180 ) | ( x832 & n20181 ) | ( n20180 & n20181 ) ;
  assign n20183 = ~n20180 & n20182 ;
  assign n20184 = ~x158 & n8793 ;
  assign n20185 = x832 | n20184 ;
  assign n20186 = ~n20183 & n20185 ;
  assign n20187 = ( n20177 & n20183 ) | ( n20177 & ~n20186 ) | ( n20183 & ~n20186 ) ;
  assign n20188 = ~x754 & x947 ;
  assign n20189 = n15644 & ~n20188 ;
  assign n20190 = x159 & ~n15653 ;
  assign n20191 = ( x38 & n20189 ) | ( x38 & n20190 ) | ( n20189 & n20190 ) ;
  assign n20192 = n20190 ^ n20189 ^ 1'b0 ;
  assign n20193 = ( x38 & n20191 ) | ( x38 & n20192 ) | ( n20191 & n20192 ) ;
  assign n20194 = ~x159 & x754 ;
  assign n20195 = ~n15486 & n20194 ;
  assign n20196 = ~x159 & n19453 ;
  assign n20197 = x159 & ~n19436 ;
  assign n20198 = ( x754 & ~n20196 ) | ( x754 & n20197 ) | ( ~n20196 & n20197 ) ;
  assign n20199 = n20196 | n20198 ;
  assign n20200 = x39 & ~n20199 ;
  assign n20201 = ( x39 & n20195 ) | ( x39 & n20200 ) | ( n20195 & n20200 ) ;
  assign n20202 = n15332 ^ x754 ^ 1'b0 ;
  assign n20203 = ( x159 & x754 ) | ( x159 & ~n20202 ) | ( x754 & ~n20202 ) ;
  assign n20204 = ( x39 & n19443 ) | ( x39 & ~n20203 ) | ( n19443 & ~n20203 ) ;
  assign n20205 = n20203 | n20204 ;
  assign n20206 = ( x38 & ~n20201 ) | ( x38 & n20205 ) | ( ~n20201 & n20205 ) ;
  assign n20207 = ~x38 & n20206 ;
  assign n20208 = ( x709 & n20193 ) | ( x709 & ~n20207 ) | ( n20193 & ~n20207 ) ;
  assign n20209 = ~n20193 & n20208 ;
  assign n20210 = x754 & x947 ;
  assign n20211 = ( x39 & n19568 ) | ( x39 & ~n20210 ) | ( n19568 & ~n20210 ) ;
  assign n20212 = ~x39 & n20211 ;
  assign n20213 = x159 | n15644 ;
  assign n20214 = x38 & n20213 ;
  assign n20215 = n20214 ^ n20212 ^ 1'b0 ;
  assign n20216 = ( n20212 & n20214 ) | ( n20212 & n20215 ) | ( n20214 & n20215 ) ;
  assign n20217 = ( x709 & ~n20212 ) | ( x709 & n20216 ) | ( ~n20212 & n20216 ) ;
  assign n20222 = x159 & ~n19410 ;
  assign n20223 = ~x159 & n19393 ;
  assign n20224 = ( x754 & n20222 ) | ( x754 & ~n20223 ) | ( n20222 & ~n20223 ) ;
  assign n20225 = ~n20222 & n20224 ;
  assign n20218 = ~x159 & n19378 ;
  assign n20219 = x159 & ~n19354 ;
  assign n20220 = ( x754 & ~n20218 ) | ( x754 & n20219 ) | ( ~n20218 & n20219 ) ;
  assign n20221 = n20218 | n20220 ;
  assign n20226 = n20225 ^ n20221 ^ 1'b0 ;
  assign n20227 = ( x39 & ~n20221 ) | ( x39 & n20225 ) | ( ~n20221 & n20225 ) ;
  assign n20228 = ( x39 & ~n20226 ) | ( x39 & n20227 ) | ( ~n20226 & n20227 ) ;
  assign n20229 = x159 & ~n15332 ;
  assign n20230 = n19394 & ~n20188 ;
  assign n20231 = ( x39 & ~n20229 ) | ( x39 & n20230 ) | ( ~n20229 & n20230 ) ;
  assign n20232 = n20229 | n20231 ;
  assign n20233 = ( x38 & ~n20228 ) | ( x38 & n20232 ) | ( ~n20228 & n20232 ) ;
  assign n20234 = ~x38 & n20233 ;
  assign n20235 = ( ~n20209 & n20217 ) | ( ~n20209 & n20234 ) | ( n20217 & n20234 ) ;
  assign n20236 = ~n20209 & n20235 ;
  assign n20237 = ( n2069 & n7318 ) | ( n2069 & ~n20236 ) | ( n7318 & ~n20236 ) ;
  assign n20238 = n20236 | n20237 ;
  assign n20239 = ~x709 & n19256 ;
  assign n20240 = n20188 | n20239 ;
  assign n20241 = n1611 & n20240 ;
  assign n20242 = x159 | n1611 ;
  assign n20243 = ( x832 & n20241 ) | ( x832 & n20242 ) | ( n20241 & n20242 ) ;
  assign n20244 = ~n20241 & n20243 ;
  assign n20245 = ~x159 & n8793 ;
  assign n20246 = x832 | n20245 ;
  assign n20247 = ~n20244 & n20246 ;
  assign n20248 = ( n20238 & n20244 ) | ( n20238 & ~n20247 ) | ( n20244 & ~n20247 ) ;
  assign n20249 = x160 | n1611 ;
  assign n20250 = x832 & n20249 ;
  assign n20252 = ~x756 & x947 ;
  assign n20270 = n15644 & ~n20252 ;
  assign n20271 = x160 & ~n15653 ;
  assign n20272 = ( x38 & n20270 ) | ( x38 & ~n20271 ) | ( n20270 & ~n20271 ) ;
  assign n20273 = ~n20270 & n20272 ;
  assign n20251 = x160 | n15332 ;
  assign n20253 = n15332 & n20252 ;
  assign n20254 = ( x39 & n20251 ) | ( x39 & ~n20253 ) | ( n20251 & ~n20253 ) ;
  assign n20255 = ~x39 & n20254 ;
  assign n20256 = ~x160 & x756 ;
  assign n20257 = ~n15486 & n20256 ;
  assign n20258 = x39 & ~n20257 ;
  assign n20259 = x160 | n15484 ;
  assign n20260 = ~n19428 & n20259 ;
  assign n20261 = x160 & n19516 ;
  assign n20262 = x299 & ~n20261 ;
  assign n20263 = x160 | n19451 ;
  assign n20264 = n20262 & n20263 ;
  assign n20265 = ( x756 & ~n20260 ) | ( x756 & n20264 ) | ( ~n20260 & n20264 ) ;
  assign n20266 = n20260 | n20265 ;
  assign n20267 = n20258 & n20266 ;
  assign n20268 = ( x38 & ~n20255 ) | ( x38 & n20267 ) | ( ~n20255 & n20267 ) ;
  assign n20269 = n20255 | n20268 ;
  assign n20274 = n20273 ^ n20269 ^ 1'b0 ;
  assign n20275 = ( x734 & ~n20269 ) | ( x734 & n20273 ) | ( ~n20269 & n20273 ) ;
  assign n20276 = ( x734 & ~n20274 ) | ( x734 & n20275 ) | ( ~n20274 & n20275 ) ;
  assign n20277 = x756 & x947 ;
  assign n20278 = ( x39 & n19568 ) | ( x39 & ~n20277 ) | ( n19568 & ~n20277 ) ;
  assign n20279 = ~x39 & n20278 ;
  assign n20280 = x160 | n15644 ;
  assign n20281 = x38 & n20280 ;
  assign n20282 = n20281 ^ n20279 ^ 1'b0 ;
  assign n20283 = ( n20279 & n20281 ) | ( n20279 & n20282 ) | ( n20281 & n20282 ) ;
  assign n20284 = ( x734 & ~n20279 ) | ( x734 & n20283 ) | ( ~n20279 & n20283 ) ;
  assign n20285 = ~x160 & n19390 ;
  assign n20286 = x756 & ~n19392 ;
  assign n20287 = x160 & ~n19407 ;
  assign n20288 = ( n20285 & n20286 ) | ( n20285 & ~n20287 ) | ( n20286 & ~n20287 ) ;
  assign n20289 = ~n20285 & n20288 ;
  assign n20290 = ~x160 & n19378 ;
  assign n20291 = x160 & ~n19354 ;
  assign n20292 = ( x756 & ~n20290 ) | ( x756 & n20291 ) | ( ~n20290 & n20291 ) ;
  assign n20293 = n20290 | n20292 ;
  assign n20294 = ( x39 & n20289 ) | ( x39 & n20293 ) | ( n20289 & n20293 ) ;
  assign n20295 = ~n20289 & n20294 ;
  assign n20296 = ~n19397 & n20255 ;
  assign n20297 = ( ~x38 & n20295 ) | ( ~x38 & n20296 ) | ( n20295 & n20296 ) ;
  assign n20298 = ~x38 & n20297 ;
  assign n20299 = ( ~n20276 & n20284 ) | ( ~n20276 & n20298 ) | ( n20284 & n20298 ) ;
  assign n20300 = ~n20276 & n20299 ;
  assign n20301 = ( n2069 & n7318 ) | ( n2069 & ~n20300 ) | ( n7318 & ~n20300 ) ;
  assign n20302 = n20300 | n20301 ;
  assign n20303 = ~x160 & n8793 ;
  assign n20304 = ( x832 & n20302 ) | ( x832 & ~n20303 ) | ( n20302 & ~n20303 ) ;
  assign n20305 = ~x832 & n20304 ;
  assign n20306 = ~x734 & n19256 ;
  assign n20307 = n20252 | n20306 ;
  assign n20308 = n1611 & n20307 ;
  assign n20309 = ~n20305 & n20308 ;
  assign n20310 = ( n20250 & n20305 ) | ( n20250 & ~n20309 ) | ( n20305 & ~n20309 ) ;
  assign n20311 = ~x161 & n8793 ;
  assign n20312 = x832 | n20311 ;
  assign n20313 = x758 & x947 ;
  assign n20314 = x39 | n20313 ;
  assign n20315 = ( x39 & n15333 ) | ( x39 & n20314 ) | ( n15333 & n20314 ) ;
  assign n20316 = n15332 & ~n20315 ;
  assign n20317 = ( x161 & n20315 ) | ( x161 & ~n20316 ) | ( n20315 & ~n20316 ) ;
  assign n20318 = n19397 | n20317 ;
  assign n20319 = x161 | n15482 ;
  assign n20320 = n19362 & n20319 ;
  assign n20321 = x299 | n20320 ;
  assign n20322 = x161 | n15337 ;
  assign n20323 = ~n19761 & n20322 ;
  assign n20324 = n1359 | n20323 ;
  assign n20325 = x161 | n15476 ;
  assign n20326 = n19766 & n20325 ;
  assign n20327 = n19769 & ~n20326 ;
  assign n20328 = ( x223 & n20324 ) | ( x223 & ~n20327 ) | ( n20324 & ~n20327 ) ;
  assign n20329 = ~x223 & n20328 ;
  assign n20330 = n19363 & n20319 ;
  assign n20331 = ( ~n20321 & n20329 ) | ( ~n20321 & n20330 ) | ( n20329 & n20330 ) ;
  assign n20332 = n20321 | n20331 ;
  assign n20333 = n2263 | n20323 ;
  assign n20334 = ~x215 & n20333 ;
  assign n20335 = x161 & ~n19371 ;
  assign n20336 = n19778 & ~n20335 ;
  assign n20337 = ~n15434 & n20336 ;
  assign n20338 = n20334 & ~n20337 ;
  assign n20339 = x161 | n15379 ;
  assign n20340 = n19368 & n20339 ;
  assign n20341 = ( x299 & n20338 ) | ( x299 & ~n20340 ) | ( n20338 & ~n20340 ) ;
  assign n20342 = ~n20338 & n20341 ;
  assign n20343 = x758 & ~n20342 ;
  assign n20344 = n20332 & n20343 ;
  assign n20345 = n19790 & n20325 ;
  assign n20346 = n20324 ^ n19792 ^ n1359 ;
  assign n20347 = ( ~x223 & n20345 ) | ( ~x223 & n20346 ) | ( n20345 & n20346 ) ;
  assign n20348 = ~x223 & n20347 ;
  assign n20349 = ( x299 & n20330 ) | ( x299 & ~n20348 ) | ( n20330 & ~n20348 ) ;
  assign n20350 = n20348 | n20349 ;
  assign n20351 = ~n19369 & n20334 ;
  assign n20352 = ~n20336 & n20351 ;
  assign n20353 = n19800 & n20340 ;
  assign n20354 = ( x299 & n20352 ) | ( x299 & ~n20353 ) | ( n20352 & ~n20353 ) ;
  assign n20355 = ~n20352 & n20354 ;
  assign n20356 = ( x758 & n20350 ) | ( x758 & ~n20355 ) | ( n20350 & ~n20355 ) ;
  assign n20357 = ~x758 & n20356 ;
  assign n20358 = ( x39 & n20344 ) | ( x39 & ~n20357 ) | ( n20344 & ~n20357 ) ;
  assign n20359 = ~n20344 & n20358 ;
  assign n20360 = ( x38 & n20318 ) | ( x38 & ~n20359 ) | ( n20318 & ~n20359 ) ;
  assign n20361 = ~x38 & n20360 ;
  assign n20362 = x161 | n15644 ;
  assign n20363 = n19811 & ~n20314 ;
  assign n20364 = x38 & ~n20363 ;
  assign n20365 = n20362 & n20364 ;
  assign n20366 = ( x736 & n20361 ) | ( x736 & ~n20365 ) | ( n20361 & ~n20365 ) ;
  assign n20367 = ~n20361 & n20366 ;
  assign n20368 = x161 | n15653 ;
  assign n20369 = n20368 ^ x736 ^ 1'b0 ;
  assign n20370 = n15644 & ~n20313 ;
  assign n20371 = x38 & ~n20370 ;
  assign n20372 = ( n20368 & ~n20369 ) | ( n20368 & n20371 ) | ( ~n20369 & n20371 ) ;
  assign n20373 = ( x736 & n20369 ) | ( x736 & n20372 ) | ( n20369 & n20372 ) ;
  assign n20374 = x161 & ~n18576 ;
  assign n20375 = ~n19825 & n20322 ;
  assign n20376 = ~n1359 & n20375 ;
  assign n20377 = n20326 | n20376 ;
  assign n20378 = x223 | n20377 ;
  assign n20379 = ( ~x223 & n20321 ) | ( ~x223 & n20378 ) | ( n20321 & n20378 ) ;
  assign n20380 = x161 & n19445 ;
  assign n20381 = n2263 | n20375 ;
  assign n20382 = ( n19399 & n19433 ) | ( n19399 & n20336 ) | ( n19433 & n20336 ) ;
  assign n20383 = ( x215 & n20381 ) | ( x215 & ~n20382 ) | ( n20381 & ~n20382 ) ;
  assign n20384 = ~x215 & n20383 ;
  assign n20385 = ( n19429 & n20380 ) | ( n19429 & ~n20384 ) | ( n20380 & ~n20384 ) ;
  assign n20386 = ~n20380 & n20385 ;
  assign n20387 = x758 & ~n20386 ;
  assign n20388 = n20379 & n20387 ;
  assign n20389 = ( x39 & n20374 ) | ( x39 & ~n20388 ) | ( n20374 & ~n20388 ) ;
  assign n20390 = ~n20374 & n20389 ;
  assign n20391 = ( x38 & n20317 ) | ( x38 & ~n20390 ) | ( n20317 & ~n20390 ) ;
  assign n20392 = ~x38 & n20391 ;
  assign n20393 = ( ~n20367 & n20373 ) | ( ~n20367 & n20392 ) | ( n20373 & n20392 ) ;
  assign n20394 = ~n20367 & n20393 ;
  assign n20395 = ( n8793 & ~n20312 ) | ( n8793 & n20394 ) | ( ~n20312 & n20394 ) ;
  assign n20396 = ~n20312 & n20395 ;
  assign n20397 = n1611 & ~n20313 ;
  assign n20398 = x736 & n19256 ;
  assign n20399 = n20397 & ~n20398 ;
  assign n20400 = x161 | n1611 ;
  assign n20401 = x832 & n20400 ;
  assign n20402 = n20401 ^ n20399 ^ 1'b0 ;
  assign n20403 = ( n20399 & n20401 ) | ( n20399 & n20402 ) | ( n20401 & n20402 ) ;
  assign n20404 = ( n20396 & ~n20399 ) | ( n20396 & n20403 ) | ( ~n20399 & n20403 ) ;
  assign n20415 = ~x761 & x947 ;
  assign n20421 = n15644 & ~n20415 ;
  assign n20422 = x162 & ~n15653 ;
  assign n20423 = ( x38 & n20421 ) | ( x38 & ~n20422 ) | ( n20421 & ~n20422 ) ;
  assign n20424 = ~n20421 & n20423 ;
  assign n20405 = n13460 & n19516 ;
  assign n20406 = ( ~x761 & n19444 ) | ( ~x761 & n20405 ) | ( n19444 & n20405 ) ;
  assign n20407 = ~x761 & n20406 ;
  assign n20408 = x761 & n15486 ;
  assign n20409 = ~x761 & n19452 ;
  assign n20410 = ( x162 & ~n20408 ) | ( x162 & n20409 ) | ( ~n20408 & n20409 ) ;
  assign n20411 = n20408 | n20410 ;
  assign n20412 = ( x39 & n20407 ) | ( x39 & n20411 ) | ( n20407 & n20411 ) ;
  assign n20413 = ~n20407 & n20412 ;
  assign n20414 = x162 | n15332 ;
  assign n20416 = n15332 & n20415 ;
  assign n20417 = ( x39 & n20414 ) | ( x39 & ~n20416 ) | ( n20414 & ~n20416 ) ;
  assign n20418 = ~x39 & n20417 ;
  assign n20419 = ( x38 & ~n20413 ) | ( x38 & n20418 ) | ( ~n20413 & n20418 ) ;
  assign n20420 = n20413 | n20419 ;
  assign n20425 = n20424 ^ n20420 ^ 1'b0 ;
  assign n20426 = ( x738 & ~n20420 ) | ( x738 & n20424 ) | ( ~n20420 & n20424 ) ;
  assign n20427 = ( x738 & ~n20425 ) | ( x738 & n20426 ) | ( ~n20425 & n20426 ) ;
  assign n20428 = x761 & x947 ;
  assign n20429 = ( x39 & n19568 ) | ( x39 & ~n20428 ) | ( n19568 & ~n20428 ) ;
  assign n20430 = ~x39 & n20429 ;
  assign n20431 = x162 | n15644 ;
  assign n20432 = x38 & n20431 ;
  assign n20433 = n20432 ^ n20430 ^ 1'b0 ;
  assign n20434 = ( n20430 & n20432 ) | ( n20430 & n20433 ) | ( n20432 & n20433 ) ;
  assign n20435 = ( x738 & ~n20430 ) | ( x738 & n20434 ) | ( ~n20430 & n20434 ) ;
  assign n20436 = ~n13460 & n19393 ;
  assign n20437 = x162 & ~n19407 ;
  assign n20438 = ( x761 & n20436 ) | ( x761 & ~n20437 ) | ( n20436 & ~n20437 ) ;
  assign n20439 = ~n20436 & n20438 ;
  assign n20440 = ~x162 & n19378 ;
  assign n20441 = x162 & ~n19354 ;
  assign n20442 = ( x761 & ~n20440 ) | ( x761 & n20441 ) | ( ~n20440 & n20441 ) ;
  assign n20443 = n20440 | n20442 ;
  assign n20444 = ( x39 & n20439 ) | ( x39 & n20443 ) | ( n20439 & n20443 ) ;
  assign n20445 = ~n20439 & n20444 ;
  assign n20446 = ~n19397 & n20418 ;
  assign n20447 = ( ~x38 & n20445 ) | ( ~x38 & n20446 ) | ( n20445 & n20446 ) ;
  assign n20448 = ~x38 & n20447 ;
  assign n20449 = ( ~n20427 & n20435 ) | ( ~n20427 & n20448 ) | ( n20435 & n20448 ) ;
  assign n20450 = ~n20427 & n20449 ;
  assign n20451 = ( n2069 & n7318 ) | ( n2069 & ~n20450 ) | ( n7318 & ~n20450 ) ;
  assign n20452 = n20450 | n20451 ;
  assign n20453 = ~x738 & n19256 ;
  assign n20454 = n20415 | n20453 ;
  assign n20455 = n1611 & n20454 ;
  assign n20456 = x162 | n1611 ;
  assign n20457 = ( x832 & n20455 ) | ( x832 & n20456 ) | ( n20455 & n20456 ) ;
  assign n20458 = ~n20455 & n20457 ;
  assign n20459 = ~x162 & n8793 ;
  assign n20460 = x832 | n20459 ;
  assign n20461 = ~n20458 & n20460 ;
  assign n20462 = ( n20452 & n20458 ) | ( n20452 & ~n20461 ) | ( n20458 & ~n20461 ) ;
  assign n20463 = x163 | n1611 ;
  assign n20464 = x832 & n20463 ;
  assign n20466 = ~x777 & x947 ;
  assign n20483 = n15644 & ~n20466 ;
  assign n20484 = x163 & ~n15653 ;
  assign n20485 = ( x38 & n20483 ) | ( x38 & ~n20484 ) | ( n20483 & ~n20484 ) ;
  assign n20486 = ~n20483 & n20485 ;
  assign n20465 = x163 | n15332 ;
  assign n20467 = n15332 & n20466 ;
  assign n20468 = ( x39 & n20465 ) | ( x39 & ~n20467 ) | ( n20465 & ~n20467 ) ;
  assign n20469 = ~x39 & n20468 ;
  assign n20470 = ~x163 & x777 ;
  assign n20471 = ~n15486 & n20470 ;
  assign n20472 = x39 & ~n20471 ;
  assign n20473 = x163 | n15484 ;
  assign n20474 = ~n19428 & n20473 ;
  assign n20475 = n13259 | n19435 ;
  assign n20476 = x163 | n19451 ;
  assign n20477 = n20475 & n20476 ;
  assign n20478 = ( x777 & ~n20474 ) | ( x777 & n20477 ) | ( ~n20474 & n20477 ) ;
  assign n20479 = n20474 | n20478 ;
  assign n20480 = n20472 & n20479 ;
  assign n20481 = ( x38 & ~n20469 ) | ( x38 & n20480 ) | ( ~n20469 & n20480 ) ;
  assign n20482 = n20469 | n20481 ;
  assign n20487 = n20486 ^ n20482 ^ 1'b0 ;
  assign n20488 = ( x737 & ~n20482 ) | ( x737 & n20486 ) | ( ~n20482 & n20486 ) ;
  assign n20489 = ( x737 & ~n20487 ) | ( x737 & n20488 ) | ( ~n20487 & n20488 ) ;
  assign n20490 = x777 & x947 ;
  assign n20491 = ( x39 & n19568 ) | ( x39 & ~n20490 ) | ( n19568 & ~n20490 ) ;
  assign n20492 = ~x39 & n20491 ;
  assign n20493 = x163 | n15644 ;
  assign n20494 = x38 & n20493 ;
  assign n20495 = n20494 ^ n20492 ^ 1'b0 ;
  assign n20496 = ( n20492 & n20494 ) | ( n20492 & n20495 ) | ( n20494 & n20495 ) ;
  assign n20497 = ( x737 & ~n20492 ) | ( x737 & n20496 ) | ( ~n20492 & n20496 ) ;
  assign n20498 = ~x163 & n19390 ;
  assign n20499 = x777 & ~n19392 ;
  assign n20500 = x163 & ~n19407 ;
  assign n20501 = ( n20498 & n20499 ) | ( n20498 & ~n20500 ) | ( n20499 & ~n20500 ) ;
  assign n20502 = ~n20498 & n20501 ;
  assign n20503 = ~x163 & n19378 ;
  assign n20504 = x163 & ~n19354 ;
  assign n20505 = ( x777 & ~n20503 ) | ( x777 & n20504 ) | ( ~n20503 & n20504 ) ;
  assign n20506 = n20503 | n20505 ;
  assign n20507 = ( x39 & n20502 ) | ( x39 & n20506 ) | ( n20502 & n20506 ) ;
  assign n20508 = ~n20502 & n20507 ;
  assign n20509 = ~n19397 & n20469 ;
  assign n20510 = ( ~x38 & n20508 ) | ( ~x38 & n20509 ) | ( n20508 & n20509 ) ;
  assign n20511 = ~x38 & n20510 ;
  assign n20512 = ( ~n20489 & n20497 ) | ( ~n20489 & n20511 ) | ( n20497 & n20511 ) ;
  assign n20513 = ~n20489 & n20512 ;
  assign n20514 = ( n2069 & n7318 ) | ( n2069 & ~n20513 ) | ( n7318 & ~n20513 ) ;
  assign n20515 = n20513 | n20514 ;
  assign n20516 = ~x163 & n8793 ;
  assign n20517 = ( x832 & n20515 ) | ( x832 & ~n20516 ) | ( n20515 & ~n20516 ) ;
  assign n20518 = ~x832 & n20517 ;
  assign n20519 = ~x737 & n19256 ;
  assign n20520 = n20466 | n20519 ;
  assign n20521 = n1611 & n20520 ;
  assign n20522 = ~n20518 & n20521 ;
  assign n20523 = ( n20464 & n20518 ) | ( n20464 & ~n20522 ) | ( n20518 & ~n20522 ) ;
  assign n20524 = x164 | n1611 ;
  assign n20525 = x832 & n20524 ;
  assign n20526 = ~x164 & n8793 ;
  assign n20527 = x832 | n20526 ;
  assign n20536 = ( x38 & x164 ) | ( x38 & n19413 ) | ( x164 & n19413 ) ;
  assign n20537 = ( x164 & n19396 ) | ( x164 & ~n20536 ) | ( n19396 & ~n20536 ) ;
  assign n20538 = ~n20536 & n20537 ;
  assign n20539 = ( x164 & n19418 ) | ( x164 & n19419 ) | ( n19418 & n19419 ) ;
  assign n20540 = ( x752 & n20538 ) | ( x752 & ~n20539 ) | ( n20538 & ~n20539 ) ;
  assign n20541 = ~n20538 & n20540 ;
  assign n20528 = x164 | n19341 ;
  assign n20529 = n19344 & n20528 ;
  assign n20530 = x164 & n19356 ;
  assign n20531 = x38 | n20530 ;
  assign n20532 = ( x164 & n19382 ) | ( x164 & ~n20531 ) | ( n19382 & ~n20531 ) ;
  assign n20533 = ~n20531 & n20532 ;
  assign n20534 = ( x752 & ~n20529 ) | ( x752 & n20533 ) | ( ~n20529 & n20533 ) ;
  assign n20535 = n20529 | n20534 ;
  assign n20542 = n20541 ^ n20535 ^ 1'b0 ;
  assign n20543 = ( x703 & ~n20535 ) | ( x703 & n20541 ) | ( ~n20535 & n20541 ) ;
  assign n20544 = ( x703 & ~n20542 ) | ( x703 & n20543 ) | ( ~n20542 & n20543 ) ;
  assign n20545 = x164 & ~n19458 ;
  assign n20546 = ( x752 & n19459 ) | ( x752 & ~n20545 ) | ( n19459 & ~n20545 ) ;
  assign n20547 = ~x752 & n20546 ;
  assign n20548 = x752 & n15655 ;
  assign n20549 = ~x752 & n19440 ;
  assign n20550 = x164 & ~n20549 ;
  assign n20551 = ( x703 & ~n20548 ) | ( x703 & n20550 ) | ( ~n20548 & n20550 ) ;
  assign n20552 = n20548 | n20551 ;
  assign n20553 = ( ~n20544 & n20547 ) | ( ~n20544 & n20552 ) | ( n20547 & n20552 ) ;
  assign n20554 = ~n20544 & n20553 ;
  assign n20555 = ( n8793 & ~n20527 ) | ( n8793 & n20554 ) | ( ~n20527 & n20554 ) ;
  assign n20556 = ~n20527 & n20555 ;
  assign n20557 = x703 & n19256 ;
  assign n20558 = ~x752 & x947 ;
  assign n20559 = ( n1611 & n20557 ) | ( n1611 & n20558 ) | ( n20557 & n20558 ) ;
  assign n20560 = n20558 ^ n20557 ^ 1'b0 ;
  assign n20561 = ( n1611 & n20559 ) | ( n1611 & n20560 ) | ( n20559 & n20560 ) ;
  assign n20562 = ~n20556 & n20561 ;
  assign n20563 = ( n20525 & n20556 ) | ( n20525 & ~n20562 ) | ( n20556 & ~n20562 ) ;
  assign n20564 = x165 | n1611 ;
  assign n20565 = x832 & n20564 ;
  assign n20566 = ~x165 & n8793 ;
  assign n20567 = x832 | n20566 ;
  assign n20576 = ( x38 & x165 ) | ( x38 & n19413 ) | ( x165 & n19413 ) ;
  assign n20577 = ( x165 & n19396 ) | ( x165 & ~n20576 ) | ( n19396 & ~n20576 ) ;
  assign n20578 = ~n20576 & n20577 ;
  assign n20579 = ( x165 & n19418 ) | ( x165 & n19419 ) | ( n19418 & n19419 ) ;
  assign n20580 = ( x774 & n20578 ) | ( x774 & ~n20579 ) | ( n20578 & ~n20579 ) ;
  assign n20581 = ~n20578 & n20580 ;
  assign n20568 = x165 | n19341 ;
  assign n20569 = n19344 & n20568 ;
  assign n20570 = x165 & n19356 ;
  assign n20571 = x38 | n20570 ;
  assign n20572 = ( x165 & n19382 ) | ( x165 & ~n20571 ) | ( n19382 & ~n20571 ) ;
  assign n20573 = ~n20571 & n20572 ;
  assign n20574 = ( x774 & ~n20569 ) | ( x774 & n20573 ) | ( ~n20569 & n20573 ) ;
  assign n20575 = n20569 | n20574 ;
  assign n20582 = n20581 ^ n20575 ^ 1'b0 ;
  assign n20583 = ( x687 & ~n20575 ) | ( x687 & n20581 ) | ( ~n20575 & n20581 ) ;
  assign n20584 = ( x687 & ~n20582 ) | ( x687 & n20583 ) | ( ~n20582 & n20583 ) ;
  assign n20585 = x165 & ~n19458 ;
  assign n20586 = ( x774 & n19459 ) | ( x774 & ~n20585 ) | ( n19459 & ~n20585 ) ;
  assign n20587 = ~x774 & n20586 ;
  assign n20588 = x774 & n15655 ;
  assign n20589 = ~x774 & n19440 ;
  assign n20590 = x165 & ~n20589 ;
  assign n20591 = ( x687 & ~n20588 ) | ( x687 & n20590 ) | ( ~n20588 & n20590 ) ;
  assign n20592 = n20588 | n20591 ;
  assign n20593 = ( ~n20584 & n20587 ) | ( ~n20584 & n20592 ) | ( n20587 & n20592 ) ;
  assign n20594 = ~n20584 & n20593 ;
  assign n20595 = ( n8793 & ~n20567 ) | ( n8793 & n20594 ) | ( ~n20567 & n20594 ) ;
  assign n20596 = ~n20567 & n20595 ;
  assign n20597 = x687 & n19256 ;
  assign n20598 = ~x774 & x947 ;
  assign n20599 = ( n1611 & n20597 ) | ( n1611 & n20598 ) | ( n20597 & n20598 ) ;
  assign n20600 = n20598 ^ n20597 ^ 1'b0 ;
  assign n20601 = ( n1611 & n20599 ) | ( n1611 & n20600 ) | ( n20599 & n20600 ) ;
  assign n20602 = ~n20596 & n20601 ;
  assign n20603 = ( n20565 & n20596 ) | ( n20565 & ~n20602 ) | ( n20596 & ~n20602 ) ;
  assign n20604 = x772 | n15486 ;
  assign n20605 = x166 & ~n20604 ;
  assign n20606 = x166 | n15476 ;
  assign n20607 = n19766 & n20606 ;
  assign n20608 = x166 | n15337 ;
  assign n20609 = ~n19825 & n20608 ;
  assign n20610 = ~n1359 & n20609 ;
  assign n20611 = ( ~x223 & n20607 ) | ( ~x223 & n20610 ) | ( n20607 & n20610 ) ;
  assign n20612 = ~x223 & n20611 ;
  assign n20613 = x166 | n15482 ;
  assign n20614 = n19362 & n20613 ;
  assign n20615 = ( x299 & ~n20612 ) | ( x299 & n20614 ) | ( ~n20612 & n20614 ) ;
  assign n20616 = n20612 | n20615 ;
  assign n20617 = x166 & n19445 ;
  assign n20618 = n2263 | n20609 ;
  assign n20619 = x166 & ~n19371 ;
  assign n20620 = n19778 & ~n20619 ;
  assign n20621 = ( n19399 & n19433 ) | ( n19399 & n20620 ) | ( n19433 & n20620 ) ;
  assign n20622 = ( x215 & n20618 ) | ( x215 & ~n20621 ) | ( n20618 & ~n20621 ) ;
  assign n20623 = ~x215 & n20622 ;
  assign n20624 = ( n19429 & n20617 ) | ( n19429 & ~n20623 ) | ( n20617 & ~n20623 ) ;
  assign n20625 = ~n20617 & n20624 ;
  assign n20626 = x772 & ~n20625 ;
  assign n20627 = n20616 & n20626 ;
  assign n20628 = ( x39 & n20605 ) | ( x39 & ~n20627 ) | ( n20605 & ~n20627 ) ;
  assign n20629 = ~n20605 & n20628 ;
  assign n20630 = x772 & x947 ;
  assign n20631 = x39 | n20630 ;
  assign n20632 = n15333 & n20631 ;
  assign n20633 = x166 & ~n15332 ;
  assign n20634 = n20632 | n20633 ;
  assign n20635 = ( x38 & ~n20629 ) | ( x38 & n20634 ) | ( ~n20629 & n20634 ) ;
  assign n20636 = ~x38 & n20635 ;
  assign n20637 = n15644 & ~n20630 ;
  assign n20638 = x166 | n15653 ;
  assign n20639 = ( x38 & n20637 ) | ( x38 & n20638 ) | ( n20637 & n20638 ) ;
  assign n20640 = ~n20637 & n20639 ;
  assign n20641 = ( x727 & ~n20636 ) | ( x727 & n20640 ) | ( ~n20636 & n20640 ) ;
  assign n20642 = n20636 | n20641 ;
  assign n20643 = x166 | n15379 ;
  assign n20644 = n19368 & n20643 ;
  assign n20645 = ~n19761 & n20608 ;
  assign n20646 = n2263 | n20645 ;
  assign n20647 = ~x215 & n20646 ;
  assign n20648 = ~n15434 & n20620 ;
  assign n20649 = n20647 & ~n20648 ;
  assign n20650 = ( x299 & n20644 ) | ( x299 & ~n20649 ) | ( n20644 & ~n20649 ) ;
  assign n20651 = ~n20644 & n20650 ;
  assign n20652 = n1359 | n20645 ;
  assign n20653 = ~x223 & n20652 ;
  assign n20654 = n15476 ^ x166 ^ 1'b0 ;
  assign n20655 = ( x166 & n19256 ) | ( x166 & n20654 ) | ( n19256 & n20654 ) ;
  assign n20656 = n19769 & ~n20655 ;
  assign n20657 = n20653 & ~n20656 ;
  assign n20658 = x299 | n20614 ;
  assign n20659 = n5055 & n15482 ;
  assign n20660 = ( x166 & n19363 ) | ( x166 & n20659 ) | ( n19363 & n20659 ) ;
  assign n20661 = n19363 & n20660 ;
  assign n20662 = ( ~n20657 & n20658 ) | ( ~n20657 & n20661 ) | ( n20658 & n20661 ) ;
  assign n20663 = n20657 | n20662 ;
  assign n20664 = ( x772 & n20651 ) | ( x772 & n20663 ) | ( n20651 & n20663 ) ;
  assign n20665 = ~n20651 & n20664 ;
  assign n20666 = n19800 & n20644 ;
  assign n20667 = ~n19369 & n20647 ;
  assign n20668 = ~n20620 & n20667 ;
  assign n20669 = ( x299 & n20666 ) | ( x299 & ~n20668 ) | ( n20666 & ~n20668 ) ;
  assign n20670 = ~n20666 & n20669 ;
  assign n20671 = n1359 & ~n20655 ;
  assign n20672 = ( n19792 & n20653 ) | ( n19792 & ~n20671 ) | ( n20653 & ~n20671 ) ;
  assign n20673 = ~n19792 & n20672 ;
  assign n20674 = ( x299 & ~n20661 ) | ( x299 & n20673 ) | ( ~n20661 & n20673 ) ;
  assign n20675 = n20661 | n20674 ;
  assign n20676 = ( x772 & ~n20670 ) | ( x772 & n20675 ) | ( ~n20670 & n20675 ) ;
  assign n20677 = ~x772 & n20676 ;
  assign n20678 = ( x39 & n20665 ) | ( x39 & ~n20677 ) | ( n20665 & ~n20677 ) ;
  assign n20679 = ~n20665 & n20678 ;
  assign n20680 = n19397 | n20634 ;
  assign n20681 = ( x38 & ~n20679 ) | ( x38 & n20680 ) | ( ~n20679 & n20680 ) ;
  assign n20682 = ~x38 & n20681 ;
  assign n20683 = x166 | n15644 ;
  assign n20684 = n19811 & ~n20631 ;
  assign n20685 = x38 & ~n20684 ;
  assign n20686 = x727 & ~n20685 ;
  assign n20687 = ( x727 & ~n20683 ) | ( x727 & n20686 ) | ( ~n20683 & n20686 ) ;
  assign n20688 = n20642 & ~n20687 ;
  assign n20689 = ( n20642 & n20682 ) | ( n20642 & n20688 ) | ( n20682 & n20688 ) ;
  assign n20690 = ( n2069 & n7318 ) | ( n2069 & ~n20689 ) | ( n7318 & ~n20689 ) ;
  assign n20691 = n20689 | n20690 ;
  assign n20692 = x166 | n1611 ;
  assign n20693 = n1611 & ~n20630 ;
  assign n20694 = x727 & n19256 ;
  assign n20695 = n20693 & ~n20694 ;
  assign n20696 = x832 & ~n20695 ;
  assign n20697 = n20692 & n20696 ;
  assign n20698 = ~x166 & n8793 ;
  assign n20699 = x832 | n20698 ;
  assign n20700 = ~n20697 & n20699 ;
  assign n20701 = ( n20691 & n20697 ) | ( n20691 & ~n20700 ) | ( n20697 & ~n20700 ) ;
  assign n20702 = x167 | n1611 ;
  assign n20703 = x832 & n20702 ;
  assign n20704 = ( x38 & x167 ) | ( x38 & n19413 ) | ( x167 & n19413 ) ;
  assign n20705 = ( x167 & n19396 ) | ( x167 & ~n20704 ) | ( n19396 & ~n20704 ) ;
  assign n20706 = ~n20704 & n20705 ;
  assign n20707 = ( x167 & n19418 ) | ( x167 & n19419 ) | ( n19418 & n19419 ) ;
  assign n20708 = ( x768 & n20706 ) | ( x768 & ~n20707 ) | ( n20706 & ~n20707 ) ;
  assign n20709 = ~n20706 & n20708 ;
  assign n20710 = x167 | n19382 ;
  assign n20711 = x167 & n19356 ;
  assign n20712 = ( x38 & n20710 ) | ( x38 & ~n20711 ) | ( n20710 & ~n20711 ) ;
  assign n20713 = ~x38 & n20712 ;
  assign n20714 = x167 | n19341 ;
  assign n20715 = n19344 & n20714 ;
  assign n20716 = ( x768 & ~n20713 ) | ( x768 & n20715 ) | ( ~n20713 & n20715 ) ;
  assign n20717 = n20713 | n20716 ;
  assign n20718 = ( x705 & n20709 ) | ( x705 & n20717 ) | ( n20709 & n20717 ) ;
  assign n20719 = ~n20709 & n20718 ;
  assign n20720 = x167 | n19455 ;
  assign n20721 = x167 & n19438 ;
  assign n20722 = ( x38 & n20720 ) | ( x38 & ~n20721 ) | ( n20720 & ~n20721 ) ;
  assign n20723 = ~x38 & n20722 ;
  assign n20724 = x167 | n15653 ;
  assign n20725 = n19425 & n20724 ;
  assign n20726 = ( x768 & ~n20723 ) | ( x768 & n20725 ) | ( ~n20723 & n20725 ) ;
  assign n20727 = n20723 | n20726 ;
  assign n20728 = x768 & ~n15655 ;
  assign n20729 = ~x167 & n20728 ;
  assign n20730 = ( x705 & n20727 ) | ( x705 & ~n20729 ) | ( n20727 & ~n20729 ) ;
  assign n20731 = ~x705 & n20730 ;
  assign n20732 = ( n8793 & ~n20719 ) | ( n8793 & n20731 ) | ( ~n20719 & n20731 ) ;
  assign n20733 = n20719 | n20732 ;
  assign n20734 = ~x167 & n8793 ;
  assign n20735 = ( x832 & n20733 ) | ( x832 & ~n20734 ) | ( n20733 & ~n20734 ) ;
  assign n20736 = ~x832 & n20735 ;
  assign n20737 = x705 & n19256 ;
  assign n20738 = ~x768 & x947 ;
  assign n20739 = ( n1611 & n20737 ) | ( n1611 & n20738 ) | ( n20737 & n20738 ) ;
  assign n20740 = n20738 ^ n20737 ^ 1'b0 ;
  assign n20741 = ( n1611 & n20739 ) | ( n1611 & n20740 ) | ( n20739 & n20740 ) ;
  assign n20742 = ~n20736 & n20741 ;
  assign n20743 = ( n20703 & n20736 ) | ( n20703 & ~n20742 ) | ( n20736 & ~n20742 ) ;
  assign n20744 = x763 & x947 ;
  assign n20745 = n1611 & ~n20744 ;
  assign n20746 = x699 & n19256 ;
  assign n20747 = n20745 & ~n20746 ;
  assign n20748 = x168 & ~n1611 ;
  assign n20749 = ( x832 & n20747 ) | ( x832 & ~n20748 ) | ( n20747 & ~n20748 ) ;
  assign n20750 = ~n20747 & n20749 ;
  assign n20751 = x57 & x168 ;
  assign n20752 = x832 | n20751 ;
  assign n20753 = ~x763 & x947 ;
  assign n20754 = ( x39 & n19568 ) | ( x39 & ~n20753 ) | ( n19568 & ~n20753 ) ;
  assign n20755 = ~x39 & n20754 ;
  assign n20756 = x168 | n15644 ;
  assign n20757 = ( x38 & n20755 ) | ( x38 & n20756 ) | ( n20755 & n20756 ) ;
  assign n20758 = ~n20755 & n20757 ;
  assign n20759 = x168 | n15484 ;
  assign n20760 = ~n19409 & n20759 ;
  assign n20761 = x168 & n2263 ;
  assign n20762 = n15434 | n20761 ;
  assign n20763 = ( ~n15434 & n15471 ) | ( ~n15434 & n20762 ) | ( n15471 & n20762 ) ;
  assign n20764 = x168 | n15337 ;
  assign n20765 = ~n19710 & n20764 ;
  assign n20766 = n19372 | n20765 ;
  assign n20767 = ( ~x215 & n20763 ) | ( ~x215 & n20766 ) | ( n20763 & n20766 ) ;
  assign n20768 = ~x215 & n20767 ;
  assign n20769 = x168 & ~n15379 ;
  assign n20770 = n19368 & ~n20769 ;
  assign n20771 = n20770 ^ n19388 ^ x215 ;
  assign n20772 = ( x299 & n20768 ) | ( x299 & n20771 ) | ( n20768 & n20771 ) ;
  assign n20773 = n20771 ^ n20768 ^ 1'b0 ;
  assign n20774 = ( x299 & n20772 ) | ( x299 & n20773 ) | ( n20772 & n20773 ) ;
  assign n20775 = ( x763 & ~n20760 ) | ( x763 & n20774 ) | ( ~n20760 & n20774 ) ;
  assign n20776 = n20760 | n20775 ;
  assign n20779 = ( n2264 & ~n19432 ) | ( n2264 & n20765 ) | ( ~n19432 & n20765 ) ;
  assign n20780 = n20763 | n20779 ;
  assign n20781 = n20780 ^ n20770 ^ 1'b0 ;
  assign n20782 = ( x299 & n20770 ) | ( x299 & ~n20780 ) | ( n20770 & ~n20780 ) ;
  assign n20783 = ( x299 & ~n20781 ) | ( x299 & n20782 ) | ( ~n20781 & n20782 ) ;
  assign n20777 = x168 & ~n19351 ;
  assign n20778 = n19367 | n20777 ;
  assign n20784 = n20783 ^ n20778 ^ 1'b0 ;
  assign n20785 = ( x763 & ~n20778 ) | ( x763 & n20783 ) | ( ~n20778 & n20783 ) ;
  assign n20786 = ( x763 & ~n20784 ) | ( x763 & n20785 ) | ( ~n20784 & n20785 ) ;
  assign n20787 = x39 & ~n20786 ;
  assign n20788 = n20776 & n20787 ;
  assign n20789 = ~x763 & n15487 ;
  assign n20790 = n19901 & ~n20789 ;
  assign n20791 = x168 | n15332 ;
  assign n20792 = ~n20790 & n20791 ;
  assign n20793 = ~n19397 & n20792 ;
  assign n20794 = ( ~x38 & n20788 ) | ( ~x38 & n20793 ) | ( n20788 & n20793 ) ;
  assign n20795 = ~x38 & n20794 ;
  assign n20796 = ( x699 & n20758 ) | ( x699 & n20795 ) | ( n20758 & n20795 ) ;
  assign n20797 = n20795 ^ n20758 ^ 1'b0 ;
  assign n20798 = ( x699 & n20796 ) | ( x699 & n20797 ) | ( n20796 & n20797 ) ;
  assign n20799 = x168 & ~n15653 ;
  assign n20800 = ~n5017 & n20745 ;
  assign n20801 = x38 & ~n20800 ;
  assign n20802 = n20801 ^ n20799 ^ 1'b0 ;
  assign n20803 = ( n20799 & n20801 ) | ( n20799 & n20802 ) | ( n20801 & n20802 ) ;
  assign n20804 = ( x699 & ~n20799 ) | ( x699 & n20803 ) | ( ~n20799 & n20803 ) ;
  assign n20805 = ~n19428 & n20759 ;
  assign n20806 = n19445 & ~n20769 ;
  assign n20807 = ~n19431 & n20764 ;
  assign n20808 = n20763 | n20807 ;
  assign n20809 = n19449 | n20808 ;
  assign n20810 = ( x299 & n20806 ) | ( x299 & n20809 ) | ( n20806 & n20809 ) ;
  assign n20811 = ~n20806 & n20810 ;
  assign n20812 = ( x763 & n20805 ) | ( x763 & ~n20811 ) | ( n20805 & ~n20811 ) ;
  assign n20813 = ~n20805 & n20812 ;
  assign n20814 = x168 | x763 ;
  assign n20815 = n15486 | n20814 ;
  assign n20816 = ( x39 & n20813 ) | ( x39 & n20815 ) | ( n20813 & n20815 ) ;
  assign n20817 = ~n20813 & n20816 ;
  assign n20818 = x38 | n20792 ;
  assign n20819 = ( ~n20804 & n20817 ) | ( ~n20804 & n20818 ) | ( n20817 & n20818 ) ;
  assign n20820 = ~n20804 & n20819 ;
  assign n20821 = ( n19509 & ~n20798 ) | ( n19509 & n20820 ) | ( ~n20798 & n20820 ) ;
  assign n20822 = n20798 | n20821 ;
  assign n20823 = ~x168 & n19509 ;
  assign n20824 = ( x57 & n20822 ) | ( x57 & ~n20823 ) | ( n20822 & ~n20823 ) ;
  assign n20825 = ~x57 & n20824 ;
  assign n20826 = ( ~n20750 & n20752 ) | ( ~n20750 & n20825 ) | ( n20752 & n20825 ) ;
  assign n20827 = ~n20750 & n20826 ;
  assign n20828 = x746 & x947 ;
  assign n20829 = n1611 & ~n20828 ;
  assign n20830 = x729 & n19256 ;
  assign n20831 = n20829 & ~n20830 ;
  assign n20832 = x169 & ~n1611 ;
  assign n20833 = ( x832 & n20831 ) | ( x832 & ~n20832 ) | ( n20831 & ~n20832 ) ;
  assign n20834 = ~n20831 & n20833 ;
  assign n20835 = x57 & x169 ;
  assign n20836 = x832 | n20835 ;
  assign n20837 = ~x746 & x947 ;
  assign n20838 = ( x39 & n19568 ) | ( x39 & ~n20837 ) | ( n19568 & ~n20837 ) ;
  assign n20839 = ~x39 & n20838 ;
  assign n20840 = x169 | n15644 ;
  assign n20841 = ( x38 & n20839 ) | ( x38 & n20840 ) | ( n20839 & n20840 ) ;
  assign n20842 = ~n20839 & n20841 ;
  assign n20843 = x169 | n15484 ;
  assign n20844 = ~n19409 & n20843 ;
  assign n20845 = x169 & n2263 ;
  assign n20846 = n15434 | n20845 ;
  assign n20847 = ( ~n15434 & n15471 ) | ( ~n15434 & n20846 ) | ( n15471 & n20846 ) ;
  assign n20848 = x169 | n15337 ;
  assign n20849 = ~n19710 & n20848 ;
  assign n20850 = n19372 | n20849 ;
  assign n20851 = ( ~x215 & n20847 ) | ( ~x215 & n20850 ) | ( n20847 & n20850 ) ;
  assign n20852 = ~x215 & n20851 ;
  assign n20853 = x169 & ~n15379 ;
  assign n20854 = n19368 & ~n20853 ;
  assign n20855 = n20854 ^ n19388 ^ x215 ;
  assign n20856 = ( x299 & n20852 ) | ( x299 & n20855 ) | ( n20852 & n20855 ) ;
  assign n20857 = n20855 ^ n20852 ^ 1'b0 ;
  assign n20858 = ( x299 & n20856 ) | ( x299 & n20857 ) | ( n20856 & n20857 ) ;
  assign n20859 = ( x746 & ~n20844 ) | ( x746 & n20858 ) | ( ~n20844 & n20858 ) ;
  assign n20860 = n20844 | n20859 ;
  assign n20863 = ( n2264 & ~n19432 ) | ( n2264 & n20849 ) | ( ~n19432 & n20849 ) ;
  assign n20864 = n20847 | n20863 ;
  assign n20865 = n20864 ^ n20854 ^ 1'b0 ;
  assign n20866 = ( x299 & n20854 ) | ( x299 & ~n20864 ) | ( n20854 & ~n20864 ) ;
  assign n20867 = ( x299 & ~n20865 ) | ( x299 & n20866 ) | ( ~n20865 & n20866 ) ;
  assign n20861 = x169 & ~n19351 ;
  assign n20862 = n19367 | n20861 ;
  assign n20868 = n20867 ^ n20862 ^ 1'b0 ;
  assign n20869 = ( x746 & ~n20862 ) | ( x746 & n20867 ) | ( ~n20862 & n20867 ) ;
  assign n20870 = ( x746 & ~n20868 ) | ( x746 & n20869 ) | ( ~n20868 & n20869 ) ;
  assign n20871 = x39 & ~n20870 ;
  assign n20872 = n20860 & n20871 ;
  assign n20873 = ~x746 & n15487 ;
  assign n20874 = n19901 & ~n20873 ;
  assign n20875 = x169 | n15332 ;
  assign n20876 = ~n20874 & n20875 ;
  assign n20877 = ~n19397 & n20876 ;
  assign n20878 = ( ~x38 & n20872 ) | ( ~x38 & n20877 ) | ( n20872 & n20877 ) ;
  assign n20879 = ~x38 & n20878 ;
  assign n20880 = ( x729 & n20842 ) | ( x729 & n20879 ) | ( n20842 & n20879 ) ;
  assign n20881 = n20879 ^ n20842 ^ 1'b0 ;
  assign n20882 = ( x729 & n20880 ) | ( x729 & n20881 ) | ( n20880 & n20881 ) ;
  assign n20883 = x169 & ~n15653 ;
  assign n20884 = ~n5017 & n20829 ;
  assign n20885 = x38 & ~n20884 ;
  assign n20886 = n20885 ^ n20883 ^ 1'b0 ;
  assign n20887 = ( n20883 & n20885 ) | ( n20883 & n20886 ) | ( n20885 & n20886 ) ;
  assign n20888 = ( x729 & ~n20883 ) | ( x729 & n20887 ) | ( ~n20883 & n20887 ) ;
  assign n20889 = ~n19428 & n20843 ;
  assign n20890 = n19445 & ~n20853 ;
  assign n20891 = ~n19431 & n20848 ;
  assign n20892 = n20847 | n20891 ;
  assign n20893 = n19449 | n20892 ;
  assign n20894 = ( x299 & n20890 ) | ( x299 & n20893 ) | ( n20890 & n20893 ) ;
  assign n20895 = ~n20890 & n20894 ;
  assign n20896 = ( x746 & n20889 ) | ( x746 & ~n20895 ) | ( n20889 & ~n20895 ) ;
  assign n20897 = ~n20889 & n20896 ;
  assign n20898 = x169 | x746 ;
  assign n20899 = n15486 | n20898 ;
  assign n20900 = ( x39 & n20897 ) | ( x39 & n20899 ) | ( n20897 & n20899 ) ;
  assign n20901 = ~n20897 & n20900 ;
  assign n20902 = x38 | n20876 ;
  assign n20903 = ( ~n20888 & n20901 ) | ( ~n20888 & n20902 ) | ( n20901 & n20902 ) ;
  assign n20904 = ~n20888 & n20903 ;
  assign n20905 = ( n19509 & ~n20882 ) | ( n19509 & n20904 ) | ( ~n20882 & n20904 ) ;
  assign n20906 = n20882 | n20905 ;
  assign n20907 = ~x169 & n19509 ;
  assign n20908 = ( x57 & n20906 ) | ( x57 & ~n20907 ) | ( n20906 & ~n20907 ) ;
  assign n20909 = ~x57 & n20908 ;
  assign n20910 = ( ~n20834 & n20836 ) | ( ~n20834 & n20909 ) | ( n20836 & n20909 ) ;
  assign n20911 = ~n20834 & n20910 ;
  assign n20912 = x748 & x947 ;
  assign n20913 = x730 & n19256 ;
  assign n20914 = ( n1611 & n20912 ) | ( n1611 & ~n20913 ) | ( n20912 & ~n20913 ) ;
  assign n20915 = ~n20912 & n20914 ;
  assign n20916 = x170 & ~n1611 ;
  assign n20917 = ( x832 & n20915 ) | ( x832 & ~n20916 ) | ( n20915 & ~n20916 ) ;
  assign n20918 = ~n20915 & n20917 ;
  assign n20919 = ~x170 & n19509 ;
  assign n20920 = x170 | n15653 ;
  assign n20921 = n19425 & n20920 ;
  assign n20922 = x170 & ~n15379 ;
  assign n20923 = n19445 & ~n20922 ;
  assign n20924 = x299 & ~n20923 ;
  assign n20925 = x170 & n2263 ;
  assign n20926 = n15434 | n20925 ;
  assign n20927 = ( ~n15434 & n15471 ) | ( ~n15434 & n20926 ) | ( n15471 & n20926 ) ;
  assign n20928 = x170 | n15337 ;
  assign n20929 = ~n19431 & n20928 ;
  assign n20930 = n20927 | n20929 ;
  assign n20931 = n19449 | n20930 ;
  assign n20932 = n20924 & n20931 ;
  assign n20933 = ( x170 & ~x299 ) | ( x170 & n19391 ) | ( ~x299 & n19391 ) ;
  assign n20934 = ~n19427 & n20933 ;
  assign n20935 = ( x39 & n20932 ) | ( x39 & n20934 ) | ( n20932 & n20934 ) ;
  assign n20936 = n20934 ^ n20932 ^ 1'b0 ;
  assign n20937 = ( x39 & n20935 ) | ( x39 & n20936 ) | ( n20935 & n20936 ) ;
  assign n20938 = x170 | n15332 ;
  assign n20939 = ~n19901 & n20938 ;
  assign n20940 = ( ~x38 & n20937 ) | ( ~x38 & n20939 ) | ( n20937 & n20939 ) ;
  assign n20941 = ~x38 & n20940 ;
  assign n20942 = ( x748 & n20921 ) | ( x748 & ~n20941 ) | ( n20921 & ~n20941 ) ;
  assign n20943 = ~n20921 & n20942 ;
  assign n20944 = x170 | x748 ;
  assign n20945 = n15655 | n20944 ;
  assign n20946 = ( x730 & ~n20943 ) | ( x730 & n20945 ) | ( ~n20943 & n20945 ) ;
  assign n20947 = ~x730 & n20946 ;
  assign n20948 = x170 | n15644 ;
  assign n20949 = n19418 & n20948 ;
  assign n20950 = ~n19710 & n20928 ;
  assign n20951 = n19372 | n20950 ;
  assign n20952 = ( ~x215 & n20927 ) | ( ~x215 & n20951 ) | ( n20927 & n20951 ) ;
  assign n20953 = ~x215 & n20952 ;
  assign n20954 = n19368 & ~n20922 ;
  assign n20955 = n20954 ^ n19388 ^ x215 ;
  assign n20956 = ( x299 & n20953 ) | ( x299 & n20955 ) | ( n20953 & n20955 ) ;
  assign n20957 = n20955 ^ n20953 ^ 1'b0 ;
  assign n20958 = ( x299 & n20956 ) | ( x299 & n20957 ) | ( n20956 & n20957 ) ;
  assign n20959 = ~n19408 & n20933 ;
  assign n20960 = ( x39 & n20958 ) | ( x39 & n20959 ) | ( n20958 & n20959 ) ;
  assign n20961 = n20959 ^ n20958 ^ 1'b0 ;
  assign n20962 = ( x39 & n20960 ) | ( x39 & n20961 ) | ( n20960 & n20961 ) ;
  assign n20963 = ~n19733 & n20938 ;
  assign n20964 = ( ~x38 & n20962 ) | ( ~x38 & n20963 ) | ( n20962 & n20963 ) ;
  assign n20965 = ~x38 & n20964 ;
  assign n20966 = ( x748 & ~n20949 ) | ( x748 & n20965 ) | ( ~n20949 & n20965 ) ;
  assign n20967 = n20949 | n20966 ;
  assign n20968 = ~n19380 & n20938 ;
  assign n20969 = x39 & ~x299 ;
  assign n20970 = ( n2264 & ~n19432 ) | ( n2264 & n20950 ) | ( ~n19432 & n20950 ) ;
  assign n20971 = n20927 | n20970 ;
  assign n20972 = ~n20954 & n20971 ;
  assign n20973 = ( x39 & n20969 ) | ( x39 & n20972 ) | ( n20969 & n20972 ) ;
  assign n20974 = x170 & ~n19351 ;
  assign n20975 = n20974 ^ n19367 ^ 1'b0 ;
  assign n20976 = ( n19367 & n20974 ) | ( n19367 & ~n20975 ) | ( n20974 & ~n20975 ) ;
  assign n20977 = ( n20973 & n20975 ) | ( n20973 & n20976 ) | ( n20975 & n20976 ) ;
  assign n20978 = ( ~x38 & n20968 ) | ( ~x38 & n20977 ) | ( n20968 & n20977 ) ;
  assign n20979 = ~x38 & n20978 ;
  assign n20980 = n19344 & n20948 ;
  assign n20981 = ( x748 & n20979 ) | ( x748 & ~n20980 ) | ( n20979 & ~n20980 ) ;
  assign n20982 = ~n20979 & n20981 ;
  assign n20983 = x730 & ~n20982 ;
  assign n20984 = n20967 & n20983 ;
  assign n20985 = ( n19509 & ~n20947 ) | ( n19509 & n20984 ) | ( ~n20947 & n20984 ) ;
  assign n20986 = n20947 | n20985 ;
  assign n20987 = ( x57 & ~n20919 ) | ( x57 & n20986 ) | ( ~n20919 & n20986 ) ;
  assign n20988 = ~x57 & n20987 ;
  assign n20989 = x57 & x170 ;
  assign n20990 = x832 | n20989 ;
  assign n20991 = ( ~n20918 & n20988 ) | ( ~n20918 & n20990 ) | ( n20988 & n20990 ) ;
  assign n20992 = ~n20918 & n20991 ;
  assign n20993 = x764 & x947 ;
  assign n20994 = n1611 & ~n20993 ;
  assign n20995 = x691 & n19256 ;
  assign n20996 = n20994 & ~n20995 ;
  assign n20997 = x171 & ~n1611 ;
  assign n20998 = ( x832 & n20996 ) | ( x832 & ~n20997 ) | ( n20996 & ~n20997 ) ;
  assign n20999 = ~n20996 & n20998 ;
  assign n21000 = x57 & x171 ;
  assign n21001 = x832 | n21000 ;
  assign n21002 = ~x764 & x947 ;
  assign n21003 = ( x39 & n19568 ) | ( x39 & ~n21002 ) | ( n19568 & ~n21002 ) ;
  assign n21004 = ~x39 & n21003 ;
  assign n21005 = x171 | n15644 ;
  assign n21006 = ( x38 & n21004 ) | ( x38 & n21005 ) | ( n21004 & n21005 ) ;
  assign n21007 = ~n21004 & n21006 ;
  assign n21008 = x171 | n15484 ;
  assign n21009 = ~n19409 & n21008 ;
  assign n21010 = x171 & n2263 ;
  assign n21011 = n15434 | n21010 ;
  assign n21012 = ( ~n15434 & n15471 ) | ( ~n15434 & n21011 ) | ( n15471 & n21011 ) ;
  assign n21013 = x171 | n15337 ;
  assign n21014 = ~n19710 & n21013 ;
  assign n21015 = n19372 | n21014 ;
  assign n21016 = ( ~x215 & n21012 ) | ( ~x215 & n21015 ) | ( n21012 & n21015 ) ;
  assign n21017 = ~x215 & n21016 ;
  assign n21018 = x171 & ~n15379 ;
  assign n21019 = n19368 & ~n21018 ;
  assign n21020 = n21019 ^ n19388 ^ x215 ;
  assign n21021 = ( x299 & n21017 ) | ( x299 & n21020 ) | ( n21017 & n21020 ) ;
  assign n21022 = n21020 ^ n21017 ^ 1'b0 ;
  assign n21023 = ( x299 & n21021 ) | ( x299 & n21022 ) | ( n21021 & n21022 ) ;
  assign n21024 = ( x764 & ~n21009 ) | ( x764 & n21023 ) | ( ~n21009 & n21023 ) ;
  assign n21025 = n21009 | n21024 ;
  assign n21028 = ( n2264 & ~n19432 ) | ( n2264 & n21014 ) | ( ~n19432 & n21014 ) ;
  assign n21029 = n21012 | n21028 ;
  assign n21030 = n21029 ^ n21019 ^ 1'b0 ;
  assign n21031 = ( x299 & n21019 ) | ( x299 & ~n21029 ) | ( n21019 & ~n21029 ) ;
  assign n21032 = ( x299 & ~n21030 ) | ( x299 & n21031 ) | ( ~n21030 & n21031 ) ;
  assign n21026 = x171 & ~n19351 ;
  assign n21027 = n19367 | n21026 ;
  assign n21033 = n21032 ^ n21027 ^ 1'b0 ;
  assign n21034 = ( x764 & ~n21027 ) | ( x764 & n21032 ) | ( ~n21027 & n21032 ) ;
  assign n21035 = ( x764 & ~n21033 ) | ( x764 & n21034 ) | ( ~n21033 & n21034 ) ;
  assign n21036 = x39 & ~n21035 ;
  assign n21037 = n21025 & n21036 ;
  assign n21038 = ~x764 & n15487 ;
  assign n21039 = n19901 & ~n21038 ;
  assign n21040 = x171 | n15332 ;
  assign n21041 = ~n21039 & n21040 ;
  assign n21042 = ~n19397 & n21041 ;
  assign n21043 = ( ~x38 & n21037 ) | ( ~x38 & n21042 ) | ( n21037 & n21042 ) ;
  assign n21044 = ~x38 & n21043 ;
  assign n21045 = ( x691 & n21007 ) | ( x691 & n21044 ) | ( n21007 & n21044 ) ;
  assign n21046 = n21044 ^ n21007 ^ 1'b0 ;
  assign n21047 = ( x691 & n21045 ) | ( x691 & n21046 ) | ( n21045 & n21046 ) ;
  assign n21048 = x171 & ~n15653 ;
  assign n21049 = ~n5017 & n20994 ;
  assign n21050 = x38 & ~n21049 ;
  assign n21051 = n21050 ^ n21048 ^ 1'b0 ;
  assign n21052 = ( n21048 & n21050 ) | ( n21048 & n21051 ) | ( n21050 & n21051 ) ;
  assign n21053 = ( x691 & ~n21048 ) | ( x691 & n21052 ) | ( ~n21048 & n21052 ) ;
  assign n21054 = ~n19428 & n21008 ;
  assign n21055 = n19445 & ~n21018 ;
  assign n21056 = ~n19431 & n21013 ;
  assign n21057 = n21012 | n21056 ;
  assign n21058 = n19449 | n21057 ;
  assign n21059 = ( x299 & n21055 ) | ( x299 & n21058 ) | ( n21055 & n21058 ) ;
  assign n21060 = ~n21055 & n21059 ;
  assign n21061 = ( x764 & n21054 ) | ( x764 & ~n21060 ) | ( n21054 & ~n21060 ) ;
  assign n21062 = ~n21054 & n21061 ;
  assign n21063 = x171 | x764 ;
  assign n21064 = n15486 | n21063 ;
  assign n21065 = ( x39 & n21062 ) | ( x39 & n21064 ) | ( n21062 & n21064 ) ;
  assign n21066 = ~n21062 & n21065 ;
  assign n21067 = x38 | n21041 ;
  assign n21068 = ( ~n21053 & n21066 ) | ( ~n21053 & n21067 ) | ( n21066 & n21067 ) ;
  assign n21069 = ~n21053 & n21068 ;
  assign n21070 = ( n19509 & ~n21047 ) | ( n19509 & n21069 ) | ( ~n21047 & n21069 ) ;
  assign n21071 = n21047 | n21070 ;
  assign n21072 = ~x171 & n19509 ;
  assign n21073 = ( x57 & n21071 ) | ( x57 & ~n21072 ) | ( n21071 & ~n21072 ) ;
  assign n21074 = ~x57 & n21073 ;
  assign n21075 = ( ~n20999 & n21001 ) | ( ~n20999 & n21074 ) | ( n21001 & n21074 ) ;
  assign n21076 = ~n20999 & n21075 ;
  assign n21077 = x739 & x947 ;
  assign n21078 = n1611 & ~n21077 ;
  assign n21079 = x690 & n19256 ;
  assign n21080 = n21078 & ~n21079 ;
  assign n21081 = x172 & ~n1611 ;
  assign n21082 = ( x832 & n21080 ) | ( x832 & ~n21081 ) | ( n21080 & ~n21081 ) ;
  assign n21083 = ~n21080 & n21082 ;
  assign n21084 = x57 & x172 ;
  assign n21085 = x832 | n21084 ;
  assign n21086 = ~x739 & x947 ;
  assign n21087 = ( x39 & n19568 ) | ( x39 & ~n21086 ) | ( n19568 & ~n21086 ) ;
  assign n21088 = ~x39 & n21087 ;
  assign n21089 = x172 | n15644 ;
  assign n21090 = ( x38 & n21088 ) | ( x38 & n21089 ) | ( n21088 & n21089 ) ;
  assign n21091 = ~n21088 & n21090 ;
  assign n21092 = x172 | n15484 ;
  assign n21093 = ~n19409 & n21092 ;
  assign n21094 = x172 & n2263 ;
  assign n21095 = n15434 | n21094 ;
  assign n21096 = ( ~n15434 & n15471 ) | ( ~n15434 & n21095 ) | ( n15471 & n21095 ) ;
  assign n21097 = x172 | n15337 ;
  assign n21098 = ~n19710 & n21097 ;
  assign n21099 = n19372 | n21098 ;
  assign n21100 = ( ~x215 & n21096 ) | ( ~x215 & n21099 ) | ( n21096 & n21099 ) ;
  assign n21101 = ~x215 & n21100 ;
  assign n21102 = x172 & ~n15379 ;
  assign n21103 = n19368 & ~n21102 ;
  assign n21104 = n21103 ^ n19388 ^ x215 ;
  assign n21105 = ( x299 & n21101 ) | ( x299 & n21104 ) | ( n21101 & n21104 ) ;
  assign n21106 = n21104 ^ n21101 ^ 1'b0 ;
  assign n21107 = ( x299 & n21105 ) | ( x299 & n21106 ) | ( n21105 & n21106 ) ;
  assign n21108 = ( x739 & ~n21093 ) | ( x739 & n21107 ) | ( ~n21093 & n21107 ) ;
  assign n21109 = n21093 | n21108 ;
  assign n21112 = ( n2264 & ~n19432 ) | ( n2264 & n21098 ) | ( ~n19432 & n21098 ) ;
  assign n21113 = n21096 | n21112 ;
  assign n21114 = n21113 ^ n21103 ^ 1'b0 ;
  assign n21115 = ( x299 & n21103 ) | ( x299 & ~n21113 ) | ( n21103 & ~n21113 ) ;
  assign n21116 = ( x299 & ~n21114 ) | ( x299 & n21115 ) | ( ~n21114 & n21115 ) ;
  assign n21110 = x172 & ~n19351 ;
  assign n21111 = n19367 | n21110 ;
  assign n21117 = n21116 ^ n21111 ^ 1'b0 ;
  assign n21118 = ( x739 & ~n21111 ) | ( x739 & n21116 ) | ( ~n21111 & n21116 ) ;
  assign n21119 = ( x739 & ~n21117 ) | ( x739 & n21118 ) | ( ~n21117 & n21118 ) ;
  assign n21120 = x39 & ~n21119 ;
  assign n21121 = n21109 & n21120 ;
  assign n21122 = x172 | n15332 ;
  assign n21123 = n15332 & n21077 ;
  assign n21124 = ( x39 & n21122 ) | ( x39 & ~n21123 ) | ( n21122 & ~n21123 ) ;
  assign n21125 = ~x39 & n21124 ;
  assign n21126 = ~n19397 & n21125 ;
  assign n21127 = ( ~x38 & n21121 ) | ( ~x38 & n21126 ) | ( n21121 & n21126 ) ;
  assign n21128 = ~x38 & n21127 ;
  assign n21129 = ( x690 & n21091 ) | ( x690 & n21128 ) | ( n21091 & n21128 ) ;
  assign n21130 = n21128 ^ n21091 ^ 1'b0 ;
  assign n21131 = ( x690 & n21129 ) | ( x690 & n21130 ) | ( n21129 & n21130 ) ;
  assign n21132 = x172 & ~n15653 ;
  assign n21133 = ~n5017 & n21078 ;
  assign n21134 = x38 & ~n21133 ;
  assign n21135 = n21134 ^ n21132 ^ 1'b0 ;
  assign n21136 = ( n21132 & n21134 ) | ( n21132 & n21135 ) | ( n21134 & n21135 ) ;
  assign n21137 = ( x690 & ~n21132 ) | ( x690 & n21136 ) | ( ~n21132 & n21136 ) ;
  assign n21138 = ~n19428 & n21092 ;
  assign n21139 = n19445 & ~n21102 ;
  assign n21140 = ~n19431 & n21097 ;
  assign n21141 = n21096 | n21140 ;
  assign n21142 = n19449 | n21141 ;
  assign n21143 = ( x299 & n21139 ) | ( x299 & n21142 ) | ( n21139 & n21142 ) ;
  assign n21144 = ~n21139 & n21143 ;
  assign n21145 = ( x739 & n21138 ) | ( x739 & ~n21144 ) | ( n21138 & ~n21144 ) ;
  assign n21146 = ~n21138 & n21145 ;
  assign n21147 = x172 | x739 ;
  assign n21148 = n15486 | n21147 ;
  assign n21149 = ( x39 & n21146 ) | ( x39 & n21148 ) | ( n21146 & n21148 ) ;
  assign n21150 = ~n21146 & n21149 ;
  assign n21151 = x38 | n21125 ;
  assign n21152 = ( ~n21137 & n21150 ) | ( ~n21137 & n21151 ) | ( n21150 & n21151 ) ;
  assign n21153 = ~n21137 & n21152 ;
  assign n21154 = ( n19509 & ~n21131 ) | ( n19509 & n21153 ) | ( ~n21131 & n21153 ) ;
  assign n21155 = n21131 | n21154 ;
  assign n21156 = ~x172 & n19509 ;
  assign n21157 = ( x57 & n21155 ) | ( x57 & ~n21156 ) | ( n21155 & ~n21156 ) ;
  assign n21158 = ~x57 & n21157 ;
  assign n21159 = ( ~n21083 & n21085 ) | ( ~n21083 & n21158 ) | ( n21085 & n21158 ) ;
  assign n21160 = ~n21083 & n21159 ;
  assign n21161 = ~x173 & n7318 ;
  assign n21162 = x832 | n21161 ;
  assign n21163 = x173 | n15656 ;
  assign n21164 = x173 | n15644 ;
  assign n21165 = x38 & n21164 ;
  assign n21166 = x173 | x745 ;
  assign n21167 = n15587 & ~n21166 ;
  assign n21168 = n15640 & ~n21167 ;
  assign n21169 = ( x173 & n21167 ) | ( x173 & ~n21168 ) | ( n21167 & ~n21168 ) ;
  assign n21170 = x173 | n15488 ;
  assign n21171 = x745 & n21170 ;
  assign n21172 = ( ~x38 & n21169 ) | ( ~x38 & n21171 ) | ( n21169 & n21171 ) ;
  assign n21173 = ~x38 & n21172 ;
  assign n21174 = ~x745 & n15646 ;
  assign n21175 = ~n21173 & n21174 ;
  assign n21176 = ( n21165 & n21173 ) | ( n21165 & ~n21175 ) | ( n21173 & ~n21175 ) ;
  assign n21177 = ~n2069 & n21176 ;
  assign n21178 = x173 & n2069 ;
  assign n21179 = n21177 | n21178 ;
  assign n21180 = n21163 ^ n15659 ^ 1'b0 ;
  assign n21181 = ( n21163 & n21179 ) | ( n21163 & ~n21180 ) | ( n21179 & ~n21180 ) ;
  assign n21182 = ~n15659 & n21179 ;
  assign n21183 = x609 & n21182 ;
  assign n21184 = ~n15668 & n21163 ;
  assign n21185 = n21183 | n21184 ;
  assign n21186 = ~x609 & n21182 ;
  assign n21187 = n15662 & n21163 ;
  assign n21188 = n21186 | n21187 ;
  assign n21189 = n21185 ^ x1155 ^ 1'b0 ;
  assign n21190 = ( n21185 & n21188 ) | ( n21185 & ~n21189 ) | ( n21188 & ~n21189 ) ;
  assign n21191 = n21181 ^ x785 ^ 1'b0 ;
  assign n21192 = ( n21181 & n21190 ) | ( n21181 & n21191 ) | ( n21190 & n21191 ) ;
  assign n21193 = x618 & ~n21192 ;
  assign n21194 = x618 | n21163 ;
  assign n21195 = ( x1154 & n21193 ) | ( x1154 & n21194 ) | ( n21193 & n21194 ) ;
  assign n21196 = ~n21193 & n21195 ;
  assign n21197 = x618 & ~n21163 ;
  assign n21198 = x1154 | n21197 ;
  assign n21199 = ( n21192 & n21193 ) | ( n21192 & ~n21198 ) | ( n21193 & ~n21198 ) ;
  assign n21200 = n21196 | n21199 ;
  assign n21201 = n21192 ^ x781 ^ 1'b0 ;
  assign n21202 = ( n21192 & n21200 ) | ( n21192 & n21201 ) | ( n21200 & n21201 ) ;
  assign n21203 = x619 & ~n21202 ;
  assign n21204 = x619 | n21163 ;
  assign n21205 = ( x1159 & n21203 ) | ( x1159 & n21204 ) | ( n21203 & n21204 ) ;
  assign n21206 = ~n21203 & n21205 ;
  assign n21207 = x619 & ~n21163 ;
  assign n21208 = x1159 | n21207 ;
  assign n21209 = ( n21202 & n21203 ) | ( n21202 & ~n21208 ) | ( n21203 & ~n21208 ) ;
  assign n21210 = n21206 | n21209 ;
  assign n21211 = n21202 ^ x789 ^ 1'b0 ;
  assign n21212 = ( n21202 & n21210 ) | ( n21202 & n21211 ) | ( n21210 & n21211 ) ;
  assign n21213 = x626 & ~n21212 ;
  assign n21214 = x626 & ~n21163 ;
  assign n21215 = x1158 | n21214 ;
  assign n21216 = ( n21212 & n21213 ) | ( n21212 & ~n21215 ) | ( n21213 & ~n21215 ) ;
  assign n21217 = n21213 & ~n21216 ;
  assign n21218 = ( x1158 & n21163 ) | ( x1158 & n21214 ) | ( n21163 & n21214 ) ;
  assign n21219 = ( n21216 & ~n21217 ) | ( n21216 & n21218 ) | ( ~n21217 & n21218 ) ;
  assign n21220 = n21212 ^ x788 ^ 1'b0 ;
  assign n21221 = ( n21212 & n21219 ) | ( n21212 & n21220 ) | ( n21219 & n21220 ) ;
  assign n21222 = n21163 ^ n16339 ^ 1'b0 ;
  assign n21223 = ( n21163 & n21221 ) | ( n21163 & ~n21222 ) | ( n21221 & ~n21222 ) ;
  assign n21224 = n21163 ^ n16376 ^ 1'b0 ;
  assign n21225 = ( n21163 & n21223 ) | ( n21163 & ~n21224 ) | ( n21223 & ~n21224 ) ;
  assign n21226 = x644 & ~n21225 ;
  assign n21227 = x644 & ~n21163 ;
  assign n21228 = ( ~x715 & n21163 ) | ( ~x715 & n21227 ) | ( n21163 & n21227 ) ;
  assign n21229 = x1160 & ~n21228 ;
  assign n21230 = ( x1160 & n21226 ) | ( x1160 & n21229 ) | ( n21226 & n21229 ) ;
  assign n21231 = n16185 & n21164 ;
  assign n21232 = ( x38 & x173 ) | ( x38 & n16700 ) | ( x173 & n16700 ) ;
  assign n21233 = ~n2069 & n21232 ;
  assign n21234 = ( x173 & n16697 ) | ( x173 & ~n21233 ) | ( n16697 & ~n21233 ) ;
  assign n21235 = ~n21233 & n21234 ;
  assign n21236 = ( x723 & ~n21231 ) | ( x723 & n21235 ) | ( ~n21231 & n21235 ) ;
  assign n21237 = n21231 | n21236 ;
  assign n21238 = n21237 ^ n21163 ^ 1'b0 ;
  assign n21239 = x723 | n2069 ;
  assign n21240 = ( n21163 & n21238 ) | ( n21163 & ~n21239 ) | ( n21238 & ~n21239 ) ;
  assign n21241 = ( n21237 & ~n21238 ) | ( n21237 & n21240 ) | ( ~n21238 & n21240 ) ;
  assign n21242 = x625 & ~n21241 ;
  assign n21243 = x625 | n21163 ;
  assign n21244 = ( x1153 & n21242 ) | ( x1153 & n21243 ) | ( n21242 & n21243 ) ;
  assign n21245 = ~n21242 & n21244 ;
  assign n21246 = x625 & ~n21163 ;
  assign n21247 = x1153 | n21246 ;
  assign n21248 = ( x625 & n21241 ) | ( x625 & ~n21247 ) | ( n21241 & ~n21247 ) ;
  assign n21249 = ~n21247 & n21248 ;
  assign n21250 = n21245 | n21249 ;
  assign n21251 = n21241 ^ x778 ^ 1'b0 ;
  assign n21252 = ( n21241 & n21250 ) | ( n21241 & n21251 ) | ( n21250 & n21251 ) ;
  assign n21253 = n21163 ^ n16234 ^ 1'b0 ;
  assign n21254 = ( n21163 & n21252 ) | ( n21163 & ~n21253 ) | ( n21252 & ~n21253 ) ;
  assign n21255 = n21163 ^ n16254 ^ 1'b0 ;
  assign n21256 = ( n21163 & n21254 ) | ( n21163 & ~n21255 ) | ( n21254 & ~n21255 ) ;
  assign n21257 = n21163 ^ n16279 ^ 1'b0 ;
  assign n21258 = ( n21163 & n21256 ) | ( n21163 & ~n21257 ) | ( n21256 & ~n21257 ) ;
  assign n21259 = n21163 ^ n16318 ^ 1'b0 ;
  assign n21260 = ( n21163 & n21258 ) | ( n21163 & ~n21259 ) | ( n21258 & ~n21259 ) ;
  assign n21261 = x628 & ~n21260 ;
  assign n21262 = x628 | n21163 ;
  assign n21263 = ( x1156 & n21261 ) | ( x1156 & n21262 ) | ( n21261 & n21262 ) ;
  assign n21264 = ~n21261 & n21263 ;
  assign n21265 = x628 & ~n21163 ;
  assign n21266 = x1156 | n21265 ;
  assign n21267 = ( n21260 & n21261 ) | ( n21260 & ~n21266 ) | ( n21261 & ~n21266 ) ;
  assign n21268 = n21264 | n21267 ;
  assign n21269 = n21260 ^ x792 ^ 1'b0 ;
  assign n21270 = ( n21260 & n21268 ) | ( n21260 & n21269 ) | ( n21268 & n21269 ) ;
  assign n21271 = n21163 ^ x647 ^ 1'b0 ;
  assign n21272 = ( n21163 & n21270 ) | ( n21163 & ~n21271 ) | ( n21270 & ~n21271 ) ;
  assign n21273 = ( n21163 & n21270 ) | ( n21163 & n21271 ) | ( n21270 & n21271 ) ;
  assign n21274 = n21272 ^ x1157 ^ 1'b0 ;
  assign n21275 = ( n21272 & n21273 ) | ( n21272 & n21274 ) | ( n21273 & n21274 ) ;
  assign n21276 = n21270 ^ x787 ^ 1'b0 ;
  assign n21277 = ( n21270 & n21275 ) | ( n21270 & n21276 ) | ( n21275 & n21276 ) ;
  assign n21278 = x644 & ~n21277 ;
  assign n21279 = ( x715 & n21277 ) | ( x715 & n21278 ) | ( n21277 & n21278 ) ;
  assign n21280 = n21230 & ~n21279 ;
  assign n21408 = x715 & ~n21227 ;
  assign n21409 = ( n21225 & n21226 ) | ( n21225 & n21408 ) | ( n21226 & n21408 ) ;
  assign n21281 = x715 | n21278 ;
  assign n21282 = x723 & ~n21176 ;
  assign n21283 = x173 & ~n16054 ;
  assign n21284 = ~x173 & n16048 ;
  assign n21285 = ( x745 & ~n21283 ) | ( x745 & n21284 ) | ( ~n21283 & n21284 ) ;
  assign n21286 = n21283 | n21285 ;
  assign n21287 = ~x173 & n16044 ;
  assign n21288 = x173 & ~n16029 ;
  assign n21289 = ( x745 & n21287 ) | ( x745 & ~n21288 ) | ( n21287 & ~n21288 ) ;
  assign n21290 = ~n21287 & n21289 ;
  assign n21291 = ( x39 & n21286 ) | ( x39 & ~n21290 ) | ( n21286 & ~n21290 ) ;
  assign n21292 = n21291 ^ n21286 ^ 1'b0 ;
  assign n21293 = ( x39 & n21291 ) | ( x39 & ~n21292 ) | ( n21291 & ~n21292 ) ;
  assign n21294 = x173 & n15795 ;
  assign n21295 = x745 & ~n21294 ;
  assign n21296 = x173 | n15876 ;
  assign n21297 = n21295 & n21296 ;
  assign n21298 = x173 & n15943 ;
  assign n21299 = x173 | n16003 ;
  assign n21300 = ( x745 & ~n21298 ) | ( x745 & n21299 ) | ( ~n21298 & n21299 ) ;
  assign n21301 = ~x745 & n21300 ;
  assign n21302 = ( x39 & n21297 ) | ( x39 & ~n21301 ) | ( n21297 & ~n21301 ) ;
  assign n21303 = ~n21297 & n21302 ;
  assign n21304 = ( x38 & n21293 ) | ( x38 & ~n21303 ) | ( n21293 & ~n21303 ) ;
  assign n21305 = ~x38 & n21304 ;
  assign n21306 = x745 | n15968 ;
  assign n21307 = n17889 & n21306 ;
  assign n21308 = x173 | n21307 ;
  assign n21309 = n21308 ^ x723 ^ 1'b0 ;
  assign n21310 = ~x745 & n15591 ;
  assign n21311 = n17156 | n21310 ;
  assign n21312 = x173 & ~n5017 ;
  assign n21313 = n21311 & n21312 ;
  assign n21314 = x38 & ~n21313 ;
  assign n21315 = ( n21308 & ~n21309 ) | ( n21308 & n21314 ) | ( ~n21309 & n21314 ) ;
  assign n21316 = ( x723 & n21309 ) | ( x723 & n21315 ) | ( n21309 & n21315 ) ;
  assign n21317 = ( ~n2069 & n21305 ) | ( ~n2069 & n21316 ) | ( n21305 & n21316 ) ;
  assign n21318 = ~n2069 & n21317 ;
  assign n21319 = n21318 ^ n21282 ^ 1'b0 ;
  assign n21320 = ( n21282 & n21318 ) | ( n21282 & n21319 ) | ( n21318 & n21319 ) ;
  assign n21321 = ( n21178 & ~n21282 ) | ( n21178 & n21320 ) | ( ~n21282 & n21320 ) ;
  assign n21322 = x625 & ~n21321 ;
  assign n21323 = x625 | n21179 ;
  assign n21324 = ( x1153 & n21322 ) | ( x1153 & n21323 ) | ( n21322 & n21323 ) ;
  assign n21325 = ~n21322 & n21324 ;
  assign n21326 = ( x608 & n21249 ) | ( x608 & ~n21325 ) | ( n21249 & ~n21325 ) ;
  assign n21327 = ~n21249 & n21326 ;
  assign n21328 = x608 | n21245 ;
  assign n21329 = x625 & ~n21179 ;
  assign n21330 = x1153 | n21329 ;
  assign n21331 = ( n21321 & n21322 ) | ( n21321 & ~n21330 ) | ( n21322 & ~n21330 ) ;
  assign n21332 = ( ~n21327 & n21328 ) | ( ~n21327 & n21331 ) | ( n21328 & n21331 ) ;
  assign n21333 = ~n21327 & n21332 ;
  assign n21334 = n21321 ^ x778 ^ 1'b0 ;
  assign n21335 = ( n21321 & n21333 ) | ( n21321 & n21334 ) | ( n21333 & n21334 ) ;
  assign n21336 = x609 & ~n21335 ;
  assign n21337 = x609 | n21252 ;
  assign n21338 = ( x1155 & n21336 ) | ( x1155 & n21337 ) | ( n21336 & n21337 ) ;
  assign n21339 = ~n21336 & n21338 ;
  assign n21340 = ~x1155 & n21188 ;
  assign n21341 = ( x660 & n21339 ) | ( x660 & ~n21340 ) | ( n21339 & ~n21340 ) ;
  assign n21342 = ~n21339 & n21341 ;
  assign n21343 = x1155 & n21185 ;
  assign n21344 = x660 | n21343 ;
  assign n21345 = x609 & ~n21252 ;
  assign n21346 = x1155 | n21345 ;
  assign n21347 = ( n21335 & n21336 ) | ( n21335 & ~n21346 ) | ( n21336 & ~n21346 ) ;
  assign n21348 = ( ~n21342 & n21344 ) | ( ~n21342 & n21347 ) | ( n21344 & n21347 ) ;
  assign n21349 = ~n21342 & n21348 ;
  assign n21350 = n21335 ^ x785 ^ 1'b0 ;
  assign n21351 = ( n21335 & n21349 ) | ( n21335 & n21350 ) | ( n21349 & n21350 ) ;
  assign n21352 = x618 & ~n21351 ;
  assign n21353 = x618 | n21254 ;
  assign n21354 = ( x1154 & n21352 ) | ( x1154 & n21353 ) | ( n21352 & n21353 ) ;
  assign n21355 = ~n21352 & n21354 ;
  assign n21356 = ( x627 & n21199 ) | ( x627 & ~n21355 ) | ( n21199 & ~n21355 ) ;
  assign n21357 = ~n21199 & n21356 ;
  assign n21358 = x627 | n21196 ;
  assign n21359 = x618 & ~n21254 ;
  assign n21360 = x1154 | n21359 ;
  assign n21361 = ( n21351 & n21352 ) | ( n21351 & ~n21360 ) | ( n21352 & ~n21360 ) ;
  assign n21362 = ( ~n21357 & n21358 ) | ( ~n21357 & n21361 ) | ( n21358 & n21361 ) ;
  assign n21363 = ~n21357 & n21362 ;
  assign n21364 = n21351 ^ x781 ^ 1'b0 ;
  assign n21365 = ( n21351 & n21363 ) | ( n21351 & n21364 ) | ( n21363 & n21364 ) ;
  assign n21366 = x619 | n21365 ;
  assign n21367 = x619 & ~n21256 ;
  assign n21368 = ( x1159 & n21366 ) | ( x1159 & ~n21367 ) | ( n21366 & ~n21367 ) ;
  assign n21369 = ~x1159 & n21368 ;
  assign n21370 = ( x648 & n21206 ) | ( x648 & ~n21369 ) | ( n21206 & ~n21369 ) ;
  assign n21371 = n21369 | n21370 ;
  assign n21372 = x619 & ~n21365 ;
  assign n21373 = x619 | n21256 ;
  assign n21374 = ( x1159 & n21372 ) | ( x1159 & n21373 ) | ( n21372 & n21373 ) ;
  assign n21375 = ~n21372 & n21374 ;
  assign n21376 = ( x648 & n21209 ) | ( x648 & ~n21375 ) | ( n21209 & ~n21375 ) ;
  assign n21377 = ~n21209 & n21376 ;
  assign n21378 = x789 & ~n21377 ;
  assign n21379 = n21371 & n21378 ;
  assign n21380 = ~x789 & n21365 ;
  assign n21381 = ( n16519 & ~n21379 ) | ( n16519 & n21380 ) | ( ~n21379 & n21380 ) ;
  assign n21382 = n21379 | n21381 ;
  assign n21383 = n16317 & ~n21219 ;
  assign n21384 = n16459 & ~n21258 ;
  assign n21385 = ( x788 & n21383 ) | ( x788 & n21384 ) | ( n21383 & n21384 ) ;
  assign n21386 = n21384 ^ n21383 ^ 1'b0 ;
  assign n21387 = ( x788 & n21385 ) | ( x788 & n21386 ) | ( n21385 & n21386 ) ;
  assign n21388 = ( n18482 & n21382 ) | ( n18482 & ~n21387 ) | ( n21382 & ~n21387 ) ;
  assign n21389 = ~n18482 & n21388 ;
  assign n21390 = n21264 ^ x629 ^ 1'b0 ;
  assign n21391 = ( n21264 & n21267 ) | ( n21264 & n21390 ) | ( n21267 & n21390 ) ;
  assign n21392 = n19046 & n21221 ;
  assign n21393 = ( x792 & n21391 ) | ( x792 & n21392 ) | ( n21391 & n21392 ) ;
  assign n21394 = n21392 ^ n21391 ^ 1'b0 ;
  assign n21395 = ( x792 & n21393 ) | ( x792 & n21394 ) | ( n21393 & n21394 ) ;
  assign n21396 = ( ~n18484 & n21389 ) | ( ~n18484 & n21395 ) | ( n21389 & n21395 ) ;
  assign n21397 = ~n18484 & n21396 ;
  assign n21398 = n16374 & n21272 ;
  assign n21399 = n19055 & n21223 ;
  assign n21400 = n16373 & n21273 ;
  assign n21401 = ( ~n21398 & n21399 ) | ( ~n21398 & n21400 ) | ( n21399 & n21400 ) ;
  assign n21402 = n21398 | n21401 ;
  assign n21403 = n21397 ^ x787 ^ 1'b0 ;
  assign n21404 = ( ~x787 & n21402 ) | ( ~x787 & n21403 ) | ( n21402 & n21403 ) ;
  assign n21405 = ( x787 & n21397 ) | ( x787 & n21404 ) | ( n21397 & n21404 ) ;
  assign n21406 = ( x644 & ~n21281 ) | ( x644 & n21405 ) | ( ~n21281 & n21405 ) ;
  assign n21407 = ~n21281 & n21406 ;
  assign n21410 = ( x1160 & n21407 ) | ( x1160 & ~n21409 ) | ( n21407 & ~n21409 ) ;
  assign n21411 = n21409 | n21410 ;
  assign n21412 = x790 & ~n21411 ;
  assign n21413 = ( x790 & n21280 ) | ( x790 & n21412 ) | ( n21280 & n21412 ) ;
  assign n21414 = x644 & n21230 ;
  assign n21415 = x790 & ~n21414 ;
  assign n21416 = ( n21405 & ~n21413 ) | ( n21405 & n21415 ) | ( ~n21413 & n21415 ) ;
  assign n21417 = ~n21413 & n21416 ;
  assign n21418 = ( n7318 & ~n21162 ) | ( n7318 & n21417 ) | ( ~n21162 & n21417 ) ;
  assign n21419 = ~n21162 & n21418 ;
  assign n21420 = x173 | n1611 ;
  assign n21421 = ~n21310 & n21420 ;
  assign n21422 = n16397 | n21421 ;
  assign n21423 = ~n15662 & n21310 ;
  assign n21424 = ~x1155 & n21420 ;
  assign n21425 = ~n21423 & n21424 ;
  assign n21426 = ( x1155 & n21422 ) | ( x1155 & n21423 ) | ( n21422 & n21423 ) ;
  assign n21427 = n21425 | n21426 ;
  assign n21428 = n21422 ^ x785 ^ 1'b0 ;
  assign n21429 = ( n21422 & n21427 ) | ( n21422 & n21428 ) | ( n21427 & n21428 ) ;
  assign n21430 = n16411 | n21429 ;
  assign n21431 = x1154 & n21430 ;
  assign n21432 = n16414 | n21429 ;
  assign n21433 = ~x1154 & n21432 ;
  assign n21434 = n21431 | n21433 ;
  assign n21435 = n21429 ^ x781 ^ 1'b0 ;
  assign n21436 = ( n21429 & n21434 ) | ( n21429 & n21435 ) | ( n21434 & n21435 ) ;
  assign n21437 = ~x619 & n1611 ;
  assign n21438 = n21436 | n21437 ;
  assign n21439 = x1159 & n21438 ;
  assign n21440 = x619 & n1611 ;
  assign n21441 = n21436 | n21440 ;
  assign n21442 = ~x1159 & n21441 ;
  assign n21443 = n21439 | n21442 ;
  assign n21444 = n21436 ^ x789 ^ 1'b0 ;
  assign n21445 = ( n21436 & n21443 ) | ( n21436 & n21444 ) | ( n21443 & n21444 ) ;
  assign n21446 = x626 & ~n21445 ;
  assign n21447 = x626 & ~n21420 ;
  assign n21448 = x1158 | n21447 ;
  assign n21449 = ( n21445 & n21446 ) | ( n21445 & ~n21448 ) | ( n21446 & ~n21448 ) ;
  assign n21450 = n21446 & ~n21449 ;
  assign n21451 = ( x1158 & n21420 ) | ( x1158 & n21447 ) | ( n21420 & n21447 ) ;
  assign n21452 = ( n21449 & ~n21450 ) | ( n21449 & n21451 ) | ( ~n21450 & n21451 ) ;
  assign n21453 = n21445 ^ x788 ^ 1'b0 ;
  assign n21454 = ( n21445 & n21452 ) | ( n21445 & n21453 ) | ( n21452 & n21453 ) ;
  assign n21455 = n21420 ^ n16339 ^ 1'b0 ;
  assign n21456 = ( n21420 & n21454 ) | ( n21420 & ~n21455 ) | ( n21454 & ~n21455 ) ;
  assign n21457 = n19055 & n21456 ;
  assign n21458 = x647 & ~n21420 ;
  assign n21459 = x1157 | n21458 ;
  assign n21460 = ~x723 & n15778 ;
  assign n21461 = ~x625 & n21460 ;
  assign n21462 = ~x1153 & n21420 ;
  assign n21463 = ~n21461 & n21462 ;
  assign n21464 = x778 & ~n21463 ;
  assign n21465 = n21420 & ~n21460 ;
  assign n21466 = ( x1153 & n21461 ) | ( x1153 & n21465 ) | ( n21461 & n21465 ) ;
  assign n21467 = n21464 & ~n21466 ;
  assign n21468 = ( x778 & n21465 ) | ( x778 & ~n21467 ) | ( n21465 & ~n21467 ) ;
  assign n21469 = ~n21467 & n21468 ;
  assign n21470 = n16447 | n21469 ;
  assign n21471 = n16449 | n21470 ;
  assign n21472 = n16451 | n21471 ;
  assign n21473 = n16530 | n21472 ;
  assign n21474 = n16560 | n21473 ;
  assign n21475 = ( x647 & ~n21459 ) | ( x647 & n21474 ) | ( ~n21459 & n21474 ) ;
  assign n21476 = ~n21459 & n21475 ;
  assign n21477 = n21420 ^ x647 ^ 1'b0 ;
  assign n21478 = ( n21420 & n21474 ) | ( n21420 & n21477 ) | ( n21474 & n21477 ) ;
  assign n21479 = x1157 & n21478 ;
  assign n21480 = ( n16375 & n21476 ) | ( n16375 & n21479 ) | ( n21476 & n21479 ) ;
  assign n21481 = ( x787 & n21457 ) | ( x787 & n21480 ) | ( n21457 & n21480 ) ;
  assign n21482 = n21480 ^ n21457 ^ 1'b0 ;
  assign n21483 = ( x787 & n21481 ) | ( x787 & n21482 ) | ( n21481 & n21482 ) ;
  assign n21484 = n16459 & ~n21472 ;
  assign n21485 = n16317 & ~n21452 ;
  assign n21486 = ( x788 & n21484 ) | ( x788 & n21485 ) | ( n21484 & n21485 ) ;
  assign n21487 = n21485 ^ n21484 ^ 1'b0 ;
  assign n21488 = ( x788 & n21486 ) | ( x788 & n21487 ) | ( n21486 & n21487 ) ;
  assign n21489 = n15524 | n21465 ;
  assign n21490 = n21421 & n21489 ;
  assign n21491 = x625 & ~n21489 ;
  assign n21492 = ( n21462 & n21490 ) | ( n21462 & n21491 ) | ( n21490 & n21491 ) ;
  assign n21493 = ( x608 & n21466 ) | ( x608 & ~n21492 ) | ( n21466 & ~n21492 ) ;
  assign n21494 = n21492 | n21493 ;
  assign n21495 = x1153 & n21421 ;
  assign n21496 = ~n21491 & n21495 ;
  assign n21497 = x608 & ~n21463 ;
  assign n21498 = n21494 & ~n21497 ;
  assign n21499 = ( n21494 & n21496 ) | ( n21494 & n21498 ) | ( n21496 & n21498 ) ;
  assign n21500 = n21490 ^ x778 ^ 1'b0 ;
  assign n21501 = ( n21490 & n21499 ) | ( n21490 & n21500 ) | ( n21499 & n21500 ) ;
  assign n21502 = x609 & ~n21501 ;
  assign n21508 = x609 | n21469 ;
  assign n21509 = ( x1155 & n21502 ) | ( x1155 & n21508 ) | ( n21502 & n21508 ) ;
  assign n21510 = ~n21502 & n21509 ;
  assign n21511 = ( x660 & n21425 ) | ( x660 & ~n21510 ) | ( n21425 & ~n21510 ) ;
  assign n21512 = ~n21425 & n21511 ;
  assign n21503 = x609 & ~n21469 ;
  assign n21504 = x1155 | n21503 ;
  assign n21505 = ( n21501 & n21502 ) | ( n21501 & ~n21504 ) | ( n21502 & ~n21504 ) ;
  assign n21506 = ( x660 & n21426 ) | ( x660 & ~n21505 ) | ( n21426 & ~n21505 ) ;
  assign n21507 = n21505 | n21506 ;
  assign n21513 = n21512 ^ n21507 ^ 1'b0 ;
  assign n21514 = ( x785 & ~n21507 ) | ( x785 & n21512 ) | ( ~n21507 & n21512 ) ;
  assign n21515 = ( x785 & ~n21513 ) | ( x785 & n21514 ) | ( ~n21513 & n21514 ) ;
  assign n21516 = ( x785 & n21501 ) | ( x785 & ~n21515 ) | ( n21501 & ~n21515 ) ;
  assign n21517 = ~n21515 & n21516 ;
  assign n21518 = x618 & ~n21517 ;
  assign n21519 = x618 | n21470 ;
  assign n21520 = ( x1154 & n21518 ) | ( x1154 & n21519 ) | ( n21518 & n21519 ) ;
  assign n21521 = ~n21518 & n21520 ;
  assign n21522 = ( x627 & n21433 ) | ( x627 & ~n21521 ) | ( n21433 & ~n21521 ) ;
  assign n21523 = ~n21433 & n21522 ;
  assign n21524 = x627 | n21431 ;
  assign n21525 = x618 & ~n21470 ;
  assign n21526 = x1154 | n21525 ;
  assign n21527 = ( n21517 & n21518 ) | ( n21517 & ~n21526 ) | ( n21518 & ~n21526 ) ;
  assign n21528 = ( ~n21523 & n21524 ) | ( ~n21523 & n21527 ) | ( n21524 & n21527 ) ;
  assign n21529 = ~n21523 & n21528 ;
  assign n21530 = n21517 ^ x781 ^ 1'b0 ;
  assign n21531 = ( n21517 & n21529 ) | ( n21517 & n21530 ) | ( n21529 & n21530 ) ;
  assign n21532 = ~x789 & n21531 ;
  assign n21533 = x619 & ~n21471 ;
  assign n21534 = x1159 | n21533 ;
  assign n21535 = x619 & ~n21531 ;
  assign n21536 = ( n21531 & ~n21534 ) | ( n21531 & n21535 ) | ( ~n21534 & n21535 ) ;
  assign n21537 = ( x648 & n21439 ) | ( x648 & ~n21536 ) | ( n21439 & ~n21536 ) ;
  assign n21538 = n21536 | n21537 ;
  assign n21539 = x619 | n21471 ;
  assign n21540 = x1159 & ~n21535 ;
  assign n21541 = n21539 & n21540 ;
  assign n21542 = ( x648 & n21442 ) | ( x648 & ~n21541 ) | ( n21442 & ~n21541 ) ;
  assign n21543 = ~n21442 & n21542 ;
  assign n21544 = x789 & ~n21543 ;
  assign n21545 = n21538 & n21544 ;
  assign n21546 = ( n16519 & ~n21532 ) | ( n16519 & n21545 ) | ( ~n21532 & n21545 ) ;
  assign n21547 = n21532 | n21546 ;
  assign n21548 = n21547 ^ n21488 ^ 1'b0 ;
  assign n21549 = ( n21488 & n21547 ) | ( n21488 & n21548 ) | ( n21547 & n21548 ) ;
  assign n21550 = ( n18482 & ~n21488 ) | ( n18482 & n21549 ) | ( ~n21488 & n21549 ) ;
  assign n21551 = n16556 & ~n21454 ;
  assign n21552 = n19208 | n21473 ;
  assign n21553 = ( x629 & n21551 ) | ( x629 & n21552 ) | ( n21551 & n21552 ) ;
  assign n21554 = ~n21551 & n21553 ;
  assign n21555 = n19212 & ~n21473 ;
  assign n21556 = n16557 & ~n21454 ;
  assign n21557 = n21555 | n21556 ;
  assign n21558 = ( x629 & ~n21554 ) | ( x629 & n21557 ) | ( ~n21554 & n21557 ) ;
  assign n21559 = ~n21554 & n21558 ;
  assign n21560 = ( x792 & ~n19206 ) | ( x792 & n21559 ) | ( ~n19206 & n21559 ) ;
  assign n21561 = ( n18484 & n19206 ) | ( n18484 & n21560 ) | ( n19206 & n21560 ) ;
  assign n21562 = ( n21483 & n21550 ) | ( n21483 & ~n21561 ) | ( n21550 & ~n21561 ) ;
  assign n21563 = n21562 ^ n21550 ^ 1'b0 ;
  assign n21564 = ( n21483 & n21562 ) | ( n21483 & ~n21563 ) | ( n21562 & ~n21563 ) ;
  assign n21565 = x790 | n21564 ;
  assign n21566 = x832 & n21565 ;
  assign n21567 = x644 & ~n21564 ;
  assign n21568 = ( x787 & n21476 ) | ( x787 & ~n21479 ) | ( n21476 & ~n21479 ) ;
  assign n21569 = ~n21476 & n21568 ;
  assign n21570 = ( x787 & n21474 ) | ( x787 & ~n21569 ) | ( n21474 & ~n21569 ) ;
  assign n21571 = ~n21569 & n21570 ;
  assign n21572 = x644 | n21571 ;
  assign n21573 = ( x715 & n21567 ) | ( x715 & n21572 ) | ( n21567 & n21572 ) ;
  assign n21574 = ~n21567 & n21573 ;
  assign n21575 = x644 | n21420 ;
  assign n21576 = n21420 ^ n16376 ^ 1'b0 ;
  assign n21577 = ( n21420 & n21456 ) | ( n21420 & ~n21576 ) | ( n21456 & ~n21576 ) ;
  assign n21578 = x644 & ~n21577 ;
  assign n21579 = ( x715 & n21575 ) | ( x715 & ~n21578 ) | ( n21575 & ~n21578 ) ;
  assign n21580 = ~x715 & n21579 ;
  assign n21581 = ( x1160 & n21574 ) | ( x1160 & ~n21580 ) | ( n21574 & ~n21580 ) ;
  assign n21582 = ~n21574 & n21581 ;
  assign n21583 = x644 & ~n21420 ;
  assign n21584 = x715 & ~n21583 ;
  assign n21585 = ( n21577 & n21578 ) | ( n21577 & n21584 ) | ( n21578 & n21584 ) ;
  assign n21586 = x644 & ~n21571 ;
  assign n21587 = x715 | n21586 ;
  assign n21588 = ( n21564 & n21567 ) | ( n21564 & ~n21587 ) | ( n21567 & ~n21587 ) ;
  assign n21589 = ( x1160 & ~n21585 ) | ( x1160 & n21588 ) | ( ~n21585 & n21588 ) ;
  assign n21590 = n21585 | n21589 ;
  assign n21591 = x790 & ~n21590 ;
  assign n21592 = ( x790 & n21582 ) | ( x790 & n21591 ) | ( n21582 & n21591 ) ;
  assign n21593 = ( n21419 & n21566 ) | ( n21419 & ~n21592 ) | ( n21566 & ~n21592 ) ;
  assign n21594 = n21593 ^ n21566 ^ 1'b0 ;
  assign n21595 = ( n21419 & n21593 ) | ( n21419 & ~n21594 ) | ( n21593 & ~n21594 ) ;
  assign n21596 = x174 & ~n1611 ;
  assign n21597 = x759 & n15591 ;
  assign n21598 = ~n18309 & n21597 ;
  assign n21599 = ~n18321 & n21598 ;
  assign n21600 = ~x626 & n21599 ;
  assign n21601 = n21596 | n21600 ;
  assign n21602 = ( x641 & x1158 ) | ( x641 & ~n21601 ) | ( x1158 & ~n21601 ) ;
  assign n21603 = ( x641 & ~n16317 ) | ( x641 & n21602 ) | ( ~n16317 & n21602 ) ;
  assign n21604 = x696 & n15778 ;
  assign n21605 = n21596 | n21604 ;
  assign n21606 = x1153 & ~n21596 ;
  assign n21607 = x625 & n21604 ;
  assign n21608 = n21606 & ~n21607 ;
  assign n21609 = n21607 ^ n21604 ^ n21596 ;
  assign n21610 = x1153 | n21609 ;
  assign n21611 = ~n21608 & n21610 ;
  assign n21612 = n21605 ^ x778 ^ 1'b0 ;
  assign n21613 = ( n21605 & n21611 ) | ( n21605 & n21612 ) | ( n21611 & n21612 ) ;
  assign n21614 = ~n17087 & n21613 ;
  assign n21615 = ~n16279 & n21614 ;
  assign n21616 = n21596 | n21615 ;
  assign n21617 = ( n16453 & ~n21603 ) | ( n16453 & n21616 ) | ( ~n21603 & n21616 ) ;
  assign n21618 = n21617 ^ n21603 ^ 1'b0 ;
  assign n21619 = ( n21603 & ~n21617 ) | ( n21603 & n21618 ) | ( ~n21617 & n21618 ) ;
  assign n21620 = x626 & n21599 ;
  assign n21621 = n21596 | n21620 ;
  assign n21622 = ( x1158 & ~n16317 ) | ( x1158 & n21621 ) | ( ~n16317 & n21621 ) ;
  assign n21623 = ( x641 & n16317 ) | ( x641 & n21622 ) | ( n16317 & n21622 ) ;
  assign n21624 = n21623 ^ n16454 ^ 1'b0 ;
  assign n21625 = ( ~n16454 & n21616 ) | ( ~n16454 & n21624 ) | ( n21616 & n21624 ) ;
  assign n21626 = ( n16454 & n21623 ) | ( n16454 & n21625 ) | ( n21623 & n21625 ) ;
  assign n21627 = ( x788 & n21619 ) | ( x788 & n21626 ) | ( n21619 & n21626 ) ;
  assign n21628 = ~n21619 & n21627 ;
  assign n21629 = ( x619 & x648 ) | ( x619 & ~x1159 ) | ( x648 & ~x1159 ) ;
  assign n21630 = n21629 ^ x648 ^ 1'b0 ;
  assign n21631 = ~n18315 & n21598 ;
  assign n21632 = n18451 & n21631 ;
  assign n21633 = n16276 & ~n21632 ;
  assign n21634 = ~n18374 & n21631 ;
  assign n21635 = ~n21633 & n21634 ;
  assign n21636 = ( n16277 & n21633 ) | ( n16277 & ~n21635 ) | ( n21633 & ~n21635 ) ;
  assign n21637 = n21614 & ~n21636 ;
  assign n21638 = ( n21630 & n21636 ) | ( n21630 & ~n21637 ) | ( n21636 & ~n21637 ) ;
  assign n21639 = n21638 ^ n16519 ^ 1'b0 ;
  assign n21640 = x789 & ~n21596 ;
  assign n21641 = ( n21638 & ~n21639 ) | ( n21638 & n21640 ) | ( ~n21639 & n21640 ) ;
  assign n21642 = ( n16519 & n21639 ) | ( n16519 & n21641 ) | ( n21639 & n21641 ) ;
  assign n21643 = x608 | n21608 ;
  assign n21644 = n21596 | n21597 ;
  assign n21645 = x696 & n17156 ;
  assign n21646 = n21644 | n21645 ;
  assign n21647 = x625 & n21645 ;
  assign n21648 = n21646 & ~n21647 ;
  assign n21649 = ( x1153 & ~n21643 ) | ( x1153 & n21648 ) | ( ~n21643 & n21648 ) ;
  assign n21650 = ~n21643 & n21649 ;
  assign n21651 = x1153 & ~n21644 ;
  assign n21652 = ~n21647 & n21651 ;
  assign n21653 = ( x608 & n21610 ) | ( x608 & n21652 ) | ( n21610 & n21652 ) ;
  assign n21654 = ~n21652 & n21653 ;
  assign n21655 = ( x778 & n21650 ) | ( x778 & ~n21654 ) | ( n21650 & ~n21654 ) ;
  assign n21656 = ~n21650 & n21655 ;
  assign n21657 = ( x778 & n21646 ) | ( x778 & ~n21656 ) | ( n21646 & ~n21656 ) ;
  assign n21658 = ~n21656 & n21657 ;
  assign n21659 = ~x609 & n21658 ;
  assign n21660 = x609 & n21613 ;
  assign n21661 = ( x1155 & ~n21659 ) | ( x1155 & n21660 ) | ( ~n21659 & n21660 ) ;
  assign n21662 = n21659 | n21661 ;
  assign n21663 = x1155 | n21596 ;
  assign n21664 = ~n15662 & n21597 ;
  assign n21665 = n21663 | n21664 ;
  assign n21666 = ~x609 & n21613 ;
  assign n21667 = x609 & n21658 ;
  assign n21668 = ( x1155 & n21666 ) | ( x1155 & ~n21667 ) | ( n21666 & ~n21667 ) ;
  assign n21669 = ~n21666 & n21668 ;
  assign n21670 = x660 & ~n21669 ;
  assign n21671 = n21665 & n21670 ;
  assign n21672 = x1155 & ~n21596 ;
  assign n21673 = n15668 & n21597 ;
  assign n21674 = ( x660 & n21672 ) | ( x660 & ~n21673 ) | ( n21672 & ~n21673 ) ;
  assign n21675 = n21674 ^ n21672 ^ 1'b0 ;
  assign n21676 = ( x660 & n21674 ) | ( x660 & ~n21675 ) | ( n21674 & ~n21675 ) ;
  assign n21677 = ~n21671 & n21676 ;
  assign n21678 = ( n21662 & n21671 ) | ( n21662 & ~n21677 ) | ( n21671 & ~n21677 ) ;
  assign n21679 = n21658 ^ x785 ^ 1'b0 ;
  assign n21680 = ( n21658 & n21678 ) | ( n21658 & n21679 ) | ( n21678 & n21679 ) ;
  assign n21681 = ~x618 & n21680 ;
  assign n21682 = ~n16234 & n21613 ;
  assign n21683 = n21596 | n21682 ;
  assign n21684 = x618 & n21683 ;
  assign n21685 = ( x1154 & ~n21681 ) | ( x1154 & n21684 ) | ( ~n21681 & n21684 ) ;
  assign n21686 = n21681 | n21685 ;
  assign n21687 = x1154 & ~n21596 ;
  assign n21688 = n18431 & n21598 ;
  assign n21689 = n21687 & ~n21688 ;
  assign n21690 = ( x627 & n21686 ) | ( x627 & ~n21689 ) | ( n21686 & ~n21689 ) ;
  assign n21691 = ~x627 & n21690 ;
  assign n21692 = x1154 | n21596 ;
  assign n21693 = ~n18378 & n21598 ;
  assign n21694 = n21692 | n21693 ;
  assign n21695 = ~x618 & n21683 ;
  assign n21696 = x618 & n21680 ;
  assign n21697 = ( x1154 & n21695 ) | ( x1154 & ~n21696 ) | ( n21695 & ~n21696 ) ;
  assign n21698 = ~n21695 & n21697 ;
  assign n21699 = x627 & ~n21698 ;
  assign n21700 = n21694 & n21699 ;
  assign n21701 = ( x781 & n21691 ) | ( x781 & n21700 ) | ( n21691 & n21700 ) ;
  assign n21702 = n21700 ^ n21691 ^ 1'b0 ;
  assign n21703 = ( x781 & n21701 ) | ( x781 & n21702 ) | ( n21701 & n21702 ) ;
  assign n21704 = n16278 | n21630 ;
  assign n21705 = x789 & n21704 ;
  assign n21706 = ~x781 & n21680 ;
  assign n21707 = n21705 | n21706 ;
  assign n21708 = ( ~n21642 & n21703 ) | ( ~n21642 & n21707 ) | ( n21703 & n21707 ) ;
  assign n21709 = ~n21642 & n21708 ;
  assign n21710 = ( n18482 & ~n21628 ) | ( n18482 & n21709 ) | ( ~n21628 & n21709 ) ;
  assign n21711 = n21628 | n21710 ;
  assign n21712 = ~n17088 & n21613 ;
  assign n21713 = x628 & n21712 ;
  assign n21714 = ~n16518 & n21599 ;
  assign n21715 = x628 | n21714 ;
  assign n21716 = x629 & n21715 ;
  assign n21717 = ( x1156 & n21713 ) | ( x1156 & ~n21716 ) | ( n21713 & ~n21716 ) ;
  assign n21718 = ~n21713 & n21717 ;
  assign n21719 = x629 & ~n21712 ;
  assign n21720 = ~x629 & n21714 ;
  assign n21721 = ~n21719 & n21720 ;
  assign n21722 = ( x628 & n21719 ) | ( x628 & ~n21721 ) | ( n21719 & ~n21721 ) ;
  assign n21723 = ( ~x1156 & n21718 ) | ( ~x1156 & n21722 ) | ( n21718 & n21722 ) ;
  assign n21724 = n21718 ^ x1156 ^ 1'b0 ;
  assign n21725 = ( n21718 & n21723 ) | ( n21718 & ~n21724 ) | ( n21723 & ~n21724 ) ;
  assign n21726 = x792 & ~n21596 ;
  assign n21727 = n21725 & n21726 ;
  assign n21728 = ( n18484 & n21711 ) | ( n18484 & ~n21727 ) | ( n21711 & ~n21727 ) ;
  assign n21729 = n21728 ^ n21711 ^ 1'b0 ;
  assign n21730 = ( n18484 & n21728 ) | ( n18484 & ~n21729 ) | ( n21728 & ~n21729 ) ;
  assign n21733 = ~n17093 & n21712 ;
  assign n21734 = x630 & ~n21733 ;
  assign n21735 = ( x647 & n21733 ) | ( x647 & n21734 ) | ( n21733 & n21734 ) ;
  assign n21731 = ~n16339 & n21714 ;
  assign n21732 = x630 & n21731 ;
  assign n21736 = ( x1157 & ~n21732 ) | ( x1157 & n21735 ) | ( ~n21732 & n21735 ) ;
  assign n21737 = ~n21735 & n21736 ;
  assign n21738 = ~x630 & n21731 ;
  assign n21739 = ~n21734 & n21738 ;
  assign n21740 = ( x647 & n21734 ) | ( x647 & ~n21739 ) | ( n21734 & ~n21739 ) ;
  assign n21741 = ( ~x1157 & n21737 ) | ( ~x1157 & n21740 ) | ( n21737 & n21740 ) ;
  assign n21742 = n21737 ^ x1157 ^ 1'b0 ;
  assign n21743 = ( n21737 & n21741 ) | ( n21737 & ~n21742 ) | ( n21741 & ~n21742 ) ;
  assign n21744 = x787 & ~n21596 ;
  assign n21745 = n21730 & ~n21744 ;
  assign n21746 = ( n21730 & ~n21743 ) | ( n21730 & n21745 ) | ( ~n21743 & n21745 ) ;
  assign n21747 = ~x790 & n21746 ;
  assign n21748 = ~x644 & n21746 ;
  assign n21749 = ~n17273 & n21733 ;
  assign n21750 = n21596 | n21749 ;
  assign n21751 = x644 & n21750 ;
  assign n21752 = ( x715 & ~n21748 ) | ( x715 & n21751 ) | ( ~n21748 & n21751 ) ;
  assign n21753 = n21748 | n21752 ;
  assign n21754 = x715 & ~n21596 ;
  assign n21755 = n16339 | n16376 ;
  assign n21756 = n21714 & ~n21755 ;
  assign n21757 = ~x644 & n21756 ;
  assign n21758 = n21754 & ~n21757 ;
  assign n21759 = ( x1160 & n21753 ) | ( x1160 & ~n21758 ) | ( n21753 & ~n21758 ) ;
  assign n21760 = ~x1160 & n21759 ;
  assign n21761 = x715 | n21596 ;
  assign n21762 = x644 & n21756 ;
  assign n21763 = n21761 | n21762 ;
  assign n21764 = ~x644 & n21750 ;
  assign n21765 = x644 & n21746 ;
  assign n21766 = ( x715 & n21764 ) | ( x715 & ~n21765 ) | ( n21764 & ~n21765 ) ;
  assign n21767 = ~n21764 & n21766 ;
  assign n21768 = x1160 & ~n21767 ;
  assign n21769 = n21763 & n21768 ;
  assign n21770 = ( x790 & n21760 ) | ( x790 & n21769 ) | ( n21760 & n21769 ) ;
  assign n21771 = n21769 ^ n21760 ^ 1'b0 ;
  assign n21772 = ( x790 & n21770 ) | ( x790 & n21771 ) | ( n21770 & n21771 ) ;
  assign n21773 = ( x832 & n21747 ) | ( x832 & ~n21772 ) | ( n21747 & ~n21772 ) ;
  assign n21774 = ~n21747 & n21773 ;
  assign n21775 = ~x174 & n5193 ;
  assign n21776 = x174 & ~n15656 ;
  assign n21821 = ~x626 & n21776 ;
  assign n21822 = n21776 ^ n15659 ^ 1'b0 ;
  assign n21823 = x174 & n2069 ;
  assign n21782 = x174 | n15644 ;
  assign n21824 = x759 & n15524 ;
  assign n21825 = n15644 & ~n21824 ;
  assign n21826 = x38 & ~n21825 ;
  assign n21827 = n21782 & n21826 ;
  assign n21828 = ~x174 & x759 ;
  assign n21829 = n15640 & n21828 ;
  assign n21830 = x759 & ~n15585 ;
  assign n21831 = x39 & ~n19823 ;
  assign n21832 = ( x39 & n21830 ) | ( x39 & n21831 ) | ( n21830 & n21831 ) ;
  assign n21833 = x759 & n15509 ;
  assign n21834 = ~x759 & n15332 ;
  assign n21835 = x39 | n21834 ;
  assign n21836 = ( ~n21832 & n21833 ) | ( ~n21832 & n21835 ) | ( n21833 & n21835 ) ;
  assign n21837 = ~n21832 & n21836 ;
  assign n21838 = ~n21829 & n21837 ;
  assign n21839 = ( x174 & n21829 ) | ( x174 & ~n21838 ) | ( n21829 & ~n21838 ) ;
  assign n21840 = ( ~x38 & n21827 ) | ( ~x38 & n21839 ) | ( n21827 & n21839 ) ;
  assign n21841 = n21827 ^ x38 ^ 1'b0 ;
  assign n21842 = ( n21827 & n21840 ) | ( n21827 & ~n21841 ) | ( n21840 & ~n21841 ) ;
  assign n21843 = ~n2069 & n21842 ;
  assign n21844 = n21823 | n21843 ;
  assign n21845 = ( n21776 & ~n21822 ) | ( n21776 & n21844 ) | ( ~n21822 & n21844 ) ;
  assign n21846 = x609 & ~n21845 ;
  assign n21847 = x609 | n21776 ;
  assign n21848 = ( x1155 & n21846 ) | ( x1155 & n21847 ) | ( n21846 & n21847 ) ;
  assign n21849 = ~n21846 & n21848 ;
  assign n21850 = x609 & ~n21776 ;
  assign n21851 = x1155 | n21850 ;
  assign n21852 = ( n21845 & n21846 ) | ( n21845 & ~n21851 ) | ( n21846 & ~n21851 ) ;
  assign n21853 = n21849 | n21852 ;
  assign n21854 = n21845 ^ x785 ^ 1'b0 ;
  assign n21855 = ( n21845 & n21853 ) | ( n21845 & n21854 ) | ( n21853 & n21854 ) ;
  assign n21856 = x618 & ~n21855 ;
  assign n21857 = x618 | n21776 ;
  assign n21858 = ( x1154 & n21856 ) | ( x1154 & n21857 ) | ( n21856 & n21857 ) ;
  assign n21859 = ~n21856 & n21858 ;
  assign n21860 = x618 & ~n21776 ;
  assign n21861 = x1154 | n21860 ;
  assign n21862 = ( n21855 & n21856 ) | ( n21855 & ~n21861 ) | ( n21856 & ~n21861 ) ;
  assign n21863 = n21859 | n21862 ;
  assign n21864 = n21855 ^ x781 ^ 1'b0 ;
  assign n21865 = ( n21855 & n21863 ) | ( n21855 & n21864 ) | ( n21863 & n21864 ) ;
  assign n21866 = x619 & ~n21865 ;
  assign n21867 = x619 | n21776 ;
  assign n21868 = ( x1159 & n21866 ) | ( x1159 & n21867 ) | ( n21866 & n21867 ) ;
  assign n21869 = ~n21866 & n21868 ;
  assign n21870 = x619 & ~n21776 ;
  assign n21871 = x1159 | n21870 ;
  assign n21872 = ( n21865 & n21866 ) | ( n21865 & ~n21871 ) | ( n21866 & ~n21871 ) ;
  assign n21873 = n21869 | n21872 ;
  assign n21874 = n21865 ^ x789 ^ 1'b0 ;
  assign n21875 = ( n21865 & n21873 ) | ( n21865 & n21874 ) | ( n21873 & n21874 ) ;
  assign n21876 = x626 & n21875 ;
  assign n21877 = ( x641 & ~n21821 ) | ( x641 & n21876 ) | ( ~n21821 & n21876 ) ;
  assign n21878 = n21821 | n21877 ;
  assign n21777 = x174 | n16699 ;
  assign n21778 = x174 & n16697 ;
  assign n21779 = ( x38 & n21777 ) | ( x38 & ~n21778 ) | ( n21777 & ~n21778 ) ;
  assign n21780 = ~x38 & n21779 ;
  assign n21781 = x696 & ~n2069 ;
  assign n21783 = n18524 & n21782 ;
  assign n21784 = ( n21780 & n21781 ) | ( n21780 & ~n21783 ) | ( n21781 & ~n21783 ) ;
  assign n21785 = ~n21780 & n21784 ;
  assign n21786 = ( n21776 & n21781 ) | ( n21776 & ~n21785 ) | ( n21781 & ~n21785 ) ;
  assign n21787 = ~n21785 & n21786 ;
  assign n21788 = x625 & ~n21787 ;
  assign n21789 = x625 | n21776 ;
  assign n21790 = ( x1153 & n21788 ) | ( x1153 & n21789 ) | ( n21788 & n21789 ) ;
  assign n21791 = ~n21788 & n21790 ;
  assign n21792 = x625 & ~n21776 ;
  assign n21793 = x1153 | n21792 ;
  assign n21794 = ( x625 & n21787 ) | ( x625 & ~n21793 ) | ( n21787 & ~n21793 ) ;
  assign n21795 = ~n21793 & n21794 ;
  assign n21796 = n21791 | n21795 ;
  assign n21797 = n21787 ^ x778 ^ 1'b0 ;
  assign n21798 = ( n21787 & n21796 ) | ( n21787 & n21797 ) | ( n21796 & n21797 ) ;
  assign n21799 = n21776 ^ n16234 ^ 1'b0 ;
  assign n21800 = ( n21776 & n21798 ) | ( n21776 & ~n21799 ) | ( n21798 & ~n21799 ) ;
  assign n21801 = n21776 ^ n16254 ^ 1'b0 ;
  assign n21802 = ( n21776 & n21800 ) | ( n21776 & ~n21801 ) | ( n21800 & ~n21801 ) ;
  assign n21803 = n21776 ^ n16279 ^ 1'b0 ;
  assign n21804 = ( n21776 & n21802 ) | ( n21776 & ~n21803 ) | ( n21802 & ~n21803 ) ;
  assign n21879 = ~x626 & n21804 ;
  assign n21880 = x174 & n16048 ;
  assign n21881 = x174 | n16054 ;
  assign n21882 = ( x759 & n21880 ) | ( x759 & n21881 ) | ( n21880 & n21881 ) ;
  assign n21883 = ~n21880 & n21882 ;
  assign n21884 = x174 | n16029 ;
  assign n21885 = x174 & n16044 ;
  assign n21886 = ( x759 & n21884 ) | ( x759 & ~n21885 ) | ( n21884 & ~n21885 ) ;
  assign n21887 = ~x759 & n21886 ;
  assign n21888 = ( x39 & ~n21883 ) | ( x39 & n21887 ) | ( ~n21883 & n21887 ) ;
  assign n21889 = n21883 | n21888 ;
  assign n21890 = x174 | n15795 ;
  assign n21891 = x174 & n15876 ;
  assign n21892 = ( x759 & n21890 ) | ( x759 & ~n21891 ) | ( n21890 & ~n21891 ) ;
  assign n21893 = ~x759 & n21892 ;
  assign n21894 = x174 & n16003 ;
  assign n21895 = x174 | n15943 ;
  assign n21896 = ( x759 & n21894 ) | ( x759 & n21895 ) | ( n21894 & n21895 ) ;
  assign n21897 = ~n21894 & n21896 ;
  assign n21898 = ( x39 & n21893 ) | ( x39 & ~n21897 ) | ( n21893 & ~n21897 ) ;
  assign n21899 = ~n21893 & n21898 ;
  assign n21900 = ( x38 & n21889 ) | ( x38 & ~n21899 ) | ( n21889 & ~n21899 ) ;
  assign n21901 = ~x38 & n21900 ;
  assign n21902 = x696 & ~n17882 ;
  assign n21903 = ( n21827 & ~n21901 ) | ( n21827 & n21902 ) | ( ~n21901 & n21902 ) ;
  assign n21904 = ~n21827 & n21903 ;
  assign n21905 = ( n2051 & n2068 ) | ( n2051 & ~n21904 ) | ( n2068 & ~n21904 ) ;
  assign n21906 = n21904 | n21905 ;
  assign n21907 = ( x696 & n21842 ) | ( x696 & ~n21906 ) | ( n21842 & ~n21906 ) ;
  assign n21908 = ~n21906 & n21907 ;
  assign n21909 = n21908 ^ x174 ^ 1'b0 ;
  assign n21910 = ( ~x174 & n2069 ) | ( ~x174 & n21909 ) | ( n2069 & n21909 ) ;
  assign n21911 = ( x174 & n21908 ) | ( x174 & n21910 ) | ( n21908 & n21910 ) ;
  assign n21912 = x625 & ~n21911 ;
  assign n21918 = x625 | n21844 ;
  assign n21919 = ( x1153 & n21912 ) | ( x1153 & n21918 ) | ( n21912 & n21918 ) ;
  assign n21920 = ~n21912 & n21919 ;
  assign n21921 = ( x608 & ~n21795 ) | ( x608 & n21920 ) | ( ~n21795 & n21920 ) ;
  assign n21922 = ~n21920 & n21921 ;
  assign n21913 = x625 & ~n21844 ;
  assign n21914 = x1153 | n21913 ;
  assign n21915 = ( n21911 & n21912 ) | ( n21911 & ~n21914 ) | ( n21912 & ~n21914 ) ;
  assign n21916 = ( x608 & ~n21791 ) | ( x608 & n21915 ) | ( ~n21791 & n21915 ) ;
  assign n21917 = n21791 | n21916 ;
  assign n21923 = n21922 ^ n21917 ^ 1'b0 ;
  assign n21924 = ( x778 & ~n21917 ) | ( x778 & n21922 ) | ( ~n21917 & n21922 ) ;
  assign n21925 = ( x778 & ~n21923 ) | ( x778 & n21924 ) | ( ~n21923 & n21924 ) ;
  assign n21926 = ( x778 & n21911 ) | ( x778 & ~n21925 ) | ( n21911 & ~n21925 ) ;
  assign n21927 = ~n21925 & n21926 ;
  assign n21928 = x609 & ~n21927 ;
  assign n21934 = x609 | n21798 ;
  assign n21935 = ( x1155 & n21928 ) | ( x1155 & n21934 ) | ( n21928 & n21934 ) ;
  assign n21936 = ~n21928 & n21935 ;
  assign n21937 = ( x660 & ~n21852 ) | ( x660 & n21936 ) | ( ~n21852 & n21936 ) ;
  assign n21938 = ~n21936 & n21937 ;
  assign n21929 = x609 & ~n21798 ;
  assign n21930 = x1155 | n21929 ;
  assign n21931 = ( n21927 & n21928 ) | ( n21927 & ~n21930 ) | ( n21928 & ~n21930 ) ;
  assign n21932 = ( x660 & ~n21849 ) | ( x660 & n21931 ) | ( ~n21849 & n21931 ) ;
  assign n21933 = n21849 | n21932 ;
  assign n21939 = n21938 ^ n21933 ^ 1'b0 ;
  assign n21940 = ( x785 & ~n21933 ) | ( x785 & n21938 ) | ( ~n21933 & n21938 ) ;
  assign n21941 = ( x785 & ~n21939 ) | ( x785 & n21940 ) | ( ~n21939 & n21940 ) ;
  assign n21942 = ( x785 & n21927 ) | ( x785 & ~n21941 ) | ( n21927 & ~n21941 ) ;
  assign n21943 = ~n21941 & n21942 ;
  assign n21944 = x618 & ~n21943 ;
  assign n21950 = x618 | n21800 ;
  assign n21951 = ( x1154 & n21944 ) | ( x1154 & n21950 ) | ( n21944 & n21950 ) ;
  assign n21952 = ~n21944 & n21951 ;
  assign n21953 = ( x627 & ~n21862 ) | ( x627 & n21952 ) | ( ~n21862 & n21952 ) ;
  assign n21954 = ~n21952 & n21953 ;
  assign n21945 = x618 & ~n21800 ;
  assign n21946 = x1154 | n21945 ;
  assign n21947 = ( n21943 & n21944 ) | ( n21943 & ~n21946 ) | ( n21944 & ~n21946 ) ;
  assign n21948 = ( x627 & ~n21859 ) | ( x627 & n21947 ) | ( ~n21859 & n21947 ) ;
  assign n21949 = n21859 | n21948 ;
  assign n21955 = n21954 ^ n21949 ^ 1'b0 ;
  assign n21956 = ( x781 & ~n21949 ) | ( x781 & n21954 ) | ( ~n21949 & n21954 ) ;
  assign n21957 = ( x781 & ~n21955 ) | ( x781 & n21956 ) | ( ~n21955 & n21956 ) ;
  assign n21958 = ( x781 & n21943 ) | ( x781 & ~n21957 ) | ( n21943 & ~n21957 ) ;
  assign n21959 = ~n21957 & n21958 ;
  assign n21960 = x619 & ~n21959 ;
  assign n21966 = x619 | n21802 ;
  assign n21967 = ( x1159 & n21960 ) | ( x1159 & n21966 ) | ( n21960 & n21966 ) ;
  assign n21968 = ~n21960 & n21967 ;
  assign n21969 = ( x648 & ~n21872 ) | ( x648 & n21968 ) | ( ~n21872 & n21968 ) ;
  assign n21970 = ~n21968 & n21969 ;
  assign n21961 = x619 & ~n21802 ;
  assign n21962 = x1159 | n21961 ;
  assign n21963 = ( n21959 & n21960 ) | ( n21959 & ~n21962 ) | ( n21960 & ~n21962 ) ;
  assign n21964 = ( x648 & ~n21869 ) | ( x648 & n21963 ) | ( ~n21869 & n21963 ) ;
  assign n21965 = n21869 | n21964 ;
  assign n21971 = n21970 ^ n21965 ^ 1'b0 ;
  assign n21972 = ( x789 & ~n21965 ) | ( x789 & n21970 ) | ( ~n21965 & n21970 ) ;
  assign n21973 = ( x789 & ~n21971 ) | ( x789 & n21972 ) | ( ~n21971 & n21972 ) ;
  assign n21974 = ( x789 & n21959 ) | ( x789 & ~n21973 ) | ( n21959 & ~n21973 ) ;
  assign n21975 = ~n21973 & n21974 ;
  assign n21976 = x626 & n21975 ;
  assign n21977 = ( x641 & n21879 ) | ( x641 & ~n21976 ) | ( n21879 & ~n21976 ) ;
  assign n21978 = ~n21879 & n21977 ;
  assign n21979 = x1158 & ~n21978 ;
  assign n21980 = n21878 & n21979 ;
  assign n21981 = ~x626 & n21975 ;
  assign n21982 = x626 & n21804 ;
  assign n21983 = ( x641 & ~n21981 ) | ( x641 & n21982 ) | ( ~n21981 & n21982 ) ;
  assign n21984 = n21981 | n21983 ;
  assign n21985 = ~x626 & n21875 ;
  assign n21986 = x626 & n21776 ;
  assign n21987 = ( x641 & n21985 ) | ( x641 & ~n21986 ) | ( n21985 & ~n21986 ) ;
  assign n21988 = ~n21985 & n21987 ;
  assign n21989 = ( x1158 & n21984 ) | ( x1158 & ~n21988 ) | ( n21984 & ~n21988 ) ;
  assign n21990 = ~x1158 & n21989 ;
  assign n21991 = ( x788 & n21980 ) | ( x788 & ~n21990 ) | ( n21980 & ~n21990 ) ;
  assign n21992 = ~n21980 & n21991 ;
  assign n21993 = ( x788 & n21975 ) | ( x788 & ~n21992 ) | ( n21975 & ~n21992 ) ;
  assign n21994 = ~n21992 & n21993 ;
  assign n21995 = x628 & ~n21994 ;
  assign n21996 = n21776 ^ n16518 ^ 1'b0 ;
  assign n21997 = ( n21776 & n21875 ) | ( n21776 & ~n21996 ) | ( n21875 & ~n21996 ) ;
  assign n22003 = x628 | n21997 ;
  assign n22004 = ( x1156 & n21995 ) | ( x1156 & n22003 ) | ( n21995 & n22003 ) ;
  assign n22005 = ~n21995 & n22004 ;
  assign n21805 = n21776 ^ n16318 ^ 1'b0 ;
  assign n21806 = ( n21776 & n21804 ) | ( n21776 & ~n21805 ) | ( n21804 & ~n21805 ) ;
  assign n21807 = x628 & ~n21806 ;
  assign n21811 = x628 & ~n21776 ;
  assign n21812 = x1156 | n21811 ;
  assign n21813 = ( n21806 & n21807 ) | ( n21806 & ~n21812 ) | ( n21807 & ~n21812 ) ;
  assign n22006 = ( x629 & ~n21813 ) | ( x629 & n22005 ) | ( ~n21813 & n22005 ) ;
  assign n22007 = ~n22005 & n22006 ;
  assign n21808 = x628 | n21776 ;
  assign n21809 = ( x1156 & n21807 ) | ( x1156 & n21808 ) | ( n21807 & n21808 ) ;
  assign n21810 = ~n21807 & n21809 ;
  assign n21998 = x628 & ~n21997 ;
  assign n21999 = x1156 | n21998 ;
  assign n22000 = ( n21994 & n21995 ) | ( n21994 & ~n21999 ) | ( n21995 & ~n21999 ) ;
  assign n22001 = ( x629 & ~n21810 ) | ( x629 & n22000 ) | ( ~n21810 & n22000 ) ;
  assign n22002 = n21810 | n22001 ;
  assign n22008 = n22007 ^ n22002 ^ 1'b0 ;
  assign n22009 = ( x792 & ~n22002 ) | ( x792 & n22007 ) | ( ~n22002 & n22007 ) ;
  assign n22010 = ( x792 & ~n22008 ) | ( x792 & n22009 ) | ( ~n22008 & n22009 ) ;
  assign n22011 = ( x792 & n21994 ) | ( x792 & ~n22010 ) | ( n21994 & ~n22010 ) ;
  assign n22012 = ~n22010 & n22011 ;
  assign n22013 = x647 & ~n22012 ;
  assign n22014 = n21776 ^ n16339 ^ 1'b0 ;
  assign n22015 = ( n21776 & n21997 ) | ( n21776 & ~n22014 ) | ( n21997 & ~n22014 ) ;
  assign n22021 = x647 | n22015 ;
  assign n22022 = ( x1157 & n22013 ) | ( x1157 & n22021 ) | ( n22013 & n22021 ) ;
  assign n22023 = ~n22013 & n22022 ;
  assign n21814 = n21810 | n21813 ;
  assign n21815 = n21806 ^ x792 ^ 1'b0 ;
  assign n21816 = ( n21806 & n21814 ) | ( n21806 & n21815 ) | ( n21814 & n21815 ) ;
  assign n21817 = x647 & ~n21816 ;
  assign n22024 = x647 & ~n21776 ;
  assign n22025 = x1157 | n22024 ;
  assign n22026 = ( n21816 & n21817 ) | ( n21816 & ~n22025 ) | ( n21817 & ~n22025 ) ;
  assign n22027 = ( x630 & n22023 ) | ( x630 & ~n22026 ) | ( n22023 & ~n22026 ) ;
  assign n22028 = ~n22023 & n22027 ;
  assign n21818 = x647 | n21776 ;
  assign n21819 = ( x1157 & n21817 ) | ( x1157 & n21818 ) | ( n21817 & n21818 ) ;
  assign n21820 = ~n21817 & n21819 ;
  assign n22016 = x647 & ~n22015 ;
  assign n22017 = x1157 | n22016 ;
  assign n22018 = ( n22012 & n22013 ) | ( n22012 & ~n22017 ) | ( n22013 & ~n22017 ) ;
  assign n22019 = ( x630 & ~n21820 ) | ( x630 & n22018 ) | ( ~n21820 & n22018 ) ;
  assign n22020 = n21820 | n22019 ;
  assign n22029 = n22028 ^ n22020 ^ 1'b0 ;
  assign n22030 = ( x787 & ~n22020 ) | ( x787 & n22028 ) | ( ~n22020 & n22028 ) ;
  assign n22031 = ( x787 & ~n22029 ) | ( x787 & n22030 ) | ( ~n22029 & n22030 ) ;
  assign n22032 = ( x787 & n22012 ) | ( x787 & ~n22031 ) | ( n22012 & ~n22031 ) ;
  assign n22033 = ~n22031 & n22032 ;
  assign n22034 = ~x790 & n22033 ;
  assign n22042 = x644 & ~n21776 ;
  assign n22043 = x715 & ~n22042 ;
  assign n22044 = n21776 ^ n16376 ^ 1'b0 ;
  assign n22045 = ( n21776 & n22015 ) | ( n21776 & ~n22044 ) | ( n22015 & ~n22044 ) ;
  assign n22046 = x644 & ~n22045 ;
  assign n22047 = ( n22043 & n22045 ) | ( n22043 & n22046 ) | ( n22045 & n22046 ) ;
  assign n22035 = x644 | n22033 ;
  assign n22036 = n21820 | n22026 ;
  assign n22037 = n21816 ^ x787 ^ 1'b0 ;
  assign n22038 = ( n21816 & n22036 ) | ( n21816 & n22037 ) | ( n22036 & n22037 ) ;
  assign n22039 = x644 & ~n22038 ;
  assign n22040 = ( x715 & n22035 ) | ( x715 & ~n22039 ) | ( n22035 & ~n22039 ) ;
  assign n22041 = ~x715 & n22040 ;
  assign n22048 = ( x1160 & n22041 ) | ( x1160 & ~n22047 ) | ( n22041 & ~n22047 ) ;
  assign n22049 = n22047 | n22048 ;
  assign n22050 = x644 & ~n22033 ;
  assign n22051 = x644 | n22038 ;
  assign n22052 = ( x715 & n22050 ) | ( x715 & n22051 ) | ( n22050 & n22051 ) ;
  assign n22053 = ~n22050 & n22052 ;
  assign n22054 = x644 | n21776 ;
  assign n22055 = ( x715 & ~n22046 ) | ( x715 & n22054 ) | ( ~n22046 & n22054 ) ;
  assign n22056 = ~x715 & n22055 ;
  assign n22057 = ( x1160 & n22053 ) | ( x1160 & ~n22056 ) | ( n22053 & ~n22056 ) ;
  assign n22058 = ~n22053 & n22057 ;
  assign n22059 = x790 & ~n22058 ;
  assign n22060 = n22049 & n22059 ;
  assign n22061 = ( n5193 & ~n22034 ) | ( n5193 & n22060 ) | ( ~n22034 & n22060 ) ;
  assign n22062 = n22034 | n22061 ;
  assign n22063 = ( x57 & ~n21775 ) | ( x57 & n22062 ) | ( ~n21775 & n22062 ) ;
  assign n22064 = ~x57 & n22063 ;
  assign n22065 = x57 & x174 ;
  assign n22066 = x832 | n22065 ;
  assign n22067 = ( ~n21774 & n22064 ) | ( ~n21774 & n22066 ) | ( n22064 & n22066 ) ;
  assign n22068 = ~n21774 & n22067 ;
  assign n22069 = x175 | n15656 ;
  assign n22070 = x175 | n15644 ;
  assign n22071 = n16185 & n22070 ;
  assign n22072 = x175 | n16697 ;
  assign n22073 = x175 & n16699 ;
  assign n22074 = ( x38 & n22072 ) | ( x38 & ~n22073 ) | ( n22072 & ~n22073 ) ;
  assign n22075 = ~x38 & n22074 ;
  assign n22076 = ( x700 & n22071 ) | ( x700 & ~n22075 ) | ( n22071 & ~n22075 ) ;
  assign n22077 = ~n22071 & n22076 ;
  assign n22078 = x175 | x700 ;
  assign n22079 = n15655 | n22078 ;
  assign n22080 = ( n2069 & ~n22077 ) | ( n2069 & n22079 ) | ( ~n22077 & n22079 ) ;
  assign n22081 = ~n2069 & n22080 ;
  assign n22082 = n22081 ^ x175 ^ 1'b0 ;
  assign n22083 = ( ~x175 & n2069 ) | ( ~x175 & n22082 ) | ( n2069 & n22082 ) ;
  assign n22084 = ( x175 & n22081 ) | ( x175 & n22083 ) | ( n22081 & n22083 ) ;
  assign n22085 = x625 & ~n22084 ;
  assign n22086 = x625 | n22069 ;
  assign n22087 = ( x1153 & n22085 ) | ( x1153 & n22086 ) | ( n22085 & n22086 ) ;
  assign n22088 = ~n22085 & n22087 ;
  assign n22089 = x625 & ~n22069 ;
  assign n22090 = x1153 | n22089 ;
  assign n22091 = ( x625 & n22084 ) | ( x625 & ~n22090 ) | ( n22084 & ~n22090 ) ;
  assign n22092 = ~n22090 & n22091 ;
  assign n22093 = n22088 | n22092 ;
  assign n22094 = n22084 ^ x778 ^ 1'b0 ;
  assign n22095 = ( n22084 & n22093 ) | ( n22084 & n22094 ) | ( n22093 & n22094 ) ;
  assign n22096 = n22069 ^ n16234 ^ 1'b0 ;
  assign n22097 = ( n22069 & n22095 ) | ( n22069 & ~n22096 ) | ( n22095 & ~n22096 ) ;
  assign n22098 = n22069 ^ n16254 ^ 1'b0 ;
  assign n22099 = ( n22069 & n22097 ) | ( n22069 & ~n22098 ) | ( n22097 & ~n22098 ) ;
  assign n22100 = n22069 ^ n16279 ^ 1'b0 ;
  assign n22101 = ( n22069 & n22099 ) | ( n22069 & ~n22100 ) | ( n22099 & ~n22100 ) ;
  assign n22102 = n22069 ^ n16318 ^ 1'b0 ;
  assign n22103 = ( n22069 & n22101 ) | ( n22069 & ~n22102 ) | ( n22101 & ~n22102 ) ;
  assign n22104 = n22069 ^ x628 ^ 1'b0 ;
  assign n22105 = ( n22069 & n22103 ) | ( n22069 & ~n22104 ) | ( n22103 & ~n22104 ) ;
  assign n22106 = ( n22069 & n22103 ) | ( n22069 & n22104 ) | ( n22103 & n22104 ) ;
  assign n22107 = n22105 ^ x1156 ^ 1'b0 ;
  assign n22108 = ( n22105 & n22106 ) | ( n22105 & n22107 ) | ( n22106 & n22107 ) ;
  assign n22109 = n22103 ^ x792 ^ 1'b0 ;
  assign n22110 = ( n22103 & n22108 ) | ( n22103 & n22109 ) | ( n22108 & n22109 ) ;
  assign n22111 = n22069 ^ x647 ^ 1'b0 ;
  assign n22112 = ( n22069 & n22110 ) | ( n22069 & ~n22111 ) | ( n22110 & ~n22111 ) ;
  assign n22113 = ( n22069 & n22110 ) | ( n22069 & n22111 ) | ( n22110 & n22111 ) ;
  assign n22114 = n22112 ^ x1157 ^ 1'b0 ;
  assign n22115 = ( n22112 & n22113 ) | ( n22112 & n22114 ) | ( n22113 & n22114 ) ;
  assign n22116 = n22110 ^ x787 ^ 1'b0 ;
  assign n22117 = ( n22110 & n22115 ) | ( n22110 & n22116 ) | ( n22115 & n22116 ) ;
  assign n22118 = x644 & ~n22117 ;
  assign n22119 = x715 | n22118 ;
  assign n22120 = x644 & ~n22069 ;
  assign n22121 = x715 & ~n22120 ;
  assign n22122 = n22121 ^ x1160 ^ 1'b0 ;
  assign n22123 = x175 & n2069 ;
  assign n22124 = x38 & n22070 ;
  assign n22125 = ~x175 & x766 ;
  assign n22126 = n15587 & n22125 ;
  assign n22127 = x766 & n15639 ;
  assign n22128 = x175 & ~n22127 ;
  assign n22129 = ( n19902 & ~n22126 ) | ( n19902 & n22128 ) | ( ~n22126 & n22128 ) ;
  assign n22130 = n22126 | n22129 ;
  assign n22131 = x175 & ~n15631 ;
  assign n22132 = ~x766 & n15486 ;
  assign n22133 = ( x39 & n22131 ) | ( x39 & n22132 ) | ( n22131 & n22132 ) ;
  assign n22134 = n22132 ^ n22131 ^ 1'b0 ;
  assign n22135 = ( x39 & n22133 ) | ( x39 & n22134 ) | ( n22133 & n22134 ) ;
  assign n22136 = ( ~x38 & n22130 ) | ( ~x38 & n22135 ) | ( n22130 & n22135 ) ;
  assign n22137 = ~x38 & n22136 ;
  assign n22138 = x766 & n15646 ;
  assign n22139 = ~n22137 & n22138 ;
  assign n22140 = ( n22124 & n22137 ) | ( n22124 & ~n22139 ) | ( n22137 & ~n22139 ) ;
  assign n22141 = ~n2069 & n22140 ;
  assign n22142 = n22123 | n22141 ;
  assign n22143 = n22069 ^ n15659 ^ 1'b0 ;
  assign n22144 = ( n22069 & n22142 ) | ( n22069 & ~n22143 ) | ( n22142 & ~n22143 ) ;
  assign n22145 = n15662 & n22069 ;
  assign n22146 = ( ~n15662 & n22123 ) | ( ~n15662 & n22141 ) | ( n22123 & n22141 ) ;
  assign n22147 = n22145 | n22146 ;
  assign n22148 = n22147 ^ n22144 ^ n22069 ;
  assign n22149 = n22148 ^ x1155 ^ 1'b0 ;
  assign n22150 = ( n22147 & n22148 ) | ( n22147 & ~n22149 ) | ( n22148 & ~n22149 ) ;
  assign n22151 = n22144 ^ x785 ^ 1'b0 ;
  assign n22152 = ( n22144 & n22150 ) | ( n22144 & n22151 ) | ( n22150 & n22151 ) ;
  assign n22153 = x618 & ~n22152 ;
  assign n22154 = x618 | n22069 ;
  assign n22155 = ( x1154 & n22153 ) | ( x1154 & n22154 ) | ( n22153 & n22154 ) ;
  assign n22156 = ~n22153 & n22155 ;
  assign n22157 = x618 & ~n22069 ;
  assign n22158 = x1154 | n22157 ;
  assign n22159 = ( n22152 & n22153 ) | ( n22152 & ~n22158 ) | ( n22153 & ~n22158 ) ;
  assign n22160 = n22156 | n22159 ;
  assign n22161 = n22152 ^ x781 ^ 1'b0 ;
  assign n22162 = ( n22152 & n22160 ) | ( n22152 & n22161 ) | ( n22160 & n22161 ) ;
  assign n22163 = x619 | n22069 ;
  assign n22164 = x619 & ~n22162 ;
  assign n22165 = x1159 & ~n22164 ;
  assign n22166 = n22163 & n22165 ;
  assign n22167 = x619 & ~n22069 ;
  assign n22168 = x1159 | n22167 ;
  assign n22169 = ( n22162 & n22164 ) | ( n22162 & ~n22168 ) | ( n22164 & ~n22168 ) ;
  assign n22170 = n22166 | n22169 ;
  assign n22171 = n22162 ^ x789 ^ 1'b0 ;
  assign n22172 = ( n22162 & n22170 ) | ( n22162 & n22171 ) | ( n22170 & n22171 ) ;
  assign n22173 = n22069 ^ n16518 ^ 1'b0 ;
  assign n22174 = ( n22069 & n22172 ) | ( n22069 & ~n22173 ) | ( n22172 & ~n22173 ) ;
  assign n22175 = n22069 ^ n16339 ^ 1'b0 ;
  assign n22176 = ( n22069 & n22174 ) | ( n22069 & ~n22175 ) | ( n22174 & ~n22175 ) ;
  assign n22177 = n22069 ^ n16376 ^ 1'b0 ;
  assign n22178 = ( n22069 & n22176 ) | ( n22069 & ~n22177 ) | ( n22176 & ~n22177 ) ;
  assign n22179 = x644 | n22178 ;
  assign n22180 = ( n22121 & ~n22122 ) | ( n22121 & n22179 ) | ( ~n22122 & n22179 ) ;
  assign n22181 = ( x1160 & n22122 ) | ( x1160 & n22180 ) | ( n22122 & n22180 ) ;
  assign n22182 = n22119 & ~n22181 ;
  assign n22183 = x644 & ~n22178 ;
  assign n22184 = ( ~x715 & n22069 ) | ( ~x715 & n22120 ) | ( n22069 & n22120 ) ;
  assign n22185 = x1160 & ~n22184 ;
  assign n22186 = ( x1160 & n22183 ) | ( x1160 & n22185 ) | ( n22183 & n22185 ) ;
  assign n22187 = ( x715 & n22117 ) | ( x715 & n22118 ) | ( n22117 & n22118 ) ;
  assign n22188 = n22186 & ~n22187 ;
  assign n22189 = ( x790 & n22182 ) | ( x790 & n22188 ) | ( n22182 & n22188 ) ;
  assign n22190 = n22188 ^ n22182 ^ 1'b0 ;
  assign n22191 = ( x790 & n22189 ) | ( x790 & n22190 ) | ( n22189 & n22190 ) ;
  assign n22192 = n16374 & n22112 ;
  assign n22193 = n19055 & n22176 ;
  assign n22194 = n22192 | n22193 ;
  assign n22195 = n16373 & n22113 ;
  assign n22196 = ( x787 & n22194 ) | ( x787 & n22195 ) | ( n22194 & n22195 ) ;
  assign n22197 = n22195 ^ n22194 ^ 1'b0 ;
  assign n22198 = ( x787 & n22196 ) | ( x787 & n22197 ) | ( n22196 & n22197 ) ;
  assign n22199 = x619 & ~n22099 ;
  assign n22200 = x1159 | n22199 ;
  assign n22249 = x625 | n22142 ;
  assign n22202 = x700 | n22140 ;
  assign n22203 = x766 & n15591 ;
  assign n22204 = n17156 | n22203 ;
  assign n22205 = x175 & ~n5017 ;
  assign n22206 = n22204 & n22205 ;
  assign n22207 = n15340 & n15690 ;
  assign n22208 = ~x766 & n22207 ;
  assign n22209 = n15968 | n22208 ;
  assign n22210 = x39 | n22209 ;
  assign n22211 = ( ~x39 & x175 ) | ( ~x39 & n22210 ) | ( x175 & n22210 ) ;
  assign n22212 = ( x38 & n22206 ) | ( x38 & n22211 ) | ( n22206 & n22211 ) ;
  assign n22213 = ~n22206 & n22212 ;
  assign n22214 = x175 & n15795 ;
  assign n22215 = x766 | n22214 ;
  assign n22216 = ( x175 & n15876 ) | ( x175 & ~n22215 ) | ( n15876 & ~n22215 ) ;
  assign n22217 = ~n22215 & n22216 ;
  assign n22218 = x175 | n16003 ;
  assign n22219 = x175 & n15943 ;
  assign n22220 = x766 & ~n22219 ;
  assign n22221 = n22218 & n22220 ;
  assign n22222 = ( x39 & n22217 ) | ( x39 & ~n22221 ) | ( n22217 & ~n22221 ) ;
  assign n22223 = ~n22217 & n22222 ;
  assign n22224 = x175 & n16054 ;
  assign n22225 = x175 | n16048 ;
  assign n22226 = ( x766 & n22224 ) | ( x766 & n22225 ) | ( n22224 & n22225 ) ;
  assign n22227 = ~n22224 & n22226 ;
  assign n22228 = x175 | n16044 ;
  assign n22229 = x175 & n16029 ;
  assign n22230 = ( x766 & n22228 ) | ( x766 & ~n22229 ) | ( n22228 & ~n22229 ) ;
  assign n22231 = ~x766 & n22230 ;
  assign n22232 = ( x39 & ~n22227 ) | ( x39 & n22231 ) | ( ~n22227 & n22231 ) ;
  assign n22233 = n22227 | n22232 ;
  assign n22234 = ( x38 & ~n22223 ) | ( x38 & n22233 ) | ( ~n22223 & n22233 ) ;
  assign n22235 = ~x38 & n22234 ;
  assign n22236 = ( x700 & n22213 ) | ( x700 & ~n22235 ) | ( n22213 & ~n22235 ) ;
  assign n22237 = ~n22213 & n22236 ;
  assign n22238 = ( n2051 & n2068 ) | ( n2051 & ~n22237 ) | ( n2068 & ~n22237 ) ;
  assign n22239 = n22237 | n22238 ;
  assign n22240 = ( n22123 & n22202 ) | ( n22123 & ~n22239 ) | ( n22202 & ~n22239 ) ;
  assign n22241 = n22240 ^ n22202 ^ 1'b0 ;
  assign n22242 = ( n22123 & n22240 ) | ( n22123 & ~n22241 ) | ( n22240 & ~n22241 ) ;
  assign n22250 = x625 & ~n22242 ;
  assign n22251 = x1153 & ~n22250 ;
  assign n22252 = n22249 & n22251 ;
  assign n22253 = ( x608 & n22092 ) | ( x608 & ~n22252 ) | ( n22092 & ~n22252 ) ;
  assign n22254 = ~n22092 & n22253 ;
  assign n22243 = x625 | n22242 ;
  assign n22244 = x625 & ~n22142 ;
  assign n22245 = ( x1153 & n22243 ) | ( x1153 & ~n22244 ) | ( n22243 & ~n22244 ) ;
  assign n22246 = ~x1153 & n22245 ;
  assign n22247 = ( x608 & n22088 ) | ( x608 & ~n22246 ) | ( n22088 & ~n22246 ) ;
  assign n22248 = n22246 | n22247 ;
  assign n22255 = n22254 ^ n22248 ^ 1'b0 ;
  assign n22256 = ( x778 & ~n22248 ) | ( x778 & n22254 ) | ( ~n22248 & n22254 ) ;
  assign n22257 = ( x778 & ~n22255 ) | ( x778 & n22256 ) | ( ~n22255 & n22256 ) ;
  assign n22258 = ( x778 & n22242 ) | ( x778 & ~n22257 ) | ( n22242 & ~n22257 ) ;
  assign n22259 = ~n22257 & n22258 ;
  assign n22260 = x609 & ~n22259 ;
  assign n22266 = x609 | n22095 ;
  assign n22267 = ( x1155 & n22260 ) | ( x1155 & n22266 ) | ( n22260 & n22266 ) ;
  assign n22268 = ~n22260 & n22267 ;
  assign n22269 = ~x1155 & n22147 ;
  assign n22270 = ( x660 & n22268 ) | ( x660 & ~n22269 ) | ( n22268 & ~n22269 ) ;
  assign n22271 = ~n22268 & n22270 ;
  assign n22201 = x1155 & n22148 ;
  assign n22261 = x609 & ~n22095 ;
  assign n22262 = x1155 | n22261 ;
  assign n22263 = ( n22259 & n22260 ) | ( n22259 & ~n22262 ) | ( n22260 & ~n22262 ) ;
  assign n22264 = ( x660 & ~n22201 ) | ( x660 & n22263 ) | ( ~n22201 & n22263 ) ;
  assign n22265 = n22201 | n22264 ;
  assign n22272 = n22271 ^ n22265 ^ 1'b0 ;
  assign n22273 = ( x785 & ~n22265 ) | ( x785 & n22271 ) | ( ~n22265 & n22271 ) ;
  assign n22274 = ( x785 & ~n22272 ) | ( x785 & n22273 ) | ( ~n22272 & n22273 ) ;
  assign n22275 = ( x785 & n22259 ) | ( x785 & ~n22274 ) | ( n22259 & ~n22274 ) ;
  assign n22276 = ~n22274 & n22275 ;
  assign n22277 = x618 & ~n22276 ;
  assign n22283 = x618 | n22097 ;
  assign n22284 = ( x1154 & n22277 ) | ( x1154 & n22283 ) | ( n22277 & n22283 ) ;
  assign n22285 = ~n22277 & n22284 ;
  assign n22286 = ( x627 & n22159 ) | ( x627 & ~n22285 ) | ( n22159 & ~n22285 ) ;
  assign n22287 = ~n22159 & n22286 ;
  assign n22278 = x618 & ~n22097 ;
  assign n22279 = x1154 | n22278 ;
  assign n22280 = ( n22276 & n22277 ) | ( n22276 & ~n22279 ) | ( n22277 & ~n22279 ) ;
  assign n22281 = ( x627 & n22156 ) | ( x627 & ~n22280 ) | ( n22156 & ~n22280 ) ;
  assign n22282 = n22280 | n22281 ;
  assign n22288 = n22287 ^ n22282 ^ 1'b0 ;
  assign n22289 = ( x781 & ~n22282 ) | ( x781 & n22287 ) | ( ~n22282 & n22287 ) ;
  assign n22290 = ( x781 & ~n22288 ) | ( x781 & n22289 ) | ( ~n22288 & n22289 ) ;
  assign n22291 = ( x781 & n22276 ) | ( x781 & ~n22290 ) | ( n22276 & ~n22290 ) ;
  assign n22292 = ~n22290 & n22291 ;
  assign n22293 = x619 & ~n22292 ;
  assign n22294 = ( ~n22200 & n22292 ) | ( ~n22200 & n22293 ) | ( n22292 & n22293 ) ;
  assign n22295 = ( x648 & n22166 ) | ( x648 & ~n22294 ) | ( n22166 & ~n22294 ) ;
  assign n22296 = n22294 | n22295 ;
  assign n22297 = x619 | n22099 ;
  assign n22298 = x1159 & ~n22293 ;
  assign n22299 = n22297 & n22298 ;
  assign n22300 = ( x648 & n22169 ) | ( x648 & ~n22299 ) | ( n22169 & ~n22299 ) ;
  assign n22301 = ~n22169 & n22300 ;
  assign n22302 = x789 & ~n22301 ;
  assign n22303 = n22296 & n22302 ;
  assign n22304 = ~x789 & n22292 ;
  assign n22305 = ( n16519 & ~n22303 ) | ( n16519 & n22304 ) | ( ~n22303 & n22304 ) ;
  assign n22306 = n22303 | n22305 ;
  assign n22307 = n16337 & n22106 ;
  assign n22308 = n16338 & n22105 ;
  assign n22309 = n22307 | n22308 ;
  assign n22310 = n19046 & n22174 ;
  assign n22311 = ( x792 & n22309 ) | ( x792 & n22310 ) | ( n22309 & n22310 ) ;
  assign n22312 = n22310 ^ n22309 ^ 1'b0 ;
  assign n22313 = ( x792 & n22311 ) | ( x792 & n22312 ) | ( n22311 & n22312 ) ;
  assign n22314 = n18482 ^ x788 ^ 1'b0 ;
  assign n22315 = n16459 & ~n22101 ;
  assign n22316 = ~x626 & n22069 ;
  assign n22317 = ~x641 & x1158 ;
  assign n22318 = x626 & n22172 ;
  assign n22319 = ( n22316 & n22317 ) | ( n22316 & ~n22318 ) | ( n22317 & ~n22318 ) ;
  assign n22320 = ~n22316 & n22319 ;
  assign n22321 = ~x626 & n22172 ;
  assign n22322 = x641 & ~x1158 ;
  assign n22323 = x626 & n22069 ;
  assign n22324 = ( n22321 & n22322 ) | ( n22321 & ~n22323 ) | ( n22322 & ~n22323 ) ;
  assign n22325 = ~n22321 & n22324 ;
  assign n22326 = ( ~n22315 & n22320 ) | ( ~n22315 & n22325 ) | ( n22320 & n22325 ) ;
  assign n22327 = n22315 | n22326 ;
  assign n22328 = ( x788 & ~n22314 ) | ( x788 & n22327 ) | ( ~n22314 & n22327 ) ;
  assign n22329 = ( n18482 & n22314 ) | ( n18482 & n22328 ) | ( n22314 & n22328 ) ;
  assign n22330 = ~n22313 & n22329 ;
  assign n22331 = ( n22306 & n22313 ) | ( n22306 & ~n22330 ) | ( n22313 & ~n22330 ) ;
  assign n22332 = ( ~n18484 & n22198 ) | ( ~n18484 & n22331 ) | ( n22198 & n22331 ) ;
  assign n22333 = n22198 ^ n18484 ^ 1'b0 ;
  assign n22334 = ( n22198 & n22332 ) | ( n22198 & ~n22333 ) | ( n22332 & ~n22333 ) ;
  assign n22335 = x644 | n22181 ;
  assign n22336 = x644 & n22186 ;
  assign n22337 = x790 & ~n22336 ;
  assign n22338 = n22335 & n22337 ;
  assign n22339 = ( ~n22191 & n22334 ) | ( ~n22191 & n22338 ) | ( n22334 & n22338 ) ;
  assign n22340 = ~n22191 & n22339 ;
  assign n22341 = ( x57 & n5193 ) | ( x57 & ~n22340 ) | ( n5193 & ~n22340 ) ;
  assign n22342 = n22340 | n22341 ;
  assign n22343 = x175 | n1611 ;
  assign n22344 = ~n22203 & n22343 ;
  assign n22345 = n16397 | n22344 ;
  assign n22346 = ~n15662 & n22203 ;
  assign n22347 = ~x1155 & n22343 ;
  assign n22348 = ~n22346 & n22347 ;
  assign n22349 = ( x1155 & n22345 ) | ( x1155 & n22346 ) | ( n22345 & n22346 ) ;
  assign n22350 = n22348 | n22349 ;
  assign n22351 = n22345 ^ x785 ^ 1'b0 ;
  assign n22352 = ( n22345 & n22350 ) | ( n22345 & n22351 ) | ( n22350 & n22351 ) ;
  assign n22353 = n16411 | n22352 ;
  assign n22354 = x1154 & n22353 ;
  assign n22355 = n16414 | n22352 ;
  assign n22356 = ~x1154 & n22355 ;
  assign n22357 = n22354 | n22356 ;
  assign n22358 = n22352 ^ x781 ^ 1'b0 ;
  assign n22359 = ( n22352 & n22357 ) | ( n22352 & n22358 ) | ( n22357 & n22358 ) ;
  assign n22360 = n21437 | n22359 ;
  assign n22361 = x1159 & n22360 ;
  assign n22362 = n21440 | n22359 ;
  assign n22363 = ~x1159 & n22362 ;
  assign n22364 = n22361 | n22363 ;
  assign n22365 = n22359 ^ x789 ^ 1'b0 ;
  assign n22366 = ( n22359 & n22364 ) | ( n22359 & n22365 ) | ( n22364 & n22365 ) ;
  assign n22367 = n22343 ^ n16518 ^ 1'b0 ;
  assign n22368 = ( n22343 & n22366 ) | ( n22343 & ~n22367 ) | ( n22366 & ~n22367 ) ;
  assign n22369 = n22343 ^ n16339 ^ 1'b0 ;
  assign n22370 = ( n22343 & n22368 ) | ( n22343 & ~n22369 ) | ( n22368 & ~n22369 ) ;
  assign n22371 = n19055 & n22370 ;
  assign n22372 = x647 & ~n22343 ;
  assign n22373 = x1157 | n22372 ;
  assign n22374 = x700 & n15778 ;
  assign n22375 = ~x625 & n22374 ;
  assign n22376 = ~x1153 & n22343 ;
  assign n22377 = ~n22375 & n22376 ;
  assign n22378 = x778 & ~n22377 ;
  assign n22379 = n22343 & ~n22374 ;
  assign n22380 = ( x1153 & n22375 ) | ( x1153 & n22379 ) | ( n22375 & n22379 ) ;
  assign n22381 = n22378 & ~n22380 ;
  assign n22382 = ( x778 & n22379 ) | ( x778 & ~n22381 ) | ( n22379 & ~n22381 ) ;
  assign n22383 = ~n22381 & n22382 ;
  assign n22384 = n16447 | n22383 ;
  assign n22385 = n16449 | n22384 ;
  assign n22386 = n16451 | n22385 ;
  assign n22387 = n16530 | n22386 ;
  assign n22388 = n16560 | n22387 ;
  assign n22389 = ( x647 & ~n22373 ) | ( x647 & n22388 ) | ( ~n22373 & n22388 ) ;
  assign n22390 = ~n22373 & n22389 ;
  assign n22391 = n22343 ^ x647 ^ 1'b0 ;
  assign n22392 = ( n22343 & n22388 ) | ( n22343 & n22391 ) | ( n22388 & n22391 ) ;
  assign n22393 = x1157 & n22392 ;
  assign n22394 = ( n16375 & n22390 ) | ( n16375 & n22393 ) | ( n22390 & n22393 ) ;
  assign n22395 = ( x787 & n22371 ) | ( x787 & n22394 ) | ( n22371 & n22394 ) ;
  assign n22396 = n22394 ^ n22371 ^ 1'b0 ;
  assign n22397 = ( x787 & n22395 ) | ( x787 & n22396 ) | ( n22395 & n22396 ) ;
  assign n22398 = ~x626 & n22343 ;
  assign n22399 = x626 & n22366 ;
  assign n22400 = ( n22317 & n22398 ) | ( n22317 & ~n22399 ) | ( n22398 & ~n22399 ) ;
  assign n22401 = ~n22398 & n22400 ;
  assign n22402 = ~x626 & n22366 ;
  assign n22403 = x626 & n22343 ;
  assign n22404 = ( n22322 & n22402 ) | ( n22322 & ~n22403 ) | ( n22402 & ~n22403 ) ;
  assign n22405 = ~n22402 & n22404 ;
  assign n22406 = n22386 & ~n22405 ;
  assign n22407 = ( n16459 & n22405 ) | ( n16459 & ~n22406 ) | ( n22405 & ~n22406 ) ;
  assign n22408 = ( x788 & n22401 ) | ( x788 & n22407 ) | ( n22401 & n22407 ) ;
  assign n22409 = n22407 ^ n22401 ^ 1'b0 ;
  assign n22410 = ( x788 & n22408 ) | ( x788 & n22409 ) | ( n22408 & n22409 ) ;
  assign n22411 = n15524 | n22379 ;
  assign n22412 = n22344 & n22411 ;
  assign n22413 = x625 & ~n22411 ;
  assign n22414 = ( n22376 & n22412 ) | ( n22376 & n22413 ) | ( n22412 & n22413 ) ;
  assign n22415 = ( x608 & n22380 ) | ( x608 & ~n22414 ) | ( n22380 & ~n22414 ) ;
  assign n22416 = n22414 | n22415 ;
  assign n22417 = x1153 & n22344 ;
  assign n22418 = ~n22413 & n22417 ;
  assign n22419 = x608 & ~n22377 ;
  assign n22420 = n22416 & ~n22419 ;
  assign n22421 = ( n22416 & n22418 ) | ( n22416 & n22420 ) | ( n22418 & n22420 ) ;
  assign n22422 = n22412 ^ x778 ^ 1'b0 ;
  assign n22423 = ( n22412 & n22421 ) | ( n22412 & n22422 ) | ( n22421 & n22422 ) ;
  assign n22424 = x609 & ~n22423 ;
  assign n22430 = x609 | n22383 ;
  assign n22431 = ( x1155 & n22424 ) | ( x1155 & n22430 ) | ( n22424 & n22430 ) ;
  assign n22432 = ~n22424 & n22431 ;
  assign n22433 = ( x660 & n22348 ) | ( x660 & ~n22432 ) | ( n22348 & ~n22432 ) ;
  assign n22434 = ~n22348 & n22433 ;
  assign n22425 = x609 & ~n22383 ;
  assign n22426 = x1155 | n22425 ;
  assign n22427 = ( n22423 & n22424 ) | ( n22423 & ~n22426 ) | ( n22424 & ~n22426 ) ;
  assign n22428 = ( x660 & n22349 ) | ( x660 & ~n22427 ) | ( n22349 & ~n22427 ) ;
  assign n22429 = n22427 | n22428 ;
  assign n22435 = n22434 ^ n22429 ^ 1'b0 ;
  assign n22436 = ( x785 & ~n22429 ) | ( x785 & n22434 ) | ( ~n22429 & n22434 ) ;
  assign n22437 = ( x785 & ~n22435 ) | ( x785 & n22436 ) | ( ~n22435 & n22436 ) ;
  assign n22438 = ( x785 & n22423 ) | ( x785 & ~n22437 ) | ( n22423 & ~n22437 ) ;
  assign n22439 = ~n22437 & n22438 ;
  assign n22440 = x618 & ~n22439 ;
  assign n22441 = x618 | n22384 ;
  assign n22442 = ( x1154 & n22440 ) | ( x1154 & n22441 ) | ( n22440 & n22441 ) ;
  assign n22443 = ~n22440 & n22442 ;
  assign n22444 = ( x627 & n22356 ) | ( x627 & ~n22443 ) | ( n22356 & ~n22443 ) ;
  assign n22445 = ~n22356 & n22444 ;
  assign n22446 = x627 | n22354 ;
  assign n22447 = x618 & ~n22384 ;
  assign n22448 = x1154 | n22447 ;
  assign n22449 = ( n22439 & n22440 ) | ( n22439 & ~n22448 ) | ( n22440 & ~n22448 ) ;
  assign n22450 = ( ~n22445 & n22446 ) | ( ~n22445 & n22449 ) | ( n22446 & n22449 ) ;
  assign n22451 = ~n22445 & n22450 ;
  assign n22452 = n22439 ^ x781 ^ 1'b0 ;
  assign n22453 = ( n22439 & n22451 ) | ( n22439 & n22452 ) | ( n22451 & n22452 ) ;
  assign n22454 = ~x789 & n22453 ;
  assign n22455 = x619 & ~n22385 ;
  assign n22456 = x1159 | n22455 ;
  assign n22457 = x619 & ~n22453 ;
  assign n22458 = ( n22453 & ~n22456 ) | ( n22453 & n22457 ) | ( ~n22456 & n22457 ) ;
  assign n22459 = ( x648 & n22361 ) | ( x648 & ~n22458 ) | ( n22361 & ~n22458 ) ;
  assign n22460 = n22458 | n22459 ;
  assign n22461 = x619 | n22385 ;
  assign n22462 = x1159 & ~n22457 ;
  assign n22463 = n22461 & n22462 ;
  assign n22464 = ( x648 & n22363 ) | ( x648 & ~n22463 ) | ( n22363 & ~n22463 ) ;
  assign n22465 = ~n22363 & n22464 ;
  assign n22466 = x789 & ~n22465 ;
  assign n22467 = n22460 & n22466 ;
  assign n22468 = ( n16519 & ~n22454 ) | ( n16519 & n22467 ) | ( ~n22454 & n22467 ) ;
  assign n22469 = n22454 | n22468 ;
  assign n22470 = n22469 ^ n22410 ^ 1'b0 ;
  assign n22471 = ( n22410 & n22469 ) | ( n22410 & n22470 ) | ( n22469 & n22470 ) ;
  assign n22472 = ( n18482 & ~n22410 ) | ( n18482 & n22471 ) | ( ~n22410 & n22471 ) ;
  assign n22473 = n19208 | n22387 ;
  assign n22474 = n16556 & ~n22368 ;
  assign n22475 = x629 & ~n22474 ;
  assign n22476 = n22473 & n22475 ;
  assign n22477 = n16557 & ~n22368 ;
  assign n22478 = n19212 & ~n22387 ;
  assign n22479 = n22477 | n22478 ;
  assign n22480 = ( x629 & ~n22476 ) | ( x629 & n22479 ) | ( ~n22476 & n22479 ) ;
  assign n22481 = ~n22476 & n22480 ;
  assign n22482 = ( x792 & ~n19206 ) | ( x792 & n22481 ) | ( ~n19206 & n22481 ) ;
  assign n22483 = ( n18484 & n19206 ) | ( n18484 & n22482 ) | ( n19206 & n22482 ) ;
  assign n22484 = ( n22397 & n22472 ) | ( n22397 & ~n22483 ) | ( n22472 & ~n22483 ) ;
  assign n22485 = n22484 ^ n22472 ^ 1'b0 ;
  assign n22486 = ( n22397 & n22484 ) | ( n22397 & ~n22485 ) | ( n22484 & ~n22485 ) ;
  assign n22487 = x790 | n22486 ;
  assign n22488 = x644 & ~n22486 ;
  assign n22489 = ( x787 & n22390 ) | ( x787 & ~n22393 ) | ( n22390 & ~n22393 ) ;
  assign n22490 = ~n22390 & n22489 ;
  assign n22491 = ( x787 & n22388 ) | ( x787 & ~n22490 ) | ( n22388 & ~n22490 ) ;
  assign n22492 = ~n22490 & n22491 ;
  assign n22493 = x644 | n22492 ;
  assign n22494 = ( x715 & n22488 ) | ( x715 & n22493 ) | ( n22488 & n22493 ) ;
  assign n22495 = ~n22488 & n22494 ;
  assign n22496 = x644 | n22343 ;
  assign n22497 = n22343 ^ n16376 ^ 1'b0 ;
  assign n22498 = ( n22343 & n22370 ) | ( n22343 & ~n22497 ) | ( n22370 & ~n22497 ) ;
  assign n22499 = x644 & ~n22498 ;
  assign n22500 = ( x715 & n22496 ) | ( x715 & ~n22499 ) | ( n22496 & ~n22499 ) ;
  assign n22501 = ~x715 & n22500 ;
  assign n22502 = ( x1160 & n22495 ) | ( x1160 & ~n22501 ) | ( n22495 & ~n22501 ) ;
  assign n22503 = ~n22495 & n22502 ;
  assign n22504 = x644 & ~n22343 ;
  assign n22505 = x715 & ~n22504 ;
  assign n22506 = ( n22498 & n22499 ) | ( n22498 & n22505 ) | ( n22499 & n22505 ) ;
  assign n22507 = x644 & ~n22492 ;
  assign n22508 = x715 | n22507 ;
  assign n22509 = ( n22486 & n22488 ) | ( n22486 & ~n22508 ) | ( n22488 & ~n22508 ) ;
  assign n22510 = ( x1160 & ~n22506 ) | ( x1160 & n22509 ) | ( ~n22506 & n22509 ) ;
  assign n22511 = n22506 | n22510 ;
  assign n22512 = x790 & ~n22511 ;
  assign n22513 = ( x790 & n22503 ) | ( x790 & n22512 ) | ( n22503 & n22512 ) ;
  assign n22514 = x832 & ~n22513 ;
  assign n22515 = n22487 & n22514 ;
  assign n22516 = ~x175 & n7318 ;
  assign n22517 = x832 | n22516 ;
  assign n22518 = ~n22515 & n22517 ;
  assign n22519 = ( n22342 & n22515 ) | ( n22342 & ~n22518 ) | ( n22515 & ~n22518 ) ;
  assign n22520 = x176 | n15656 ;
  assign n22521 = x38 | n16697 ;
  assign n22522 = ~n18524 & n22521 ;
  assign n22523 = ~x176 & n22522 ;
  assign n22524 = x704 | n22523 ;
  assign n22525 = x176 | n15655 ;
  assign n22526 = x704 & ~n22525 ;
  assign n22527 = ( n2069 & n22524 ) | ( n2069 & ~n22526 ) | ( n22524 & ~n22526 ) ;
  assign n22528 = ~n2069 & n22527 ;
  assign n22529 = n2069 | n16185 ;
  assign n22530 = n16700 & ~n22529 ;
  assign n22531 = ~n22528 & n22530 ;
  assign n22532 = ( x176 & n22528 ) | ( x176 & ~n22531 ) | ( n22528 & ~n22531 ) ;
  assign n22533 = x625 & ~n22532 ;
  assign n22534 = x625 | n22520 ;
  assign n22535 = ( x1153 & n22533 ) | ( x1153 & n22534 ) | ( n22533 & n22534 ) ;
  assign n22536 = ~n22533 & n22535 ;
  assign n22537 = x625 & ~n22520 ;
  assign n22538 = x1153 | n22537 ;
  assign n22539 = ( x625 & n22532 ) | ( x625 & ~n22538 ) | ( n22532 & ~n22538 ) ;
  assign n22540 = ~n22538 & n22539 ;
  assign n22541 = n22536 | n22540 ;
  assign n22542 = n22532 ^ x778 ^ 1'b0 ;
  assign n22543 = ( n22532 & n22541 ) | ( n22532 & n22542 ) | ( n22541 & n22542 ) ;
  assign n22544 = n22520 ^ n16234 ^ 1'b0 ;
  assign n22545 = ( n22520 & n22543 ) | ( n22520 & ~n22544 ) | ( n22543 & ~n22544 ) ;
  assign n22546 = n22520 ^ n16254 ^ 1'b0 ;
  assign n22547 = ( n22520 & n22545 ) | ( n22520 & ~n22546 ) | ( n22545 & ~n22546 ) ;
  assign n22548 = n22520 ^ n16279 ^ 1'b0 ;
  assign n22549 = ( n22520 & n22547 ) | ( n22520 & ~n22548 ) | ( n22547 & ~n22548 ) ;
  assign n22550 = n22520 ^ n16318 ^ 1'b0 ;
  assign n22551 = ( n22520 & n22549 ) | ( n22520 & ~n22550 ) | ( n22549 & ~n22550 ) ;
  assign n22552 = n22520 ^ x628 ^ 1'b0 ;
  assign n22553 = ( n22520 & n22551 ) | ( n22520 & ~n22552 ) | ( n22551 & ~n22552 ) ;
  assign n22554 = ( n22520 & n22551 ) | ( n22520 & n22552 ) | ( n22551 & n22552 ) ;
  assign n22555 = n22553 ^ x1156 ^ 1'b0 ;
  assign n22556 = ( n22553 & n22554 ) | ( n22553 & n22555 ) | ( n22554 & n22555 ) ;
  assign n22557 = n22551 ^ x792 ^ 1'b0 ;
  assign n22558 = ( n22551 & n22556 ) | ( n22551 & n22557 ) | ( n22556 & n22557 ) ;
  assign n22559 = n22520 ^ x647 ^ 1'b0 ;
  assign n22560 = ( n22520 & n22558 ) | ( n22520 & ~n22559 ) | ( n22558 & ~n22559 ) ;
  assign n22561 = ( n22520 & n22558 ) | ( n22520 & n22559 ) | ( n22558 & n22559 ) ;
  assign n22562 = n22560 ^ x1157 ^ 1'b0 ;
  assign n22563 = ( n22560 & n22561 ) | ( n22560 & n22562 ) | ( n22561 & n22562 ) ;
  assign n22564 = n22558 ^ x787 ^ 1'b0 ;
  assign n22565 = ( n22558 & n22563 ) | ( n22558 & n22564 ) | ( n22563 & n22564 ) ;
  assign n22566 = x644 & ~n22565 ;
  assign n22567 = x715 | n22566 ;
  assign n22568 = x644 & ~n22520 ;
  assign n22569 = x715 & ~n22568 ;
  assign n22570 = n22569 ^ x1160 ^ 1'b0 ;
  assign n22571 = n15640 ^ x38 ^ 1'b0 ;
  assign n22572 = ( n15640 & n17838 ) | ( n15640 & n22571 ) | ( n17838 & n22571 ) ;
  assign n22573 = n17843 ^ x176 ^ 1'b0 ;
  assign n22574 = ( n17843 & ~n22572 ) | ( n17843 & n22573 ) | ( ~n22572 & n22573 ) ;
  assign n22575 = n22525 ^ x742 ^ 1'b0 ;
  assign n22576 = ( n22525 & n22574 ) | ( n22525 & ~n22575 ) | ( n22574 & ~n22575 ) ;
  assign n22577 = n22576 ^ n2069 ^ 1'b0 ;
  assign n22578 = ( x176 & n22576 ) | ( x176 & n22577 ) | ( n22576 & n22577 ) ;
  assign n22579 = n22520 ^ n15659 ^ 1'b0 ;
  assign n22580 = ( n22520 & n22578 ) | ( n22520 & ~n22579 ) | ( n22578 & ~n22579 ) ;
  assign n22581 = ~n15659 & n22578 ;
  assign n22582 = x609 & n22581 ;
  assign n22583 = ~n15668 & n22520 ;
  assign n22584 = ( x1155 & n22582 ) | ( x1155 & n22583 ) | ( n22582 & n22583 ) ;
  assign n22585 = n22583 ^ n22582 ^ 1'b0 ;
  assign n22586 = ( x1155 & n22584 ) | ( x1155 & n22585 ) | ( n22584 & n22585 ) ;
  assign n22587 = ~x609 & n22581 ;
  assign n22588 = n15662 & n22520 ;
  assign n22589 = ( ~x1155 & n22587 ) | ( ~x1155 & n22588 ) | ( n22587 & n22588 ) ;
  assign n22590 = ~x1155 & n22589 ;
  assign n22591 = n22586 | n22590 ;
  assign n22592 = n22580 ^ x785 ^ 1'b0 ;
  assign n22593 = ( n22580 & n22591 ) | ( n22580 & n22592 ) | ( n22591 & n22592 ) ;
  assign n22594 = x618 & ~n22593 ;
  assign n22595 = x618 | n22520 ;
  assign n22596 = ( x1154 & n22594 ) | ( x1154 & n22595 ) | ( n22594 & n22595 ) ;
  assign n22597 = ~n22594 & n22596 ;
  assign n22598 = x618 & ~n22520 ;
  assign n22599 = x1154 | n22598 ;
  assign n22600 = ( n22593 & n22594 ) | ( n22593 & ~n22599 ) | ( n22594 & ~n22599 ) ;
  assign n22601 = n22597 | n22600 ;
  assign n22602 = n22593 ^ x781 ^ 1'b0 ;
  assign n22603 = ( n22593 & n22601 ) | ( n22593 & n22602 ) | ( n22601 & n22602 ) ;
  assign n22604 = x619 & ~n22603 ;
  assign n22605 = x619 | n22520 ;
  assign n22606 = ( x1159 & n22604 ) | ( x1159 & n22605 ) | ( n22604 & n22605 ) ;
  assign n22607 = ~n22604 & n22606 ;
  assign n22608 = x619 & ~n22520 ;
  assign n22609 = x1159 | n22608 ;
  assign n22610 = ( n22603 & n22604 ) | ( n22603 & ~n22609 ) | ( n22604 & ~n22609 ) ;
  assign n22611 = n22607 | n22610 ;
  assign n22612 = n22603 ^ x789 ^ 1'b0 ;
  assign n22613 = ( n22603 & n22611 ) | ( n22603 & n22612 ) | ( n22611 & n22612 ) ;
  assign n22614 = n22520 ^ n16518 ^ 1'b0 ;
  assign n22615 = ( n22520 & n22613 ) | ( n22520 & ~n22614 ) | ( n22613 & ~n22614 ) ;
  assign n22616 = n22520 ^ n16339 ^ 1'b0 ;
  assign n22617 = ( n22520 & n22615 ) | ( n22520 & ~n22616 ) | ( n22615 & ~n22616 ) ;
  assign n22618 = n22520 ^ n16376 ^ 1'b0 ;
  assign n22619 = ( n22520 & n22617 ) | ( n22520 & ~n22618 ) | ( n22617 & ~n22618 ) ;
  assign n22620 = x644 | n22619 ;
  assign n22621 = ( n22569 & ~n22570 ) | ( n22569 & n22620 ) | ( ~n22570 & n22620 ) ;
  assign n22622 = ( x1160 & n22570 ) | ( x1160 & n22621 ) | ( n22570 & n22621 ) ;
  assign n22623 = n22567 & ~n22622 ;
  assign n22624 = x644 & ~n22619 ;
  assign n22625 = ( ~x715 & n22520 ) | ( ~x715 & n22568 ) | ( n22520 & n22568 ) ;
  assign n22626 = x1160 & ~n22625 ;
  assign n22627 = ( x1160 & n22624 ) | ( x1160 & n22626 ) | ( n22624 & n22626 ) ;
  assign n22628 = ( x715 & n22565 ) | ( x715 & n22566 ) | ( n22565 & n22566 ) ;
  assign n22629 = n22627 & ~n22628 ;
  assign n22630 = ( x790 & n22623 ) | ( x790 & n22629 ) | ( n22623 & n22629 ) ;
  assign n22631 = n22629 ^ n22623 ^ 1'b0 ;
  assign n22632 = ( x790 & n22630 ) | ( x790 & n22631 ) | ( n22630 & n22631 ) ;
  assign n22633 = x626 & n22613 ;
  assign n22634 = ~x626 & n22520 ;
  assign n22635 = ( n22317 & n22633 ) | ( n22317 & ~n22634 ) | ( n22633 & ~n22634 ) ;
  assign n22636 = ~n22633 & n22635 ;
  assign n22637 = ~x626 & n22613 ;
  assign n22638 = x626 & n22520 ;
  assign n22639 = ( n22322 & n22637 ) | ( n22322 & ~n22638 ) | ( n22637 & ~n22638 ) ;
  assign n22640 = ~n22637 & n22639 ;
  assign n22641 = n22549 & ~n22640 ;
  assign n22642 = ( n16459 & n22640 ) | ( n16459 & ~n22641 ) | ( n22640 & ~n22641 ) ;
  assign n22643 = ( x788 & n22636 ) | ( x788 & n22642 ) | ( n22636 & n22642 ) ;
  assign n22644 = n22642 ^ n22636 ^ 1'b0 ;
  assign n22645 = ( x788 & n22643 ) | ( x788 & n22644 ) | ( n22643 & n22644 ) ;
  assign n22646 = x704 & ~n22576 ;
  assign n22647 = x176 | n17902 ;
  assign n22648 = x176 & n17910 ;
  assign n22649 = ( x742 & n22647 ) | ( x742 & ~n22648 ) | ( n22647 & ~n22648 ) ;
  assign n22650 = ~x742 & n22649 ;
  assign n22651 = n17886 ^ n16659 ^ x38 ;
  assign n22652 = x176 & n22651 ;
  assign n22653 = x176 | n17893 ;
  assign n22654 = ( x742 & n22652 ) | ( x742 & n22653 ) | ( n22652 & n22653 ) ;
  assign n22655 = ~n22652 & n22654 ;
  assign n22656 = ( x704 & ~n22650 ) | ( x704 & n22655 ) | ( ~n22650 & n22655 ) ;
  assign n22657 = n22650 | n22656 ;
  assign n22658 = ( n2069 & ~n22646 ) | ( n2069 & n22657 ) | ( ~n22646 & n22657 ) ;
  assign n22659 = ~n2069 & n22658 ;
  assign n22660 = n22659 ^ x176 ^ 1'b0 ;
  assign n22661 = ( ~x176 & n2069 ) | ( ~x176 & n22660 ) | ( n2069 & n22660 ) ;
  assign n22662 = ( x176 & n22659 ) | ( x176 & n22661 ) | ( n22659 & n22661 ) ;
  assign n22663 = x625 & ~n22662 ;
  assign n22664 = x625 | n22578 ;
  assign n22665 = ( x1153 & n22663 ) | ( x1153 & n22664 ) | ( n22663 & n22664 ) ;
  assign n22666 = ~n22663 & n22665 ;
  assign n22667 = ( x608 & n22540 ) | ( x608 & ~n22666 ) | ( n22540 & ~n22666 ) ;
  assign n22668 = ~n22540 & n22667 ;
  assign n22669 = x608 | n22536 ;
  assign n22670 = x625 & ~n22578 ;
  assign n22671 = x1153 | n22670 ;
  assign n22672 = ( n22662 & n22663 ) | ( n22662 & ~n22671 ) | ( n22663 & ~n22671 ) ;
  assign n22673 = ( ~n22668 & n22669 ) | ( ~n22668 & n22672 ) | ( n22669 & n22672 ) ;
  assign n22674 = ~n22668 & n22673 ;
  assign n22675 = n22662 ^ x778 ^ 1'b0 ;
  assign n22676 = ( n22662 & n22674 ) | ( n22662 & n22675 ) | ( n22674 & n22675 ) ;
  assign n22677 = x609 & ~n22676 ;
  assign n22678 = x609 | n22543 ;
  assign n22679 = ( x1155 & n22677 ) | ( x1155 & n22678 ) | ( n22677 & n22678 ) ;
  assign n22680 = ~n22677 & n22679 ;
  assign n22681 = ( x660 & n22590 ) | ( x660 & ~n22680 ) | ( n22590 & ~n22680 ) ;
  assign n22682 = ~n22590 & n22681 ;
  assign n22683 = x660 | n22586 ;
  assign n22684 = x609 & ~n22543 ;
  assign n22685 = x1155 | n22684 ;
  assign n22686 = ( n22676 & n22677 ) | ( n22676 & ~n22685 ) | ( n22677 & ~n22685 ) ;
  assign n22687 = ( ~n22682 & n22683 ) | ( ~n22682 & n22686 ) | ( n22683 & n22686 ) ;
  assign n22688 = ~n22682 & n22687 ;
  assign n22689 = n22676 ^ x785 ^ 1'b0 ;
  assign n22690 = ( n22676 & n22688 ) | ( n22676 & n22689 ) | ( n22688 & n22689 ) ;
  assign n22691 = x618 & ~n22690 ;
  assign n22692 = x618 | n22545 ;
  assign n22693 = ( x1154 & n22691 ) | ( x1154 & n22692 ) | ( n22691 & n22692 ) ;
  assign n22694 = ~n22691 & n22693 ;
  assign n22695 = ( x627 & n22600 ) | ( x627 & ~n22694 ) | ( n22600 & ~n22694 ) ;
  assign n22696 = ~n22600 & n22695 ;
  assign n22697 = x627 | n22597 ;
  assign n22698 = x618 & ~n22545 ;
  assign n22699 = x1154 | n22698 ;
  assign n22700 = ( n22690 & n22691 ) | ( n22690 & ~n22699 ) | ( n22691 & ~n22699 ) ;
  assign n22701 = ( ~n22696 & n22697 ) | ( ~n22696 & n22700 ) | ( n22697 & n22700 ) ;
  assign n22702 = ~n22696 & n22701 ;
  assign n22703 = n22690 ^ x781 ^ 1'b0 ;
  assign n22704 = ( n22690 & n22702 ) | ( n22690 & n22703 ) | ( n22702 & n22703 ) ;
  assign n22705 = ~x789 & n22704 ;
  assign n22706 = n16519 | n22705 ;
  assign n22707 = x619 | n22704 ;
  assign n22708 = x619 & ~n22547 ;
  assign n22709 = ( x1159 & n22707 ) | ( x1159 & ~n22708 ) | ( n22707 & ~n22708 ) ;
  assign n22710 = ~x1159 & n22709 ;
  assign n22711 = ( x648 & n22607 ) | ( x648 & ~n22710 ) | ( n22607 & ~n22710 ) ;
  assign n22712 = n22710 | n22711 ;
  assign n22713 = x619 & ~n22704 ;
  assign n22714 = x619 | n22547 ;
  assign n22715 = ( x1159 & n22713 ) | ( x1159 & n22714 ) | ( n22713 & n22714 ) ;
  assign n22716 = ~n22713 & n22715 ;
  assign n22717 = ( x648 & n22610 ) | ( x648 & ~n22716 ) | ( n22610 & ~n22716 ) ;
  assign n22718 = ~n22610 & n22717 ;
  assign n22719 = x789 & ~n22718 ;
  assign n22720 = n22712 & n22719 ;
  assign n22721 = ( ~n22645 & n22706 ) | ( ~n22645 & n22720 ) | ( n22706 & n22720 ) ;
  assign n22722 = ~n22645 & n22721 ;
  assign n22723 = n19046 & n22615 ;
  assign n22724 = n16337 & n22554 ;
  assign n22725 = n16338 & n22553 ;
  assign n22726 = ( ~n22723 & n22724 ) | ( ~n22723 & n22725 ) | ( n22724 & n22725 ) ;
  assign n22727 = n22723 | n22726 ;
  assign n22728 = n22722 ^ x792 ^ 1'b0 ;
  assign n22729 = ( ~x792 & n22727 ) | ( ~x792 & n22728 ) | ( n22727 & n22728 ) ;
  assign n22730 = ( x792 & n22722 ) | ( x792 & n22729 ) | ( n22722 & n22729 ) ;
  assign n22731 = n16374 & n22560 ;
  assign n22732 = n19055 & n22617 ;
  assign n22733 = n22731 | n22732 ;
  assign n22734 = n16373 & n22561 ;
  assign n22735 = ( x787 & n22733 ) | ( x787 & n22734 ) | ( n22733 & n22734 ) ;
  assign n22736 = n22734 ^ n22733 ^ 1'b0 ;
  assign n22737 = ( x787 & n22735 ) | ( x787 & n22736 ) | ( n22735 & n22736 ) ;
  assign n22738 = n18482 & ~n22727 ;
  assign n22739 = n18484 | n22738 ;
  assign n22740 = ~n22737 & n22739 ;
  assign n22741 = ( n22730 & n22737 ) | ( n22730 & ~n22740 ) | ( n22737 & ~n22740 ) ;
  assign n22742 = x644 | n22622 ;
  assign n22743 = x644 & n22627 ;
  assign n22744 = x790 & ~n22743 ;
  assign n22745 = n22742 & n22744 ;
  assign n22746 = ( ~n22632 & n22741 ) | ( ~n22632 & n22745 ) | ( n22741 & n22745 ) ;
  assign n22747 = ~n22632 & n22746 ;
  assign n22748 = ( x57 & n5193 ) | ( x57 & ~n22747 ) | ( n5193 & ~n22747 ) ;
  assign n22749 = n22747 | n22748 ;
  assign n22750 = x176 | n1611 ;
  assign n22751 = ~x742 & n15591 ;
  assign n22752 = n22750 & ~n22751 ;
  assign n22753 = n16397 | n22752 ;
  assign n22754 = n16402 | n22752 ;
  assign n22755 = x1155 & n22754 ;
  assign n22756 = n16405 | n22753 ;
  assign n22757 = ~x1155 & n22756 ;
  assign n22758 = n22755 | n22757 ;
  assign n22759 = n22753 ^ x785 ^ 1'b0 ;
  assign n22760 = ( n22753 & n22758 ) | ( n22753 & n22759 ) | ( n22758 & n22759 ) ;
  assign n22761 = n16411 | n22760 ;
  assign n22762 = x1154 & n22761 ;
  assign n22763 = n16414 | n22760 ;
  assign n22764 = ~x1154 & n22763 ;
  assign n22765 = n22762 | n22764 ;
  assign n22766 = n22760 ^ x781 ^ 1'b0 ;
  assign n22767 = ( n22760 & n22765 ) | ( n22760 & n22766 ) | ( n22765 & n22766 ) ;
  assign n22768 = x619 & ~n22767 ;
  assign n22769 = x619 | n22750 ;
  assign n22770 = ( x1159 & n22768 ) | ( x1159 & n22769 ) | ( n22768 & n22769 ) ;
  assign n22771 = ~n22768 & n22770 ;
  assign n22772 = x619 & ~n22750 ;
  assign n22773 = x1159 | n22772 ;
  assign n22774 = ( n22767 & n22768 ) | ( n22767 & ~n22773 ) | ( n22768 & ~n22773 ) ;
  assign n22775 = n22771 | n22774 ;
  assign n22776 = n22767 ^ x789 ^ 1'b0 ;
  assign n22777 = ( n22767 & n22775 ) | ( n22767 & n22776 ) | ( n22775 & n22776 ) ;
  assign n22778 = n22750 ^ n16518 ^ 1'b0 ;
  assign n22779 = ( n22750 & n22777 ) | ( n22750 & ~n22778 ) | ( n22777 & ~n22778 ) ;
  assign n22780 = n22750 ^ n16339 ^ 1'b0 ;
  assign n22781 = ( n22750 & n22779 ) | ( n22750 & ~n22780 ) | ( n22779 & ~n22780 ) ;
  assign n22782 = n19055 & n22781 ;
  assign n22783 = x647 & ~n22750 ;
  assign n22784 = x1157 | n22783 ;
  assign n22785 = ~x704 & n15778 ;
  assign n22786 = n22750 & ~n22785 ;
  assign n22787 = ~x1153 & n22750 ;
  assign n22788 = ~x625 & n22785 ;
  assign n22789 = n22787 & ~n22788 ;
  assign n22790 = ( x1153 & n22786 ) | ( x1153 & n22788 ) | ( n22786 & n22788 ) ;
  assign n22791 = n22789 | n22790 ;
  assign n22792 = n22786 ^ x778 ^ 1'b0 ;
  assign n22793 = ( n22786 & n22791 ) | ( n22786 & n22792 ) | ( n22791 & n22792 ) ;
  assign n22794 = n16447 | n22793 ;
  assign n22795 = n16449 | n22794 ;
  assign n22796 = n16451 | n22795 ;
  assign n22797 = n16530 | n22796 ;
  assign n22798 = n16560 | n22797 ;
  assign n22799 = ( x647 & ~n22784 ) | ( x647 & n22798 ) | ( ~n22784 & n22798 ) ;
  assign n22800 = ~n22784 & n22799 ;
  assign n22801 = n22750 ^ x647 ^ 1'b0 ;
  assign n22802 = ( n22750 & n22798 ) | ( n22750 & n22801 ) | ( n22798 & n22801 ) ;
  assign n22803 = x1157 & n22802 ;
  assign n22804 = ( n16375 & n22800 ) | ( n16375 & n22803 ) | ( n22800 & n22803 ) ;
  assign n22805 = ( x787 & n22782 ) | ( x787 & n22804 ) | ( n22782 & n22804 ) ;
  assign n22806 = n22804 ^ n22782 ^ 1'b0 ;
  assign n22807 = ( x787 & n22805 ) | ( x787 & n22806 ) | ( n22805 & n22806 ) ;
  assign n22808 = ~x626 & n22750 ;
  assign n22809 = x626 & n22777 ;
  assign n22810 = ( n22317 & n22808 ) | ( n22317 & ~n22809 ) | ( n22808 & ~n22809 ) ;
  assign n22811 = ~n22808 & n22810 ;
  assign n22812 = ~x626 & n22777 ;
  assign n22813 = x626 & n22750 ;
  assign n22814 = ( n22322 & n22812 ) | ( n22322 & ~n22813 ) | ( n22812 & ~n22813 ) ;
  assign n22815 = ~n22812 & n22814 ;
  assign n22816 = n22796 & ~n22815 ;
  assign n22817 = ( n16459 & n22815 ) | ( n16459 & ~n22816 ) | ( n22815 & ~n22816 ) ;
  assign n22818 = ( x788 & n22811 ) | ( x788 & n22817 ) | ( n22811 & n22817 ) ;
  assign n22819 = n22817 ^ n22811 ^ 1'b0 ;
  assign n22820 = ( x788 & n22818 ) | ( x788 & n22819 ) | ( n22818 & n22819 ) ;
  assign n22821 = n15524 | n22786 ;
  assign n22822 = n22752 & n22821 ;
  assign n22823 = x625 & ~n22821 ;
  assign n22824 = ( n22787 & n22822 ) | ( n22787 & n22823 ) | ( n22822 & n22823 ) ;
  assign n22825 = ( x608 & n22790 ) | ( x608 & ~n22824 ) | ( n22790 & ~n22824 ) ;
  assign n22826 = n22824 | n22825 ;
  assign n22827 = x1153 & n22752 ;
  assign n22828 = ~n22823 & n22827 ;
  assign n22829 = x608 & ~n22789 ;
  assign n22830 = n22826 & ~n22829 ;
  assign n22831 = ( n22826 & n22828 ) | ( n22826 & n22830 ) | ( n22828 & n22830 ) ;
  assign n22832 = n22822 ^ x778 ^ 1'b0 ;
  assign n22833 = ( n22822 & n22831 ) | ( n22822 & n22832 ) | ( n22831 & n22832 ) ;
  assign n22834 = x609 & ~n22833 ;
  assign n22835 = x609 | n22793 ;
  assign n22836 = ( x1155 & n22834 ) | ( x1155 & n22835 ) | ( n22834 & n22835 ) ;
  assign n22837 = ~n22834 & n22836 ;
  assign n22838 = ( x660 & n22757 ) | ( x660 & ~n22837 ) | ( n22757 & ~n22837 ) ;
  assign n22839 = ~n22757 & n22838 ;
  assign n22840 = x660 | n22755 ;
  assign n22841 = x609 & ~n22793 ;
  assign n22842 = x1155 | n22841 ;
  assign n22843 = ( n22833 & n22834 ) | ( n22833 & ~n22842 ) | ( n22834 & ~n22842 ) ;
  assign n22844 = ( ~n22839 & n22840 ) | ( ~n22839 & n22843 ) | ( n22840 & n22843 ) ;
  assign n22845 = ~n22839 & n22844 ;
  assign n22846 = n22833 ^ x785 ^ 1'b0 ;
  assign n22847 = ( n22833 & n22845 ) | ( n22833 & n22846 ) | ( n22845 & n22846 ) ;
  assign n22848 = x618 & ~n22847 ;
  assign n22849 = x618 | n22794 ;
  assign n22850 = ( x1154 & n22848 ) | ( x1154 & n22849 ) | ( n22848 & n22849 ) ;
  assign n22851 = ~n22848 & n22850 ;
  assign n22852 = ( x627 & n22764 ) | ( x627 & ~n22851 ) | ( n22764 & ~n22851 ) ;
  assign n22853 = ~n22764 & n22852 ;
  assign n22854 = x627 | n22762 ;
  assign n22855 = x618 & ~n22794 ;
  assign n22856 = x1154 | n22855 ;
  assign n22857 = ( n22847 & n22848 ) | ( n22847 & ~n22856 ) | ( n22848 & ~n22856 ) ;
  assign n22858 = ( ~n22853 & n22854 ) | ( ~n22853 & n22857 ) | ( n22854 & n22857 ) ;
  assign n22859 = ~n22853 & n22858 ;
  assign n22860 = n22847 ^ x781 ^ 1'b0 ;
  assign n22861 = ( n22847 & n22859 ) | ( n22847 & n22860 ) | ( n22859 & n22860 ) ;
  assign n22862 = ~x789 & n22861 ;
  assign n22863 = x619 & ~n22795 ;
  assign n22864 = x1159 | n22863 ;
  assign n22865 = x619 & ~n22861 ;
  assign n22866 = ( n22861 & ~n22864 ) | ( n22861 & n22865 ) | ( ~n22864 & n22865 ) ;
  assign n22867 = ( x648 & n22771 ) | ( x648 & ~n22866 ) | ( n22771 & ~n22866 ) ;
  assign n22868 = n22866 | n22867 ;
  assign n22869 = x619 | n22795 ;
  assign n22870 = x1159 & ~n22865 ;
  assign n22871 = n22869 & n22870 ;
  assign n22872 = ( x648 & n22774 ) | ( x648 & ~n22871 ) | ( n22774 & ~n22871 ) ;
  assign n22873 = ~n22774 & n22872 ;
  assign n22874 = x789 & ~n22873 ;
  assign n22875 = n22868 & n22874 ;
  assign n22876 = ( n16519 & ~n22862 ) | ( n16519 & n22875 ) | ( ~n22862 & n22875 ) ;
  assign n22877 = n22862 | n22876 ;
  assign n22878 = n22877 ^ n22820 ^ 1'b0 ;
  assign n22879 = ( n22820 & n22877 ) | ( n22820 & n22878 ) | ( n22877 & n22878 ) ;
  assign n22880 = ( n18482 & ~n22820 ) | ( n18482 & n22879 ) | ( ~n22820 & n22879 ) ;
  assign n22881 = n19208 | n22797 ;
  assign n22882 = n16556 & ~n22779 ;
  assign n22883 = x629 & ~n22882 ;
  assign n22884 = n22881 & n22883 ;
  assign n22885 = n16557 & ~n22779 ;
  assign n22886 = n19212 & ~n22797 ;
  assign n22887 = n22885 | n22886 ;
  assign n22888 = ( x629 & ~n22884 ) | ( x629 & n22887 ) | ( ~n22884 & n22887 ) ;
  assign n22889 = ~n22884 & n22888 ;
  assign n22890 = ( x792 & ~n19206 ) | ( x792 & n22889 ) | ( ~n19206 & n22889 ) ;
  assign n22891 = ( n18484 & n19206 ) | ( n18484 & n22890 ) | ( n19206 & n22890 ) ;
  assign n22892 = ( n22807 & n22880 ) | ( n22807 & ~n22891 ) | ( n22880 & ~n22891 ) ;
  assign n22893 = n22892 ^ n22880 ^ 1'b0 ;
  assign n22894 = ( n22807 & n22892 ) | ( n22807 & ~n22893 ) | ( n22892 & ~n22893 ) ;
  assign n22895 = x790 | n22894 ;
  assign n22896 = x644 & ~n22894 ;
  assign n22897 = ( x787 & n22800 ) | ( x787 & ~n22803 ) | ( n22800 & ~n22803 ) ;
  assign n22898 = ~n22800 & n22897 ;
  assign n22899 = ( x787 & n22798 ) | ( x787 & ~n22898 ) | ( n22798 & ~n22898 ) ;
  assign n22900 = ~n22898 & n22899 ;
  assign n22901 = x644 | n22900 ;
  assign n22902 = ( x715 & n22896 ) | ( x715 & n22901 ) | ( n22896 & n22901 ) ;
  assign n22903 = ~n22896 & n22902 ;
  assign n22904 = x644 | n22750 ;
  assign n22905 = n22750 ^ n16376 ^ 1'b0 ;
  assign n22906 = ( n22750 & n22781 ) | ( n22750 & ~n22905 ) | ( n22781 & ~n22905 ) ;
  assign n22907 = x644 & ~n22906 ;
  assign n22908 = ( x715 & n22904 ) | ( x715 & ~n22907 ) | ( n22904 & ~n22907 ) ;
  assign n22909 = ~x715 & n22908 ;
  assign n22910 = ( x1160 & n22903 ) | ( x1160 & ~n22909 ) | ( n22903 & ~n22909 ) ;
  assign n22911 = ~n22903 & n22910 ;
  assign n22912 = x644 & ~n22750 ;
  assign n22913 = x715 & ~n22912 ;
  assign n22914 = ( n22906 & n22907 ) | ( n22906 & n22913 ) | ( n22907 & n22913 ) ;
  assign n22915 = x644 & ~n22900 ;
  assign n22916 = x715 | n22915 ;
  assign n22917 = ( n22894 & n22896 ) | ( n22894 & ~n22916 ) | ( n22896 & ~n22916 ) ;
  assign n22918 = ( x1160 & ~n22914 ) | ( x1160 & n22917 ) | ( ~n22914 & n22917 ) ;
  assign n22919 = n22914 | n22918 ;
  assign n22920 = x790 & ~n22919 ;
  assign n22921 = ( x790 & n22911 ) | ( x790 & n22920 ) | ( n22911 & n22920 ) ;
  assign n22922 = x832 & ~n22921 ;
  assign n22923 = n22895 & n22922 ;
  assign n22924 = ~x176 & n7318 ;
  assign n22925 = x832 | n22924 ;
  assign n22926 = ~n22923 & n22925 ;
  assign n22927 = ( n22749 & n22923 ) | ( n22749 & ~n22926 ) | ( n22923 & ~n22926 ) ;
  assign n22928 = x177 | n17839 ;
  assign n22929 = ( x757 & n22572 ) | ( x757 & n22928 ) | ( n22572 & n22928 ) ;
  assign n22930 = ~x757 & n22929 ;
  assign n22931 = n17843 ^ x757 ^ 1'b0 ;
  assign n22932 = ( n15655 & n17843 ) | ( n15655 & n22931 ) | ( n17843 & n22931 ) ;
  assign n22933 = ( x177 & ~n22930 ) | ( x177 & n22932 ) | ( ~n22930 & n22932 ) ;
  assign n22934 = ~n22930 & n22933 ;
  assign n22963 = x686 & ~n22934 ;
  assign n22964 = x177 | n17897 ;
  assign n22965 = ( x38 & ~x177 ) | ( x38 & n17905 ) | ( ~x177 & n17905 ) ;
  assign n22966 = n22964 & n22965 ;
  assign n22967 = x177 & n17908 ;
  assign n22968 = n16048 ^ x39 ^ 1'b0 ;
  assign n22969 = ( n16003 & n16048 ) | ( n16003 & n22968 ) | ( n16048 & n22968 ) ;
  assign n22970 = x177 | n22969 ;
  assign n22971 = ( x38 & ~n22967 ) | ( x38 & n22970 ) | ( ~n22967 & n22970 ) ;
  assign n22972 = ~x38 & n22971 ;
  assign n22973 = ( x757 & ~n22966 ) | ( x757 & n22972 ) | ( ~n22966 & n22972 ) ;
  assign n22974 = n22966 | n22973 ;
  assign n22975 = x177 | n17891 ;
  assign n22976 = x177 & n17885 ;
  assign n22977 = ( x38 & n22975 ) | ( x38 & ~n22976 ) | ( n22975 & ~n22976 ) ;
  assign n22978 = ~x38 & n22977 ;
  assign n22979 = x177 | n15644 ;
  assign n22980 = n16659 & n22979 ;
  assign n22981 = ( x757 & n22978 ) | ( x757 & ~n22980 ) | ( n22978 & ~n22980 ) ;
  assign n22982 = ~n22978 & n22981 ;
  assign n22983 = ( x686 & n22974 ) | ( x686 & ~n22982 ) | ( n22974 & ~n22982 ) ;
  assign n22984 = n22983 ^ n22974 ^ 1'b0 ;
  assign n22985 = ( x686 & n22983 ) | ( x686 & ~n22984 ) | ( n22983 & ~n22984 ) ;
  assign n22986 = ( n2069 & ~n22963 ) | ( n2069 & n22985 ) | ( ~n22963 & n22985 ) ;
  assign n22987 = ~n2069 & n22986 ;
  assign n22988 = n22987 ^ x177 ^ 1'b0 ;
  assign n22989 = ( ~x177 & n2069 ) | ( ~x177 & n22988 ) | ( n2069 & n22988 ) ;
  assign n22990 = ( x177 & n22987 ) | ( x177 & n22989 ) | ( n22987 & n22989 ) ;
  assign n22991 = x625 & ~n22990 ;
  assign n22935 = n22934 ^ n2069 ^ 1'b0 ;
  assign n22936 = ( x177 & n22934 ) | ( x177 & n22935 ) | ( n22934 & n22935 ) ;
  assign n22992 = x625 | n22936 ;
  assign n22993 = ( x1153 & n22991 ) | ( x1153 & n22992 ) | ( n22991 & n22992 ) ;
  assign n22994 = ~n22991 & n22993 ;
  assign n22937 = x177 | n15656 ;
  assign n22995 = x625 & ~n22937 ;
  assign n22996 = x1153 | n22995 ;
  assign n22997 = n16185 & n22979 ;
  assign n22998 = ( x38 & x177 ) | ( x38 & n16700 ) | ( x177 & n16700 ) ;
  assign n22999 = ( x177 & n16697 ) | ( x177 & ~n22998 ) | ( n16697 & ~n22998 ) ;
  assign n23000 = ~n22998 & n22999 ;
  assign n23001 = ( x686 & ~n22997 ) | ( x686 & n23000 ) | ( ~n22997 & n23000 ) ;
  assign n23002 = n22997 | n23001 ;
  assign n23003 = ~x177 & x686 ;
  assign n23004 = ~n15655 & n23003 ;
  assign n23005 = ( n2069 & n23002 ) | ( n2069 & ~n23004 ) | ( n23002 & ~n23004 ) ;
  assign n23006 = ~n2069 & n23005 ;
  assign n23007 = n23006 ^ x177 ^ 1'b0 ;
  assign n23008 = ( ~x177 & n2069 ) | ( ~x177 & n23007 ) | ( n2069 & n23007 ) ;
  assign n23009 = ( x177 & n23006 ) | ( x177 & n23008 ) | ( n23006 & n23008 ) ;
  assign n23010 = ( x625 & ~n22996 ) | ( x625 & n23009 ) | ( ~n22996 & n23009 ) ;
  assign n23011 = ~n22996 & n23010 ;
  assign n23012 = ( x608 & n22994 ) | ( x608 & ~n23011 ) | ( n22994 & ~n23011 ) ;
  assign n23013 = ~n22994 & n23012 ;
  assign n23014 = x625 & ~n23009 ;
  assign n23015 = x625 | n22937 ;
  assign n23016 = ( x1153 & n23014 ) | ( x1153 & n23015 ) | ( n23014 & n23015 ) ;
  assign n23017 = ~n23014 & n23016 ;
  assign n23018 = x608 | n23017 ;
  assign n23019 = x625 & ~n22936 ;
  assign n23020 = x1153 | n23019 ;
  assign n23021 = ( n22990 & n22991 ) | ( n22990 & ~n23020 ) | ( n22991 & ~n23020 ) ;
  assign n23022 = ( ~n23013 & n23018 ) | ( ~n23013 & n23021 ) | ( n23018 & n23021 ) ;
  assign n23023 = ~n23013 & n23022 ;
  assign n23024 = n22990 ^ x778 ^ 1'b0 ;
  assign n23025 = ( n22990 & n23023 ) | ( n22990 & n23024 ) | ( n23023 & n23024 ) ;
  assign n23026 = x609 & ~n23025 ;
  assign n23027 = n23011 | n23017 ;
  assign n23028 = n23009 ^ x778 ^ 1'b0 ;
  assign n23029 = ( n23009 & n23027 ) | ( n23009 & n23028 ) | ( n23027 & n23028 ) ;
  assign n23030 = x609 | n23029 ;
  assign n23031 = ( x1155 & n23026 ) | ( x1155 & n23030 ) | ( n23026 & n23030 ) ;
  assign n23032 = ~n23026 & n23031 ;
  assign n22940 = ~n15659 & n22936 ;
  assign n22941 = x609 & n22940 ;
  assign n22942 = ~n15668 & n22937 ;
  assign n22943 = n22941 | n22942 ;
  assign n22938 = n22936 ^ n15659 ^ 1'b0 ;
  assign n22939 = ( n22936 & n22937 ) | ( n22936 & n22938 ) | ( n22937 & n22938 ) ;
  assign n22945 = n22943 ^ n22939 ^ n22937 ;
  assign n23033 = ~x1155 & n22945 ;
  assign n23034 = ( x660 & n23032 ) | ( x660 & ~n23033 ) | ( n23032 & ~n23033 ) ;
  assign n23035 = ~n23032 & n23034 ;
  assign n23036 = x1155 & n22943 ;
  assign n23037 = x660 | n23036 ;
  assign n23038 = x609 & ~n23029 ;
  assign n23039 = x1155 | n23038 ;
  assign n23040 = ( n23025 & n23026 ) | ( n23025 & ~n23039 ) | ( n23026 & ~n23039 ) ;
  assign n23041 = ( ~n23035 & n23037 ) | ( ~n23035 & n23040 ) | ( n23037 & n23040 ) ;
  assign n23042 = ~n23035 & n23041 ;
  assign n23043 = n23025 ^ x785 ^ 1'b0 ;
  assign n23044 = ( n23025 & n23042 ) | ( n23025 & n23043 ) | ( n23042 & n23043 ) ;
  assign n23045 = x618 & ~n23044 ;
  assign n23046 = n22937 ^ n16234 ^ 1'b0 ;
  assign n23047 = ( n22937 & n23029 ) | ( n22937 & ~n23046 ) | ( n23029 & ~n23046 ) ;
  assign n23048 = x618 | n23047 ;
  assign n23049 = ( x1154 & n23045 ) | ( x1154 & n23048 ) | ( n23045 & n23048 ) ;
  assign n23050 = ~n23045 & n23049 ;
  assign n22944 = n22943 ^ x1155 ^ 1'b0 ;
  assign n22946 = ( n22943 & ~n22944 ) | ( n22943 & n22945 ) | ( ~n22944 & n22945 ) ;
  assign n22947 = n22939 ^ x785 ^ 1'b0 ;
  assign n22948 = ( n22939 & n22946 ) | ( n22939 & n22947 ) | ( n22946 & n22947 ) ;
  assign n22949 = x618 & ~n22948 ;
  assign n22953 = x618 & ~n22937 ;
  assign n22954 = x1154 | n22953 ;
  assign n22955 = ( n22948 & n22949 ) | ( n22948 & ~n22954 ) | ( n22949 & ~n22954 ) ;
  assign n23051 = ( x627 & ~n22955 ) | ( x627 & n23050 ) | ( ~n22955 & n23050 ) ;
  assign n23052 = ~n23050 & n23051 ;
  assign n22950 = x618 | n22937 ;
  assign n22951 = ( x1154 & n22949 ) | ( x1154 & n22950 ) | ( n22949 & n22950 ) ;
  assign n22952 = ~n22949 & n22951 ;
  assign n23053 = x627 | n22952 ;
  assign n23054 = x618 & ~n23047 ;
  assign n23055 = x1154 | n23054 ;
  assign n23056 = ( n23044 & n23045 ) | ( n23044 & ~n23055 ) | ( n23045 & ~n23055 ) ;
  assign n23057 = ( ~n23052 & n23053 ) | ( ~n23052 & n23056 ) | ( n23053 & n23056 ) ;
  assign n23058 = ~n23052 & n23057 ;
  assign n23059 = n23044 ^ x781 ^ 1'b0 ;
  assign n23060 = ( n23044 & n23058 ) | ( n23044 & n23059 ) | ( n23058 & n23059 ) ;
  assign n23061 = x619 & ~n23060 ;
  assign n23062 = n22937 ^ n16254 ^ 1'b0 ;
  assign n23063 = ( n22937 & n23047 ) | ( n22937 & ~n23062 ) | ( n23047 & ~n23062 ) ;
  assign n23069 = x619 | n23063 ;
  assign n23070 = ( x1159 & n23061 ) | ( x1159 & n23069 ) | ( n23061 & n23069 ) ;
  assign n23071 = ~n23061 & n23070 ;
  assign n22956 = n22952 | n22955 ;
  assign n22957 = n22948 ^ x781 ^ 1'b0 ;
  assign n22958 = ( n22948 & n22956 ) | ( n22948 & n22957 ) | ( n22956 & n22957 ) ;
  assign n22959 = x619 & ~n22958 ;
  assign n23072 = x619 & ~n22937 ;
  assign n23073 = x1159 | n23072 ;
  assign n23074 = ( n22958 & n22959 ) | ( n22958 & ~n23073 ) | ( n22959 & ~n23073 ) ;
  assign n23075 = ( x648 & n23071 ) | ( x648 & ~n23074 ) | ( n23071 & ~n23074 ) ;
  assign n23076 = ~n23071 & n23075 ;
  assign n22960 = x619 | n22937 ;
  assign n22961 = ( x1159 & n22959 ) | ( x1159 & n22960 ) | ( n22959 & n22960 ) ;
  assign n22962 = ~n22959 & n22961 ;
  assign n23064 = x619 & ~n23063 ;
  assign n23065 = x1159 | n23064 ;
  assign n23066 = ( n23060 & n23061 ) | ( n23060 & ~n23065 ) | ( n23061 & ~n23065 ) ;
  assign n23067 = ( x648 & ~n22962 ) | ( x648 & n23066 ) | ( ~n22962 & n23066 ) ;
  assign n23068 = n22962 | n23067 ;
  assign n23077 = n23076 ^ n23068 ^ 1'b0 ;
  assign n23078 = ( x789 & ~n23068 ) | ( x789 & n23076 ) | ( ~n23068 & n23076 ) ;
  assign n23079 = ( x789 & ~n23077 ) | ( x789 & n23078 ) | ( ~n23077 & n23078 ) ;
  assign n23080 = ( x789 & n23060 ) | ( x789 & ~n23079 ) | ( n23060 & ~n23079 ) ;
  assign n23081 = ~n23079 & n23080 ;
  assign n23082 = ~x626 & n23081 ;
  assign n23083 = n22937 ^ n16279 ^ 1'b0 ;
  assign n23084 = ( n22937 & n23063 ) | ( n22937 & ~n23083 ) | ( n23063 & ~n23083 ) ;
  assign n23085 = x626 & n23084 ;
  assign n23086 = ( x641 & ~n23082 ) | ( x641 & n23085 ) | ( ~n23082 & n23085 ) ;
  assign n23087 = n23082 | n23086 ;
  assign n23088 = ~x626 & n22937 ;
  assign n23089 = n22962 | n23074 ;
  assign n23090 = n22958 ^ x789 ^ 1'b0 ;
  assign n23091 = ( n22958 & n23089 ) | ( n22958 & n23090 ) | ( n23089 & n23090 ) ;
  assign n23092 = x626 & n23091 ;
  assign n23093 = ( x641 & ~n23088 ) | ( x641 & n23092 ) | ( ~n23088 & n23092 ) ;
  assign n23094 = n23088 | n23093 ;
  assign n23095 = ~x626 & n23084 ;
  assign n23096 = x626 & n23081 ;
  assign n23097 = ( x641 & n23095 ) | ( x641 & ~n23096 ) | ( n23095 & ~n23096 ) ;
  assign n23098 = ~n23095 & n23097 ;
  assign n23099 = x1158 & ~n23098 ;
  assign n23100 = n23094 & n23099 ;
  assign n23101 = ~x626 & n23091 ;
  assign n23102 = x626 & n22937 ;
  assign n23103 = x641 & ~n23102 ;
  assign n23104 = n23103 ^ n23101 ^ 1'b0 ;
  assign n23105 = ( n23101 & n23103 ) | ( n23101 & n23104 ) | ( n23103 & n23104 ) ;
  assign n23106 = ( x1158 & ~n23101 ) | ( x1158 & n23105 ) | ( ~n23101 & n23105 ) ;
  assign n23107 = ~n23100 & n23106 ;
  assign n23108 = ( n23087 & n23100 ) | ( n23087 & ~n23107 ) | ( n23100 & ~n23107 ) ;
  assign n23109 = n23081 ^ x788 ^ 1'b0 ;
  assign n23110 = ( n23081 & n23108 ) | ( n23081 & n23109 ) | ( n23108 & n23109 ) ;
  assign n23111 = x628 & ~n23110 ;
  assign n23112 = n22937 ^ n16518 ^ 1'b0 ;
  assign n23113 = ( n22937 & n23091 ) | ( n22937 & ~n23112 ) | ( n23091 & ~n23112 ) ;
  assign n23114 = x628 | n23113 ;
  assign n23115 = ( x1156 & n23111 ) | ( x1156 & n23114 ) | ( n23111 & n23114 ) ;
  assign n23116 = ~n23111 & n23115 ;
  assign n23117 = x628 & ~n22937 ;
  assign n23118 = x1156 | n23117 ;
  assign n23119 = n22937 ^ n16318 ^ 1'b0 ;
  assign n23120 = ( n22937 & n23084 ) | ( n22937 & ~n23119 ) | ( n23084 & ~n23119 ) ;
  assign n23121 = x628 & ~n23120 ;
  assign n23122 = ( ~n23118 & n23120 ) | ( ~n23118 & n23121 ) | ( n23120 & n23121 ) ;
  assign n23123 = ( x629 & n23116 ) | ( x629 & ~n23122 ) | ( n23116 & ~n23122 ) ;
  assign n23124 = ~n23116 & n23123 ;
  assign n23125 = x628 | n22937 ;
  assign n23126 = ( x1156 & n23121 ) | ( x1156 & n23125 ) | ( n23121 & n23125 ) ;
  assign n23127 = ~n23121 & n23126 ;
  assign n23128 = x629 | n23127 ;
  assign n23129 = x628 & ~n23113 ;
  assign n23130 = x1156 | n23129 ;
  assign n23131 = ( n23110 & n23111 ) | ( n23110 & ~n23130 ) | ( n23111 & ~n23130 ) ;
  assign n23132 = ( ~n23124 & n23128 ) | ( ~n23124 & n23131 ) | ( n23128 & n23131 ) ;
  assign n23133 = ~n23124 & n23132 ;
  assign n23134 = n23110 ^ x792 ^ 1'b0 ;
  assign n23135 = ( n23110 & n23133 ) | ( n23110 & n23134 ) | ( n23133 & n23134 ) ;
  assign n23136 = x647 & ~n23135 ;
  assign n23137 = n22937 ^ n16339 ^ 1'b0 ;
  assign n23138 = ( n22937 & n23113 ) | ( n22937 & ~n23137 ) | ( n23113 & ~n23137 ) ;
  assign n23139 = x647 | n23138 ;
  assign n23140 = ( x1157 & n23136 ) | ( x1157 & n23139 ) | ( n23136 & n23139 ) ;
  assign n23141 = ~n23136 & n23140 ;
  assign n23142 = x647 & ~n22937 ;
  assign n23143 = x1157 | n23142 ;
  assign n23144 = n23122 | n23127 ;
  assign n23145 = n23120 ^ x792 ^ 1'b0 ;
  assign n23146 = ( n23120 & n23144 ) | ( n23120 & n23145 ) | ( n23144 & n23145 ) ;
  assign n23147 = x647 & ~n23146 ;
  assign n23148 = ( ~n23143 & n23146 ) | ( ~n23143 & n23147 ) | ( n23146 & n23147 ) ;
  assign n23149 = ( x630 & n23141 ) | ( x630 & ~n23148 ) | ( n23141 & ~n23148 ) ;
  assign n23150 = ~n23141 & n23149 ;
  assign n23151 = x647 | n22937 ;
  assign n23152 = ( x1157 & n23147 ) | ( x1157 & n23151 ) | ( n23147 & n23151 ) ;
  assign n23153 = ~n23147 & n23152 ;
  assign n23154 = x630 | n23153 ;
  assign n23155 = x647 & ~n23138 ;
  assign n23156 = x1157 | n23155 ;
  assign n23157 = ( n23135 & n23136 ) | ( n23135 & ~n23156 ) | ( n23136 & ~n23156 ) ;
  assign n23158 = ( ~n23150 & n23154 ) | ( ~n23150 & n23157 ) | ( n23154 & n23157 ) ;
  assign n23159 = ~n23150 & n23158 ;
  assign n23160 = n23135 ^ x787 ^ 1'b0 ;
  assign n23161 = ( n23135 & n23159 ) | ( n23135 & n23160 ) | ( n23159 & n23160 ) ;
  assign n23162 = x644 & ~n23161 ;
  assign n23163 = n23148 | n23153 ;
  assign n23164 = n23146 ^ x787 ^ 1'b0 ;
  assign n23165 = ( n23146 & n23163 ) | ( n23146 & n23164 ) | ( n23163 & n23164 ) ;
  assign n23166 = x644 | n23165 ;
  assign n23167 = ( x715 & n23162 ) | ( x715 & n23166 ) | ( n23162 & n23166 ) ;
  assign n23168 = ~n23162 & n23167 ;
  assign n23169 = x644 | n22937 ;
  assign n23170 = n22937 ^ n16376 ^ 1'b0 ;
  assign n23171 = ( n22937 & n23138 ) | ( n22937 & ~n23170 ) | ( n23138 & ~n23170 ) ;
  assign n23172 = x644 & ~n23171 ;
  assign n23173 = ( x715 & n23169 ) | ( x715 & ~n23172 ) | ( n23169 & ~n23172 ) ;
  assign n23174 = ~x715 & n23173 ;
  assign n23175 = ( x1160 & n23168 ) | ( x1160 & ~n23174 ) | ( n23168 & ~n23174 ) ;
  assign n23176 = ~n23168 & n23175 ;
  assign n23177 = x644 & ~n22937 ;
  assign n23178 = x715 & ~n23177 ;
  assign n23179 = ( n23171 & n23172 ) | ( n23171 & n23178 ) | ( n23172 & n23178 ) ;
  assign n23180 = x644 & ~n23165 ;
  assign n23181 = x715 | n23180 ;
  assign n23182 = ( n23161 & n23162 ) | ( n23161 & ~n23181 ) | ( n23162 & ~n23181 ) ;
  assign n23183 = ( x1160 & ~n23179 ) | ( x1160 & n23182 ) | ( ~n23179 & n23182 ) ;
  assign n23184 = n23179 | n23183 ;
  assign n23185 = ( x790 & n23176 ) | ( x790 & n23184 ) | ( n23176 & n23184 ) ;
  assign n23186 = ~n23176 & n23185 ;
  assign n23187 = ~x790 & n23161 ;
  assign n23188 = ( n7318 & ~n23186 ) | ( n7318 & n23187 ) | ( ~n23186 & n23187 ) ;
  assign n23189 = n23186 | n23188 ;
  assign n23190 = x177 | n1611 ;
  assign n23191 = ~x757 & n15591 ;
  assign n23192 = n23190 & ~n23191 ;
  assign n23193 = n16397 | n23192 ;
  assign n23194 = n16402 | n23192 ;
  assign n23195 = x1155 & n23194 ;
  assign n23196 = n16405 | n23193 ;
  assign n23197 = ~x1155 & n23196 ;
  assign n23198 = n23195 | n23197 ;
  assign n23199 = n23193 ^ x785 ^ 1'b0 ;
  assign n23200 = ( n23193 & n23198 ) | ( n23193 & n23199 ) | ( n23198 & n23199 ) ;
  assign n23201 = n16411 | n23200 ;
  assign n23202 = x1154 & n23201 ;
  assign n23203 = n16414 | n23200 ;
  assign n23204 = ~x1154 & n23203 ;
  assign n23205 = n23202 | n23204 ;
  assign n23206 = n23200 ^ x781 ^ 1'b0 ;
  assign n23207 = ( n23200 & n23205 ) | ( n23200 & n23206 ) | ( n23205 & n23206 ) ;
  assign n23208 = x619 & ~n23207 ;
  assign n23209 = x619 | n23190 ;
  assign n23210 = ( x1159 & n23208 ) | ( x1159 & n23209 ) | ( n23208 & n23209 ) ;
  assign n23211 = ~n23208 & n23210 ;
  assign n23212 = x619 & ~n23190 ;
  assign n23213 = x1159 | n23212 ;
  assign n23214 = ( n23207 & n23208 ) | ( n23207 & ~n23213 ) | ( n23208 & ~n23213 ) ;
  assign n23215 = n23211 | n23214 ;
  assign n23216 = n23207 ^ x789 ^ 1'b0 ;
  assign n23217 = ( n23207 & n23215 ) | ( n23207 & n23216 ) | ( n23215 & n23216 ) ;
  assign n23218 = n23190 ^ n16518 ^ 1'b0 ;
  assign n23219 = ( n23190 & n23217 ) | ( n23190 & ~n23218 ) | ( n23217 & ~n23218 ) ;
  assign n23220 = n23190 ^ n16339 ^ 1'b0 ;
  assign n23221 = ( n23190 & n23219 ) | ( n23190 & ~n23220 ) | ( n23219 & ~n23220 ) ;
  assign n23222 = n19055 & n23221 ;
  assign n23223 = x647 & ~n23190 ;
  assign n23224 = x1157 | n23223 ;
  assign n23225 = ~x686 & n15778 ;
  assign n23226 = n23190 & ~n23225 ;
  assign n23227 = ~x1153 & n23190 ;
  assign n23228 = ~x625 & n23225 ;
  assign n23229 = n23227 & ~n23228 ;
  assign n23230 = ( x1153 & n23226 ) | ( x1153 & n23228 ) | ( n23226 & n23228 ) ;
  assign n23231 = n23229 | n23230 ;
  assign n23232 = n23226 ^ x778 ^ 1'b0 ;
  assign n23233 = ( n23226 & n23231 ) | ( n23226 & n23232 ) | ( n23231 & n23232 ) ;
  assign n23234 = n16447 | n23233 ;
  assign n23235 = n16449 | n23234 ;
  assign n23236 = n16451 | n23235 ;
  assign n23237 = n16530 | n23236 ;
  assign n23238 = n16560 | n23237 ;
  assign n23239 = ( x647 & ~n23224 ) | ( x647 & n23238 ) | ( ~n23224 & n23238 ) ;
  assign n23240 = ~n23224 & n23239 ;
  assign n23241 = n23190 ^ x647 ^ 1'b0 ;
  assign n23242 = ( n23190 & n23238 ) | ( n23190 & n23241 ) | ( n23238 & n23241 ) ;
  assign n23243 = x1157 & n23242 ;
  assign n23244 = ( n16375 & n23240 ) | ( n16375 & n23243 ) | ( n23240 & n23243 ) ;
  assign n23245 = ( x787 & n23222 ) | ( x787 & n23244 ) | ( n23222 & n23244 ) ;
  assign n23246 = n23244 ^ n23222 ^ 1'b0 ;
  assign n23247 = ( x787 & n23245 ) | ( x787 & n23246 ) | ( n23245 & n23246 ) ;
  assign n23248 = ~x626 & n23190 ;
  assign n23249 = x626 & n23217 ;
  assign n23250 = ( n22317 & n23248 ) | ( n22317 & ~n23249 ) | ( n23248 & ~n23249 ) ;
  assign n23251 = ~n23248 & n23250 ;
  assign n23252 = ~x626 & n23217 ;
  assign n23253 = x626 & n23190 ;
  assign n23254 = ( n22322 & n23252 ) | ( n22322 & ~n23253 ) | ( n23252 & ~n23253 ) ;
  assign n23255 = ~n23252 & n23254 ;
  assign n23256 = n23236 & ~n23255 ;
  assign n23257 = ( n16459 & n23255 ) | ( n16459 & ~n23256 ) | ( n23255 & ~n23256 ) ;
  assign n23258 = ( x788 & n23251 ) | ( x788 & n23257 ) | ( n23251 & n23257 ) ;
  assign n23259 = n23257 ^ n23251 ^ 1'b0 ;
  assign n23260 = ( x788 & n23258 ) | ( x788 & n23259 ) | ( n23258 & n23259 ) ;
  assign n23261 = n15524 | n23226 ;
  assign n23262 = n23192 & n23261 ;
  assign n23263 = x625 & ~n23261 ;
  assign n23264 = ( n23227 & n23262 ) | ( n23227 & n23263 ) | ( n23262 & n23263 ) ;
  assign n23265 = ( x608 & n23230 ) | ( x608 & ~n23264 ) | ( n23230 & ~n23264 ) ;
  assign n23266 = n23264 | n23265 ;
  assign n23267 = x1153 & n23192 ;
  assign n23268 = ~n23263 & n23267 ;
  assign n23269 = x608 & ~n23229 ;
  assign n23270 = n23266 & ~n23269 ;
  assign n23271 = ( n23266 & n23268 ) | ( n23266 & n23270 ) | ( n23268 & n23270 ) ;
  assign n23272 = n23262 ^ x778 ^ 1'b0 ;
  assign n23273 = ( n23262 & n23271 ) | ( n23262 & n23272 ) | ( n23271 & n23272 ) ;
  assign n23274 = x609 & ~n23273 ;
  assign n23275 = x609 | n23233 ;
  assign n23276 = ( x1155 & n23274 ) | ( x1155 & n23275 ) | ( n23274 & n23275 ) ;
  assign n23277 = ~n23274 & n23276 ;
  assign n23278 = ( x660 & n23197 ) | ( x660 & ~n23277 ) | ( n23197 & ~n23277 ) ;
  assign n23279 = ~n23197 & n23278 ;
  assign n23280 = x660 | n23195 ;
  assign n23281 = x609 & ~n23233 ;
  assign n23282 = x1155 | n23281 ;
  assign n23283 = ( n23273 & n23274 ) | ( n23273 & ~n23282 ) | ( n23274 & ~n23282 ) ;
  assign n23284 = ( ~n23279 & n23280 ) | ( ~n23279 & n23283 ) | ( n23280 & n23283 ) ;
  assign n23285 = ~n23279 & n23284 ;
  assign n23286 = n23273 ^ x785 ^ 1'b0 ;
  assign n23287 = ( n23273 & n23285 ) | ( n23273 & n23286 ) | ( n23285 & n23286 ) ;
  assign n23288 = x618 & ~n23287 ;
  assign n23289 = x618 | n23234 ;
  assign n23290 = ( x1154 & n23288 ) | ( x1154 & n23289 ) | ( n23288 & n23289 ) ;
  assign n23291 = ~n23288 & n23290 ;
  assign n23292 = ( x627 & n23204 ) | ( x627 & ~n23291 ) | ( n23204 & ~n23291 ) ;
  assign n23293 = ~n23204 & n23292 ;
  assign n23294 = x627 | n23202 ;
  assign n23295 = x618 & ~n23234 ;
  assign n23296 = x1154 | n23295 ;
  assign n23297 = ( n23287 & n23288 ) | ( n23287 & ~n23296 ) | ( n23288 & ~n23296 ) ;
  assign n23298 = ( ~n23293 & n23294 ) | ( ~n23293 & n23297 ) | ( n23294 & n23297 ) ;
  assign n23299 = ~n23293 & n23298 ;
  assign n23300 = n23287 ^ x781 ^ 1'b0 ;
  assign n23301 = ( n23287 & n23299 ) | ( n23287 & n23300 ) | ( n23299 & n23300 ) ;
  assign n23302 = ~x789 & n23301 ;
  assign n23303 = x619 & ~n23235 ;
  assign n23304 = x1159 | n23303 ;
  assign n23305 = x619 & ~n23301 ;
  assign n23306 = ( n23301 & ~n23304 ) | ( n23301 & n23305 ) | ( ~n23304 & n23305 ) ;
  assign n23307 = ( x648 & n23211 ) | ( x648 & ~n23306 ) | ( n23211 & ~n23306 ) ;
  assign n23308 = n23306 | n23307 ;
  assign n23309 = x619 | n23235 ;
  assign n23310 = x1159 & ~n23305 ;
  assign n23311 = n23309 & n23310 ;
  assign n23312 = ( x648 & n23214 ) | ( x648 & ~n23311 ) | ( n23214 & ~n23311 ) ;
  assign n23313 = ~n23214 & n23312 ;
  assign n23314 = x789 & ~n23313 ;
  assign n23315 = n23308 & n23314 ;
  assign n23316 = ( n16519 & ~n23302 ) | ( n16519 & n23315 ) | ( ~n23302 & n23315 ) ;
  assign n23317 = n23302 | n23316 ;
  assign n23318 = n23317 ^ n23260 ^ 1'b0 ;
  assign n23319 = ( n23260 & n23317 ) | ( n23260 & n23318 ) | ( n23317 & n23318 ) ;
  assign n23320 = ( n18482 & ~n23260 ) | ( n18482 & n23319 ) | ( ~n23260 & n23319 ) ;
  assign n23321 = n19208 | n23237 ;
  assign n23322 = n16556 & ~n23219 ;
  assign n23323 = x629 & ~n23322 ;
  assign n23324 = n23321 & n23323 ;
  assign n23325 = n16557 & ~n23219 ;
  assign n23326 = n19212 & ~n23237 ;
  assign n23327 = n23325 | n23326 ;
  assign n23328 = ( x629 & ~n23324 ) | ( x629 & n23327 ) | ( ~n23324 & n23327 ) ;
  assign n23329 = ~n23324 & n23328 ;
  assign n23330 = ( x792 & ~n19206 ) | ( x792 & n23329 ) | ( ~n19206 & n23329 ) ;
  assign n23331 = ( n18484 & n19206 ) | ( n18484 & n23330 ) | ( n19206 & n23330 ) ;
  assign n23332 = ( n23247 & n23320 ) | ( n23247 & ~n23331 ) | ( n23320 & ~n23331 ) ;
  assign n23333 = n23332 ^ n23320 ^ 1'b0 ;
  assign n23334 = ( n23247 & n23332 ) | ( n23247 & ~n23333 ) | ( n23332 & ~n23333 ) ;
  assign n23335 = x790 | n23334 ;
  assign n23336 = x644 & ~n23334 ;
  assign n23337 = ( x787 & n23240 ) | ( x787 & ~n23243 ) | ( n23240 & ~n23243 ) ;
  assign n23338 = ~n23240 & n23337 ;
  assign n23339 = ( x787 & n23238 ) | ( x787 & ~n23338 ) | ( n23238 & ~n23338 ) ;
  assign n23340 = ~n23338 & n23339 ;
  assign n23341 = x644 | n23340 ;
  assign n23342 = ( x715 & n23336 ) | ( x715 & n23341 ) | ( n23336 & n23341 ) ;
  assign n23343 = ~n23336 & n23342 ;
  assign n23344 = x644 | n23190 ;
  assign n23345 = n23190 ^ n16376 ^ 1'b0 ;
  assign n23346 = ( n23190 & n23221 ) | ( n23190 & ~n23345 ) | ( n23221 & ~n23345 ) ;
  assign n23347 = x644 & ~n23346 ;
  assign n23348 = ( x715 & n23344 ) | ( x715 & ~n23347 ) | ( n23344 & ~n23347 ) ;
  assign n23349 = ~x715 & n23348 ;
  assign n23350 = ( x1160 & n23343 ) | ( x1160 & ~n23349 ) | ( n23343 & ~n23349 ) ;
  assign n23351 = ~n23343 & n23350 ;
  assign n23352 = x644 & ~n23190 ;
  assign n23353 = x715 & ~n23352 ;
  assign n23354 = ( n23346 & n23347 ) | ( n23346 & n23353 ) | ( n23347 & n23353 ) ;
  assign n23355 = x644 & ~n23340 ;
  assign n23356 = x715 | n23355 ;
  assign n23357 = ( n23334 & n23336 ) | ( n23334 & ~n23356 ) | ( n23336 & ~n23356 ) ;
  assign n23358 = ( x1160 & ~n23354 ) | ( x1160 & n23357 ) | ( ~n23354 & n23357 ) ;
  assign n23359 = n23354 | n23358 ;
  assign n23360 = x790 & ~n23359 ;
  assign n23361 = ( x790 & n23351 ) | ( x790 & n23360 ) | ( n23351 & n23360 ) ;
  assign n23362 = x832 & ~n23361 ;
  assign n23363 = n23335 & n23362 ;
  assign n23364 = ~x177 & n7318 ;
  assign n23365 = x832 | n23364 ;
  assign n23366 = ~n23363 & n23365 ;
  assign n23367 = ( n23189 & n23363 ) | ( n23189 & ~n23366 ) | ( n23363 & ~n23366 ) ;
  assign n23368 = x178 | n15656 ;
  assign n23369 = x688 | n2069 ;
  assign n23370 = ~n23368 & n23369 ;
  assign n23371 = ( x38 & x178 ) | ( x38 & n16700 ) | ( x178 & n16700 ) ;
  assign n23372 = ~n2069 & n23371 ;
  assign n23373 = ( x178 & n16697 ) | ( x178 & ~n23372 ) | ( n16697 & ~n23372 ) ;
  assign n23374 = ~n23372 & n23373 ;
  assign n23375 = x178 | n15644 ;
  assign n23376 = n16185 & n23375 ;
  assign n23377 = x688 | n23376 ;
  assign n23378 = ( ~n23370 & n23374 ) | ( ~n23370 & n23377 ) | ( n23374 & n23377 ) ;
  assign n23379 = ~n23370 & n23378 ;
  assign n23380 = x625 & ~n23379 ;
  assign n23381 = x625 | n23368 ;
  assign n23382 = ( x1153 & n23380 ) | ( x1153 & n23381 ) | ( n23380 & n23381 ) ;
  assign n23383 = ~n23380 & n23382 ;
  assign n23384 = x625 & ~n23368 ;
  assign n23385 = x1153 | n23384 ;
  assign n23386 = ( x625 & n23379 ) | ( x625 & ~n23385 ) | ( n23379 & ~n23385 ) ;
  assign n23387 = ~n23385 & n23386 ;
  assign n23388 = n23383 | n23387 ;
  assign n23389 = n23379 ^ x778 ^ 1'b0 ;
  assign n23390 = ( n23379 & n23388 ) | ( n23379 & n23389 ) | ( n23388 & n23389 ) ;
  assign n23391 = n23368 ^ n16234 ^ 1'b0 ;
  assign n23392 = ( n23368 & n23390 ) | ( n23368 & ~n23391 ) | ( n23390 & ~n23391 ) ;
  assign n23393 = n23368 ^ n16254 ^ 1'b0 ;
  assign n23394 = ( n23368 & n23392 ) | ( n23368 & ~n23393 ) | ( n23392 & ~n23393 ) ;
  assign n23395 = n23368 ^ n16279 ^ 1'b0 ;
  assign n23396 = ( n23368 & n23394 ) | ( n23368 & ~n23395 ) | ( n23394 & ~n23395 ) ;
  assign n23397 = n23368 ^ n16318 ^ 1'b0 ;
  assign n23398 = ( n23368 & n23396 ) | ( n23368 & ~n23397 ) | ( n23396 & ~n23397 ) ;
  assign n23399 = x628 & ~n23398 ;
  assign n23400 = x628 | n23368 ;
  assign n23401 = ( x1156 & n23399 ) | ( x1156 & n23400 ) | ( n23399 & n23400 ) ;
  assign n23402 = ~n23399 & n23401 ;
  assign n23403 = x628 & ~n23368 ;
  assign n23404 = x1156 | n23403 ;
  assign n23405 = ( n23398 & n23399 ) | ( n23398 & ~n23404 ) | ( n23399 & ~n23404 ) ;
  assign n23406 = n23402 | n23405 ;
  assign n23407 = n23398 ^ x792 ^ 1'b0 ;
  assign n23408 = ( n23398 & n23406 ) | ( n23398 & n23407 ) | ( n23406 & n23407 ) ;
  assign n23409 = n23368 ^ x647 ^ 1'b0 ;
  assign n23410 = ( n23368 & n23408 ) | ( n23368 & ~n23409 ) | ( n23408 & ~n23409 ) ;
  assign n23411 = ( n23368 & n23408 ) | ( n23368 & n23409 ) | ( n23408 & n23409 ) ;
  assign n23412 = n23410 ^ x1157 ^ 1'b0 ;
  assign n23413 = ( n23410 & n23411 ) | ( n23410 & n23412 ) | ( n23411 & n23412 ) ;
  assign n23414 = n23408 ^ x787 ^ 1'b0 ;
  assign n23415 = ( n23408 & n23413 ) | ( n23408 & n23414 ) | ( n23413 & n23414 ) ;
  assign n23416 = x644 & ~n23415 ;
  assign n23417 = x715 | n23416 ;
  assign n23418 = x644 & ~n23368 ;
  assign n23419 = x715 & ~n23418 ;
  assign n23420 = n23419 ^ x1160 ^ 1'b0 ;
  assign n23421 = ~x760 & n15646 ;
  assign n23422 = n23375 & ~n23421 ;
  assign n23423 = ~x178 & x760 ;
  assign n23424 = ~n15488 & n23423 ;
  assign n23425 = ~x178 & n15587 ;
  assign n23426 = x178 & ~n15640 ;
  assign n23427 = x760 | n23426 ;
  assign n23428 = ( ~n23424 & n23425 ) | ( ~n23424 & n23427 ) | ( n23425 & n23427 ) ;
  assign n23429 = ~n23424 & n23428 ;
  assign n23430 = n23422 ^ x38 ^ 1'b0 ;
  assign n23431 = ( n23422 & n23429 ) | ( n23422 & ~n23430 ) | ( n23429 & ~n23430 ) ;
  assign n23432 = ~n2069 & n23431 ;
  assign n23433 = x178 & n2069 ;
  assign n23434 = n23432 | n23433 ;
  assign n23435 = n23368 ^ n15659 ^ 1'b0 ;
  assign n23436 = ( n23368 & n23434 ) | ( n23368 & ~n23435 ) | ( n23434 & ~n23435 ) ;
  assign n23437 = n15662 & n23368 ;
  assign n23438 = ( ~n15662 & n23432 ) | ( ~n15662 & n23433 ) | ( n23432 & n23433 ) ;
  assign n23439 = n23437 | n23438 ;
  assign n23440 = n23439 ^ n23436 ^ n23368 ;
  assign n23441 = n23440 ^ x1155 ^ 1'b0 ;
  assign n23442 = ( n23439 & n23440 ) | ( n23439 & ~n23441 ) | ( n23440 & ~n23441 ) ;
  assign n23443 = n23436 ^ x785 ^ 1'b0 ;
  assign n23444 = ( n23436 & n23442 ) | ( n23436 & n23443 ) | ( n23442 & n23443 ) ;
  assign n23445 = x618 & ~n23444 ;
  assign n23446 = x618 | n23368 ;
  assign n23447 = ( x1154 & n23445 ) | ( x1154 & n23446 ) | ( n23445 & n23446 ) ;
  assign n23448 = ~n23445 & n23447 ;
  assign n23449 = x618 & ~n23368 ;
  assign n23450 = x1154 | n23449 ;
  assign n23451 = ( n23444 & n23445 ) | ( n23444 & ~n23450 ) | ( n23445 & ~n23450 ) ;
  assign n23452 = n23448 | n23451 ;
  assign n23453 = n23444 ^ x781 ^ 1'b0 ;
  assign n23454 = ( n23444 & n23452 ) | ( n23444 & n23453 ) | ( n23452 & n23453 ) ;
  assign n23455 = x619 & ~n23454 ;
  assign n23456 = x619 | n23368 ;
  assign n23457 = ( x1159 & n23455 ) | ( x1159 & n23456 ) | ( n23455 & n23456 ) ;
  assign n23458 = ~n23455 & n23457 ;
  assign n23459 = x619 & ~n23368 ;
  assign n23460 = x1159 | n23459 ;
  assign n23461 = ( n23454 & n23455 ) | ( n23454 & ~n23460 ) | ( n23455 & ~n23460 ) ;
  assign n23462 = n23458 | n23461 ;
  assign n23463 = n23454 ^ x789 ^ 1'b0 ;
  assign n23464 = ( n23454 & n23462 ) | ( n23454 & n23463 ) | ( n23462 & n23463 ) ;
  assign n23465 = n23368 ^ n16518 ^ 1'b0 ;
  assign n23466 = ( n23368 & n23464 ) | ( n23368 & ~n23465 ) | ( n23464 & ~n23465 ) ;
  assign n23467 = n23368 ^ n16339 ^ 1'b0 ;
  assign n23468 = ( n23368 & n23466 ) | ( n23368 & ~n23467 ) | ( n23466 & ~n23467 ) ;
  assign n23469 = n23368 ^ n16376 ^ 1'b0 ;
  assign n23470 = ( n23368 & n23468 ) | ( n23368 & ~n23469 ) | ( n23468 & ~n23469 ) ;
  assign n23471 = x644 | n23470 ;
  assign n23472 = ( n23419 & ~n23420 ) | ( n23419 & n23471 ) | ( ~n23420 & n23471 ) ;
  assign n23473 = ( x1160 & n23420 ) | ( x1160 & n23472 ) | ( n23420 & n23472 ) ;
  assign n23474 = n23417 & ~n23473 ;
  assign n23475 = x644 & ~n23470 ;
  assign n23476 = ( ~x715 & n23368 ) | ( ~x715 & n23418 ) | ( n23368 & n23418 ) ;
  assign n23477 = x1160 & ~n23476 ;
  assign n23478 = ( x1160 & n23475 ) | ( x1160 & n23477 ) | ( n23475 & n23477 ) ;
  assign n23479 = ( x715 & n23415 ) | ( x715 & n23416 ) | ( n23415 & n23416 ) ;
  assign n23480 = n23478 & ~n23479 ;
  assign n23481 = ( x790 & n23474 ) | ( x790 & n23480 ) | ( n23474 & n23480 ) ;
  assign n23482 = n23480 ^ n23474 ^ 1'b0 ;
  assign n23483 = ( x790 & n23481 ) | ( x790 & n23482 ) | ( n23481 & n23482 ) ;
  assign n23484 = n19055 & n23468 ;
  assign n23485 = n16374 & n23410 ;
  assign n23486 = n16373 & n23411 ;
  assign n23487 = n23485 | n23486 ;
  assign n23488 = ( x787 & n23484 ) | ( x787 & n23487 ) | ( n23484 & n23487 ) ;
  assign n23489 = n23487 ^ n23484 ^ 1'b0 ;
  assign n23490 = ( x787 & n23488 ) | ( x787 & n23489 ) | ( n23488 & n23489 ) ;
  assign n23491 = x688 & ~n23431 ;
  assign n23492 = x178 & ~n16054 ;
  assign n23493 = ~x178 & n16048 ;
  assign n23494 = ( x760 & ~n23492 ) | ( x760 & n23493 ) | ( ~n23492 & n23493 ) ;
  assign n23495 = n23492 | n23494 ;
  assign n23496 = ~x178 & n16044 ;
  assign n23497 = x178 & ~n16029 ;
  assign n23498 = ( x760 & n23496 ) | ( x760 & ~n23497 ) | ( n23496 & ~n23497 ) ;
  assign n23499 = ~n23496 & n23498 ;
  assign n23500 = ( x39 & n23495 ) | ( x39 & ~n23499 ) | ( n23495 & ~n23499 ) ;
  assign n23501 = n23500 ^ n23495 ^ 1'b0 ;
  assign n23502 = ( x39 & n23500 ) | ( x39 & ~n23501 ) | ( n23500 & ~n23501 ) ;
  assign n23503 = x178 & n15795 ;
  assign n23504 = x760 & ~n23503 ;
  assign n23505 = x178 | n15876 ;
  assign n23506 = n23504 & n23505 ;
  assign n23507 = x178 & n15943 ;
  assign n23508 = x178 | n16003 ;
  assign n23509 = ( x760 & ~n23507 ) | ( x760 & n23508 ) | ( ~n23507 & n23508 ) ;
  assign n23510 = ~x760 & n23509 ;
  assign n23511 = ( x39 & n23506 ) | ( x39 & ~n23510 ) | ( n23506 & ~n23510 ) ;
  assign n23512 = ~n23506 & n23511 ;
  assign n23513 = ( x38 & n23502 ) | ( x38 & ~n23512 ) | ( n23502 & ~n23512 ) ;
  assign n23514 = ~x38 & n23513 ;
  assign n23515 = ~x760 & n15591 ;
  assign n23516 = n17156 | n23515 ;
  assign n23517 = x178 & ~n5017 ;
  assign n23518 = n23516 & n23517 ;
  assign n23519 = x38 & ~n23518 ;
  assign n23520 = n23519 ^ x688 ^ 1'b0 ;
  assign n23521 = x760 | n15968 ;
  assign n23522 = n17889 & n23521 ;
  assign n23523 = x178 | n23522 ;
  assign n23524 = ( n23519 & ~n23520 ) | ( n23519 & n23523 ) | ( ~n23520 & n23523 ) ;
  assign n23525 = ( x688 & n23520 ) | ( x688 & n23524 ) | ( n23520 & n23524 ) ;
  assign n23526 = ( ~n2069 & n23514 ) | ( ~n2069 & n23525 ) | ( n23514 & n23525 ) ;
  assign n23527 = ~n2069 & n23526 ;
  assign n23528 = n23527 ^ n23491 ^ 1'b0 ;
  assign n23529 = ( n23491 & n23527 ) | ( n23491 & n23528 ) | ( n23527 & n23528 ) ;
  assign n23530 = ( n23433 & ~n23491 ) | ( n23433 & n23529 ) | ( ~n23491 & n23529 ) ;
  assign n23531 = x625 & ~n23530 ;
  assign n23532 = x625 | n23434 ;
  assign n23533 = ( x1153 & n23531 ) | ( x1153 & n23532 ) | ( n23531 & n23532 ) ;
  assign n23534 = ~n23531 & n23533 ;
  assign n23535 = ( x608 & n23387 ) | ( x608 & ~n23534 ) | ( n23387 & ~n23534 ) ;
  assign n23536 = ~n23387 & n23535 ;
  assign n23537 = x608 | n23383 ;
  assign n23538 = x625 & ~n23434 ;
  assign n23539 = x1153 | n23538 ;
  assign n23540 = ( n23530 & n23531 ) | ( n23530 & ~n23539 ) | ( n23531 & ~n23539 ) ;
  assign n23541 = ( ~n23536 & n23537 ) | ( ~n23536 & n23540 ) | ( n23537 & n23540 ) ;
  assign n23542 = ~n23536 & n23541 ;
  assign n23543 = n23530 ^ x778 ^ 1'b0 ;
  assign n23544 = ( n23530 & n23542 ) | ( n23530 & n23543 ) | ( n23542 & n23543 ) ;
  assign n23545 = x609 & ~n23544 ;
  assign n23546 = x609 | n23390 ;
  assign n23547 = ( x1155 & n23545 ) | ( x1155 & n23546 ) | ( n23545 & n23546 ) ;
  assign n23548 = ~n23545 & n23547 ;
  assign n23549 = ~x1155 & n23439 ;
  assign n23550 = ( x660 & n23548 ) | ( x660 & ~n23549 ) | ( n23548 & ~n23549 ) ;
  assign n23551 = ~n23548 & n23550 ;
  assign n23552 = x1155 & n23440 ;
  assign n23553 = x660 | n23552 ;
  assign n23554 = x609 & ~n23390 ;
  assign n23555 = x1155 | n23554 ;
  assign n23556 = ( n23544 & n23545 ) | ( n23544 & ~n23555 ) | ( n23545 & ~n23555 ) ;
  assign n23557 = ( ~n23551 & n23553 ) | ( ~n23551 & n23556 ) | ( n23553 & n23556 ) ;
  assign n23558 = ~n23551 & n23557 ;
  assign n23559 = n23544 ^ x785 ^ 1'b0 ;
  assign n23560 = ( n23544 & n23558 ) | ( n23544 & n23559 ) | ( n23558 & n23559 ) ;
  assign n23561 = x618 & ~n23560 ;
  assign n23562 = x618 | n23392 ;
  assign n23563 = ( x1154 & n23561 ) | ( x1154 & n23562 ) | ( n23561 & n23562 ) ;
  assign n23564 = ~n23561 & n23563 ;
  assign n23565 = ( x627 & n23451 ) | ( x627 & ~n23564 ) | ( n23451 & ~n23564 ) ;
  assign n23566 = ~n23451 & n23565 ;
  assign n23567 = x627 | n23448 ;
  assign n23568 = x618 & ~n23392 ;
  assign n23569 = x1154 | n23568 ;
  assign n23570 = ( n23560 & n23561 ) | ( n23560 & ~n23569 ) | ( n23561 & ~n23569 ) ;
  assign n23571 = ( ~n23566 & n23567 ) | ( ~n23566 & n23570 ) | ( n23567 & n23570 ) ;
  assign n23572 = ~n23566 & n23571 ;
  assign n23573 = n23560 ^ x781 ^ 1'b0 ;
  assign n23574 = ( n23560 & n23572 ) | ( n23560 & n23573 ) | ( n23572 & n23573 ) ;
  assign n23575 = x619 | n23574 ;
  assign n23576 = x619 & ~n23394 ;
  assign n23577 = ( x1159 & n23575 ) | ( x1159 & ~n23576 ) | ( n23575 & ~n23576 ) ;
  assign n23578 = ~x1159 & n23577 ;
  assign n23579 = ( x648 & n23458 ) | ( x648 & ~n23578 ) | ( n23458 & ~n23578 ) ;
  assign n23580 = n23578 | n23579 ;
  assign n23581 = x619 & ~n23574 ;
  assign n23582 = x619 | n23394 ;
  assign n23583 = ( x1159 & n23581 ) | ( x1159 & n23582 ) | ( n23581 & n23582 ) ;
  assign n23584 = ~n23581 & n23583 ;
  assign n23585 = ( x648 & n23461 ) | ( x648 & ~n23584 ) | ( n23461 & ~n23584 ) ;
  assign n23586 = ~n23461 & n23585 ;
  assign n23587 = x789 & ~n23586 ;
  assign n23588 = n23580 & n23587 ;
  assign n23589 = ~x789 & n23574 ;
  assign n23590 = ( n16519 & ~n23588 ) | ( n16519 & n23589 ) | ( ~n23588 & n23589 ) ;
  assign n23591 = n23588 | n23590 ;
  assign n23592 = n23402 ^ x629 ^ 1'b0 ;
  assign n23593 = ( n23402 & n23405 ) | ( n23402 & n23592 ) | ( n23405 & n23592 ) ;
  assign n23594 = n19046 & n23466 ;
  assign n23595 = ( x792 & n23593 ) | ( x792 & n23594 ) | ( n23593 & n23594 ) ;
  assign n23596 = n23594 ^ n23593 ^ 1'b0 ;
  assign n23597 = ( x792 & n23595 ) | ( x792 & n23596 ) | ( n23595 & n23596 ) ;
  assign n23598 = n16459 & ~n23396 ;
  assign n23599 = ~x626 & n23368 ;
  assign n23600 = x626 & n23464 ;
  assign n23601 = ( n22317 & n23599 ) | ( n22317 & ~n23600 ) | ( n23599 & ~n23600 ) ;
  assign n23602 = ~n23599 & n23601 ;
  assign n23603 = ~x626 & n23464 ;
  assign n23604 = x626 & n23368 ;
  assign n23605 = ( n22322 & n23603 ) | ( n22322 & ~n23604 ) | ( n23603 & ~n23604 ) ;
  assign n23606 = ~n23603 & n23605 ;
  assign n23607 = ( ~n23598 & n23602 ) | ( ~n23598 & n23606 ) | ( n23602 & n23606 ) ;
  assign n23608 = n23598 | n23607 ;
  assign n23609 = ( x788 & ~n22314 ) | ( x788 & n23608 ) | ( ~n22314 & n23608 ) ;
  assign n23610 = ( n18482 & n22314 ) | ( n18482 & n23609 ) | ( n22314 & n23609 ) ;
  assign n23611 = ~n23597 & n23610 ;
  assign n23612 = ( n23591 & n23597 ) | ( n23591 & ~n23611 ) | ( n23597 & ~n23611 ) ;
  assign n23613 = ( ~n18484 & n23490 ) | ( ~n18484 & n23612 ) | ( n23490 & n23612 ) ;
  assign n23614 = n23490 ^ n18484 ^ 1'b0 ;
  assign n23615 = ( n23490 & n23613 ) | ( n23490 & ~n23614 ) | ( n23613 & ~n23614 ) ;
  assign n23616 = x644 | n23473 ;
  assign n23617 = x644 & n23478 ;
  assign n23618 = x790 & ~n23617 ;
  assign n23619 = n23616 & n23618 ;
  assign n23620 = ( ~n23483 & n23615 ) | ( ~n23483 & n23619 ) | ( n23615 & n23619 ) ;
  assign n23621 = ~n23483 & n23620 ;
  assign n23622 = ( x57 & n5193 ) | ( x57 & ~n23621 ) | ( n5193 & ~n23621 ) ;
  assign n23623 = n23621 | n23622 ;
  assign n23624 = x178 | n1611 ;
  assign n23625 = ~n23515 & n23624 ;
  assign n23626 = n16397 | n23625 ;
  assign n23627 = ~n15662 & n23515 ;
  assign n23628 = ~x1155 & n23624 ;
  assign n23629 = ~n23627 & n23628 ;
  assign n23630 = ( x1155 & n23626 ) | ( x1155 & n23627 ) | ( n23626 & n23627 ) ;
  assign n23631 = n23629 | n23630 ;
  assign n23632 = n23626 ^ x785 ^ 1'b0 ;
  assign n23633 = ( n23626 & n23631 ) | ( n23626 & n23632 ) | ( n23631 & n23632 ) ;
  assign n23634 = n16411 | n23633 ;
  assign n23635 = x1154 & n23634 ;
  assign n23636 = n16414 | n23633 ;
  assign n23637 = ~x1154 & n23636 ;
  assign n23638 = n23635 | n23637 ;
  assign n23639 = n23633 ^ x781 ^ 1'b0 ;
  assign n23640 = ( n23633 & n23638 ) | ( n23633 & n23639 ) | ( n23638 & n23639 ) ;
  assign n23641 = n21437 | n23640 ;
  assign n23642 = x1159 & n23641 ;
  assign n23643 = n21440 | n23640 ;
  assign n23644 = ~x1159 & n23643 ;
  assign n23645 = n23642 | n23644 ;
  assign n23646 = n23640 ^ x789 ^ 1'b0 ;
  assign n23647 = ( n23640 & n23645 ) | ( n23640 & n23646 ) | ( n23645 & n23646 ) ;
  assign n23648 = n23624 ^ n16518 ^ 1'b0 ;
  assign n23649 = ( n23624 & n23647 ) | ( n23624 & ~n23648 ) | ( n23647 & ~n23648 ) ;
  assign n23650 = n23624 ^ n16339 ^ 1'b0 ;
  assign n23651 = ( n23624 & n23649 ) | ( n23624 & ~n23650 ) | ( n23649 & ~n23650 ) ;
  assign n23652 = n19055 & n23651 ;
  assign n23653 = x647 & ~n23624 ;
  assign n23654 = x1157 | n23653 ;
  assign n23655 = ~x688 & n15778 ;
  assign n23656 = ~x625 & n23655 ;
  assign n23657 = ~x1153 & n23624 ;
  assign n23658 = ~n23656 & n23657 ;
  assign n23659 = x778 & ~n23658 ;
  assign n23660 = n23624 & ~n23655 ;
  assign n23661 = ( x1153 & n23656 ) | ( x1153 & n23660 ) | ( n23656 & n23660 ) ;
  assign n23662 = n23659 & ~n23661 ;
  assign n23663 = ( x778 & n23660 ) | ( x778 & ~n23662 ) | ( n23660 & ~n23662 ) ;
  assign n23664 = ~n23662 & n23663 ;
  assign n23665 = n16447 | n23664 ;
  assign n23666 = n16449 | n23665 ;
  assign n23667 = n16451 | n23666 ;
  assign n23668 = n16530 | n23667 ;
  assign n23669 = n16560 | n23668 ;
  assign n23670 = ( x647 & ~n23654 ) | ( x647 & n23669 ) | ( ~n23654 & n23669 ) ;
  assign n23671 = ~n23654 & n23670 ;
  assign n23672 = n23624 ^ x647 ^ 1'b0 ;
  assign n23673 = ( n23624 & n23669 ) | ( n23624 & n23672 ) | ( n23669 & n23672 ) ;
  assign n23674 = x1157 & n23673 ;
  assign n23675 = ( n16375 & n23671 ) | ( n16375 & n23674 ) | ( n23671 & n23674 ) ;
  assign n23676 = ( x787 & n23652 ) | ( x787 & n23675 ) | ( n23652 & n23675 ) ;
  assign n23677 = n23675 ^ n23652 ^ 1'b0 ;
  assign n23678 = ( x787 & n23676 ) | ( x787 & n23677 ) | ( n23676 & n23677 ) ;
  assign n23679 = ~x626 & n23624 ;
  assign n23680 = x626 & n23647 ;
  assign n23681 = ( n22317 & n23679 ) | ( n22317 & ~n23680 ) | ( n23679 & ~n23680 ) ;
  assign n23682 = ~n23679 & n23681 ;
  assign n23683 = ~x626 & n23647 ;
  assign n23684 = x626 & n23624 ;
  assign n23685 = ( n22322 & n23683 ) | ( n22322 & ~n23684 ) | ( n23683 & ~n23684 ) ;
  assign n23686 = ~n23683 & n23685 ;
  assign n23687 = n23667 & ~n23686 ;
  assign n23688 = ( n16459 & n23686 ) | ( n16459 & ~n23687 ) | ( n23686 & ~n23687 ) ;
  assign n23689 = ( x788 & n23682 ) | ( x788 & n23688 ) | ( n23682 & n23688 ) ;
  assign n23690 = n23688 ^ n23682 ^ 1'b0 ;
  assign n23691 = ( x788 & n23689 ) | ( x788 & n23690 ) | ( n23689 & n23690 ) ;
  assign n23692 = n15524 | n23660 ;
  assign n23693 = n23625 & n23692 ;
  assign n23694 = x625 & ~n23692 ;
  assign n23695 = ( n23657 & n23693 ) | ( n23657 & n23694 ) | ( n23693 & n23694 ) ;
  assign n23696 = ( x608 & n23661 ) | ( x608 & ~n23695 ) | ( n23661 & ~n23695 ) ;
  assign n23697 = n23695 | n23696 ;
  assign n23698 = x1153 & n23625 ;
  assign n23699 = ~n23694 & n23698 ;
  assign n23700 = x608 & ~n23658 ;
  assign n23701 = n23697 & ~n23700 ;
  assign n23702 = ( n23697 & n23699 ) | ( n23697 & n23701 ) | ( n23699 & n23701 ) ;
  assign n23703 = n23693 ^ x778 ^ 1'b0 ;
  assign n23704 = ( n23693 & n23702 ) | ( n23693 & n23703 ) | ( n23702 & n23703 ) ;
  assign n23705 = x609 & ~n23704 ;
  assign n23711 = x609 | n23664 ;
  assign n23712 = ( x1155 & n23705 ) | ( x1155 & n23711 ) | ( n23705 & n23711 ) ;
  assign n23713 = ~n23705 & n23712 ;
  assign n23714 = ( x660 & n23629 ) | ( x660 & ~n23713 ) | ( n23629 & ~n23713 ) ;
  assign n23715 = ~n23629 & n23714 ;
  assign n23706 = x609 & ~n23664 ;
  assign n23707 = x1155 | n23706 ;
  assign n23708 = ( n23704 & n23705 ) | ( n23704 & ~n23707 ) | ( n23705 & ~n23707 ) ;
  assign n23709 = ( x660 & n23630 ) | ( x660 & ~n23708 ) | ( n23630 & ~n23708 ) ;
  assign n23710 = n23708 | n23709 ;
  assign n23716 = n23715 ^ n23710 ^ 1'b0 ;
  assign n23717 = ( x785 & ~n23710 ) | ( x785 & n23715 ) | ( ~n23710 & n23715 ) ;
  assign n23718 = ( x785 & ~n23716 ) | ( x785 & n23717 ) | ( ~n23716 & n23717 ) ;
  assign n23719 = ( x785 & n23704 ) | ( x785 & ~n23718 ) | ( n23704 & ~n23718 ) ;
  assign n23720 = ~n23718 & n23719 ;
  assign n23721 = x618 & ~n23720 ;
  assign n23722 = x618 | n23665 ;
  assign n23723 = ( x1154 & n23721 ) | ( x1154 & n23722 ) | ( n23721 & n23722 ) ;
  assign n23724 = ~n23721 & n23723 ;
  assign n23725 = ( x627 & n23637 ) | ( x627 & ~n23724 ) | ( n23637 & ~n23724 ) ;
  assign n23726 = ~n23637 & n23725 ;
  assign n23727 = x627 | n23635 ;
  assign n23728 = x618 & ~n23665 ;
  assign n23729 = x1154 | n23728 ;
  assign n23730 = ( n23720 & n23721 ) | ( n23720 & ~n23729 ) | ( n23721 & ~n23729 ) ;
  assign n23731 = ( ~n23726 & n23727 ) | ( ~n23726 & n23730 ) | ( n23727 & n23730 ) ;
  assign n23732 = ~n23726 & n23731 ;
  assign n23733 = n23720 ^ x781 ^ 1'b0 ;
  assign n23734 = ( n23720 & n23732 ) | ( n23720 & n23733 ) | ( n23732 & n23733 ) ;
  assign n23735 = ~x789 & n23734 ;
  assign n23736 = x619 & ~n23666 ;
  assign n23737 = x1159 | n23736 ;
  assign n23738 = x619 & ~n23734 ;
  assign n23739 = ( n23734 & ~n23737 ) | ( n23734 & n23738 ) | ( ~n23737 & n23738 ) ;
  assign n23740 = ( x648 & n23642 ) | ( x648 & ~n23739 ) | ( n23642 & ~n23739 ) ;
  assign n23741 = n23739 | n23740 ;
  assign n23742 = x619 | n23666 ;
  assign n23743 = x1159 & ~n23738 ;
  assign n23744 = n23742 & n23743 ;
  assign n23745 = ( x648 & n23644 ) | ( x648 & ~n23744 ) | ( n23644 & ~n23744 ) ;
  assign n23746 = ~n23644 & n23745 ;
  assign n23747 = x789 & ~n23746 ;
  assign n23748 = n23741 & n23747 ;
  assign n23749 = ( n16519 & ~n23735 ) | ( n16519 & n23748 ) | ( ~n23735 & n23748 ) ;
  assign n23750 = n23735 | n23749 ;
  assign n23751 = n23750 ^ n23691 ^ 1'b0 ;
  assign n23752 = ( n23691 & n23750 ) | ( n23691 & n23751 ) | ( n23750 & n23751 ) ;
  assign n23753 = ( n18482 & ~n23691 ) | ( n18482 & n23752 ) | ( ~n23691 & n23752 ) ;
  assign n23754 = n19208 | n23668 ;
  assign n23755 = n16556 & ~n23649 ;
  assign n23756 = x629 & ~n23755 ;
  assign n23757 = n23754 & n23756 ;
  assign n23758 = n16557 & ~n23649 ;
  assign n23759 = n19212 & ~n23668 ;
  assign n23760 = n23758 | n23759 ;
  assign n23761 = ( x629 & ~n23757 ) | ( x629 & n23760 ) | ( ~n23757 & n23760 ) ;
  assign n23762 = ~n23757 & n23761 ;
  assign n23763 = ( x792 & ~n19206 ) | ( x792 & n23762 ) | ( ~n19206 & n23762 ) ;
  assign n23764 = ( n18484 & n19206 ) | ( n18484 & n23763 ) | ( n19206 & n23763 ) ;
  assign n23765 = ( n23678 & n23753 ) | ( n23678 & ~n23764 ) | ( n23753 & ~n23764 ) ;
  assign n23766 = n23765 ^ n23753 ^ 1'b0 ;
  assign n23767 = ( n23678 & n23765 ) | ( n23678 & ~n23766 ) | ( n23765 & ~n23766 ) ;
  assign n23768 = x790 | n23767 ;
  assign n23769 = x644 & ~n23767 ;
  assign n23770 = ( x787 & n23671 ) | ( x787 & ~n23674 ) | ( n23671 & ~n23674 ) ;
  assign n23771 = ~n23671 & n23770 ;
  assign n23772 = ( x787 & n23669 ) | ( x787 & ~n23771 ) | ( n23669 & ~n23771 ) ;
  assign n23773 = ~n23771 & n23772 ;
  assign n23774 = x644 | n23773 ;
  assign n23775 = ( x715 & n23769 ) | ( x715 & n23774 ) | ( n23769 & n23774 ) ;
  assign n23776 = ~n23769 & n23775 ;
  assign n23777 = x644 | n23624 ;
  assign n23778 = n23624 ^ n16376 ^ 1'b0 ;
  assign n23779 = ( n23624 & n23651 ) | ( n23624 & ~n23778 ) | ( n23651 & ~n23778 ) ;
  assign n23780 = x644 & ~n23779 ;
  assign n23781 = ( x715 & n23777 ) | ( x715 & ~n23780 ) | ( n23777 & ~n23780 ) ;
  assign n23782 = ~x715 & n23781 ;
  assign n23783 = ( x1160 & n23776 ) | ( x1160 & ~n23782 ) | ( n23776 & ~n23782 ) ;
  assign n23784 = ~n23776 & n23783 ;
  assign n23785 = x644 & ~n23624 ;
  assign n23786 = x715 & ~n23785 ;
  assign n23787 = ( n23779 & n23780 ) | ( n23779 & n23786 ) | ( n23780 & n23786 ) ;
  assign n23788 = x644 & ~n23773 ;
  assign n23789 = x715 | n23788 ;
  assign n23790 = ( n23767 & n23769 ) | ( n23767 & ~n23789 ) | ( n23769 & ~n23789 ) ;
  assign n23791 = ( x1160 & ~n23787 ) | ( x1160 & n23790 ) | ( ~n23787 & n23790 ) ;
  assign n23792 = n23787 | n23791 ;
  assign n23793 = x790 & ~n23792 ;
  assign n23794 = ( x790 & n23784 ) | ( x790 & n23793 ) | ( n23784 & n23793 ) ;
  assign n23795 = x832 & ~n23794 ;
  assign n23796 = n23768 & n23795 ;
  assign n23797 = ~x178 & n7318 ;
  assign n23798 = x832 | n23797 ;
  assign n23799 = ~n23796 & n23798 ;
  assign n23800 = ( n23623 & n23796 ) | ( n23623 & ~n23799 ) | ( n23796 & ~n23799 ) ;
  assign n23836 = x179 & n15795 ;
  assign n23837 = x39 & ~n23836 ;
  assign n23838 = x179 | n15876 ;
  assign n23839 = n23837 & n23838 ;
  assign n23840 = x179 | n16044 ;
  assign n23841 = x179 & n16029 ;
  assign n23842 = ( x39 & n23840 ) | ( x39 & ~n23841 ) | ( n23840 & ~n23841 ) ;
  assign n23843 = ~x39 & n23842 ;
  assign n23844 = ( ~x38 & n23839 ) | ( ~x38 & n23843 ) | ( n23839 & n23843 ) ;
  assign n23845 = ~x38 & n23844 ;
  assign n23846 = x179 | n15644 ;
  assign n23847 = n16659 & n23846 ;
  assign n23848 = ( x741 & n23845 ) | ( x741 & n23847 ) | ( n23845 & n23847 ) ;
  assign n23849 = n23847 ^ n23845 ^ 1'b0 ;
  assign n23850 = ( x741 & n23848 ) | ( x741 & n23849 ) | ( n23848 & n23849 ) ;
  assign n23851 = x179 | n17902 ;
  assign n23852 = x179 & n17910 ;
  assign n23853 = ( x741 & n23851 ) | ( x741 & ~n23852 ) | ( n23851 & ~n23852 ) ;
  assign n23854 = ~x741 & n23853 ;
  assign n23855 = ( x724 & ~n23850 ) | ( x724 & n23854 ) | ( ~n23850 & n23854 ) ;
  assign n23856 = n23850 | n23855 ;
  assign n23801 = x179 | x741 ;
  assign n23802 = ( n17839 & n17843 ) | ( n17839 & ~n23801 ) | ( n17843 & ~n23801 ) ;
  assign n23803 = ~n17839 & n23802 ;
  assign n23804 = ~x741 & n22572 ;
  assign n23805 = x179 & ~n23804 ;
  assign n23806 = ( n20040 & ~n23803 ) | ( n20040 & n23805 ) | ( ~n23803 & n23805 ) ;
  assign n23807 = n23803 | n23806 ;
  assign n23857 = x724 & ~n23807 ;
  assign n23858 = ( n2069 & n23856 ) | ( n2069 & ~n23857 ) | ( n23856 & ~n23857 ) ;
  assign n23859 = ~n2069 & n23858 ;
  assign n23860 = n23859 ^ x179 ^ 1'b0 ;
  assign n23861 = ( ~x179 & n2069 ) | ( ~x179 & n23860 ) | ( n2069 & n23860 ) ;
  assign n23862 = ( x179 & n23859 ) | ( x179 & n23861 ) | ( n23859 & n23861 ) ;
  assign n23863 = x625 & ~n23862 ;
  assign n23808 = n23807 ^ n2069 ^ 1'b0 ;
  assign n23809 = ( x179 & n23807 ) | ( x179 & n23808 ) | ( n23807 & n23808 ) ;
  assign n23864 = x625 | n23809 ;
  assign n23865 = ( x1153 & n23863 ) | ( x1153 & n23864 ) | ( n23863 & n23864 ) ;
  assign n23866 = ~n23863 & n23865 ;
  assign n23810 = x179 | n15656 ;
  assign n23867 = x625 & ~n23810 ;
  assign n23868 = x1153 | n23867 ;
  assign n23869 = n16185 & n23846 ;
  assign n23870 = ( x38 & x179 ) | ( x38 & n16700 ) | ( x179 & n16700 ) ;
  assign n23871 = ~n2069 & n23870 ;
  assign n23872 = ( x179 & n16697 ) | ( x179 & ~n23871 ) | ( n16697 & ~n23871 ) ;
  assign n23873 = ~n23871 & n23872 ;
  assign n23874 = ( x724 & ~n23869 ) | ( x724 & n23873 ) | ( ~n23869 & n23873 ) ;
  assign n23875 = n23869 | n23874 ;
  assign n23876 = n23875 ^ n23810 ^ 1'b0 ;
  assign n23877 = x724 | n2069 ;
  assign n23878 = ( n23810 & n23876 ) | ( n23810 & ~n23877 ) | ( n23876 & ~n23877 ) ;
  assign n23879 = ( n23875 & ~n23876 ) | ( n23875 & n23878 ) | ( ~n23876 & n23878 ) ;
  assign n23880 = ( x625 & ~n23868 ) | ( x625 & n23879 ) | ( ~n23868 & n23879 ) ;
  assign n23881 = ~n23868 & n23880 ;
  assign n23882 = ( x608 & n23866 ) | ( x608 & ~n23881 ) | ( n23866 & ~n23881 ) ;
  assign n23883 = ~n23866 & n23882 ;
  assign n23884 = x625 & ~n23879 ;
  assign n23885 = x625 | n23810 ;
  assign n23886 = ( x1153 & n23884 ) | ( x1153 & n23885 ) | ( n23884 & n23885 ) ;
  assign n23887 = ~n23884 & n23886 ;
  assign n23888 = x608 | n23887 ;
  assign n23889 = x625 & ~n23809 ;
  assign n23890 = x1153 | n23889 ;
  assign n23891 = ( n23862 & n23863 ) | ( n23862 & ~n23890 ) | ( n23863 & ~n23890 ) ;
  assign n23892 = ( ~n23883 & n23888 ) | ( ~n23883 & n23891 ) | ( n23888 & n23891 ) ;
  assign n23893 = ~n23883 & n23892 ;
  assign n23894 = n23862 ^ x778 ^ 1'b0 ;
  assign n23895 = ( n23862 & n23893 ) | ( n23862 & n23894 ) | ( n23893 & n23894 ) ;
  assign n23896 = x609 & ~n23895 ;
  assign n23897 = n23881 | n23887 ;
  assign n23898 = n23879 ^ x778 ^ 1'b0 ;
  assign n23899 = ( n23879 & n23897 ) | ( n23879 & n23898 ) | ( n23897 & n23898 ) ;
  assign n23900 = x609 | n23899 ;
  assign n23901 = ( x1155 & n23896 ) | ( x1155 & n23900 ) | ( n23896 & n23900 ) ;
  assign n23902 = ~n23896 & n23901 ;
  assign n23813 = ~n15659 & n23809 ;
  assign n23814 = x609 & n23813 ;
  assign n23815 = ~n15668 & n23810 ;
  assign n23816 = n23814 | n23815 ;
  assign n23811 = n23809 ^ n15659 ^ 1'b0 ;
  assign n23812 = ( n23809 & n23810 ) | ( n23809 & n23811 ) | ( n23810 & n23811 ) ;
  assign n23818 = n23816 ^ n23812 ^ n23810 ;
  assign n23903 = ~x1155 & n23818 ;
  assign n23904 = ( x660 & n23902 ) | ( x660 & ~n23903 ) | ( n23902 & ~n23903 ) ;
  assign n23905 = ~n23902 & n23904 ;
  assign n23906 = x1155 & n23816 ;
  assign n23907 = x660 | n23906 ;
  assign n23908 = x609 & ~n23899 ;
  assign n23909 = x1155 | n23908 ;
  assign n23910 = ( n23895 & n23896 ) | ( n23895 & ~n23909 ) | ( n23896 & ~n23909 ) ;
  assign n23911 = ( ~n23905 & n23907 ) | ( ~n23905 & n23910 ) | ( n23907 & n23910 ) ;
  assign n23912 = ~n23905 & n23911 ;
  assign n23913 = n23895 ^ x785 ^ 1'b0 ;
  assign n23914 = ( n23895 & n23912 ) | ( n23895 & n23913 ) | ( n23912 & n23913 ) ;
  assign n23915 = x618 & ~n23914 ;
  assign n23916 = n23810 ^ n16234 ^ 1'b0 ;
  assign n23917 = ( n23810 & n23899 ) | ( n23810 & ~n23916 ) | ( n23899 & ~n23916 ) ;
  assign n23918 = x618 | n23917 ;
  assign n23919 = ( x1154 & n23915 ) | ( x1154 & n23918 ) | ( n23915 & n23918 ) ;
  assign n23920 = ~n23915 & n23919 ;
  assign n23817 = n23816 ^ x1155 ^ 1'b0 ;
  assign n23819 = ( n23816 & ~n23817 ) | ( n23816 & n23818 ) | ( ~n23817 & n23818 ) ;
  assign n23820 = n23812 ^ x785 ^ 1'b0 ;
  assign n23821 = ( n23812 & n23819 ) | ( n23812 & n23820 ) | ( n23819 & n23820 ) ;
  assign n23822 = x618 & ~n23821 ;
  assign n23826 = x618 & ~n23810 ;
  assign n23827 = x1154 | n23826 ;
  assign n23828 = ( n23821 & n23822 ) | ( n23821 & ~n23827 ) | ( n23822 & ~n23827 ) ;
  assign n23921 = ( x627 & ~n23828 ) | ( x627 & n23920 ) | ( ~n23828 & n23920 ) ;
  assign n23922 = ~n23920 & n23921 ;
  assign n23823 = x618 | n23810 ;
  assign n23824 = ( x1154 & n23822 ) | ( x1154 & n23823 ) | ( n23822 & n23823 ) ;
  assign n23825 = ~n23822 & n23824 ;
  assign n23923 = x627 | n23825 ;
  assign n23924 = x618 & ~n23917 ;
  assign n23925 = x1154 | n23924 ;
  assign n23926 = ( n23914 & n23915 ) | ( n23914 & ~n23925 ) | ( n23915 & ~n23925 ) ;
  assign n23927 = ( ~n23922 & n23923 ) | ( ~n23922 & n23926 ) | ( n23923 & n23926 ) ;
  assign n23928 = ~n23922 & n23927 ;
  assign n23929 = n23914 ^ x781 ^ 1'b0 ;
  assign n23930 = ( n23914 & n23928 ) | ( n23914 & n23929 ) | ( n23928 & n23929 ) ;
  assign n23931 = x619 & ~n23930 ;
  assign n23932 = n23810 ^ n16254 ^ 1'b0 ;
  assign n23933 = ( n23810 & n23917 ) | ( n23810 & ~n23932 ) | ( n23917 & ~n23932 ) ;
  assign n23939 = x619 | n23933 ;
  assign n23940 = ( x1159 & n23931 ) | ( x1159 & n23939 ) | ( n23931 & n23939 ) ;
  assign n23941 = ~n23931 & n23940 ;
  assign n23829 = n23825 | n23828 ;
  assign n23830 = n23821 ^ x781 ^ 1'b0 ;
  assign n23831 = ( n23821 & n23829 ) | ( n23821 & n23830 ) | ( n23829 & n23830 ) ;
  assign n23832 = x619 & ~n23831 ;
  assign n23942 = x619 & ~n23810 ;
  assign n23943 = x1159 | n23942 ;
  assign n23944 = ( n23831 & n23832 ) | ( n23831 & ~n23943 ) | ( n23832 & ~n23943 ) ;
  assign n23945 = ( x648 & n23941 ) | ( x648 & ~n23944 ) | ( n23941 & ~n23944 ) ;
  assign n23946 = ~n23941 & n23945 ;
  assign n23833 = x619 | n23810 ;
  assign n23834 = ( x1159 & n23832 ) | ( x1159 & n23833 ) | ( n23832 & n23833 ) ;
  assign n23835 = ~n23832 & n23834 ;
  assign n23934 = x619 & ~n23933 ;
  assign n23935 = x1159 | n23934 ;
  assign n23936 = ( n23930 & n23931 ) | ( n23930 & ~n23935 ) | ( n23931 & ~n23935 ) ;
  assign n23937 = ( x648 & ~n23835 ) | ( x648 & n23936 ) | ( ~n23835 & n23936 ) ;
  assign n23938 = n23835 | n23937 ;
  assign n23947 = n23946 ^ n23938 ^ 1'b0 ;
  assign n23948 = ( x789 & ~n23938 ) | ( x789 & n23946 ) | ( ~n23938 & n23946 ) ;
  assign n23949 = ( x789 & ~n23947 ) | ( x789 & n23948 ) | ( ~n23947 & n23948 ) ;
  assign n23950 = ( x789 & n23930 ) | ( x789 & ~n23949 ) | ( n23930 & ~n23949 ) ;
  assign n23951 = ~n23949 & n23950 ;
  assign n23952 = ~x626 & n23951 ;
  assign n23953 = n23810 ^ n16279 ^ 1'b0 ;
  assign n23954 = ( n23810 & n23933 ) | ( n23810 & ~n23953 ) | ( n23933 & ~n23953 ) ;
  assign n23955 = x626 & n23954 ;
  assign n23956 = ( x641 & ~n23952 ) | ( x641 & n23955 ) | ( ~n23952 & n23955 ) ;
  assign n23957 = n23952 | n23956 ;
  assign n23958 = ~x626 & n23810 ;
  assign n23959 = n23835 | n23944 ;
  assign n23960 = n23831 ^ x789 ^ 1'b0 ;
  assign n23961 = ( n23831 & n23959 ) | ( n23831 & n23960 ) | ( n23959 & n23960 ) ;
  assign n23962 = x626 & n23961 ;
  assign n23963 = ( x641 & ~n23958 ) | ( x641 & n23962 ) | ( ~n23958 & n23962 ) ;
  assign n23964 = n23958 | n23963 ;
  assign n23965 = ~x626 & n23954 ;
  assign n23966 = x626 & n23951 ;
  assign n23967 = ( x641 & n23965 ) | ( x641 & ~n23966 ) | ( n23965 & ~n23966 ) ;
  assign n23968 = ~n23965 & n23967 ;
  assign n23969 = x1158 & ~n23968 ;
  assign n23970 = n23964 & n23969 ;
  assign n23971 = ~x626 & n23961 ;
  assign n23972 = x626 & n23810 ;
  assign n23973 = x641 & ~n23972 ;
  assign n23974 = n23973 ^ n23971 ^ 1'b0 ;
  assign n23975 = ( n23971 & n23973 ) | ( n23971 & n23974 ) | ( n23973 & n23974 ) ;
  assign n23976 = ( x1158 & ~n23971 ) | ( x1158 & n23975 ) | ( ~n23971 & n23975 ) ;
  assign n23977 = ~n23970 & n23976 ;
  assign n23978 = ( n23957 & n23970 ) | ( n23957 & ~n23977 ) | ( n23970 & ~n23977 ) ;
  assign n23979 = n23951 ^ x788 ^ 1'b0 ;
  assign n23980 = ( n23951 & n23978 ) | ( n23951 & n23979 ) | ( n23978 & n23979 ) ;
  assign n23981 = x628 & ~n23980 ;
  assign n23982 = n23810 ^ n16518 ^ 1'b0 ;
  assign n23983 = ( n23810 & n23961 ) | ( n23810 & ~n23982 ) | ( n23961 & ~n23982 ) ;
  assign n23984 = x628 | n23983 ;
  assign n23985 = ( x1156 & n23981 ) | ( x1156 & n23984 ) | ( n23981 & n23984 ) ;
  assign n23986 = ~n23981 & n23985 ;
  assign n23987 = x628 & ~n23810 ;
  assign n23988 = x1156 | n23987 ;
  assign n23989 = n23810 ^ n16318 ^ 1'b0 ;
  assign n23990 = ( n23810 & n23954 ) | ( n23810 & ~n23989 ) | ( n23954 & ~n23989 ) ;
  assign n23991 = x628 & ~n23990 ;
  assign n23992 = ( ~n23988 & n23990 ) | ( ~n23988 & n23991 ) | ( n23990 & n23991 ) ;
  assign n23993 = ( x629 & n23986 ) | ( x629 & ~n23992 ) | ( n23986 & ~n23992 ) ;
  assign n23994 = ~n23986 & n23993 ;
  assign n23995 = x628 | n23810 ;
  assign n23996 = ( x1156 & n23991 ) | ( x1156 & n23995 ) | ( n23991 & n23995 ) ;
  assign n23997 = ~n23991 & n23996 ;
  assign n23998 = x629 | n23997 ;
  assign n23999 = x628 & ~n23983 ;
  assign n24000 = x1156 | n23999 ;
  assign n24001 = ( n23980 & n23981 ) | ( n23980 & ~n24000 ) | ( n23981 & ~n24000 ) ;
  assign n24002 = ( ~n23994 & n23998 ) | ( ~n23994 & n24001 ) | ( n23998 & n24001 ) ;
  assign n24003 = ~n23994 & n24002 ;
  assign n24004 = n23980 ^ x792 ^ 1'b0 ;
  assign n24005 = ( n23980 & n24003 ) | ( n23980 & n24004 ) | ( n24003 & n24004 ) ;
  assign n24006 = x647 & ~n24005 ;
  assign n24007 = n23810 ^ n16339 ^ 1'b0 ;
  assign n24008 = ( n23810 & n23983 ) | ( n23810 & ~n24007 ) | ( n23983 & ~n24007 ) ;
  assign n24009 = x647 | n24008 ;
  assign n24010 = ( x1157 & n24006 ) | ( x1157 & n24009 ) | ( n24006 & n24009 ) ;
  assign n24011 = ~n24006 & n24010 ;
  assign n24012 = x647 & ~n23810 ;
  assign n24013 = x1157 | n24012 ;
  assign n24014 = n23992 | n23997 ;
  assign n24015 = n23990 ^ x792 ^ 1'b0 ;
  assign n24016 = ( n23990 & n24014 ) | ( n23990 & n24015 ) | ( n24014 & n24015 ) ;
  assign n24017 = x647 & ~n24016 ;
  assign n24018 = ( ~n24013 & n24016 ) | ( ~n24013 & n24017 ) | ( n24016 & n24017 ) ;
  assign n24019 = ( x630 & n24011 ) | ( x630 & ~n24018 ) | ( n24011 & ~n24018 ) ;
  assign n24020 = ~n24011 & n24019 ;
  assign n24021 = x647 | n23810 ;
  assign n24022 = ( x1157 & n24017 ) | ( x1157 & n24021 ) | ( n24017 & n24021 ) ;
  assign n24023 = ~n24017 & n24022 ;
  assign n24024 = x630 | n24023 ;
  assign n24025 = x647 & ~n24008 ;
  assign n24026 = x1157 | n24025 ;
  assign n24027 = ( n24005 & n24006 ) | ( n24005 & ~n24026 ) | ( n24006 & ~n24026 ) ;
  assign n24028 = ( ~n24020 & n24024 ) | ( ~n24020 & n24027 ) | ( n24024 & n24027 ) ;
  assign n24029 = ~n24020 & n24028 ;
  assign n24030 = n24005 ^ x787 ^ 1'b0 ;
  assign n24031 = ( n24005 & n24029 ) | ( n24005 & n24030 ) | ( n24029 & n24030 ) ;
  assign n24032 = x644 & ~n24031 ;
  assign n24033 = n24018 | n24023 ;
  assign n24034 = n24016 ^ x787 ^ 1'b0 ;
  assign n24035 = ( n24016 & n24033 ) | ( n24016 & n24034 ) | ( n24033 & n24034 ) ;
  assign n24036 = x644 | n24035 ;
  assign n24037 = ( x715 & n24032 ) | ( x715 & n24036 ) | ( n24032 & n24036 ) ;
  assign n24038 = ~n24032 & n24037 ;
  assign n24039 = x644 | n23810 ;
  assign n24040 = n23810 ^ n16376 ^ 1'b0 ;
  assign n24041 = ( n23810 & n24008 ) | ( n23810 & ~n24040 ) | ( n24008 & ~n24040 ) ;
  assign n24042 = x644 & ~n24041 ;
  assign n24043 = ( x715 & n24039 ) | ( x715 & ~n24042 ) | ( n24039 & ~n24042 ) ;
  assign n24044 = ~x715 & n24043 ;
  assign n24045 = ( x1160 & n24038 ) | ( x1160 & ~n24044 ) | ( n24038 & ~n24044 ) ;
  assign n24046 = ~n24038 & n24045 ;
  assign n24047 = x644 & ~n23810 ;
  assign n24048 = x715 & ~n24047 ;
  assign n24049 = ( n24041 & n24042 ) | ( n24041 & n24048 ) | ( n24042 & n24048 ) ;
  assign n24050 = x644 & ~n24035 ;
  assign n24051 = x715 | n24050 ;
  assign n24052 = ( n24031 & n24032 ) | ( n24031 & ~n24051 ) | ( n24032 & ~n24051 ) ;
  assign n24053 = ( x1160 & ~n24049 ) | ( x1160 & n24052 ) | ( ~n24049 & n24052 ) ;
  assign n24054 = n24049 | n24053 ;
  assign n24055 = ( x790 & n24046 ) | ( x790 & n24054 ) | ( n24046 & n24054 ) ;
  assign n24056 = ~n24046 & n24055 ;
  assign n24057 = ~x790 & n24031 ;
  assign n24058 = ( n7318 & ~n24056 ) | ( n7318 & n24057 ) | ( ~n24056 & n24057 ) ;
  assign n24059 = n24056 | n24058 ;
  assign n24060 = x179 | n1611 ;
  assign n24061 = ~x741 & n15591 ;
  assign n24062 = n24060 & ~n24061 ;
  assign n24063 = n16397 | n24062 ;
  assign n24064 = n16402 | n24062 ;
  assign n24065 = x1155 & n24064 ;
  assign n24066 = n16405 | n24063 ;
  assign n24067 = ~x1155 & n24066 ;
  assign n24068 = n24065 | n24067 ;
  assign n24069 = n24063 ^ x785 ^ 1'b0 ;
  assign n24070 = ( n24063 & n24068 ) | ( n24063 & n24069 ) | ( n24068 & n24069 ) ;
  assign n24071 = n16411 | n24070 ;
  assign n24072 = x1154 & n24071 ;
  assign n24073 = n16414 | n24070 ;
  assign n24074 = ~x1154 & n24073 ;
  assign n24075 = n24072 | n24074 ;
  assign n24076 = n24070 ^ x781 ^ 1'b0 ;
  assign n24077 = ( n24070 & n24075 ) | ( n24070 & n24076 ) | ( n24075 & n24076 ) ;
  assign n24078 = x619 & ~n24077 ;
  assign n24079 = x619 | n24060 ;
  assign n24080 = ( x1159 & n24078 ) | ( x1159 & n24079 ) | ( n24078 & n24079 ) ;
  assign n24081 = ~n24078 & n24080 ;
  assign n24082 = x619 & ~n24060 ;
  assign n24083 = x1159 | n24082 ;
  assign n24084 = ( n24077 & n24078 ) | ( n24077 & ~n24083 ) | ( n24078 & ~n24083 ) ;
  assign n24085 = n24081 | n24084 ;
  assign n24086 = n24077 ^ x789 ^ 1'b0 ;
  assign n24087 = ( n24077 & n24085 ) | ( n24077 & n24086 ) | ( n24085 & n24086 ) ;
  assign n24088 = n24060 ^ n16518 ^ 1'b0 ;
  assign n24089 = ( n24060 & n24087 ) | ( n24060 & ~n24088 ) | ( n24087 & ~n24088 ) ;
  assign n24090 = n24060 ^ n16339 ^ 1'b0 ;
  assign n24091 = ( n24060 & n24089 ) | ( n24060 & ~n24090 ) | ( n24089 & ~n24090 ) ;
  assign n24092 = n19055 & n24091 ;
  assign n24093 = x647 & ~n24060 ;
  assign n24094 = x1157 | n24093 ;
  assign n24095 = ~x724 & n15778 ;
  assign n24096 = n24060 & ~n24095 ;
  assign n24097 = ~x1153 & n24060 ;
  assign n24098 = ~x625 & n24095 ;
  assign n24099 = n24097 & ~n24098 ;
  assign n24100 = ( x1153 & n24096 ) | ( x1153 & n24098 ) | ( n24096 & n24098 ) ;
  assign n24101 = n24099 | n24100 ;
  assign n24102 = n24096 ^ x778 ^ 1'b0 ;
  assign n24103 = ( n24096 & n24101 ) | ( n24096 & n24102 ) | ( n24101 & n24102 ) ;
  assign n24104 = n16447 | n24103 ;
  assign n24105 = n16449 | n24104 ;
  assign n24106 = n16451 | n24105 ;
  assign n24107 = n16530 | n24106 ;
  assign n24108 = n16560 | n24107 ;
  assign n24109 = ( x647 & ~n24094 ) | ( x647 & n24108 ) | ( ~n24094 & n24108 ) ;
  assign n24110 = ~n24094 & n24109 ;
  assign n24111 = n24060 ^ x647 ^ 1'b0 ;
  assign n24112 = ( n24060 & n24108 ) | ( n24060 & n24111 ) | ( n24108 & n24111 ) ;
  assign n24113 = x1157 & n24112 ;
  assign n24114 = ( n16375 & n24110 ) | ( n16375 & n24113 ) | ( n24110 & n24113 ) ;
  assign n24115 = ( x787 & n24092 ) | ( x787 & n24114 ) | ( n24092 & n24114 ) ;
  assign n24116 = n24114 ^ n24092 ^ 1'b0 ;
  assign n24117 = ( x787 & n24115 ) | ( x787 & n24116 ) | ( n24115 & n24116 ) ;
  assign n24118 = ~x626 & n24060 ;
  assign n24119 = x626 & n24087 ;
  assign n24120 = ( n22317 & n24118 ) | ( n22317 & ~n24119 ) | ( n24118 & ~n24119 ) ;
  assign n24121 = ~n24118 & n24120 ;
  assign n24122 = ~x626 & n24087 ;
  assign n24123 = x626 & n24060 ;
  assign n24124 = ( n22322 & n24122 ) | ( n22322 & ~n24123 ) | ( n24122 & ~n24123 ) ;
  assign n24125 = ~n24122 & n24124 ;
  assign n24126 = n24106 & ~n24125 ;
  assign n24127 = ( n16459 & n24125 ) | ( n16459 & ~n24126 ) | ( n24125 & ~n24126 ) ;
  assign n24128 = ( x788 & n24121 ) | ( x788 & n24127 ) | ( n24121 & n24127 ) ;
  assign n24129 = n24127 ^ n24121 ^ 1'b0 ;
  assign n24130 = ( x788 & n24128 ) | ( x788 & n24129 ) | ( n24128 & n24129 ) ;
  assign n24131 = n15524 | n24096 ;
  assign n24132 = n24062 & n24131 ;
  assign n24133 = x625 & ~n24131 ;
  assign n24134 = ( n24097 & n24132 ) | ( n24097 & n24133 ) | ( n24132 & n24133 ) ;
  assign n24135 = ( x608 & n24100 ) | ( x608 & ~n24134 ) | ( n24100 & ~n24134 ) ;
  assign n24136 = n24134 | n24135 ;
  assign n24137 = x1153 & n24062 ;
  assign n24138 = ~n24133 & n24137 ;
  assign n24139 = x608 & ~n24099 ;
  assign n24140 = n24136 & ~n24139 ;
  assign n24141 = ( n24136 & n24138 ) | ( n24136 & n24140 ) | ( n24138 & n24140 ) ;
  assign n24142 = n24132 ^ x778 ^ 1'b0 ;
  assign n24143 = ( n24132 & n24141 ) | ( n24132 & n24142 ) | ( n24141 & n24142 ) ;
  assign n24144 = x609 & ~n24143 ;
  assign n24145 = x609 | n24103 ;
  assign n24146 = ( x1155 & n24144 ) | ( x1155 & n24145 ) | ( n24144 & n24145 ) ;
  assign n24147 = ~n24144 & n24146 ;
  assign n24148 = ( x660 & n24067 ) | ( x660 & ~n24147 ) | ( n24067 & ~n24147 ) ;
  assign n24149 = ~n24067 & n24148 ;
  assign n24150 = x660 | n24065 ;
  assign n24151 = x609 & ~n24103 ;
  assign n24152 = x1155 | n24151 ;
  assign n24153 = ( n24143 & n24144 ) | ( n24143 & ~n24152 ) | ( n24144 & ~n24152 ) ;
  assign n24154 = ( ~n24149 & n24150 ) | ( ~n24149 & n24153 ) | ( n24150 & n24153 ) ;
  assign n24155 = ~n24149 & n24154 ;
  assign n24156 = n24143 ^ x785 ^ 1'b0 ;
  assign n24157 = ( n24143 & n24155 ) | ( n24143 & n24156 ) | ( n24155 & n24156 ) ;
  assign n24158 = x618 & ~n24157 ;
  assign n24159 = x618 | n24104 ;
  assign n24160 = ( x1154 & n24158 ) | ( x1154 & n24159 ) | ( n24158 & n24159 ) ;
  assign n24161 = ~n24158 & n24160 ;
  assign n24162 = ( x627 & n24074 ) | ( x627 & ~n24161 ) | ( n24074 & ~n24161 ) ;
  assign n24163 = ~n24074 & n24162 ;
  assign n24164 = x627 | n24072 ;
  assign n24165 = x618 & ~n24104 ;
  assign n24166 = x1154 | n24165 ;
  assign n24167 = ( n24157 & n24158 ) | ( n24157 & ~n24166 ) | ( n24158 & ~n24166 ) ;
  assign n24168 = ( ~n24163 & n24164 ) | ( ~n24163 & n24167 ) | ( n24164 & n24167 ) ;
  assign n24169 = ~n24163 & n24168 ;
  assign n24170 = n24157 ^ x781 ^ 1'b0 ;
  assign n24171 = ( n24157 & n24169 ) | ( n24157 & n24170 ) | ( n24169 & n24170 ) ;
  assign n24172 = ~x789 & n24171 ;
  assign n24173 = x619 & ~n24105 ;
  assign n24174 = x1159 | n24173 ;
  assign n24175 = x619 & ~n24171 ;
  assign n24176 = ( n24171 & ~n24174 ) | ( n24171 & n24175 ) | ( ~n24174 & n24175 ) ;
  assign n24177 = ( x648 & n24081 ) | ( x648 & ~n24176 ) | ( n24081 & ~n24176 ) ;
  assign n24178 = n24176 | n24177 ;
  assign n24179 = x619 | n24105 ;
  assign n24180 = x1159 & ~n24175 ;
  assign n24181 = n24179 & n24180 ;
  assign n24182 = ( x648 & n24084 ) | ( x648 & ~n24181 ) | ( n24084 & ~n24181 ) ;
  assign n24183 = ~n24084 & n24182 ;
  assign n24184 = x789 & ~n24183 ;
  assign n24185 = n24178 & n24184 ;
  assign n24186 = ( n16519 & ~n24172 ) | ( n16519 & n24185 ) | ( ~n24172 & n24185 ) ;
  assign n24187 = n24172 | n24186 ;
  assign n24188 = n24187 ^ n24130 ^ 1'b0 ;
  assign n24189 = ( n24130 & n24187 ) | ( n24130 & n24188 ) | ( n24187 & n24188 ) ;
  assign n24190 = ( n18482 & ~n24130 ) | ( n18482 & n24189 ) | ( ~n24130 & n24189 ) ;
  assign n24191 = n19208 | n24107 ;
  assign n24192 = n16556 & ~n24089 ;
  assign n24193 = x629 & ~n24192 ;
  assign n24194 = n24191 & n24193 ;
  assign n24195 = n16557 & ~n24089 ;
  assign n24196 = n19212 & ~n24107 ;
  assign n24197 = n24195 | n24196 ;
  assign n24198 = ( x629 & ~n24194 ) | ( x629 & n24197 ) | ( ~n24194 & n24197 ) ;
  assign n24199 = ~n24194 & n24198 ;
  assign n24200 = ( x792 & ~n19206 ) | ( x792 & n24199 ) | ( ~n19206 & n24199 ) ;
  assign n24201 = ( n18484 & n19206 ) | ( n18484 & n24200 ) | ( n19206 & n24200 ) ;
  assign n24202 = ( n24117 & n24190 ) | ( n24117 & ~n24201 ) | ( n24190 & ~n24201 ) ;
  assign n24203 = n24202 ^ n24190 ^ 1'b0 ;
  assign n24204 = ( n24117 & n24202 ) | ( n24117 & ~n24203 ) | ( n24202 & ~n24203 ) ;
  assign n24205 = x790 | n24204 ;
  assign n24206 = x644 & ~n24204 ;
  assign n24207 = ( x787 & n24110 ) | ( x787 & ~n24113 ) | ( n24110 & ~n24113 ) ;
  assign n24208 = ~n24110 & n24207 ;
  assign n24209 = ( x787 & n24108 ) | ( x787 & ~n24208 ) | ( n24108 & ~n24208 ) ;
  assign n24210 = ~n24208 & n24209 ;
  assign n24211 = x644 | n24210 ;
  assign n24212 = ( x715 & n24206 ) | ( x715 & n24211 ) | ( n24206 & n24211 ) ;
  assign n24213 = ~n24206 & n24212 ;
  assign n24214 = x644 | n24060 ;
  assign n24215 = n24060 ^ n16376 ^ 1'b0 ;
  assign n24216 = ( n24060 & n24091 ) | ( n24060 & ~n24215 ) | ( n24091 & ~n24215 ) ;
  assign n24217 = x644 & ~n24216 ;
  assign n24218 = ( x715 & n24214 ) | ( x715 & ~n24217 ) | ( n24214 & ~n24217 ) ;
  assign n24219 = ~x715 & n24218 ;
  assign n24220 = ( x1160 & n24213 ) | ( x1160 & ~n24219 ) | ( n24213 & ~n24219 ) ;
  assign n24221 = ~n24213 & n24220 ;
  assign n24222 = x644 & ~n24060 ;
  assign n24223 = x715 & ~n24222 ;
  assign n24224 = ( n24216 & n24217 ) | ( n24216 & n24223 ) | ( n24217 & n24223 ) ;
  assign n24225 = x644 & ~n24210 ;
  assign n24226 = x715 | n24225 ;
  assign n24227 = ( n24204 & n24206 ) | ( n24204 & ~n24226 ) | ( n24206 & ~n24226 ) ;
  assign n24228 = ( x1160 & ~n24224 ) | ( x1160 & n24227 ) | ( ~n24224 & n24227 ) ;
  assign n24229 = n24224 | n24228 ;
  assign n24230 = x790 & ~n24229 ;
  assign n24231 = ( x790 & n24221 ) | ( x790 & n24230 ) | ( n24221 & n24230 ) ;
  assign n24232 = x832 & ~n24231 ;
  assign n24233 = n24205 & n24232 ;
  assign n24234 = ~x179 & n7318 ;
  assign n24235 = x832 | n24234 ;
  assign n24236 = ~n24233 & n24235 ;
  assign n24237 = ( n24059 & n24233 ) | ( n24059 & ~n24236 ) | ( n24233 & ~n24236 ) ;
  assign n24238 = x180 | n15656 ;
  assign n24239 = x702 | n2069 ;
  assign n24240 = ~n24238 & n24239 ;
  assign n24241 = ( x38 & x180 ) | ( x38 & n16700 ) | ( x180 & n16700 ) ;
  assign n24242 = ~n2069 & n24241 ;
  assign n24243 = ( x180 & n16697 ) | ( x180 & ~n24242 ) | ( n16697 & ~n24242 ) ;
  assign n24244 = ~n24242 & n24243 ;
  assign n24245 = x180 | n15644 ;
  assign n24246 = n16185 & n24245 ;
  assign n24247 = x702 | n24246 ;
  assign n24248 = ( ~n24240 & n24244 ) | ( ~n24240 & n24247 ) | ( n24244 & n24247 ) ;
  assign n24249 = ~n24240 & n24248 ;
  assign n24250 = x625 & ~n24249 ;
  assign n24251 = x625 | n24238 ;
  assign n24252 = ( x1153 & n24250 ) | ( x1153 & n24251 ) | ( n24250 & n24251 ) ;
  assign n24253 = ~n24250 & n24252 ;
  assign n24254 = x625 & ~n24238 ;
  assign n24255 = x1153 | n24254 ;
  assign n24256 = ( x625 & n24249 ) | ( x625 & ~n24255 ) | ( n24249 & ~n24255 ) ;
  assign n24257 = ~n24255 & n24256 ;
  assign n24258 = n24253 | n24257 ;
  assign n24259 = n24249 ^ x778 ^ 1'b0 ;
  assign n24260 = ( n24249 & n24258 ) | ( n24249 & n24259 ) | ( n24258 & n24259 ) ;
  assign n24261 = n24238 ^ n16234 ^ 1'b0 ;
  assign n24262 = ( n24238 & n24260 ) | ( n24238 & ~n24261 ) | ( n24260 & ~n24261 ) ;
  assign n24263 = n24238 ^ n16254 ^ 1'b0 ;
  assign n24264 = ( n24238 & n24262 ) | ( n24238 & ~n24263 ) | ( n24262 & ~n24263 ) ;
  assign n24265 = n24238 ^ n16279 ^ 1'b0 ;
  assign n24266 = ( n24238 & n24264 ) | ( n24238 & ~n24265 ) | ( n24264 & ~n24265 ) ;
  assign n24267 = n24238 ^ n16318 ^ 1'b0 ;
  assign n24268 = ( n24238 & n24266 ) | ( n24238 & ~n24267 ) | ( n24266 & ~n24267 ) ;
  assign n24269 = x628 & ~n24268 ;
  assign n24270 = x628 | n24238 ;
  assign n24271 = ( x1156 & n24269 ) | ( x1156 & n24270 ) | ( n24269 & n24270 ) ;
  assign n24272 = ~n24269 & n24271 ;
  assign n24273 = x628 & ~n24238 ;
  assign n24274 = x1156 | n24273 ;
  assign n24275 = ( n24268 & n24269 ) | ( n24268 & ~n24274 ) | ( n24269 & ~n24274 ) ;
  assign n24276 = n24272 | n24275 ;
  assign n24277 = n24268 ^ x792 ^ 1'b0 ;
  assign n24278 = ( n24268 & n24276 ) | ( n24268 & n24277 ) | ( n24276 & n24277 ) ;
  assign n24279 = n24238 ^ x647 ^ 1'b0 ;
  assign n24280 = ( n24238 & n24278 ) | ( n24238 & ~n24279 ) | ( n24278 & ~n24279 ) ;
  assign n24281 = ( n24238 & n24278 ) | ( n24238 & n24279 ) | ( n24278 & n24279 ) ;
  assign n24282 = n24280 ^ x1157 ^ 1'b0 ;
  assign n24283 = ( n24280 & n24281 ) | ( n24280 & n24282 ) | ( n24281 & n24282 ) ;
  assign n24284 = n24278 ^ x787 ^ 1'b0 ;
  assign n24285 = ( n24278 & n24283 ) | ( n24278 & n24284 ) | ( n24283 & n24284 ) ;
  assign n24286 = x644 & ~n24285 ;
  assign n24287 = x715 | n24286 ;
  assign n24288 = x644 & ~n24238 ;
  assign n24289 = x715 & ~n24288 ;
  assign n24290 = n24289 ^ x1160 ^ 1'b0 ;
  assign n24291 = x38 & n24245 ;
  assign n24292 = x753 & n15332 ;
  assign n24293 = x180 & ~n15638 ;
  assign n24294 = ( ~x39 & n24292 ) | ( ~x39 & n24293 ) | ( n24292 & n24293 ) ;
  assign n24295 = ~x39 & n24294 ;
  assign n24296 = n24295 ^ x180 ^ 1'b0 ;
  assign n24297 = ( ~x180 & x753 ) | ( ~x180 & n24296 ) | ( x753 & n24296 ) ;
  assign n24298 = ( x180 & n24295 ) | ( x180 & n24297 ) | ( n24295 & n24297 ) ;
  assign n24299 = n24297 ^ n24295 ^ x180 ;
  assign n24300 = ( n15587 & n24298 ) | ( n15587 & ~n24299 ) | ( n24298 & ~n24299 ) ;
  assign n24301 = x180 & ~n15631 ;
  assign n24302 = x753 & n15486 ;
  assign n24303 = ( x39 & n24301 ) | ( x39 & n24302 ) | ( n24301 & n24302 ) ;
  assign n24304 = n24302 ^ n24301 ^ 1'b0 ;
  assign n24305 = ( x39 & n24303 ) | ( x39 & n24304 ) | ( n24303 & n24304 ) ;
  assign n24306 = ( ~x38 & n24300 ) | ( ~x38 & n24305 ) | ( n24300 & n24305 ) ;
  assign n24307 = ~x38 & n24306 ;
  assign n24308 = ~x753 & n15646 ;
  assign n24309 = ~n24307 & n24308 ;
  assign n24310 = ( n24291 & n24307 ) | ( n24291 & ~n24309 ) | ( n24307 & ~n24309 ) ;
  assign n24311 = ~n2069 & n24310 ;
  assign n24312 = x180 & n2069 ;
  assign n24313 = n24311 | n24312 ;
  assign n24314 = n24238 ^ n15659 ^ 1'b0 ;
  assign n24315 = ( n24238 & n24313 ) | ( n24238 & ~n24314 ) | ( n24313 & ~n24314 ) ;
  assign n24316 = n15662 & n24238 ;
  assign n24317 = ( ~n15662 & n24311 ) | ( ~n15662 & n24312 ) | ( n24311 & n24312 ) ;
  assign n24318 = n24316 | n24317 ;
  assign n24319 = n24318 ^ n24315 ^ n24238 ;
  assign n24320 = n24319 ^ x1155 ^ 1'b0 ;
  assign n24321 = ( n24318 & n24319 ) | ( n24318 & ~n24320 ) | ( n24319 & ~n24320 ) ;
  assign n24322 = n24315 ^ x785 ^ 1'b0 ;
  assign n24323 = ( n24315 & n24321 ) | ( n24315 & n24322 ) | ( n24321 & n24322 ) ;
  assign n24324 = x618 & ~n24323 ;
  assign n24325 = x618 | n24238 ;
  assign n24326 = ( x1154 & n24324 ) | ( x1154 & n24325 ) | ( n24324 & n24325 ) ;
  assign n24327 = ~n24324 & n24326 ;
  assign n24328 = x618 & ~n24238 ;
  assign n24329 = x1154 | n24328 ;
  assign n24330 = ( n24323 & n24324 ) | ( n24323 & ~n24329 ) | ( n24324 & ~n24329 ) ;
  assign n24331 = n24327 | n24330 ;
  assign n24332 = n24323 ^ x781 ^ 1'b0 ;
  assign n24333 = ( n24323 & n24331 ) | ( n24323 & n24332 ) | ( n24331 & n24332 ) ;
  assign n24334 = x619 & ~n24333 ;
  assign n24335 = x619 | n24238 ;
  assign n24336 = ( x1159 & n24334 ) | ( x1159 & n24335 ) | ( n24334 & n24335 ) ;
  assign n24337 = ~n24334 & n24336 ;
  assign n24338 = x619 & ~n24238 ;
  assign n24339 = x1159 | n24338 ;
  assign n24340 = ( n24333 & n24334 ) | ( n24333 & ~n24339 ) | ( n24334 & ~n24339 ) ;
  assign n24341 = n24337 | n24340 ;
  assign n24342 = n24333 ^ x789 ^ 1'b0 ;
  assign n24343 = ( n24333 & n24341 ) | ( n24333 & n24342 ) | ( n24341 & n24342 ) ;
  assign n24344 = n24238 ^ n16518 ^ 1'b0 ;
  assign n24345 = ( n24238 & n24343 ) | ( n24238 & ~n24344 ) | ( n24343 & ~n24344 ) ;
  assign n24346 = n24238 ^ n16339 ^ 1'b0 ;
  assign n24347 = ( n24238 & n24345 ) | ( n24238 & ~n24346 ) | ( n24345 & ~n24346 ) ;
  assign n24348 = n24238 ^ n16376 ^ 1'b0 ;
  assign n24349 = ( n24238 & n24347 ) | ( n24238 & ~n24348 ) | ( n24347 & ~n24348 ) ;
  assign n24350 = x644 | n24349 ;
  assign n24351 = ( n24289 & ~n24290 ) | ( n24289 & n24350 ) | ( ~n24290 & n24350 ) ;
  assign n24352 = ( x1160 & n24290 ) | ( x1160 & n24351 ) | ( n24290 & n24351 ) ;
  assign n24353 = n24287 & ~n24352 ;
  assign n24354 = x644 & ~n24349 ;
  assign n24355 = ( ~x715 & n24238 ) | ( ~x715 & n24288 ) | ( n24238 & n24288 ) ;
  assign n24356 = x1160 & ~n24355 ;
  assign n24357 = ( x1160 & n24354 ) | ( x1160 & n24356 ) | ( n24354 & n24356 ) ;
  assign n24358 = ( x715 & n24285 ) | ( x715 & n24286 ) | ( n24285 & n24286 ) ;
  assign n24359 = n24357 & ~n24358 ;
  assign n24360 = ( x790 & n24353 ) | ( x790 & n24359 ) | ( n24353 & n24359 ) ;
  assign n24361 = n24359 ^ n24353 ^ 1'b0 ;
  assign n24362 = ( x790 & n24360 ) | ( x790 & n24361 ) | ( n24360 & n24361 ) ;
  assign n24363 = n19055 & n24347 ;
  assign n24364 = n16374 & n24280 ;
  assign n24365 = n16373 & n24281 ;
  assign n24366 = n24364 | n24365 ;
  assign n24367 = ( x787 & n24363 ) | ( x787 & n24366 ) | ( n24363 & n24366 ) ;
  assign n24368 = n24366 ^ n24363 ^ 1'b0 ;
  assign n24369 = ( x787 & n24367 ) | ( x787 & n24368 ) | ( n24367 & n24368 ) ;
  assign n24370 = x702 & ~n24310 ;
  assign n24371 = x180 & ~n16054 ;
  assign n24372 = ~x180 & n16048 ;
  assign n24373 = ( x753 & ~n24371 ) | ( x753 & n24372 ) | ( ~n24371 & n24372 ) ;
  assign n24374 = n24371 | n24373 ;
  assign n24375 = ~x180 & n16044 ;
  assign n24376 = x180 & ~n16029 ;
  assign n24377 = ( x753 & n24375 ) | ( x753 & ~n24376 ) | ( n24375 & ~n24376 ) ;
  assign n24378 = ~n24375 & n24377 ;
  assign n24379 = ( x39 & n24374 ) | ( x39 & ~n24378 ) | ( n24374 & ~n24378 ) ;
  assign n24380 = n24379 ^ n24374 ^ 1'b0 ;
  assign n24381 = ( x39 & n24379 ) | ( x39 & ~n24380 ) | ( n24379 & ~n24380 ) ;
  assign n24382 = x180 & n15795 ;
  assign n24383 = x753 & ~n24382 ;
  assign n24384 = x180 | n15876 ;
  assign n24385 = n24383 & n24384 ;
  assign n24386 = x180 & n15943 ;
  assign n24387 = x180 | n16003 ;
  assign n24388 = ( x753 & ~n24386 ) | ( x753 & n24387 ) | ( ~n24386 & n24387 ) ;
  assign n24389 = ~x753 & n24388 ;
  assign n24390 = ( x39 & n24385 ) | ( x39 & ~n24389 ) | ( n24385 & ~n24389 ) ;
  assign n24391 = ~n24385 & n24390 ;
  assign n24392 = ( x38 & n24381 ) | ( x38 & ~n24391 ) | ( n24381 & ~n24391 ) ;
  assign n24393 = ~x38 & n24392 ;
  assign n24394 = ~x753 & n15591 ;
  assign n24395 = n17156 | n24394 ;
  assign n24396 = x180 & ~n5017 ;
  assign n24397 = n24395 & n24396 ;
  assign n24398 = x38 & ~n24397 ;
  assign n24399 = n24398 ^ x702 ^ 1'b0 ;
  assign n24400 = x753 | n15968 ;
  assign n24401 = n17889 & n24400 ;
  assign n24402 = x180 | n24401 ;
  assign n24403 = ( n24398 & ~n24399 ) | ( n24398 & n24402 ) | ( ~n24399 & n24402 ) ;
  assign n24404 = ( x702 & n24399 ) | ( x702 & n24403 ) | ( n24399 & n24403 ) ;
  assign n24405 = ( ~n2069 & n24393 ) | ( ~n2069 & n24404 ) | ( n24393 & n24404 ) ;
  assign n24406 = ~n2069 & n24405 ;
  assign n24407 = n24406 ^ n24370 ^ 1'b0 ;
  assign n24408 = ( n24370 & n24406 ) | ( n24370 & n24407 ) | ( n24406 & n24407 ) ;
  assign n24409 = ( n24312 & ~n24370 ) | ( n24312 & n24408 ) | ( ~n24370 & n24408 ) ;
  assign n24410 = x625 & ~n24409 ;
  assign n24411 = x625 | n24313 ;
  assign n24412 = ( x1153 & n24410 ) | ( x1153 & n24411 ) | ( n24410 & n24411 ) ;
  assign n24413 = ~n24410 & n24412 ;
  assign n24414 = ( x608 & n24257 ) | ( x608 & ~n24413 ) | ( n24257 & ~n24413 ) ;
  assign n24415 = ~n24257 & n24414 ;
  assign n24416 = x608 | n24253 ;
  assign n24417 = x625 & ~n24313 ;
  assign n24418 = x1153 | n24417 ;
  assign n24419 = ( n24409 & n24410 ) | ( n24409 & ~n24418 ) | ( n24410 & ~n24418 ) ;
  assign n24420 = ( ~n24415 & n24416 ) | ( ~n24415 & n24419 ) | ( n24416 & n24419 ) ;
  assign n24421 = ~n24415 & n24420 ;
  assign n24422 = n24409 ^ x778 ^ 1'b0 ;
  assign n24423 = ( n24409 & n24421 ) | ( n24409 & n24422 ) | ( n24421 & n24422 ) ;
  assign n24424 = x609 & ~n24423 ;
  assign n24425 = x609 | n24260 ;
  assign n24426 = ( x1155 & n24424 ) | ( x1155 & n24425 ) | ( n24424 & n24425 ) ;
  assign n24427 = ~n24424 & n24426 ;
  assign n24428 = ~x1155 & n24318 ;
  assign n24429 = ( x660 & n24427 ) | ( x660 & ~n24428 ) | ( n24427 & ~n24428 ) ;
  assign n24430 = ~n24427 & n24429 ;
  assign n24431 = x1155 & n24319 ;
  assign n24432 = x660 | n24431 ;
  assign n24433 = x609 & ~n24260 ;
  assign n24434 = x1155 | n24433 ;
  assign n24435 = ( n24423 & n24424 ) | ( n24423 & ~n24434 ) | ( n24424 & ~n24434 ) ;
  assign n24436 = ( ~n24430 & n24432 ) | ( ~n24430 & n24435 ) | ( n24432 & n24435 ) ;
  assign n24437 = ~n24430 & n24436 ;
  assign n24438 = n24423 ^ x785 ^ 1'b0 ;
  assign n24439 = ( n24423 & n24437 ) | ( n24423 & n24438 ) | ( n24437 & n24438 ) ;
  assign n24440 = x618 & ~n24439 ;
  assign n24441 = x618 | n24262 ;
  assign n24442 = ( x1154 & n24440 ) | ( x1154 & n24441 ) | ( n24440 & n24441 ) ;
  assign n24443 = ~n24440 & n24442 ;
  assign n24444 = ( x627 & n24330 ) | ( x627 & ~n24443 ) | ( n24330 & ~n24443 ) ;
  assign n24445 = ~n24330 & n24444 ;
  assign n24446 = x627 | n24327 ;
  assign n24447 = x618 & ~n24262 ;
  assign n24448 = x1154 | n24447 ;
  assign n24449 = ( n24439 & n24440 ) | ( n24439 & ~n24448 ) | ( n24440 & ~n24448 ) ;
  assign n24450 = ( ~n24445 & n24446 ) | ( ~n24445 & n24449 ) | ( n24446 & n24449 ) ;
  assign n24451 = ~n24445 & n24450 ;
  assign n24452 = n24439 ^ x781 ^ 1'b0 ;
  assign n24453 = ( n24439 & n24451 ) | ( n24439 & n24452 ) | ( n24451 & n24452 ) ;
  assign n24454 = x619 | n24453 ;
  assign n24455 = x619 & ~n24264 ;
  assign n24456 = ( x1159 & n24454 ) | ( x1159 & ~n24455 ) | ( n24454 & ~n24455 ) ;
  assign n24457 = ~x1159 & n24456 ;
  assign n24458 = ( x648 & n24337 ) | ( x648 & ~n24457 ) | ( n24337 & ~n24457 ) ;
  assign n24459 = n24457 | n24458 ;
  assign n24460 = x619 & ~n24453 ;
  assign n24461 = x619 | n24264 ;
  assign n24462 = ( x1159 & n24460 ) | ( x1159 & n24461 ) | ( n24460 & n24461 ) ;
  assign n24463 = ~n24460 & n24462 ;
  assign n24464 = ( x648 & n24340 ) | ( x648 & ~n24463 ) | ( n24340 & ~n24463 ) ;
  assign n24465 = ~n24340 & n24464 ;
  assign n24466 = x789 & ~n24465 ;
  assign n24467 = n24459 & n24466 ;
  assign n24468 = ~x789 & n24453 ;
  assign n24469 = ( n16519 & ~n24467 ) | ( n16519 & n24468 ) | ( ~n24467 & n24468 ) ;
  assign n24470 = n24467 | n24469 ;
  assign n24471 = n24272 ^ x629 ^ 1'b0 ;
  assign n24472 = ( n24272 & n24275 ) | ( n24272 & n24471 ) | ( n24275 & n24471 ) ;
  assign n24473 = n19046 & n24345 ;
  assign n24474 = ( x792 & n24472 ) | ( x792 & n24473 ) | ( n24472 & n24473 ) ;
  assign n24475 = n24473 ^ n24472 ^ 1'b0 ;
  assign n24476 = ( x792 & n24474 ) | ( x792 & n24475 ) | ( n24474 & n24475 ) ;
  assign n24477 = n16459 & ~n24266 ;
  assign n24478 = ~x626 & n24238 ;
  assign n24479 = x626 & n24343 ;
  assign n24480 = ( n22317 & n24478 ) | ( n22317 & ~n24479 ) | ( n24478 & ~n24479 ) ;
  assign n24481 = ~n24478 & n24480 ;
  assign n24482 = ~x626 & n24343 ;
  assign n24483 = x626 & n24238 ;
  assign n24484 = ( n22322 & n24482 ) | ( n22322 & ~n24483 ) | ( n24482 & ~n24483 ) ;
  assign n24485 = ~n24482 & n24484 ;
  assign n24486 = ( ~n24477 & n24481 ) | ( ~n24477 & n24485 ) | ( n24481 & n24485 ) ;
  assign n24487 = n24477 | n24486 ;
  assign n24488 = ( x788 & ~n22314 ) | ( x788 & n24487 ) | ( ~n22314 & n24487 ) ;
  assign n24489 = ( n18482 & n22314 ) | ( n18482 & n24488 ) | ( n22314 & n24488 ) ;
  assign n24490 = ~n24476 & n24489 ;
  assign n24491 = ( n24470 & n24476 ) | ( n24470 & ~n24490 ) | ( n24476 & ~n24490 ) ;
  assign n24492 = ( ~n18484 & n24369 ) | ( ~n18484 & n24491 ) | ( n24369 & n24491 ) ;
  assign n24493 = n24369 ^ n18484 ^ 1'b0 ;
  assign n24494 = ( n24369 & n24492 ) | ( n24369 & ~n24493 ) | ( n24492 & ~n24493 ) ;
  assign n24495 = x644 | n24352 ;
  assign n24496 = x644 & n24357 ;
  assign n24497 = x790 & ~n24496 ;
  assign n24498 = n24495 & n24497 ;
  assign n24499 = ( ~n24362 & n24494 ) | ( ~n24362 & n24498 ) | ( n24494 & n24498 ) ;
  assign n24500 = ~n24362 & n24499 ;
  assign n24501 = ( x57 & n5193 ) | ( x57 & ~n24500 ) | ( n5193 & ~n24500 ) ;
  assign n24502 = n24500 | n24501 ;
  assign n24503 = x180 | n1611 ;
  assign n24504 = ~n24394 & n24503 ;
  assign n24505 = n16397 | n24504 ;
  assign n24506 = ~n15662 & n24394 ;
  assign n24507 = ~x1155 & n24503 ;
  assign n24508 = ~n24506 & n24507 ;
  assign n24509 = ( x1155 & n24505 ) | ( x1155 & n24506 ) | ( n24505 & n24506 ) ;
  assign n24510 = n24508 | n24509 ;
  assign n24511 = n24505 ^ x785 ^ 1'b0 ;
  assign n24512 = ( n24505 & n24510 ) | ( n24505 & n24511 ) | ( n24510 & n24511 ) ;
  assign n24513 = n16411 | n24512 ;
  assign n24514 = x1154 & n24513 ;
  assign n24515 = n16414 | n24512 ;
  assign n24516 = ~x1154 & n24515 ;
  assign n24517 = n24514 | n24516 ;
  assign n24518 = n24512 ^ x781 ^ 1'b0 ;
  assign n24519 = ( n24512 & n24517 ) | ( n24512 & n24518 ) | ( n24517 & n24518 ) ;
  assign n24520 = n21437 | n24519 ;
  assign n24521 = x1159 & n24520 ;
  assign n24522 = n21440 | n24519 ;
  assign n24523 = ~x1159 & n24522 ;
  assign n24524 = n24521 | n24523 ;
  assign n24525 = n24519 ^ x789 ^ 1'b0 ;
  assign n24526 = ( n24519 & n24524 ) | ( n24519 & n24525 ) | ( n24524 & n24525 ) ;
  assign n24527 = n24503 ^ n16518 ^ 1'b0 ;
  assign n24528 = ( n24503 & n24526 ) | ( n24503 & ~n24527 ) | ( n24526 & ~n24527 ) ;
  assign n24529 = n24503 ^ n16339 ^ 1'b0 ;
  assign n24530 = ( n24503 & n24528 ) | ( n24503 & ~n24529 ) | ( n24528 & ~n24529 ) ;
  assign n24531 = n19055 & n24530 ;
  assign n24532 = x647 & ~n24503 ;
  assign n24533 = x1157 | n24532 ;
  assign n24534 = ~x702 & n15778 ;
  assign n24535 = ~x625 & n24534 ;
  assign n24536 = ~x1153 & n24503 ;
  assign n24537 = ~n24535 & n24536 ;
  assign n24538 = x778 & ~n24537 ;
  assign n24539 = n24503 & ~n24534 ;
  assign n24540 = ( x1153 & n24535 ) | ( x1153 & n24539 ) | ( n24535 & n24539 ) ;
  assign n24541 = n24538 & ~n24540 ;
  assign n24542 = ( x778 & n24539 ) | ( x778 & ~n24541 ) | ( n24539 & ~n24541 ) ;
  assign n24543 = ~n24541 & n24542 ;
  assign n24544 = n16447 | n24543 ;
  assign n24545 = n16449 | n24544 ;
  assign n24546 = n16451 | n24545 ;
  assign n24547 = n16530 | n24546 ;
  assign n24548 = n16560 | n24547 ;
  assign n24549 = ( x647 & ~n24533 ) | ( x647 & n24548 ) | ( ~n24533 & n24548 ) ;
  assign n24550 = ~n24533 & n24549 ;
  assign n24551 = n24503 ^ x647 ^ 1'b0 ;
  assign n24552 = ( n24503 & n24548 ) | ( n24503 & n24551 ) | ( n24548 & n24551 ) ;
  assign n24553 = x1157 & n24552 ;
  assign n24554 = ( n16375 & n24550 ) | ( n16375 & n24553 ) | ( n24550 & n24553 ) ;
  assign n24555 = ( x787 & n24531 ) | ( x787 & n24554 ) | ( n24531 & n24554 ) ;
  assign n24556 = n24554 ^ n24531 ^ 1'b0 ;
  assign n24557 = ( x787 & n24555 ) | ( x787 & n24556 ) | ( n24555 & n24556 ) ;
  assign n24558 = ~x626 & n24503 ;
  assign n24559 = x626 & n24526 ;
  assign n24560 = ( n22317 & n24558 ) | ( n22317 & ~n24559 ) | ( n24558 & ~n24559 ) ;
  assign n24561 = ~n24558 & n24560 ;
  assign n24562 = ~x626 & n24526 ;
  assign n24563 = x626 & n24503 ;
  assign n24564 = ( n22322 & n24562 ) | ( n22322 & ~n24563 ) | ( n24562 & ~n24563 ) ;
  assign n24565 = ~n24562 & n24564 ;
  assign n24566 = n24546 & ~n24565 ;
  assign n24567 = ( n16459 & n24565 ) | ( n16459 & ~n24566 ) | ( n24565 & ~n24566 ) ;
  assign n24568 = ( x788 & n24561 ) | ( x788 & n24567 ) | ( n24561 & n24567 ) ;
  assign n24569 = n24567 ^ n24561 ^ 1'b0 ;
  assign n24570 = ( x788 & n24568 ) | ( x788 & n24569 ) | ( n24568 & n24569 ) ;
  assign n24571 = n15524 | n24539 ;
  assign n24572 = n24504 & n24571 ;
  assign n24573 = x625 & ~n24571 ;
  assign n24574 = ( n24536 & n24572 ) | ( n24536 & n24573 ) | ( n24572 & n24573 ) ;
  assign n24575 = ( x608 & n24540 ) | ( x608 & ~n24574 ) | ( n24540 & ~n24574 ) ;
  assign n24576 = n24574 | n24575 ;
  assign n24577 = x1153 & n24504 ;
  assign n24578 = ~n24573 & n24577 ;
  assign n24579 = x608 & ~n24537 ;
  assign n24580 = n24576 & ~n24579 ;
  assign n24581 = ( n24576 & n24578 ) | ( n24576 & n24580 ) | ( n24578 & n24580 ) ;
  assign n24582 = n24572 ^ x778 ^ 1'b0 ;
  assign n24583 = ( n24572 & n24581 ) | ( n24572 & n24582 ) | ( n24581 & n24582 ) ;
  assign n24584 = x609 & ~n24583 ;
  assign n24590 = x609 | n24543 ;
  assign n24591 = ( x1155 & n24584 ) | ( x1155 & n24590 ) | ( n24584 & n24590 ) ;
  assign n24592 = ~n24584 & n24591 ;
  assign n24593 = ( x660 & n24508 ) | ( x660 & ~n24592 ) | ( n24508 & ~n24592 ) ;
  assign n24594 = ~n24508 & n24593 ;
  assign n24585 = x609 & ~n24543 ;
  assign n24586 = x1155 | n24585 ;
  assign n24587 = ( n24583 & n24584 ) | ( n24583 & ~n24586 ) | ( n24584 & ~n24586 ) ;
  assign n24588 = ( x660 & n24509 ) | ( x660 & ~n24587 ) | ( n24509 & ~n24587 ) ;
  assign n24589 = n24587 | n24588 ;
  assign n24595 = n24594 ^ n24589 ^ 1'b0 ;
  assign n24596 = ( x785 & ~n24589 ) | ( x785 & n24594 ) | ( ~n24589 & n24594 ) ;
  assign n24597 = ( x785 & ~n24595 ) | ( x785 & n24596 ) | ( ~n24595 & n24596 ) ;
  assign n24598 = ( x785 & n24583 ) | ( x785 & ~n24597 ) | ( n24583 & ~n24597 ) ;
  assign n24599 = ~n24597 & n24598 ;
  assign n24600 = x618 & ~n24599 ;
  assign n24601 = x618 | n24544 ;
  assign n24602 = ( x1154 & n24600 ) | ( x1154 & n24601 ) | ( n24600 & n24601 ) ;
  assign n24603 = ~n24600 & n24602 ;
  assign n24604 = ( x627 & n24516 ) | ( x627 & ~n24603 ) | ( n24516 & ~n24603 ) ;
  assign n24605 = ~n24516 & n24604 ;
  assign n24606 = x627 | n24514 ;
  assign n24607 = x618 & ~n24544 ;
  assign n24608 = x1154 | n24607 ;
  assign n24609 = ( n24599 & n24600 ) | ( n24599 & ~n24608 ) | ( n24600 & ~n24608 ) ;
  assign n24610 = ( ~n24605 & n24606 ) | ( ~n24605 & n24609 ) | ( n24606 & n24609 ) ;
  assign n24611 = ~n24605 & n24610 ;
  assign n24612 = n24599 ^ x781 ^ 1'b0 ;
  assign n24613 = ( n24599 & n24611 ) | ( n24599 & n24612 ) | ( n24611 & n24612 ) ;
  assign n24614 = ~x789 & n24613 ;
  assign n24615 = x619 & ~n24545 ;
  assign n24616 = x1159 | n24615 ;
  assign n24617 = x619 & ~n24613 ;
  assign n24618 = ( n24613 & ~n24616 ) | ( n24613 & n24617 ) | ( ~n24616 & n24617 ) ;
  assign n24619 = ( x648 & n24521 ) | ( x648 & ~n24618 ) | ( n24521 & ~n24618 ) ;
  assign n24620 = n24618 | n24619 ;
  assign n24621 = x619 | n24545 ;
  assign n24622 = x1159 & ~n24617 ;
  assign n24623 = n24621 & n24622 ;
  assign n24624 = ( x648 & n24523 ) | ( x648 & ~n24623 ) | ( n24523 & ~n24623 ) ;
  assign n24625 = ~n24523 & n24624 ;
  assign n24626 = x789 & ~n24625 ;
  assign n24627 = n24620 & n24626 ;
  assign n24628 = ( n16519 & ~n24614 ) | ( n16519 & n24627 ) | ( ~n24614 & n24627 ) ;
  assign n24629 = n24614 | n24628 ;
  assign n24630 = n24629 ^ n24570 ^ 1'b0 ;
  assign n24631 = ( n24570 & n24629 ) | ( n24570 & n24630 ) | ( n24629 & n24630 ) ;
  assign n24632 = ( n18482 & ~n24570 ) | ( n18482 & n24631 ) | ( ~n24570 & n24631 ) ;
  assign n24633 = n19208 | n24547 ;
  assign n24634 = n16556 & ~n24528 ;
  assign n24635 = x629 & ~n24634 ;
  assign n24636 = n24633 & n24635 ;
  assign n24637 = n16557 & ~n24528 ;
  assign n24638 = n19212 & ~n24547 ;
  assign n24639 = n24637 | n24638 ;
  assign n24640 = ( x629 & ~n24636 ) | ( x629 & n24639 ) | ( ~n24636 & n24639 ) ;
  assign n24641 = ~n24636 & n24640 ;
  assign n24642 = ( x792 & ~n19206 ) | ( x792 & n24641 ) | ( ~n19206 & n24641 ) ;
  assign n24643 = ( n18484 & n19206 ) | ( n18484 & n24642 ) | ( n19206 & n24642 ) ;
  assign n24644 = ( n24557 & n24632 ) | ( n24557 & ~n24643 ) | ( n24632 & ~n24643 ) ;
  assign n24645 = n24644 ^ n24632 ^ 1'b0 ;
  assign n24646 = ( n24557 & n24644 ) | ( n24557 & ~n24645 ) | ( n24644 & ~n24645 ) ;
  assign n24647 = x790 | n24646 ;
  assign n24648 = x644 & ~n24646 ;
  assign n24649 = ( x787 & n24550 ) | ( x787 & ~n24553 ) | ( n24550 & ~n24553 ) ;
  assign n24650 = ~n24550 & n24649 ;
  assign n24651 = ( x787 & n24548 ) | ( x787 & ~n24650 ) | ( n24548 & ~n24650 ) ;
  assign n24652 = ~n24650 & n24651 ;
  assign n24653 = x644 | n24652 ;
  assign n24654 = ( x715 & n24648 ) | ( x715 & n24653 ) | ( n24648 & n24653 ) ;
  assign n24655 = ~n24648 & n24654 ;
  assign n24656 = x644 | n24503 ;
  assign n24657 = n24503 ^ n16376 ^ 1'b0 ;
  assign n24658 = ( n24503 & n24530 ) | ( n24503 & ~n24657 ) | ( n24530 & ~n24657 ) ;
  assign n24659 = x644 & ~n24658 ;
  assign n24660 = ( x715 & n24656 ) | ( x715 & ~n24659 ) | ( n24656 & ~n24659 ) ;
  assign n24661 = ~x715 & n24660 ;
  assign n24662 = ( x1160 & n24655 ) | ( x1160 & ~n24661 ) | ( n24655 & ~n24661 ) ;
  assign n24663 = ~n24655 & n24662 ;
  assign n24664 = x644 & ~n24503 ;
  assign n24665 = x715 & ~n24664 ;
  assign n24666 = ( n24658 & n24659 ) | ( n24658 & n24665 ) | ( n24659 & n24665 ) ;
  assign n24667 = x644 & ~n24652 ;
  assign n24668 = x715 | n24667 ;
  assign n24669 = ( n24646 & n24648 ) | ( n24646 & ~n24668 ) | ( n24648 & ~n24668 ) ;
  assign n24670 = ( x1160 & ~n24666 ) | ( x1160 & n24669 ) | ( ~n24666 & n24669 ) ;
  assign n24671 = n24666 | n24670 ;
  assign n24672 = x790 & ~n24671 ;
  assign n24673 = ( x790 & n24663 ) | ( x790 & n24672 ) | ( n24663 & n24672 ) ;
  assign n24674 = x832 & ~n24673 ;
  assign n24675 = n24647 & n24674 ;
  assign n24676 = ~x180 & n7318 ;
  assign n24677 = x832 | n24676 ;
  assign n24678 = ~n24675 & n24677 ;
  assign n24679 = ( n24502 & n24675 ) | ( n24502 & ~n24678 ) | ( n24675 & ~n24678 ) ;
  assign n24680 = x181 | n15656 ;
  assign n24681 = x709 | n2069 ;
  assign n24682 = ~n24680 & n24681 ;
  assign n24683 = ( x38 & x181 ) | ( x38 & n16700 ) | ( x181 & n16700 ) ;
  assign n24684 = ~n2069 & n24683 ;
  assign n24685 = ( x181 & n16697 ) | ( x181 & ~n24684 ) | ( n16697 & ~n24684 ) ;
  assign n24686 = ~n24684 & n24685 ;
  assign n24687 = x181 | n15644 ;
  assign n24688 = n16185 & n24687 ;
  assign n24689 = x709 | n24688 ;
  assign n24690 = ( ~n24682 & n24686 ) | ( ~n24682 & n24689 ) | ( n24686 & n24689 ) ;
  assign n24691 = ~n24682 & n24690 ;
  assign n24692 = x625 & ~n24691 ;
  assign n24693 = x625 | n24680 ;
  assign n24694 = ( x1153 & n24692 ) | ( x1153 & n24693 ) | ( n24692 & n24693 ) ;
  assign n24695 = ~n24692 & n24694 ;
  assign n24696 = x625 & ~n24680 ;
  assign n24697 = x1153 | n24696 ;
  assign n24698 = ( x625 & n24691 ) | ( x625 & ~n24697 ) | ( n24691 & ~n24697 ) ;
  assign n24699 = ~n24697 & n24698 ;
  assign n24700 = n24695 | n24699 ;
  assign n24701 = n24691 ^ x778 ^ 1'b0 ;
  assign n24702 = ( n24691 & n24700 ) | ( n24691 & n24701 ) | ( n24700 & n24701 ) ;
  assign n24703 = n24680 ^ n16234 ^ 1'b0 ;
  assign n24704 = ( n24680 & n24702 ) | ( n24680 & ~n24703 ) | ( n24702 & ~n24703 ) ;
  assign n24705 = n24680 ^ n16254 ^ 1'b0 ;
  assign n24706 = ( n24680 & n24704 ) | ( n24680 & ~n24705 ) | ( n24704 & ~n24705 ) ;
  assign n24707 = n24680 ^ n16279 ^ 1'b0 ;
  assign n24708 = ( n24680 & n24706 ) | ( n24680 & ~n24707 ) | ( n24706 & ~n24707 ) ;
  assign n24709 = n24680 ^ n16318 ^ 1'b0 ;
  assign n24710 = ( n24680 & n24708 ) | ( n24680 & ~n24709 ) | ( n24708 & ~n24709 ) ;
  assign n24711 = x628 & ~n24710 ;
  assign n24712 = x628 | n24680 ;
  assign n24713 = ( x1156 & n24711 ) | ( x1156 & n24712 ) | ( n24711 & n24712 ) ;
  assign n24714 = ~n24711 & n24713 ;
  assign n24715 = x628 & ~n24680 ;
  assign n24716 = x1156 | n24715 ;
  assign n24717 = ( n24710 & n24711 ) | ( n24710 & ~n24716 ) | ( n24711 & ~n24716 ) ;
  assign n24718 = n24714 | n24717 ;
  assign n24719 = n24710 ^ x792 ^ 1'b0 ;
  assign n24720 = ( n24710 & n24718 ) | ( n24710 & n24719 ) | ( n24718 & n24719 ) ;
  assign n24721 = n24680 ^ x647 ^ 1'b0 ;
  assign n24722 = ( n24680 & n24720 ) | ( n24680 & ~n24721 ) | ( n24720 & ~n24721 ) ;
  assign n24723 = ( n24680 & n24720 ) | ( n24680 & n24721 ) | ( n24720 & n24721 ) ;
  assign n24724 = n24722 ^ x1157 ^ 1'b0 ;
  assign n24725 = ( n24722 & n24723 ) | ( n24722 & n24724 ) | ( n24723 & n24724 ) ;
  assign n24726 = n24720 ^ x787 ^ 1'b0 ;
  assign n24727 = ( n24720 & n24725 ) | ( n24720 & n24726 ) | ( n24725 & n24726 ) ;
  assign n24728 = x644 & ~n24727 ;
  assign n24729 = x715 | n24728 ;
  assign n24730 = x644 & ~n24680 ;
  assign n24731 = x715 & ~n24730 ;
  assign n24732 = n24731 ^ x1160 ^ 1'b0 ;
  assign n24733 = x38 & n24687 ;
  assign n24734 = x754 & n15332 ;
  assign n24735 = x181 & ~n15638 ;
  assign n24736 = ( ~x39 & n24734 ) | ( ~x39 & n24735 ) | ( n24734 & n24735 ) ;
  assign n24737 = ~x39 & n24736 ;
  assign n24738 = n24737 ^ x181 ^ 1'b0 ;
  assign n24739 = ( ~x181 & x754 ) | ( ~x181 & n24738 ) | ( x754 & n24738 ) ;
  assign n24740 = ( x181 & n24737 ) | ( x181 & n24739 ) | ( n24737 & n24739 ) ;
  assign n24741 = n24739 ^ n24737 ^ x181 ;
  assign n24742 = ( n15587 & n24740 ) | ( n15587 & ~n24741 ) | ( n24740 & ~n24741 ) ;
  assign n24743 = x181 & ~n15631 ;
  assign n24744 = x754 & n15486 ;
  assign n24745 = ( x39 & n24743 ) | ( x39 & n24744 ) | ( n24743 & n24744 ) ;
  assign n24746 = n24744 ^ n24743 ^ 1'b0 ;
  assign n24747 = ( x39 & n24745 ) | ( x39 & n24746 ) | ( n24745 & n24746 ) ;
  assign n24748 = ( ~x38 & n24742 ) | ( ~x38 & n24747 ) | ( n24742 & n24747 ) ;
  assign n24749 = ~x38 & n24748 ;
  assign n24750 = ~x754 & n15646 ;
  assign n24751 = ~n24749 & n24750 ;
  assign n24752 = ( n24733 & n24749 ) | ( n24733 & ~n24751 ) | ( n24749 & ~n24751 ) ;
  assign n24753 = ~n2069 & n24752 ;
  assign n24754 = x181 & n2069 ;
  assign n24755 = n24753 | n24754 ;
  assign n24756 = n24680 ^ n15659 ^ 1'b0 ;
  assign n24757 = ( n24680 & n24755 ) | ( n24680 & ~n24756 ) | ( n24755 & ~n24756 ) ;
  assign n24758 = n15662 & n24680 ;
  assign n24759 = ( ~n15662 & n24753 ) | ( ~n15662 & n24754 ) | ( n24753 & n24754 ) ;
  assign n24760 = n24758 | n24759 ;
  assign n24761 = n24760 ^ n24757 ^ n24680 ;
  assign n24762 = n24761 ^ x1155 ^ 1'b0 ;
  assign n24763 = ( n24760 & n24761 ) | ( n24760 & ~n24762 ) | ( n24761 & ~n24762 ) ;
  assign n24764 = n24757 ^ x785 ^ 1'b0 ;
  assign n24765 = ( n24757 & n24763 ) | ( n24757 & n24764 ) | ( n24763 & n24764 ) ;
  assign n24766 = x618 & ~n24765 ;
  assign n24767 = x618 | n24680 ;
  assign n24768 = ( x1154 & n24766 ) | ( x1154 & n24767 ) | ( n24766 & n24767 ) ;
  assign n24769 = ~n24766 & n24768 ;
  assign n24770 = x618 & ~n24680 ;
  assign n24771 = x1154 | n24770 ;
  assign n24772 = ( n24765 & n24766 ) | ( n24765 & ~n24771 ) | ( n24766 & ~n24771 ) ;
  assign n24773 = n24769 | n24772 ;
  assign n24774 = n24765 ^ x781 ^ 1'b0 ;
  assign n24775 = ( n24765 & n24773 ) | ( n24765 & n24774 ) | ( n24773 & n24774 ) ;
  assign n24776 = x619 & ~n24775 ;
  assign n24777 = x619 | n24680 ;
  assign n24778 = ( x1159 & n24776 ) | ( x1159 & n24777 ) | ( n24776 & n24777 ) ;
  assign n24779 = ~n24776 & n24778 ;
  assign n24780 = x619 & ~n24680 ;
  assign n24781 = x1159 | n24780 ;
  assign n24782 = ( n24775 & n24776 ) | ( n24775 & ~n24781 ) | ( n24776 & ~n24781 ) ;
  assign n24783 = n24779 | n24782 ;
  assign n24784 = n24775 ^ x789 ^ 1'b0 ;
  assign n24785 = ( n24775 & n24783 ) | ( n24775 & n24784 ) | ( n24783 & n24784 ) ;
  assign n24786 = n24680 ^ n16518 ^ 1'b0 ;
  assign n24787 = ( n24680 & n24785 ) | ( n24680 & ~n24786 ) | ( n24785 & ~n24786 ) ;
  assign n24788 = n24680 ^ n16339 ^ 1'b0 ;
  assign n24789 = ( n24680 & n24787 ) | ( n24680 & ~n24788 ) | ( n24787 & ~n24788 ) ;
  assign n24790 = n24680 ^ n16376 ^ 1'b0 ;
  assign n24791 = ( n24680 & n24789 ) | ( n24680 & ~n24790 ) | ( n24789 & ~n24790 ) ;
  assign n24792 = x644 | n24791 ;
  assign n24793 = ( n24731 & ~n24732 ) | ( n24731 & n24792 ) | ( ~n24732 & n24792 ) ;
  assign n24794 = ( x1160 & n24732 ) | ( x1160 & n24793 ) | ( n24732 & n24793 ) ;
  assign n24795 = n24729 & ~n24794 ;
  assign n24796 = x644 & ~n24791 ;
  assign n24797 = ( ~x715 & n24680 ) | ( ~x715 & n24730 ) | ( n24680 & n24730 ) ;
  assign n24798 = x1160 & ~n24797 ;
  assign n24799 = ( x1160 & n24796 ) | ( x1160 & n24798 ) | ( n24796 & n24798 ) ;
  assign n24800 = ( x715 & n24727 ) | ( x715 & n24728 ) | ( n24727 & n24728 ) ;
  assign n24801 = n24799 & ~n24800 ;
  assign n24802 = ( x790 & n24795 ) | ( x790 & n24801 ) | ( n24795 & n24801 ) ;
  assign n24803 = n24801 ^ n24795 ^ 1'b0 ;
  assign n24804 = ( x790 & n24802 ) | ( x790 & n24803 ) | ( n24802 & n24803 ) ;
  assign n24805 = n19055 & n24789 ;
  assign n24806 = n16374 & n24722 ;
  assign n24807 = n16373 & n24723 ;
  assign n24808 = n24806 | n24807 ;
  assign n24809 = ( x787 & n24805 ) | ( x787 & n24808 ) | ( n24805 & n24808 ) ;
  assign n24810 = n24808 ^ n24805 ^ 1'b0 ;
  assign n24811 = ( x787 & n24809 ) | ( x787 & n24810 ) | ( n24809 & n24810 ) ;
  assign n24812 = x709 & ~n24752 ;
  assign n24813 = x181 & ~n16054 ;
  assign n24814 = ~x181 & n16048 ;
  assign n24815 = ( x754 & ~n24813 ) | ( x754 & n24814 ) | ( ~n24813 & n24814 ) ;
  assign n24816 = n24813 | n24815 ;
  assign n24817 = ~x181 & n16044 ;
  assign n24818 = x181 & ~n16029 ;
  assign n24819 = ( x754 & n24817 ) | ( x754 & ~n24818 ) | ( n24817 & ~n24818 ) ;
  assign n24820 = ~n24817 & n24819 ;
  assign n24821 = ( x39 & n24816 ) | ( x39 & ~n24820 ) | ( n24816 & ~n24820 ) ;
  assign n24822 = n24821 ^ n24816 ^ 1'b0 ;
  assign n24823 = ( x39 & n24821 ) | ( x39 & ~n24822 ) | ( n24821 & ~n24822 ) ;
  assign n24824 = x181 & n15795 ;
  assign n24825 = x754 & ~n24824 ;
  assign n24826 = x181 | n15876 ;
  assign n24827 = n24825 & n24826 ;
  assign n24828 = x181 & n15943 ;
  assign n24829 = x181 | n16003 ;
  assign n24830 = ( x754 & ~n24828 ) | ( x754 & n24829 ) | ( ~n24828 & n24829 ) ;
  assign n24831 = ~x754 & n24830 ;
  assign n24832 = ( x39 & n24827 ) | ( x39 & ~n24831 ) | ( n24827 & ~n24831 ) ;
  assign n24833 = ~n24827 & n24832 ;
  assign n24834 = ( x38 & n24823 ) | ( x38 & ~n24833 ) | ( n24823 & ~n24833 ) ;
  assign n24835 = ~x38 & n24834 ;
  assign n24836 = ~x754 & n15591 ;
  assign n24837 = n17156 | n24836 ;
  assign n24838 = x181 & ~n5017 ;
  assign n24839 = n24837 & n24838 ;
  assign n24840 = x38 & ~n24839 ;
  assign n24841 = n24840 ^ x709 ^ 1'b0 ;
  assign n24842 = x754 | n15968 ;
  assign n24843 = n17889 & n24842 ;
  assign n24844 = x181 | n24843 ;
  assign n24845 = ( n24840 & ~n24841 ) | ( n24840 & n24844 ) | ( ~n24841 & n24844 ) ;
  assign n24846 = ( x709 & n24841 ) | ( x709 & n24845 ) | ( n24841 & n24845 ) ;
  assign n24847 = ( ~n2069 & n24835 ) | ( ~n2069 & n24846 ) | ( n24835 & n24846 ) ;
  assign n24848 = ~n2069 & n24847 ;
  assign n24849 = n24848 ^ n24812 ^ 1'b0 ;
  assign n24850 = ( n24812 & n24848 ) | ( n24812 & n24849 ) | ( n24848 & n24849 ) ;
  assign n24851 = ( n24754 & ~n24812 ) | ( n24754 & n24850 ) | ( ~n24812 & n24850 ) ;
  assign n24852 = x625 & ~n24851 ;
  assign n24853 = x625 | n24755 ;
  assign n24854 = ( x1153 & n24852 ) | ( x1153 & n24853 ) | ( n24852 & n24853 ) ;
  assign n24855 = ~n24852 & n24854 ;
  assign n24856 = ( x608 & n24699 ) | ( x608 & ~n24855 ) | ( n24699 & ~n24855 ) ;
  assign n24857 = ~n24699 & n24856 ;
  assign n24858 = x608 | n24695 ;
  assign n24859 = x625 & ~n24755 ;
  assign n24860 = x1153 | n24859 ;
  assign n24861 = ( n24851 & n24852 ) | ( n24851 & ~n24860 ) | ( n24852 & ~n24860 ) ;
  assign n24862 = ( ~n24857 & n24858 ) | ( ~n24857 & n24861 ) | ( n24858 & n24861 ) ;
  assign n24863 = ~n24857 & n24862 ;
  assign n24864 = n24851 ^ x778 ^ 1'b0 ;
  assign n24865 = ( n24851 & n24863 ) | ( n24851 & n24864 ) | ( n24863 & n24864 ) ;
  assign n24866 = x609 & ~n24865 ;
  assign n24867 = x609 | n24702 ;
  assign n24868 = ( x1155 & n24866 ) | ( x1155 & n24867 ) | ( n24866 & n24867 ) ;
  assign n24869 = ~n24866 & n24868 ;
  assign n24870 = ~x1155 & n24760 ;
  assign n24871 = ( x660 & n24869 ) | ( x660 & ~n24870 ) | ( n24869 & ~n24870 ) ;
  assign n24872 = ~n24869 & n24871 ;
  assign n24873 = x1155 & n24761 ;
  assign n24874 = x660 | n24873 ;
  assign n24875 = x609 & ~n24702 ;
  assign n24876 = x1155 | n24875 ;
  assign n24877 = ( n24865 & n24866 ) | ( n24865 & ~n24876 ) | ( n24866 & ~n24876 ) ;
  assign n24878 = ( ~n24872 & n24874 ) | ( ~n24872 & n24877 ) | ( n24874 & n24877 ) ;
  assign n24879 = ~n24872 & n24878 ;
  assign n24880 = n24865 ^ x785 ^ 1'b0 ;
  assign n24881 = ( n24865 & n24879 ) | ( n24865 & n24880 ) | ( n24879 & n24880 ) ;
  assign n24882 = x618 & ~n24881 ;
  assign n24883 = x618 | n24704 ;
  assign n24884 = ( x1154 & n24882 ) | ( x1154 & n24883 ) | ( n24882 & n24883 ) ;
  assign n24885 = ~n24882 & n24884 ;
  assign n24886 = ( x627 & n24772 ) | ( x627 & ~n24885 ) | ( n24772 & ~n24885 ) ;
  assign n24887 = ~n24772 & n24886 ;
  assign n24888 = x627 | n24769 ;
  assign n24889 = x618 & ~n24704 ;
  assign n24890 = x1154 | n24889 ;
  assign n24891 = ( n24881 & n24882 ) | ( n24881 & ~n24890 ) | ( n24882 & ~n24890 ) ;
  assign n24892 = ( ~n24887 & n24888 ) | ( ~n24887 & n24891 ) | ( n24888 & n24891 ) ;
  assign n24893 = ~n24887 & n24892 ;
  assign n24894 = n24881 ^ x781 ^ 1'b0 ;
  assign n24895 = ( n24881 & n24893 ) | ( n24881 & n24894 ) | ( n24893 & n24894 ) ;
  assign n24896 = x619 | n24895 ;
  assign n24897 = x619 & ~n24706 ;
  assign n24898 = ( x1159 & n24896 ) | ( x1159 & ~n24897 ) | ( n24896 & ~n24897 ) ;
  assign n24899 = ~x1159 & n24898 ;
  assign n24900 = ( x648 & n24779 ) | ( x648 & ~n24899 ) | ( n24779 & ~n24899 ) ;
  assign n24901 = n24899 | n24900 ;
  assign n24902 = x619 & ~n24895 ;
  assign n24903 = x619 | n24706 ;
  assign n24904 = ( x1159 & n24902 ) | ( x1159 & n24903 ) | ( n24902 & n24903 ) ;
  assign n24905 = ~n24902 & n24904 ;
  assign n24906 = ( x648 & n24782 ) | ( x648 & ~n24905 ) | ( n24782 & ~n24905 ) ;
  assign n24907 = ~n24782 & n24906 ;
  assign n24908 = x789 & ~n24907 ;
  assign n24909 = n24901 & n24908 ;
  assign n24910 = ~x789 & n24895 ;
  assign n24911 = ( n16519 & ~n24909 ) | ( n16519 & n24910 ) | ( ~n24909 & n24910 ) ;
  assign n24912 = n24909 | n24911 ;
  assign n24913 = n24714 ^ x629 ^ 1'b0 ;
  assign n24914 = ( n24714 & n24717 ) | ( n24714 & n24913 ) | ( n24717 & n24913 ) ;
  assign n24915 = n19046 & n24787 ;
  assign n24916 = ( x792 & n24914 ) | ( x792 & n24915 ) | ( n24914 & n24915 ) ;
  assign n24917 = n24915 ^ n24914 ^ 1'b0 ;
  assign n24918 = ( x792 & n24916 ) | ( x792 & n24917 ) | ( n24916 & n24917 ) ;
  assign n24919 = n16459 & ~n24708 ;
  assign n24920 = ~x626 & n24680 ;
  assign n24921 = x626 & n24785 ;
  assign n24922 = ( n22317 & n24920 ) | ( n22317 & ~n24921 ) | ( n24920 & ~n24921 ) ;
  assign n24923 = ~n24920 & n24922 ;
  assign n24924 = ~x626 & n24785 ;
  assign n24925 = x626 & n24680 ;
  assign n24926 = ( n22322 & n24924 ) | ( n22322 & ~n24925 ) | ( n24924 & ~n24925 ) ;
  assign n24927 = ~n24924 & n24926 ;
  assign n24928 = ( ~n24919 & n24923 ) | ( ~n24919 & n24927 ) | ( n24923 & n24927 ) ;
  assign n24929 = n24919 | n24928 ;
  assign n24930 = ( x788 & ~n22314 ) | ( x788 & n24929 ) | ( ~n22314 & n24929 ) ;
  assign n24931 = ( n18482 & n22314 ) | ( n18482 & n24930 ) | ( n22314 & n24930 ) ;
  assign n24932 = ~n24918 & n24931 ;
  assign n24933 = ( n24912 & n24918 ) | ( n24912 & ~n24932 ) | ( n24918 & ~n24932 ) ;
  assign n24934 = ( ~n18484 & n24811 ) | ( ~n18484 & n24933 ) | ( n24811 & n24933 ) ;
  assign n24935 = n24811 ^ n18484 ^ 1'b0 ;
  assign n24936 = ( n24811 & n24934 ) | ( n24811 & ~n24935 ) | ( n24934 & ~n24935 ) ;
  assign n24937 = x644 | n24794 ;
  assign n24938 = x644 & n24799 ;
  assign n24939 = x790 & ~n24938 ;
  assign n24940 = n24937 & n24939 ;
  assign n24941 = ( ~n24804 & n24936 ) | ( ~n24804 & n24940 ) | ( n24936 & n24940 ) ;
  assign n24942 = ~n24804 & n24941 ;
  assign n24943 = ( x57 & n5193 ) | ( x57 & ~n24942 ) | ( n5193 & ~n24942 ) ;
  assign n24944 = n24942 | n24943 ;
  assign n24945 = x181 | n1611 ;
  assign n24946 = ~n24836 & n24945 ;
  assign n24947 = n16397 | n24946 ;
  assign n24948 = ~n15662 & n24836 ;
  assign n24949 = ~x1155 & n24945 ;
  assign n24950 = ~n24948 & n24949 ;
  assign n24951 = ( x1155 & n24947 ) | ( x1155 & n24948 ) | ( n24947 & n24948 ) ;
  assign n24952 = n24950 | n24951 ;
  assign n24953 = n24947 ^ x785 ^ 1'b0 ;
  assign n24954 = ( n24947 & n24952 ) | ( n24947 & n24953 ) | ( n24952 & n24953 ) ;
  assign n24955 = n16411 | n24954 ;
  assign n24956 = x1154 & n24955 ;
  assign n24957 = n16414 | n24954 ;
  assign n24958 = ~x1154 & n24957 ;
  assign n24959 = n24956 | n24958 ;
  assign n24960 = n24954 ^ x781 ^ 1'b0 ;
  assign n24961 = ( n24954 & n24959 ) | ( n24954 & n24960 ) | ( n24959 & n24960 ) ;
  assign n24962 = n21437 | n24961 ;
  assign n24963 = x1159 & n24962 ;
  assign n24964 = n21440 | n24961 ;
  assign n24965 = ~x1159 & n24964 ;
  assign n24966 = n24963 | n24965 ;
  assign n24967 = n24961 ^ x789 ^ 1'b0 ;
  assign n24968 = ( n24961 & n24966 ) | ( n24961 & n24967 ) | ( n24966 & n24967 ) ;
  assign n24969 = n24945 ^ n16518 ^ 1'b0 ;
  assign n24970 = ( n24945 & n24968 ) | ( n24945 & ~n24969 ) | ( n24968 & ~n24969 ) ;
  assign n24971 = n24945 ^ n16339 ^ 1'b0 ;
  assign n24972 = ( n24945 & n24970 ) | ( n24945 & ~n24971 ) | ( n24970 & ~n24971 ) ;
  assign n24973 = n19055 & n24972 ;
  assign n24974 = x647 & ~n24945 ;
  assign n24975 = x1157 | n24974 ;
  assign n24976 = ~x709 & n15778 ;
  assign n24977 = ~x625 & n24976 ;
  assign n24978 = ~x1153 & n24945 ;
  assign n24979 = ~n24977 & n24978 ;
  assign n24980 = x778 & ~n24979 ;
  assign n24981 = n24945 & ~n24976 ;
  assign n24982 = ( x1153 & n24977 ) | ( x1153 & n24981 ) | ( n24977 & n24981 ) ;
  assign n24983 = n24980 & ~n24982 ;
  assign n24984 = ( x778 & n24981 ) | ( x778 & ~n24983 ) | ( n24981 & ~n24983 ) ;
  assign n24985 = ~n24983 & n24984 ;
  assign n24986 = n16447 | n24985 ;
  assign n24987 = n16449 | n24986 ;
  assign n24988 = n16451 | n24987 ;
  assign n24989 = n16530 | n24988 ;
  assign n24990 = n16560 | n24989 ;
  assign n24991 = ( x647 & ~n24975 ) | ( x647 & n24990 ) | ( ~n24975 & n24990 ) ;
  assign n24992 = ~n24975 & n24991 ;
  assign n24993 = n24945 ^ x647 ^ 1'b0 ;
  assign n24994 = ( n24945 & n24990 ) | ( n24945 & n24993 ) | ( n24990 & n24993 ) ;
  assign n24995 = x1157 & n24994 ;
  assign n24996 = ( n16375 & n24992 ) | ( n16375 & n24995 ) | ( n24992 & n24995 ) ;
  assign n24997 = ( x787 & n24973 ) | ( x787 & n24996 ) | ( n24973 & n24996 ) ;
  assign n24998 = n24996 ^ n24973 ^ 1'b0 ;
  assign n24999 = ( x787 & n24997 ) | ( x787 & n24998 ) | ( n24997 & n24998 ) ;
  assign n25000 = ~x626 & n24945 ;
  assign n25001 = x626 & n24968 ;
  assign n25002 = ( n22317 & n25000 ) | ( n22317 & ~n25001 ) | ( n25000 & ~n25001 ) ;
  assign n25003 = ~n25000 & n25002 ;
  assign n25004 = ~x626 & n24968 ;
  assign n25005 = x626 & n24945 ;
  assign n25006 = ( n22322 & n25004 ) | ( n22322 & ~n25005 ) | ( n25004 & ~n25005 ) ;
  assign n25007 = ~n25004 & n25006 ;
  assign n25008 = n24988 & ~n25007 ;
  assign n25009 = ( n16459 & n25007 ) | ( n16459 & ~n25008 ) | ( n25007 & ~n25008 ) ;
  assign n25010 = ( x788 & n25003 ) | ( x788 & n25009 ) | ( n25003 & n25009 ) ;
  assign n25011 = n25009 ^ n25003 ^ 1'b0 ;
  assign n25012 = ( x788 & n25010 ) | ( x788 & n25011 ) | ( n25010 & n25011 ) ;
  assign n25013 = n15524 | n24981 ;
  assign n25014 = n24946 & n25013 ;
  assign n25015 = x625 & ~n25013 ;
  assign n25016 = ( n24978 & n25014 ) | ( n24978 & n25015 ) | ( n25014 & n25015 ) ;
  assign n25017 = ( x608 & n24982 ) | ( x608 & ~n25016 ) | ( n24982 & ~n25016 ) ;
  assign n25018 = n25016 | n25017 ;
  assign n25019 = x1153 & n24946 ;
  assign n25020 = ~n25015 & n25019 ;
  assign n25021 = x608 & ~n24979 ;
  assign n25022 = n25018 & ~n25021 ;
  assign n25023 = ( n25018 & n25020 ) | ( n25018 & n25022 ) | ( n25020 & n25022 ) ;
  assign n25024 = n25014 ^ x778 ^ 1'b0 ;
  assign n25025 = ( n25014 & n25023 ) | ( n25014 & n25024 ) | ( n25023 & n25024 ) ;
  assign n25026 = x609 & ~n25025 ;
  assign n25032 = x609 | n24985 ;
  assign n25033 = ( x1155 & n25026 ) | ( x1155 & n25032 ) | ( n25026 & n25032 ) ;
  assign n25034 = ~n25026 & n25033 ;
  assign n25035 = ( x660 & n24950 ) | ( x660 & ~n25034 ) | ( n24950 & ~n25034 ) ;
  assign n25036 = ~n24950 & n25035 ;
  assign n25027 = x609 & ~n24985 ;
  assign n25028 = x1155 | n25027 ;
  assign n25029 = ( n25025 & n25026 ) | ( n25025 & ~n25028 ) | ( n25026 & ~n25028 ) ;
  assign n25030 = ( x660 & n24951 ) | ( x660 & ~n25029 ) | ( n24951 & ~n25029 ) ;
  assign n25031 = n25029 | n25030 ;
  assign n25037 = n25036 ^ n25031 ^ 1'b0 ;
  assign n25038 = ( x785 & ~n25031 ) | ( x785 & n25036 ) | ( ~n25031 & n25036 ) ;
  assign n25039 = ( x785 & ~n25037 ) | ( x785 & n25038 ) | ( ~n25037 & n25038 ) ;
  assign n25040 = ( x785 & n25025 ) | ( x785 & ~n25039 ) | ( n25025 & ~n25039 ) ;
  assign n25041 = ~n25039 & n25040 ;
  assign n25042 = x618 & ~n25041 ;
  assign n25043 = x618 | n24986 ;
  assign n25044 = ( x1154 & n25042 ) | ( x1154 & n25043 ) | ( n25042 & n25043 ) ;
  assign n25045 = ~n25042 & n25044 ;
  assign n25046 = ( x627 & n24958 ) | ( x627 & ~n25045 ) | ( n24958 & ~n25045 ) ;
  assign n25047 = ~n24958 & n25046 ;
  assign n25048 = x627 | n24956 ;
  assign n25049 = x618 & ~n24986 ;
  assign n25050 = x1154 | n25049 ;
  assign n25051 = ( n25041 & n25042 ) | ( n25041 & ~n25050 ) | ( n25042 & ~n25050 ) ;
  assign n25052 = ( ~n25047 & n25048 ) | ( ~n25047 & n25051 ) | ( n25048 & n25051 ) ;
  assign n25053 = ~n25047 & n25052 ;
  assign n25054 = n25041 ^ x781 ^ 1'b0 ;
  assign n25055 = ( n25041 & n25053 ) | ( n25041 & n25054 ) | ( n25053 & n25054 ) ;
  assign n25056 = ~x789 & n25055 ;
  assign n25057 = x619 & ~n24987 ;
  assign n25058 = x1159 | n25057 ;
  assign n25059 = x619 & ~n25055 ;
  assign n25060 = ( n25055 & ~n25058 ) | ( n25055 & n25059 ) | ( ~n25058 & n25059 ) ;
  assign n25061 = ( x648 & n24963 ) | ( x648 & ~n25060 ) | ( n24963 & ~n25060 ) ;
  assign n25062 = n25060 | n25061 ;
  assign n25063 = x619 | n24987 ;
  assign n25064 = x1159 & ~n25059 ;
  assign n25065 = n25063 & n25064 ;
  assign n25066 = ( x648 & n24965 ) | ( x648 & ~n25065 ) | ( n24965 & ~n25065 ) ;
  assign n25067 = ~n24965 & n25066 ;
  assign n25068 = x789 & ~n25067 ;
  assign n25069 = n25062 & n25068 ;
  assign n25070 = ( n16519 & ~n25056 ) | ( n16519 & n25069 ) | ( ~n25056 & n25069 ) ;
  assign n25071 = n25056 | n25070 ;
  assign n25072 = n25071 ^ n25012 ^ 1'b0 ;
  assign n25073 = ( n25012 & n25071 ) | ( n25012 & n25072 ) | ( n25071 & n25072 ) ;
  assign n25074 = ( n18482 & ~n25012 ) | ( n18482 & n25073 ) | ( ~n25012 & n25073 ) ;
  assign n25075 = n19208 | n24989 ;
  assign n25076 = n16556 & ~n24970 ;
  assign n25077 = x629 & ~n25076 ;
  assign n25078 = n25075 & n25077 ;
  assign n25079 = n16557 & ~n24970 ;
  assign n25080 = n19212 & ~n24989 ;
  assign n25081 = n25079 | n25080 ;
  assign n25082 = ( x629 & ~n25078 ) | ( x629 & n25081 ) | ( ~n25078 & n25081 ) ;
  assign n25083 = ~n25078 & n25082 ;
  assign n25084 = ( x792 & ~n19206 ) | ( x792 & n25083 ) | ( ~n19206 & n25083 ) ;
  assign n25085 = ( n18484 & n19206 ) | ( n18484 & n25084 ) | ( n19206 & n25084 ) ;
  assign n25086 = ( n24999 & n25074 ) | ( n24999 & ~n25085 ) | ( n25074 & ~n25085 ) ;
  assign n25087 = n25086 ^ n25074 ^ 1'b0 ;
  assign n25088 = ( n24999 & n25086 ) | ( n24999 & ~n25087 ) | ( n25086 & ~n25087 ) ;
  assign n25089 = x790 | n25088 ;
  assign n25090 = x644 & ~n25088 ;
  assign n25091 = ( x787 & n24992 ) | ( x787 & ~n24995 ) | ( n24992 & ~n24995 ) ;
  assign n25092 = ~n24992 & n25091 ;
  assign n25093 = ( x787 & n24990 ) | ( x787 & ~n25092 ) | ( n24990 & ~n25092 ) ;
  assign n25094 = ~n25092 & n25093 ;
  assign n25095 = x644 | n25094 ;
  assign n25096 = ( x715 & n25090 ) | ( x715 & n25095 ) | ( n25090 & n25095 ) ;
  assign n25097 = ~n25090 & n25096 ;
  assign n25098 = x644 | n24945 ;
  assign n25099 = n24945 ^ n16376 ^ 1'b0 ;
  assign n25100 = ( n24945 & n24972 ) | ( n24945 & ~n25099 ) | ( n24972 & ~n25099 ) ;
  assign n25101 = x644 & ~n25100 ;
  assign n25102 = ( x715 & n25098 ) | ( x715 & ~n25101 ) | ( n25098 & ~n25101 ) ;
  assign n25103 = ~x715 & n25102 ;
  assign n25104 = ( x1160 & n25097 ) | ( x1160 & ~n25103 ) | ( n25097 & ~n25103 ) ;
  assign n25105 = ~n25097 & n25104 ;
  assign n25106 = x644 & ~n24945 ;
  assign n25107 = x715 & ~n25106 ;
  assign n25108 = ( n25100 & n25101 ) | ( n25100 & n25107 ) | ( n25101 & n25107 ) ;
  assign n25109 = x644 & ~n25094 ;
  assign n25110 = x715 | n25109 ;
  assign n25111 = ( n25088 & n25090 ) | ( n25088 & ~n25110 ) | ( n25090 & ~n25110 ) ;
  assign n25112 = ( x1160 & ~n25108 ) | ( x1160 & n25111 ) | ( ~n25108 & n25111 ) ;
  assign n25113 = n25108 | n25112 ;
  assign n25114 = x790 & ~n25113 ;
  assign n25115 = ( x790 & n25105 ) | ( x790 & n25114 ) | ( n25105 & n25114 ) ;
  assign n25116 = x832 & ~n25115 ;
  assign n25117 = n25089 & n25116 ;
  assign n25118 = ~x181 & n7318 ;
  assign n25119 = x832 | n25118 ;
  assign n25120 = ~n25117 & n25119 ;
  assign n25121 = ( n24944 & n25117 ) | ( n24944 & ~n25120 ) | ( n25117 & ~n25120 ) ;
  assign n25122 = x182 | n15656 ;
  assign n25123 = x734 | n2069 ;
  assign n25124 = ~n25122 & n25123 ;
  assign n25125 = ( x38 & x182 ) | ( x38 & n16700 ) | ( x182 & n16700 ) ;
  assign n25126 = ~n2069 & n25125 ;
  assign n25127 = ( x182 & n16697 ) | ( x182 & ~n25126 ) | ( n16697 & ~n25126 ) ;
  assign n25128 = ~n25126 & n25127 ;
  assign n25129 = x182 | n15644 ;
  assign n25130 = n16185 & n25129 ;
  assign n25131 = x734 | n25130 ;
  assign n25132 = ( ~n25124 & n25128 ) | ( ~n25124 & n25131 ) | ( n25128 & n25131 ) ;
  assign n25133 = ~n25124 & n25132 ;
  assign n25134 = x625 & ~n25133 ;
  assign n25135 = x625 | n25122 ;
  assign n25136 = ( x1153 & n25134 ) | ( x1153 & n25135 ) | ( n25134 & n25135 ) ;
  assign n25137 = ~n25134 & n25136 ;
  assign n25138 = x625 & ~n25122 ;
  assign n25139 = x1153 | n25138 ;
  assign n25140 = ( x625 & n25133 ) | ( x625 & ~n25139 ) | ( n25133 & ~n25139 ) ;
  assign n25141 = ~n25139 & n25140 ;
  assign n25142 = n25137 | n25141 ;
  assign n25143 = n25133 ^ x778 ^ 1'b0 ;
  assign n25144 = ( n25133 & n25142 ) | ( n25133 & n25143 ) | ( n25142 & n25143 ) ;
  assign n25145 = n25122 ^ n16234 ^ 1'b0 ;
  assign n25146 = ( n25122 & n25144 ) | ( n25122 & ~n25145 ) | ( n25144 & ~n25145 ) ;
  assign n25147 = n25122 ^ n16254 ^ 1'b0 ;
  assign n25148 = ( n25122 & n25146 ) | ( n25122 & ~n25147 ) | ( n25146 & ~n25147 ) ;
  assign n25149 = n25122 ^ n16279 ^ 1'b0 ;
  assign n25150 = ( n25122 & n25148 ) | ( n25122 & ~n25149 ) | ( n25148 & ~n25149 ) ;
  assign n25151 = n25122 ^ n16318 ^ 1'b0 ;
  assign n25152 = ( n25122 & n25150 ) | ( n25122 & ~n25151 ) | ( n25150 & ~n25151 ) ;
  assign n25153 = x628 & ~n25152 ;
  assign n25154 = x628 | n25122 ;
  assign n25155 = ( x1156 & n25153 ) | ( x1156 & n25154 ) | ( n25153 & n25154 ) ;
  assign n25156 = ~n25153 & n25155 ;
  assign n25157 = x628 & ~n25122 ;
  assign n25158 = x1156 | n25157 ;
  assign n25159 = ( n25152 & n25153 ) | ( n25152 & ~n25158 ) | ( n25153 & ~n25158 ) ;
  assign n25160 = n25156 | n25159 ;
  assign n25161 = n25152 ^ x792 ^ 1'b0 ;
  assign n25162 = ( n25152 & n25160 ) | ( n25152 & n25161 ) | ( n25160 & n25161 ) ;
  assign n25163 = n25122 ^ x647 ^ 1'b0 ;
  assign n25164 = ( n25122 & n25162 ) | ( n25122 & ~n25163 ) | ( n25162 & ~n25163 ) ;
  assign n25165 = ( n25122 & n25162 ) | ( n25122 & n25163 ) | ( n25162 & n25163 ) ;
  assign n25166 = n25164 ^ x1157 ^ 1'b0 ;
  assign n25167 = ( n25164 & n25165 ) | ( n25164 & n25166 ) | ( n25165 & n25166 ) ;
  assign n25168 = n25162 ^ x787 ^ 1'b0 ;
  assign n25169 = ( n25162 & n25167 ) | ( n25162 & n25168 ) | ( n25167 & n25168 ) ;
  assign n25170 = x644 & ~n25169 ;
  assign n25171 = x715 | n25170 ;
  assign n25172 = x644 & ~n25122 ;
  assign n25173 = x715 & ~n25172 ;
  assign n25174 = n25173 ^ x1160 ^ 1'b0 ;
  assign n25175 = ~x756 & n15646 ;
  assign n25176 = n25129 & ~n25175 ;
  assign n25177 = ~x182 & x756 ;
  assign n25178 = ~n15488 & n25177 ;
  assign n25179 = ~x182 & n15587 ;
  assign n25180 = x182 & ~n15640 ;
  assign n25181 = x756 | n25180 ;
  assign n25182 = ( ~n25178 & n25179 ) | ( ~n25178 & n25181 ) | ( n25179 & n25181 ) ;
  assign n25183 = ~n25178 & n25182 ;
  assign n25184 = n25176 ^ x38 ^ 1'b0 ;
  assign n25185 = ( n25176 & n25183 ) | ( n25176 & ~n25184 ) | ( n25183 & ~n25184 ) ;
  assign n25186 = ~n2069 & n25185 ;
  assign n25187 = x182 & n2069 ;
  assign n25188 = n25186 | n25187 ;
  assign n25189 = n25122 ^ n15659 ^ 1'b0 ;
  assign n25190 = ( n25122 & n25188 ) | ( n25122 & ~n25189 ) | ( n25188 & ~n25189 ) ;
  assign n25191 = n15662 & n25122 ;
  assign n25192 = ( ~n15662 & n25186 ) | ( ~n15662 & n25187 ) | ( n25186 & n25187 ) ;
  assign n25193 = n25191 | n25192 ;
  assign n25194 = n25193 ^ n25190 ^ n25122 ;
  assign n25195 = n25194 ^ x1155 ^ 1'b0 ;
  assign n25196 = ( n25193 & n25194 ) | ( n25193 & ~n25195 ) | ( n25194 & ~n25195 ) ;
  assign n25197 = n25190 ^ x785 ^ 1'b0 ;
  assign n25198 = ( n25190 & n25196 ) | ( n25190 & n25197 ) | ( n25196 & n25197 ) ;
  assign n25199 = x618 & ~n25198 ;
  assign n25200 = x618 | n25122 ;
  assign n25201 = ( x1154 & n25199 ) | ( x1154 & n25200 ) | ( n25199 & n25200 ) ;
  assign n25202 = ~n25199 & n25201 ;
  assign n25203 = x618 & ~n25122 ;
  assign n25204 = x1154 | n25203 ;
  assign n25205 = ( n25198 & n25199 ) | ( n25198 & ~n25204 ) | ( n25199 & ~n25204 ) ;
  assign n25206 = n25202 | n25205 ;
  assign n25207 = n25198 ^ x781 ^ 1'b0 ;
  assign n25208 = ( n25198 & n25206 ) | ( n25198 & n25207 ) | ( n25206 & n25207 ) ;
  assign n25209 = x619 & ~n25208 ;
  assign n25210 = x619 | n25122 ;
  assign n25211 = ( x1159 & n25209 ) | ( x1159 & n25210 ) | ( n25209 & n25210 ) ;
  assign n25212 = ~n25209 & n25211 ;
  assign n25213 = x619 & ~n25122 ;
  assign n25214 = x1159 | n25213 ;
  assign n25215 = ( n25208 & n25209 ) | ( n25208 & ~n25214 ) | ( n25209 & ~n25214 ) ;
  assign n25216 = n25212 | n25215 ;
  assign n25217 = n25208 ^ x789 ^ 1'b0 ;
  assign n25218 = ( n25208 & n25216 ) | ( n25208 & n25217 ) | ( n25216 & n25217 ) ;
  assign n25219 = n25122 ^ n16518 ^ 1'b0 ;
  assign n25220 = ( n25122 & n25218 ) | ( n25122 & ~n25219 ) | ( n25218 & ~n25219 ) ;
  assign n25221 = n25122 ^ n16339 ^ 1'b0 ;
  assign n25222 = ( n25122 & n25220 ) | ( n25122 & ~n25221 ) | ( n25220 & ~n25221 ) ;
  assign n25223 = n25122 ^ n16376 ^ 1'b0 ;
  assign n25224 = ( n25122 & n25222 ) | ( n25122 & ~n25223 ) | ( n25222 & ~n25223 ) ;
  assign n25225 = x644 | n25224 ;
  assign n25226 = ( n25173 & ~n25174 ) | ( n25173 & n25225 ) | ( ~n25174 & n25225 ) ;
  assign n25227 = ( x1160 & n25174 ) | ( x1160 & n25226 ) | ( n25174 & n25226 ) ;
  assign n25228 = n25171 & ~n25227 ;
  assign n25229 = x644 & ~n25224 ;
  assign n25230 = ( ~x715 & n25122 ) | ( ~x715 & n25172 ) | ( n25122 & n25172 ) ;
  assign n25231 = x1160 & ~n25230 ;
  assign n25232 = ( x1160 & n25229 ) | ( x1160 & n25231 ) | ( n25229 & n25231 ) ;
  assign n25233 = ( x715 & n25169 ) | ( x715 & n25170 ) | ( n25169 & n25170 ) ;
  assign n25234 = n25232 & ~n25233 ;
  assign n25235 = ( x790 & n25228 ) | ( x790 & n25234 ) | ( n25228 & n25234 ) ;
  assign n25236 = n25234 ^ n25228 ^ 1'b0 ;
  assign n25237 = ( x790 & n25235 ) | ( x790 & n25236 ) | ( n25235 & n25236 ) ;
  assign n25238 = n19055 & n25222 ;
  assign n25239 = n16374 & n25164 ;
  assign n25240 = n16373 & n25165 ;
  assign n25241 = n25239 | n25240 ;
  assign n25242 = ( x787 & n25238 ) | ( x787 & n25241 ) | ( n25238 & n25241 ) ;
  assign n25243 = n25241 ^ n25238 ^ 1'b0 ;
  assign n25244 = ( x787 & n25242 ) | ( x787 & n25243 ) | ( n25242 & n25243 ) ;
  assign n25245 = x734 & ~n25185 ;
  assign n25246 = x182 & ~n16054 ;
  assign n25247 = ~x182 & n16048 ;
  assign n25248 = ( x756 & ~n25246 ) | ( x756 & n25247 ) | ( ~n25246 & n25247 ) ;
  assign n25249 = n25246 | n25248 ;
  assign n25250 = ~x182 & n16044 ;
  assign n25251 = x182 & ~n16029 ;
  assign n25252 = ( x756 & n25250 ) | ( x756 & ~n25251 ) | ( n25250 & ~n25251 ) ;
  assign n25253 = ~n25250 & n25252 ;
  assign n25254 = ( x39 & n25249 ) | ( x39 & ~n25253 ) | ( n25249 & ~n25253 ) ;
  assign n25255 = n25254 ^ n25249 ^ 1'b0 ;
  assign n25256 = ( x39 & n25254 ) | ( x39 & ~n25255 ) | ( n25254 & ~n25255 ) ;
  assign n25257 = x182 & n15795 ;
  assign n25258 = x756 & ~n25257 ;
  assign n25259 = x182 | n15876 ;
  assign n25260 = n25258 & n25259 ;
  assign n25261 = x182 & n15943 ;
  assign n25262 = x182 | n16003 ;
  assign n25263 = ( x756 & ~n25261 ) | ( x756 & n25262 ) | ( ~n25261 & n25262 ) ;
  assign n25264 = ~x756 & n25263 ;
  assign n25265 = ( x39 & n25260 ) | ( x39 & ~n25264 ) | ( n25260 & ~n25264 ) ;
  assign n25266 = ~n25260 & n25265 ;
  assign n25267 = ( x38 & n25256 ) | ( x38 & ~n25266 ) | ( n25256 & ~n25266 ) ;
  assign n25268 = ~x38 & n25267 ;
  assign n25269 = ~x756 & n15591 ;
  assign n25270 = n17156 | n25269 ;
  assign n25271 = x182 & ~n5017 ;
  assign n25272 = n25270 & n25271 ;
  assign n25273 = x38 & ~n25272 ;
  assign n25274 = n25273 ^ x734 ^ 1'b0 ;
  assign n25275 = x756 | n15968 ;
  assign n25276 = n17889 & n25275 ;
  assign n25277 = x182 | n25276 ;
  assign n25278 = ( n25273 & ~n25274 ) | ( n25273 & n25277 ) | ( ~n25274 & n25277 ) ;
  assign n25279 = ( x734 & n25274 ) | ( x734 & n25278 ) | ( n25274 & n25278 ) ;
  assign n25280 = ( ~n2069 & n25268 ) | ( ~n2069 & n25279 ) | ( n25268 & n25279 ) ;
  assign n25281 = ~n2069 & n25280 ;
  assign n25282 = n25281 ^ n25245 ^ 1'b0 ;
  assign n25283 = ( n25245 & n25281 ) | ( n25245 & n25282 ) | ( n25281 & n25282 ) ;
  assign n25284 = ( n25187 & ~n25245 ) | ( n25187 & n25283 ) | ( ~n25245 & n25283 ) ;
  assign n25285 = x625 & ~n25284 ;
  assign n25286 = x625 | n25188 ;
  assign n25287 = ( x1153 & n25285 ) | ( x1153 & n25286 ) | ( n25285 & n25286 ) ;
  assign n25288 = ~n25285 & n25287 ;
  assign n25289 = ( x608 & n25141 ) | ( x608 & ~n25288 ) | ( n25141 & ~n25288 ) ;
  assign n25290 = ~n25141 & n25289 ;
  assign n25291 = x608 | n25137 ;
  assign n25292 = x625 & ~n25188 ;
  assign n25293 = x1153 | n25292 ;
  assign n25294 = ( n25284 & n25285 ) | ( n25284 & ~n25293 ) | ( n25285 & ~n25293 ) ;
  assign n25295 = ( ~n25290 & n25291 ) | ( ~n25290 & n25294 ) | ( n25291 & n25294 ) ;
  assign n25296 = ~n25290 & n25295 ;
  assign n25297 = n25284 ^ x778 ^ 1'b0 ;
  assign n25298 = ( n25284 & n25296 ) | ( n25284 & n25297 ) | ( n25296 & n25297 ) ;
  assign n25299 = x609 & ~n25298 ;
  assign n25300 = x609 | n25144 ;
  assign n25301 = ( x1155 & n25299 ) | ( x1155 & n25300 ) | ( n25299 & n25300 ) ;
  assign n25302 = ~n25299 & n25301 ;
  assign n25303 = ~x1155 & n25193 ;
  assign n25304 = ( x660 & n25302 ) | ( x660 & ~n25303 ) | ( n25302 & ~n25303 ) ;
  assign n25305 = ~n25302 & n25304 ;
  assign n25306 = x1155 & n25194 ;
  assign n25307 = x660 | n25306 ;
  assign n25308 = x609 & ~n25144 ;
  assign n25309 = x1155 | n25308 ;
  assign n25310 = ( n25298 & n25299 ) | ( n25298 & ~n25309 ) | ( n25299 & ~n25309 ) ;
  assign n25311 = ( ~n25305 & n25307 ) | ( ~n25305 & n25310 ) | ( n25307 & n25310 ) ;
  assign n25312 = ~n25305 & n25311 ;
  assign n25313 = n25298 ^ x785 ^ 1'b0 ;
  assign n25314 = ( n25298 & n25312 ) | ( n25298 & n25313 ) | ( n25312 & n25313 ) ;
  assign n25315 = x618 & ~n25314 ;
  assign n25316 = x618 | n25146 ;
  assign n25317 = ( x1154 & n25315 ) | ( x1154 & n25316 ) | ( n25315 & n25316 ) ;
  assign n25318 = ~n25315 & n25317 ;
  assign n25319 = ( x627 & n25205 ) | ( x627 & ~n25318 ) | ( n25205 & ~n25318 ) ;
  assign n25320 = ~n25205 & n25319 ;
  assign n25321 = x627 | n25202 ;
  assign n25322 = x618 & ~n25146 ;
  assign n25323 = x1154 | n25322 ;
  assign n25324 = ( n25314 & n25315 ) | ( n25314 & ~n25323 ) | ( n25315 & ~n25323 ) ;
  assign n25325 = ( ~n25320 & n25321 ) | ( ~n25320 & n25324 ) | ( n25321 & n25324 ) ;
  assign n25326 = ~n25320 & n25325 ;
  assign n25327 = n25314 ^ x781 ^ 1'b0 ;
  assign n25328 = ( n25314 & n25326 ) | ( n25314 & n25327 ) | ( n25326 & n25327 ) ;
  assign n25329 = x619 | n25328 ;
  assign n25330 = x619 & ~n25148 ;
  assign n25331 = ( x1159 & n25329 ) | ( x1159 & ~n25330 ) | ( n25329 & ~n25330 ) ;
  assign n25332 = ~x1159 & n25331 ;
  assign n25333 = ( x648 & n25212 ) | ( x648 & ~n25332 ) | ( n25212 & ~n25332 ) ;
  assign n25334 = n25332 | n25333 ;
  assign n25335 = x619 & ~n25328 ;
  assign n25336 = x619 | n25148 ;
  assign n25337 = ( x1159 & n25335 ) | ( x1159 & n25336 ) | ( n25335 & n25336 ) ;
  assign n25338 = ~n25335 & n25337 ;
  assign n25339 = ( x648 & n25215 ) | ( x648 & ~n25338 ) | ( n25215 & ~n25338 ) ;
  assign n25340 = ~n25215 & n25339 ;
  assign n25341 = x789 & ~n25340 ;
  assign n25342 = n25334 & n25341 ;
  assign n25343 = ~x789 & n25328 ;
  assign n25344 = ( n16519 & ~n25342 ) | ( n16519 & n25343 ) | ( ~n25342 & n25343 ) ;
  assign n25345 = n25342 | n25344 ;
  assign n25346 = n25156 ^ x629 ^ 1'b0 ;
  assign n25347 = ( n25156 & n25159 ) | ( n25156 & n25346 ) | ( n25159 & n25346 ) ;
  assign n25348 = n19046 & n25220 ;
  assign n25349 = ( x792 & n25347 ) | ( x792 & n25348 ) | ( n25347 & n25348 ) ;
  assign n25350 = n25348 ^ n25347 ^ 1'b0 ;
  assign n25351 = ( x792 & n25349 ) | ( x792 & n25350 ) | ( n25349 & n25350 ) ;
  assign n25352 = n16459 & ~n25150 ;
  assign n25353 = ~x626 & n25122 ;
  assign n25354 = x626 & n25218 ;
  assign n25355 = ( n22317 & n25353 ) | ( n22317 & ~n25354 ) | ( n25353 & ~n25354 ) ;
  assign n25356 = ~n25353 & n25355 ;
  assign n25357 = ~x626 & n25218 ;
  assign n25358 = x626 & n25122 ;
  assign n25359 = ( n22322 & n25357 ) | ( n22322 & ~n25358 ) | ( n25357 & ~n25358 ) ;
  assign n25360 = ~n25357 & n25359 ;
  assign n25361 = ( ~n25352 & n25356 ) | ( ~n25352 & n25360 ) | ( n25356 & n25360 ) ;
  assign n25362 = n25352 | n25361 ;
  assign n25363 = ( x788 & ~n22314 ) | ( x788 & n25362 ) | ( ~n22314 & n25362 ) ;
  assign n25364 = ( n18482 & n22314 ) | ( n18482 & n25363 ) | ( n22314 & n25363 ) ;
  assign n25365 = ~n25351 & n25364 ;
  assign n25366 = ( n25345 & n25351 ) | ( n25345 & ~n25365 ) | ( n25351 & ~n25365 ) ;
  assign n25367 = ( ~n18484 & n25244 ) | ( ~n18484 & n25366 ) | ( n25244 & n25366 ) ;
  assign n25368 = n25244 ^ n18484 ^ 1'b0 ;
  assign n25369 = ( n25244 & n25367 ) | ( n25244 & ~n25368 ) | ( n25367 & ~n25368 ) ;
  assign n25370 = x644 | n25227 ;
  assign n25371 = x644 & n25232 ;
  assign n25372 = x790 & ~n25371 ;
  assign n25373 = n25370 & n25372 ;
  assign n25374 = ( ~n25237 & n25369 ) | ( ~n25237 & n25373 ) | ( n25369 & n25373 ) ;
  assign n25375 = ~n25237 & n25374 ;
  assign n25376 = ( x57 & n5193 ) | ( x57 & ~n25375 ) | ( n5193 & ~n25375 ) ;
  assign n25377 = n25375 | n25376 ;
  assign n25378 = x182 | n1611 ;
  assign n25379 = ~n25269 & n25378 ;
  assign n25380 = n16397 | n25379 ;
  assign n25381 = ~n15662 & n25269 ;
  assign n25382 = ~x1155 & n25378 ;
  assign n25383 = ~n25381 & n25382 ;
  assign n25384 = ( x1155 & n25380 ) | ( x1155 & n25381 ) | ( n25380 & n25381 ) ;
  assign n25385 = n25383 | n25384 ;
  assign n25386 = n25380 ^ x785 ^ 1'b0 ;
  assign n25387 = ( n25380 & n25385 ) | ( n25380 & n25386 ) | ( n25385 & n25386 ) ;
  assign n25388 = n16411 | n25387 ;
  assign n25389 = x1154 & n25388 ;
  assign n25390 = n16414 | n25387 ;
  assign n25391 = ~x1154 & n25390 ;
  assign n25392 = n25389 | n25391 ;
  assign n25393 = n25387 ^ x781 ^ 1'b0 ;
  assign n25394 = ( n25387 & n25392 ) | ( n25387 & n25393 ) | ( n25392 & n25393 ) ;
  assign n25395 = n21437 | n25394 ;
  assign n25396 = x1159 & n25395 ;
  assign n25397 = n21440 | n25394 ;
  assign n25398 = ~x1159 & n25397 ;
  assign n25399 = n25396 | n25398 ;
  assign n25400 = n25394 ^ x789 ^ 1'b0 ;
  assign n25401 = ( n25394 & n25399 ) | ( n25394 & n25400 ) | ( n25399 & n25400 ) ;
  assign n25402 = n25378 ^ n16518 ^ 1'b0 ;
  assign n25403 = ( n25378 & n25401 ) | ( n25378 & ~n25402 ) | ( n25401 & ~n25402 ) ;
  assign n25404 = n25378 ^ n16339 ^ 1'b0 ;
  assign n25405 = ( n25378 & n25403 ) | ( n25378 & ~n25404 ) | ( n25403 & ~n25404 ) ;
  assign n25406 = n19055 & n25405 ;
  assign n25407 = x647 & ~n25378 ;
  assign n25408 = x1157 | n25407 ;
  assign n25409 = ~x734 & n15778 ;
  assign n25410 = ~x625 & n25409 ;
  assign n25411 = ~x1153 & n25378 ;
  assign n25412 = ~n25410 & n25411 ;
  assign n25413 = x778 & ~n25412 ;
  assign n25414 = n25378 & ~n25409 ;
  assign n25415 = ( x1153 & n25410 ) | ( x1153 & n25414 ) | ( n25410 & n25414 ) ;
  assign n25416 = n25413 & ~n25415 ;
  assign n25417 = ( x778 & n25414 ) | ( x778 & ~n25416 ) | ( n25414 & ~n25416 ) ;
  assign n25418 = ~n25416 & n25417 ;
  assign n25419 = n16447 | n25418 ;
  assign n25420 = n16449 | n25419 ;
  assign n25421 = n16451 | n25420 ;
  assign n25422 = n16530 | n25421 ;
  assign n25423 = n16560 | n25422 ;
  assign n25424 = ( x647 & ~n25408 ) | ( x647 & n25423 ) | ( ~n25408 & n25423 ) ;
  assign n25425 = ~n25408 & n25424 ;
  assign n25426 = n25378 ^ x647 ^ 1'b0 ;
  assign n25427 = ( n25378 & n25423 ) | ( n25378 & n25426 ) | ( n25423 & n25426 ) ;
  assign n25428 = x1157 & n25427 ;
  assign n25429 = ( n16375 & n25425 ) | ( n16375 & n25428 ) | ( n25425 & n25428 ) ;
  assign n25430 = ( x787 & n25406 ) | ( x787 & n25429 ) | ( n25406 & n25429 ) ;
  assign n25431 = n25429 ^ n25406 ^ 1'b0 ;
  assign n25432 = ( x787 & n25430 ) | ( x787 & n25431 ) | ( n25430 & n25431 ) ;
  assign n25433 = ~x626 & n25378 ;
  assign n25434 = x626 & n25401 ;
  assign n25435 = ( n22317 & n25433 ) | ( n22317 & ~n25434 ) | ( n25433 & ~n25434 ) ;
  assign n25436 = ~n25433 & n25435 ;
  assign n25437 = ~x626 & n25401 ;
  assign n25438 = x626 & n25378 ;
  assign n25439 = ( n22322 & n25437 ) | ( n22322 & ~n25438 ) | ( n25437 & ~n25438 ) ;
  assign n25440 = ~n25437 & n25439 ;
  assign n25441 = n25421 & ~n25440 ;
  assign n25442 = ( n16459 & n25440 ) | ( n16459 & ~n25441 ) | ( n25440 & ~n25441 ) ;
  assign n25443 = ( x788 & n25436 ) | ( x788 & n25442 ) | ( n25436 & n25442 ) ;
  assign n25444 = n25442 ^ n25436 ^ 1'b0 ;
  assign n25445 = ( x788 & n25443 ) | ( x788 & n25444 ) | ( n25443 & n25444 ) ;
  assign n25446 = n15524 | n25414 ;
  assign n25447 = n25379 & n25446 ;
  assign n25448 = x625 & ~n25446 ;
  assign n25449 = ( n25411 & n25447 ) | ( n25411 & n25448 ) | ( n25447 & n25448 ) ;
  assign n25450 = ( x608 & n25415 ) | ( x608 & ~n25449 ) | ( n25415 & ~n25449 ) ;
  assign n25451 = n25449 | n25450 ;
  assign n25452 = x1153 & n25379 ;
  assign n25453 = ~n25448 & n25452 ;
  assign n25454 = x608 & ~n25412 ;
  assign n25455 = n25451 & ~n25454 ;
  assign n25456 = ( n25451 & n25453 ) | ( n25451 & n25455 ) | ( n25453 & n25455 ) ;
  assign n25457 = n25447 ^ x778 ^ 1'b0 ;
  assign n25458 = ( n25447 & n25456 ) | ( n25447 & n25457 ) | ( n25456 & n25457 ) ;
  assign n25459 = x609 & ~n25458 ;
  assign n25465 = x609 | n25418 ;
  assign n25466 = ( x1155 & n25459 ) | ( x1155 & n25465 ) | ( n25459 & n25465 ) ;
  assign n25467 = ~n25459 & n25466 ;
  assign n25468 = ( x660 & n25383 ) | ( x660 & ~n25467 ) | ( n25383 & ~n25467 ) ;
  assign n25469 = ~n25383 & n25468 ;
  assign n25460 = x609 & ~n25418 ;
  assign n25461 = x1155 | n25460 ;
  assign n25462 = ( n25458 & n25459 ) | ( n25458 & ~n25461 ) | ( n25459 & ~n25461 ) ;
  assign n25463 = ( x660 & n25384 ) | ( x660 & ~n25462 ) | ( n25384 & ~n25462 ) ;
  assign n25464 = n25462 | n25463 ;
  assign n25470 = n25469 ^ n25464 ^ 1'b0 ;
  assign n25471 = ( x785 & ~n25464 ) | ( x785 & n25469 ) | ( ~n25464 & n25469 ) ;
  assign n25472 = ( x785 & ~n25470 ) | ( x785 & n25471 ) | ( ~n25470 & n25471 ) ;
  assign n25473 = ( x785 & n25458 ) | ( x785 & ~n25472 ) | ( n25458 & ~n25472 ) ;
  assign n25474 = ~n25472 & n25473 ;
  assign n25475 = x618 & ~n25474 ;
  assign n25476 = x618 | n25419 ;
  assign n25477 = ( x1154 & n25475 ) | ( x1154 & n25476 ) | ( n25475 & n25476 ) ;
  assign n25478 = ~n25475 & n25477 ;
  assign n25479 = ( x627 & n25391 ) | ( x627 & ~n25478 ) | ( n25391 & ~n25478 ) ;
  assign n25480 = ~n25391 & n25479 ;
  assign n25481 = x627 | n25389 ;
  assign n25482 = x618 & ~n25419 ;
  assign n25483 = x1154 | n25482 ;
  assign n25484 = ( n25474 & n25475 ) | ( n25474 & ~n25483 ) | ( n25475 & ~n25483 ) ;
  assign n25485 = ( ~n25480 & n25481 ) | ( ~n25480 & n25484 ) | ( n25481 & n25484 ) ;
  assign n25486 = ~n25480 & n25485 ;
  assign n25487 = n25474 ^ x781 ^ 1'b0 ;
  assign n25488 = ( n25474 & n25486 ) | ( n25474 & n25487 ) | ( n25486 & n25487 ) ;
  assign n25489 = ~x789 & n25488 ;
  assign n25490 = x619 & ~n25420 ;
  assign n25491 = x1159 | n25490 ;
  assign n25492 = x619 & ~n25488 ;
  assign n25493 = ( n25488 & ~n25491 ) | ( n25488 & n25492 ) | ( ~n25491 & n25492 ) ;
  assign n25494 = ( x648 & n25396 ) | ( x648 & ~n25493 ) | ( n25396 & ~n25493 ) ;
  assign n25495 = n25493 | n25494 ;
  assign n25496 = x619 | n25420 ;
  assign n25497 = x1159 & ~n25492 ;
  assign n25498 = n25496 & n25497 ;
  assign n25499 = ( x648 & n25398 ) | ( x648 & ~n25498 ) | ( n25398 & ~n25498 ) ;
  assign n25500 = ~n25398 & n25499 ;
  assign n25501 = x789 & ~n25500 ;
  assign n25502 = n25495 & n25501 ;
  assign n25503 = ( n16519 & ~n25489 ) | ( n16519 & n25502 ) | ( ~n25489 & n25502 ) ;
  assign n25504 = n25489 | n25503 ;
  assign n25505 = n25504 ^ n25445 ^ 1'b0 ;
  assign n25506 = ( n25445 & n25504 ) | ( n25445 & n25505 ) | ( n25504 & n25505 ) ;
  assign n25507 = ( n18482 & ~n25445 ) | ( n18482 & n25506 ) | ( ~n25445 & n25506 ) ;
  assign n25508 = n19208 | n25422 ;
  assign n25509 = n16556 & ~n25403 ;
  assign n25510 = x629 & ~n25509 ;
  assign n25511 = n25508 & n25510 ;
  assign n25512 = n16557 & ~n25403 ;
  assign n25513 = n19212 & ~n25422 ;
  assign n25514 = n25512 | n25513 ;
  assign n25515 = ( x629 & ~n25511 ) | ( x629 & n25514 ) | ( ~n25511 & n25514 ) ;
  assign n25516 = ~n25511 & n25515 ;
  assign n25517 = ( x792 & ~n19206 ) | ( x792 & n25516 ) | ( ~n19206 & n25516 ) ;
  assign n25518 = ( n18484 & n19206 ) | ( n18484 & n25517 ) | ( n19206 & n25517 ) ;
  assign n25519 = ( n25432 & n25507 ) | ( n25432 & ~n25518 ) | ( n25507 & ~n25518 ) ;
  assign n25520 = n25519 ^ n25507 ^ 1'b0 ;
  assign n25521 = ( n25432 & n25519 ) | ( n25432 & ~n25520 ) | ( n25519 & ~n25520 ) ;
  assign n25522 = x790 | n25521 ;
  assign n25523 = x644 & ~n25521 ;
  assign n25524 = ( x787 & n25425 ) | ( x787 & ~n25428 ) | ( n25425 & ~n25428 ) ;
  assign n25525 = ~n25425 & n25524 ;
  assign n25526 = ( x787 & n25423 ) | ( x787 & ~n25525 ) | ( n25423 & ~n25525 ) ;
  assign n25527 = ~n25525 & n25526 ;
  assign n25528 = x644 | n25527 ;
  assign n25529 = ( x715 & n25523 ) | ( x715 & n25528 ) | ( n25523 & n25528 ) ;
  assign n25530 = ~n25523 & n25529 ;
  assign n25531 = x644 | n25378 ;
  assign n25532 = n25378 ^ n16376 ^ 1'b0 ;
  assign n25533 = ( n25378 & n25405 ) | ( n25378 & ~n25532 ) | ( n25405 & ~n25532 ) ;
  assign n25534 = x644 & ~n25533 ;
  assign n25535 = ( x715 & n25531 ) | ( x715 & ~n25534 ) | ( n25531 & ~n25534 ) ;
  assign n25536 = ~x715 & n25535 ;
  assign n25537 = ( x1160 & n25530 ) | ( x1160 & ~n25536 ) | ( n25530 & ~n25536 ) ;
  assign n25538 = ~n25530 & n25537 ;
  assign n25539 = x644 & ~n25378 ;
  assign n25540 = x715 & ~n25539 ;
  assign n25541 = ( n25533 & n25534 ) | ( n25533 & n25540 ) | ( n25534 & n25540 ) ;
  assign n25542 = x644 & ~n25527 ;
  assign n25543 = x715 | n25542 ;
  assign n25544 = ( n25521 & n25523 ) | ( n25521 & ~n25543 ) | ( n25523 & ~n25543 ) ;
  assign n25545 = ( x1160 & ~n25541 ) | ( x1160 & n25544 ) | ( ~n25541 & n25544 ) ;
  assign n25546 = n25541 | n25545 ;
  assign n25547 = x790 & ~n25546 ;
  assign n25548 = ( x790 & n25538 ) | ( x790 & n25547 ) | ( n25538 & n25547 ) ;
  assign n25549 = x832 & ~n25548 ;
  assign n25550 = n25522 & n25549 ;
  assign n25551 = ~x182 & n7318 ;
  assign n25552 = x832 | n25551 ;
  assign n25553 = ~n25550 & n25552 ;
  assign n25554 = ( n25377 & n25550 ) | ( n25377 & ~n25553 ) | ( n25550 & ~n25553 ) ;
  assign n25555 = x183 | n15656 ;
  assign n25556 = x725 | n2069 ;
  assign n25557 = ~n25555 & n25556 ;
  assign n25558 = ( x38 & x183 ) | ( x38 & n16700 ) | ( x183 & n16700 ) ;
  assign n25559 = ~n2069 & n25558 ;
  assign n25560 = ( x183 & n16697 ) | ( x183 & ~n25559 ) | ( n16697 & ~n25559 ) ;
  assign n25561 = ~n25559 & n25560 ;
  assign n25562 = x183 | n15644 ;
  assign n25563 = n16185 & n25562 ;
  assign n25564 = x725 | n25563 ;
  assign n25565 = ( ~n25557 & n25561 ) | ( ~n25557 & n25564 ) | ( n25561 & n25564 ) ;
  assign n25566 = ~n25557 & n25565 ;
  assign n25567 = x625 & ~n25566 ;
  assign n25568 = x625 | n25555 ;
  assign n25569 = ( x1153 & n25567 ) | ( x1153 & n25568 ) | ( n25567 & n25568 ) ;
  assign n25570 = ~n25567 & n25569 ;
  assign n25571 = x625 & ~n25555 ;
  assign n25572 = x1153 | n25571 ;
  assign n25573 = ( x625 & n25566 ) | ( x625 & ~n25572 ) | ( n25566 & ~n25572 ) ;
  assign n25574 = ~n25572 & n25573 ;
  assign n25575 = n25570 | n25574 ;
  assign n25576 = n25566 ^ x778 ^ 1'b0 ;
  assign n25577 = ( n25566 & n25575 ) | ( n25566 & n25576 ) | ( n25575 & n25576 ) ;
  assign n25578 = n25555 ^ n16234 ^ 1'b0 ;
  assign n25579 = ( n25555 & n25577 ) | ( n25555 & ~n25578 ) | ( n25577 & ~n25578 ) ;
  assign n25580 = n25555 ^ n16254 ^ 1'b0 ;
  assign n25581 = ( n25555 & n25579 ) | ( n25555 & ~n25580 ) | ( n25579 & ~n25580 ) ;
  assign n25582 = n25555 ^ n16279 ^ 1'b0 ;
  assign n25583 = ( n25555 & n25581 ) | ( n25555 & ~n25582 ) | ( n25581 & ~n25582 ) ;
  assign n25584 = n25555 ^ n16318 ^ 1'b0 ;
  assign n25585 = ( n25555 & n25583 ) | ( n25555 & ~n25584 ) | ( n25583 & ~n25584 ) ;
  assign n25586 = x628 & ~n25585 ;
  assign n25587 = x628 | n25555 ;
  assign n25588 = ( x1156 & n25586 ) | ( x1156 & n25587 ) | ( n25586 & n25587 ) ;
  assign n25589 = ~n25586 & n25588 ;
  assign n25590 = x628 & ~n25555 ;
  assign n25591 = x1156 | n25590 ;
  assign n25592 = ( n25585 & n25586 ) | ( n25585 & ~n25591 ) | ( n25586 & ~n25591 ) ;
  assign n25593 = n25589 | n25592 ;
  assign n25594 = n25585 ^ x792 ^ 1'b0 ;
  assign n25595 = ( n25585 & n25593 ) | ( n25585 & n25594 ) | ( n25593 & n25594 ) ;
  assign n25596 = n25555 ^ x647 ^ 1'b0 ;
  assign n25597 = ( n25555 & n25595 ) | ( n25555 & ~n25596 ) | ( n25595 & ~n25596 ) ;
  assign n25598 = ( n25555 & n25595 ) | ( n25555 & n25596 ) | ( n25595 & n25596 ) ;
  assign n25599 = n25597 ^ x1157 ^ 1'b0 ;
  assign n25600 = ( n25597 & n25598 ) | ( n25597 & n25599 ) | ( n25598 & n25599 ) ;
  assign n25601 = n25595 ^ x787 ^ 1'b0 ;
  assign n25602 = ( n25595 & n25600 ) | ( n25595 & n25601 ) | ( n25600 & n25601 ) ;
  assign n25603 = x644 & ~n25602 ;
  assign n25604 = x715 | n25603 ;
  assign n25605 = x644 & ~n25555 ;
  assign n25606 = x715 & ~n25605 ;
  assign n25607 = n25606 ^ x1160 ^ 1'b0 ;
  assign n25608 = ~x755 & n15646 ;
  assign n25609 = n25562 & ~n25608 ;
  assign n25610 = ~x183 & x755 ;
  assign n25611 = ~n15488 & n25610 ;
  assign n25612 = ~x183 & n15587 ;
  assign n25613 = x183 & ~n15640 ;
  assign n25614 = x755 | n25613 ;
  assign n25615 = ( ~n25611 & n25612 ) | ( ~n25611 & n25614 ) | ( n25612 & n25614 ) ;
  assign n25616 = ~n25611 & n25615 ;
  assign n25617 = n25609 ^ x38 ^ 1'b0 ;
  assign n25618 = ( n25609 & n25616 ) | ( n25609 & ~n25617 ) | ( n25616 & ~n25617 ) ;
  assign n25619 = ~n2069 & n25618 ;
  assign n25620 = x183 & n2069 ;
  assign n25621 = n25619 | n25620 ;
  assign n25622 = n25555 ^ n15659 ^ 1'b0 ;
  assign n25623 = ( n25555 & n25621 ) | ( n25555 & ~n25622 ) | ( n25621 & ~n25622 ) ;
  assign n25624 = n15662 & n25555 ;
  assign n25625 = ( ~n15662 & n25619 ) | ( ~n15662 & n25620 ) | ( n25619 & n25620 ) ;
  assign n25626 = n25624 | n25625 ;
  assign n25627 = n25626 ^ n25623 ^ n25555 ;
  assign n25628 = n25627 ^ x1155 ^ 1'b0 ;
  assign n25629 = ( n25626 & n25627 ) | ( n25626 & ~n25628 ) | ( n25627 & ~n25628 ) ;
  assign n25630 = n25623 ^ x785 ^ 1'b0 ;
  assign n25631 = ( n25623 & n25629 ) | ( n25623 & n25630 ) | ( n25629 & n25630 ) ;
  assign n25632 = x618 & ~n25631 ;
  assign n25633 = x618 | n25555 ;
  assign n25634 = ( x1154 & n25632 ) | ( x1154 & n25633 ) | ( n25632 & n25633 ) ;
  assign n25635 = ~n25632 & n25634 ;
  assign n25636 = x618 & ~n25555 ;
  assign n25637 = x1154 | n25636 ;
  assign n25638 = ( n25631 & n25632 ) | ( n25631 & ~n25637 ) | ( n25632 & ~n25637 ) ;
  assign n25639 = n25635 | n25638 ;
  assign n25640 = n25631 ^ x781 ^ 1'b0 ;
  assign n25641 = ( n25631 & n25639 ) | ( n25631 & n25640 ) | ( n25639 & n25640 ) ;
  assign n25642 = x619 & ~n25641 ;
  assign n25643 = x619 | n25555 ;
  assign n25644 = ( x1159 & n25642 ) | ( x1159 & n25643 ) | ( n25642 & n25643 ) ;
  assign n25645 = ~n25642 & n25644 ;
  assign n25646 = x619 & ~n25555 ;
  assign n25647 = x1159 | n25646 ;
  assign n25648 = ( n25641 & n25642 ) | ( n25641 & ~n25647 ) | ( n25642 & ~n25647 ) ;
  assign n25649 = n25645 | n25648 ;
  assign n25650 = n25641 ^ x789 ^ 1'b0 ;
  assign n25651 = ( n25641 & n25649 ) | ( n25641 & n25650 ) | ( n25649 & n25650 ) ;
  assign n25652 = n25555 ^ n16518 ^ 1'b0 ;
  assign n25653 = ( n25555 & n25651 ) | ( n25555 & ~n25652 ) | ( n25651 & ~n25652 ) ;
  assign n25654 = n25555 ^ n16339 ^ 1'b0 ;
  assign n25655 = ( n25555 & n25653 ) | ( n25555 & ~n25654 ) | ( n25653 & ~n25654 ) ;
  assign n25656 = n25555 ^ n16376 ^ 1'b0 ;
  assign n25657 = ( n25555 & n25655 ) | ( n25555 & ~n25656 ) | ( n25655 & ~n25656 ) ;
  assign n25658 = x644 | n25657 ;
  assign n25659 = ( n25606 & ~n25607 ) | ( n25606 & n25658 ) | ( ~n25607 & n25658 ) ;
  assign n25660 = ( x1160 & n25607 ) | ( x1160 & n25659 ) | ( n25607 & n25659 ) ;
  assign n25661 = n25604 & ~n25660 ;
  assign n25662 = x644 & ~n25657 ;
  assign n25663 = ( ~x715 & n25555 ) | ( ~x715 & n25605 ) | ( n25555 & n25605 ) ;
  assign n25664 = x1160 & ~n25663 ;
  assign n25665 = ( x1160 & n25662 ) | ( x1160 & n25664 ) | ( n25662 & n25664 ) ;
  assign n25666 = ( x715 & n25602 ) | ( x715 & n25603 ) | ( n25602 & n25603 ) ;
  assign n25667 = n25665 & ~n25666 ;
  assign n25668 = ( x790 & n25661 ) | ( x790 & n25667 ) | ( n25661 & n25667 ) ;
  assign n25669 = n25667 ^ n25661 ^ 1'b0 ;
  assign n25670 = ( x790 & n25668 ) | ( x790 & n25669 ) | ( n25668 & n25669 ) ;
  assign n25671 = n19055 & n25655 ;
  assign n25672 = n16374 & n25597 ;
  assign n25673 = n16373 & n25598 ;
  assign n25674 = n25672 | n25673 ;
  assign n25675 = ( x787 & n25671 ) | ( x787 & n25674 ) | ( n25671 & n25674 ) ;
  assign n25676 = n25674 ^ n25671 ^ 1'b0 ;
  assign n25677 = ( x787 & n25675 ) | ( x787 & n25676 ) | ( n25675 & n25676 ) ;
  assign n25678 = x725 & ~n25618 ;
  assign n25679 = x183 & ~n16054 ;
  assign n25680 = ~x183 & n16048 ;
  assign n25681 = ( x755 & ~n25679 ) | ( x755 & n25680 ) | ( ~n25679 & n25680 ) ;
  assign n25682 = n25679 | n25681 ;
  assign n25683 = ~x183 & n16044 ;
  assign n25684 = x183 & ~n16029 ;
  assign n25685 = ( x755 & n25683 ) | ( x755 & ~n25684 ) | ( n25683 & ~n25684 ) ;
  assign n25686 = ~n25683 & n25685 ;
  assign n25687 = ( x39 & n25682 ) | ( x39 & ~n25686 ) | ( n25682 & ~n25686 ) ;
  assign n25688 = n25687 ^ n25682 ^ 1'b0 ;
  assign n25689 = ( x39 & n25687 ) | ( x39 & ~n25688 ) | ( n25687 & ~n25688 ) ;
  assign n25690 = x183 & n15795 ;
  assign n25691 = x755 & ~n25690 ;
  assign n25692 = x183 | n15876 ;
  assign n25693 = n25691 & n25692 ;
  assign n25694 = x183 & n15943 ;
  assign n25695 = x183 | n16003 ;
  assign n25696 = ( x755 & ~n25694 ) | ( x755 & n25695 ) | ( ~n25694 & n25695 ) ;
  assign n25697 = ~x755 & n25696 ;
  assign n25698 = ( x39 & n25693 ) | ( x39 & ~n25697 ) | ( n25693 & ~n25697 ) ;
  assign n25699 = ~n25693 & n25698 ;
  assign n25700 = ( x38 & n25689 ) | ( x38 & ~n25699 ) | ( n25689 & ~n25699 ) ;
  assign n25701 = ~x38 & n25700 ;
  assign n25702 = ~x755 & n15591 ;
  assign n25703 = n17156 | n25702 ;
  assign n25704 = x183 & ~n5017 ;
  assign n25705 = n25703 & n25704 ;
  assign n25706 = x38 & ~n25705 ;
  assign n25707 = n25706 ^ x725 ^ 1'b0 ;
  assign n25708 = x755 | n15968 ;
  assign n25709 = n17889 & n25708 ;
  assign n25710 = x183 | n25709 ;
  assign n25711 = ( n25706 & ~n25707 ) | ( n25706 & n25710 ) | ( ~n25707 & n25710 ) ;
  assign n25712 = ( x725 & n25707 ) | ( x725 & n25711 ) | ( n25707 & n25711 ) ;
  assign n25713 = ( ~n2069 & n25701 ) | ( ~n2069 & n25712 ) | ( n25701 & n25712 ) ;
  assign n25714 = ~n2069 & n25713 ;
  assign n25715 = n25714 ^ n25678 ^ 1'b0 ;
  assign n25716 = ( n25678 & n25714 ) | ( n25678 & n25715 ) | ( n25714 & n25715 ) ;
  assign n25717 = ( n25620 & ~n25678 ) | ( n25620 & n25716 ) | ( ~n25678 & n25716 ) ;
  assign n25718 = x625 & ~n25717 ;
  assign n25719 = x625 | n25621 ;
  assign n25720 = ( x1153 & n25718 ) | ( x1153 & n25719 ) | ( n25718 & n25719 ) ;
  assign n25721 = ~n25718 & n25720 ;
  assign n25722 = ( x608 & n25574 ) | ( x608 & ~n25721 ) | ( n25574 & ~n25721 ) ;
  assign n25723 = ~n25574 & n25722 ;
  assign n25724 = x608 | n25570 ;
  assign n25725 = x625 & ~n25621 ;
  assign n25726 = x1153 | n25725 ;
  assign n25727 = ( n25717 & n25718 ) | ( n25717 & ~n25726 ) | ( n25718 & ~n25726 ) ;
  assign n25728 = ( ~n25723 & n25724 ) | ( ~n25723 & n25727 ) | ( n25724 & n25727 ) ;
  assign n25729 = ~n25723 & n25728 ;
  assign n25730 = n25717 ^ x778 ^ 1'b0 ;
  assign n25731 = ( n25717 & n25729 ) | ( n25717 & n25730 ) | ( n25729 & n25730 ) ;
  assign n25732 = x609 & ~n25731 ;
  assign n25733 = x609 | n25577 ;
  assign n25734 = ( x1155 & n25732 ) | ( x1155 & n25733 ) | ( n25732 & n25733 ) ;
  assign n25735 = ~n25732 & n25734 ;
  assign n25736 = ~x1155 & n25626 ;
  assign n25737 = ( x660 & n25735 ) | ( x660 & ~n25736 ) | ( n25735 & ~n25736 ) ;
  assign n25738 = ~n25735 & n25737 ;
  assign n25739 = x1155 & n25627 ;
  assign n25740 = x660 | n25739 ;
  assign n25741 = x609 & ~n25577 ;
  assign n25742 = x1155 | n25741 ;
  assign n25743 = ( n25731 & n25732 ) | ( n25731 & ~n25742 ) | ( n25732 & ~n25742 ) ;
  assign n25744 = ( ~n25738 & n25740 ) | ( ~n25738 & n25743 ) | ( n25740 & n25743 ) ;
  assign n25745 = ~n25738 & n25744 ;
  assign n25746 = n25731 ^ x785 ^ 1'b0 ;
  assign n25747 = ( n25731 & n25745 ) | ( n25731 & n25746 ) | ( n25745 & n25746 ) ;
  assign n25748 = x618 & ~n25747 ;
  assign n25749 = x618 | n25579 ;
  assign n25750 = ( x1154 & n25748 ) | ( x1154 & n25749 ) | ( n25748 & n25749 ) ;
  assign n25751 = ~n25748 & n25750 ;
  assign n25752 = ( x627 & n25638 ) | ( x627 & ~n25751 ) | ( n25638 & ~n25751 ) ;
  assign n25753 = ~n25638 & n25752 ;
  assign n25754 = x627 | n25635 ;
  assign n25755 = x618 & ~n25579 ;
  assign n25756 = x1154 | n25755 ;
  assign n25757 = ( n25747 & n25748 ) | ( n25747 & ~n25756 ) | ( n25748 & ~n25756 ) ;
  assign n25758 = ( ~n25753 & n25754 ) | ( ~n25753 & n25757 ) | ( n25754 & n25757 ) ;
  assign n25759 = ~n25753 & n25758 ;
  assign n25760 = n25747 ^ x781 ^ 1'b0 ;
  assign n25761 = ( n25747 & n25759 ) | ( n25747 & n25760 ) | ( n25759 & n25760 ) ;
  assign n25762 = x619 | n25761 ;
  assign n25763 = x619 & ~n25581 ;
  assign n25764 = ( x1159 & n25762 ) | ( x1159 & ~n25763 ) | ( n25762 & ~n25763 ) ;
  assign n25765 = ~x1159 & n25764 ;
  assign n25766 = ( x648 & n25645 ) | ( x648 & ~n25765 ) | ( n25645 & ~n25765 ) ;
  assign n25767 = n25765 | n25766 ;
  assign n25768 = x619 & ~n25761 ;
  assign n25769 = x619 | n25581 ;
  assign n25770 = ( x1159 & n25768 ) | ( x1159 & n25769 ) | ( n25768 & n25769 ) ;
  assign n25771 = ~n25768 & n25770 ;
  assign n25772 = ( x648 & n25648 ) | ( x648 & ~n25771 ) | ( n25648 & ~n25771 ) ;
  assign n25773 = ~n25648 & n25772 ;
  assign n25774 = x789 & ~n25773 ;
  assign n25775 = n25767 & n25774 ;
  assign n25776 = ~x789 & n25761 ;
  assign n25777 = ( n16519 & ~n25775 ) | ( n16519 & n25776 ) | ( ~n25775 & n25776 ) ;
  assign n25778 = n25775 | n25777 ;
  assign n25779 = n25589 ^ x629 ^ 1'b0 ;
  assign n25780 = ( n25589 & n25592 ) | ( n25589 & n25779 ) | ( n25592 & n25779 ) ;
  assign n25781 = n19046 & n25653 ;
  assign n25782 = ( x792 & n25780 ) | ( x792 & n25781 ) | ( n25780 & n25781 ) ;
  assign n25783 = n25781 ^ n25780 ^ 1'b0 ;
  assign n25784 = ( x792 & n25782 ) | ( x792 & n25783 ) | ( n25782 & n25783 ) ;
  assign n25785 = n16459 & ~n25583 ;
  assign n25786 = ~x626 & n25555 ;
  assign n25787 = x626 & n25651 ;
  assign n25788 = ( n22317 & n25786 ) | ( n22317 & ~n25787 ) | ( n25786 & ~n25787 ) ;
  assign n25789 = ~n25786 & n25788 ;
  assign n25790 = ~x626 & n25651 ;
  assign n25791 = x626 & n25555 ;
  assign n25792 = ( n22322 & n25790 ) | ( n22322 & ~n25791 ) | ( n25790 & ~n25791 ) ;
  assign n25793 = ~n25790 & n25792 ;
  assign n25794 = ( ~n25785 & n25789 ) | ( ~n25785 & n25793 ) | ( n25789 & n25793 ) ;
  assign n25795 = n25785 | n25794 ;
  assign n25796 = ( x788 & ~n22314 ) | ( x788 & n25795 ) | ( ~n22314 & n25795 ) ;
  assign n25797 = ( n18482 & n22314 ) | ( n18482 & n25796 ) | ( n22314 & n25796 ) ;
  assign n25798 = ~n25784 & n25797 ;
  assign n25799 = ( n25778 & n25784 ) | ( n25778 & ~n25798 ) | ( n25784 & ~n25798 ) ;
  assign n25800 = ( ~n18484 & n25677 ) | ( ~n18484 & n25799 ) | ( n25677 & n25799 ) ;
  assign n25801 = n25677 ^ n18484 ^ 1'b0 ;
  assign n25802 = ( n25677 & n25800 ) | ( n25677 & ~n25801 ) | ( n25800 & ~n25801 ) ;
  assign n25803 = x644 | n25660 ;
  assign n25804 = x644 & n25665 ;
  assign n25805 = x790 & ~n25804 ;
  assign n25806 = n25803 & n25805 ;
  assign n25807 = ( ~n25670 & n25802 ) | ( ~n25670 & n25806 ) | ( n25802 & n25806 ) ;
  assign n25808 = ~n25670 & n25807 ;
  assign n25809 = ( x57 & n5193 ) | ( x57 & ~n25808 ) | ( n5193 & ~n25808 ) ;
  assign n25810 = n25808 | n25809 ;
  assign n25811 = x183 | n1611 ;
  assign n25812 = ~n25702 & n25811 ;
  assign n25813 = n16397 | n25812 ;
  assign n25814 = ~n15662 & n25702 ;
  assign n25815 = ~x1155 & n25811 ;
  assign n25816 = ~n25814 & n25815 ;
  assign n25817 = ( x1155 & n25813 ) | ( x1155 & n25814 ) | ( n25813 & n25814 ) ;
  assign n25818 = n25816 | n25817 ;
  assign n25819 = n25813 ^ x785 ^ 1'b0 ;
  assign n25820 = ( n25813 & n25818 ) | ( n25813 & n25819 ) | ( n25818 & n25819 ) ;
  assign n25821 = n16411 | n25820 ;
  assign n25822 = x1154 & n25821 ;
  assign n25823 = n16414 | n25820 ;
  assign n25824 = ~x1154 & n25823 ;
  assign n25825 = n25822 | n25824 ;
  assign n25826 = n25820 ^ x781 ^ 1'b0 ;
  assign n25827 = ( n25820 & n25825 ) | ( n25820 & n25826 ) | ( n25825 & n25826 ) ;
  assign n25828 = n21437 | n25827 ;
  assign n25829 = x1159 & n25828 ;
  assign n25830 = n21440 | n25827 ;
  assign n25831 = ~x1159 & n25830 ;
  assign n25832 = n25829 | n25831 ;
  assign n25833 = n25827 ^ x789 ^ 1'b0 ;
  assign n25834 = ( n25827 & n25832 ) | ( n25827 & n25833 ) | ( n25832 & n25833 ) ;
  assign n25835 = n25811 ^ n16518 ^ 1'b0 ;
  assign n25836 = ( n25811 & n25834 ) | ( n25811 & ~n25835 ) | ( n25834 & ~n25835 ) ;
  assign n25837 = n25811 ^ n16339 ^ 1'b0 ;
  assign n25838 = ( n25811 & n25836 ) | ( n25811 & ~n25837 ) | ( n25836 & ~n25837 ) ;
  assign n25839 = n19055 & n25838 ;
  assign n25840 = x647 & ~n25811 ;
  assign n25841 = x1157 | n25840 ;
  assign n25842 = ~x725 & n15778 ;
  assign n25843 = ~x625 & n25842 ;
  assign n25844 = ~x1153 & n25811 ;
  assign n25845 = ~n25843 & n25844 ;
  assign n25846 = x778 & ~n25845 ;
  assign n25847 = n25811 & ~n25842 ;
  assign n25848 = ( x1153 & n25843 ) | ( x1153 & n25847 ) | ( n25843 & n25847 ) ;
  assign n25849 = n25846 & ~n25848 ;
  assign n25850 = ( x778 & n25847 ) | ( x778 & ~n25849 ) | ( n25847 & ~n25849 ) ;
  assign n25851 = ~n25849 & n25850 ;
  assign n25852 = n16447 | n25851 ;
  assign n25853 = n16449 | n25852 ;
  assign n25854 = n16451 | n25853 ;
  assign n25855 = n16530 | n25854 ;
  assign n25856 = n16560 | n25855 ;
  assign n25857 = ( x647 & ~n25841 ) | ( x647 & n25856 ) | ( ~n25841 & n25856 ) ;
  assign n25858 = ~n25841 & n25857 ;
  assign n25859 = n25811 ^ x647 ^ 1'b0 ;
  assign n25860 = ( n25811 & n25856 ) | ( n25811 & n25859 ) | ( n25856 & n25859 ) ;
  assign n25861 = x1157 & n25860 ;
  assign n25862 = ( n16375 & n25858 ) | ( n16375 & n25861 ) | ( n25858 & n25861 ) ;
  assign n25863 = ( x787 & n25839 ) | ( x787 & n25862 ) | ( n25839 & n25862 ) ;
  assign n25864 = n25862 ^ n25839 ^ 1'b0 ;
  assign n25865 = ( x787 & n25863 ) | ( x787 & n25864 ) | ( n25863 & n25864 ) ;
  assign n25866 = ~x626 & n25811 ;
  assign n25867 = x626 & n25834 ;
  assign n25868 = ( n22317 & n25866 ) | ( n22317 & ~n25867 ) | ( n25866 & ~n25867 ) ;
  assign n25869 = ~n25866 & n25868 ;
  assign n25870 = ~x626 & n25834 ;
  assign n25871 = x626 & n25811 ;
  assign n25872 = ( n22322 & n25870 ) | ( n22322 & ~n25871 ) | ( n25870 & ~n25871 ) ;
  assign n25873 = ~n25870 & n25872 ;
  assign n25874 = n25854 & ~n25873 ;
  assign n25875 = ( n16459 & n25873 ) | ( n16459 & ~n25874 ) | ( n25873 & ~n25874 ) ;
  assign n25876 = ( x788 & n25869 ) | ( x788 & n25875 ) | ( n25869 & n25875 ) ;
  assign n25877 = n25875 ^ n25869 ^ 1'b0 ;
  assign n25878 = ( x788 & n25876 ) | ( x788 & n25877 ) | ( n25876 & n25877 ) ;
  assign n25879 = n15524 | n25847 ;
  assign n25880 = n25812 & n25879 ;
  assign n25881 = x625 & ~n25879 ;
  assign n25882 = ( n25844 & n25880 ) | ( n25844 & n25881 ) | ( n25880 & n25881 ) ;
  assign n25883 = ( x608 & n25848 ) | ( x608 & ~n25882 ) | ( n25848 & ~n25882 ) ;
  assign n25884 = n25882 | n25883 ;
  assign n25885 = x1153 & n25812 ;
  assign n25886 = ~n25881 & n25885 ;
  assign n25887 = x608 & ~n25845 ;
  assign n25888 = n25884 & ~n25887 ;
  assign n25889 = ( n25884 & n25886 ) | ( n25884 & n25888 ) | ( n25886 & n25888 ) ;
  assign n25890 = n25880 ^ x778 ^ 1'b0 ;
  assign n25891 = ( n25880 & n25889 ) | ( n25880 & n25890 ) | ( n25889 & n25890 ) ;
  assign n25892 = x609 & ~n25891 ;
  assign n25898 = x609 | n25851 ;
  assign n25899 = ( x1155 & n25892 ) | ( x1155 & n25898 ) | ( n25892 & n25898 ) ;
  assign n25900 = ~n25892 & n25899 ;
  assign n25901 = ( x660 & n25816 ) | ( x660 & ~n25900 ) | ( n25816 & ~n25900 ) ;
  assign n25902 = ~n25816 & n25901 ;
  assign n25893 = x609 & ~n25851 ;
  assign n25894 = x1155 | n25893 ;
  assign n25895 = ( n25891 & n25892 ) | ( n25891 & ~n25894 ) | ( n25892 & ~n25894 ) ;
  assign n25896 = ( x660 & n25817 ) | ( x660 & ~n25895 ) | ( n25817 & ~n25895 ) ;
  assign n25897 = n25895 | n25896 ;
  assign n25903 = n25902 ^ n25897 ^ 1'b0 ;
  assign n25904 = ( x785 & ~n25897 ) | ( x785 & n25902 ) | ( ~n25897 & n25902 ) ;
  assign n25905 = ( x785 & ~n25903 ) | ( x785 & n25904 ) | ( ~n25903 & n25904 ) ;
  assign n25906 = ( x785 & n25891 ) | ( x785 & ~n25905 ) | ( n25891 & ~n25905 ) ;
  assign n25907 = ~n25905 & n25906 ;
  assign n25908 = x618 & ~n25907 ;
  assign n25909 = x618 | n25852 ;
  assign n25910 = ( x1154 & n25908 ) | ( x1154 & n25909 ) | ( n25908 & n25909 ) ;
  assign n25911 = ~n25908 & n25910 ;
  assign n25912 = ( x627 & n25824 ) | ( x627 & ~n25911 ) | ( n25824 & ~n25911 ) ;
  assign n25913 = ~n25824 & n25912 ;
  assign n25914 = x627 | n25822 ;
  assign n25915 = x618 & ~n25852 ;
  assign n25916 = x1154 | n25915 ;
  assign n25917 = ( n25907 & n25908 ) | ( n25907 & ~n25916 ) | ( n25908 & ~n25916 ) ;
  assign n25918 = ( ~n25913 & n25914 ) | ( ~n25913 & n25917 ) | ( n25914 & n25917 ) ;
  assign n25919 = ~n25913 & n25918 ;
  assign n25920 = n25907 ^ x781 ^ 1'b0 ;
  assign n25921 = ( n25907 & n25919 ) | ( n25907 & n25920 ) | ( n25919 & n25920 ) ;
  assign n25922 = ~x789 & n25921 ;
  assign n25923 = x619 & ~n25853 ;
  assign n25924 = x1159 | n25923 ;
  assign n25925 = x619 & ~n25921 ;
  assign n25926 = ( n25921 & ~n25924 ) | ( n25921 & n25925 ) | ( ~n25924 & n25925 ) ;
  assign n25927 = ( x648 & n25829 ) | ( x648 & ~n25926 ) | ( n25829 & ~n25926 ) ;
  assign n25928 = n25926 | n25927 ;
  assign n25929 = x619 | n25853 ;
  assign n25930 = x1159 & ~n25925 ;
  assign n25931 = n25929 & n25930 ;
  assign n25932 = ( x648 & n25831 ) | ( x648 & ~n25931 ) | ( n25831 & ~n25931 ) ;
  assign n25933 = ~n25831 & n25932 ;
  assign n25934 = x789 & ~n25933 ;
  assign n25935 = n25928 & n25934 ;
  assign n25936 = ( n16519 & ~n25922 ) | ( n16519 & n25935 ) | ( ~n25922 & n25935 ) ;
  assign n25937 = n25922 | n25936 ;
  assign n25938 = n25937 ^ n25878 ^ 1'b0 ;
  assign n25939 = ( n25878 & n25937 ) | ( n25878 & n25938 ) | ( n25937 & n25938 ) ;
  assign n25940 = ( n18482 & ~n25878 ) | ( n18482 & n25939 ) | ( ~n25878 & n25939 ) ;
  assign n25941 = n19208 | n25855 ;
  assign n25942 = n16556 & ~n25836 ;
  assign n25943 = x629 & ~n25942 ;
  assign n25944 = n25941 & n25943 ;
  assign n25945 = n16557 & ~n25836 ;
  assign n25946 = n19212 & ~n25855 ;
  assign n25947 = n25945 | n25946 ;
  assign n25948 = ( x629 & ~n25944 ) | ( x629 & n25947 ) | ( ~n25944 & n25947 ) ;
  assign n25949 = ~n25944 & n25948 ;
  assign n25950 = ( x792 & ~n19206 ) | ( x792 & n25949 ) | ( ~n19206 & n25949 ) ;
  assign n25951 = ( n18484 & n19206 ) | ( n18484 & n25950 ) | ( n19206 & n25950 ) ;
  assign n25952 = ( n25865 & n25940 ) | ( n25865 & ~n25951 ) | ( n25940 & ~n25951 ) ;
  assign n25953 = n25952 ^ n25940 ^ 1'b0 ;
  assign n25954 = ( n25865 & n25952 ) | ( n25865 & ~n25953 ) | ( n25952 & ~n25953 ) ;
  assign n25955 = x790 | n25954 ;
  assign n25956 = x644 & ~n25954 ;
  assign n25957 = ( x787 & n25858 ) | ( x787 & ~n25861 ) | ( n25858 & ~n25861 ) ;
  assign n25958 = ~n25858 & n25957 ;
  assign n25959 = ( x787 & n25856 ) | ( x787 & ~n25958 ) | ( n25856 & ~n25958 ) ;
  assign n25960 = ~n25958 & n25959 ;
  assign n25961 = x644 | n25960 ;
  assign n25962 = ( x715 & n25956 ) | ( x715 & n25961 ) | ( n25956 & n25961 ) ;
  assign n25963 = ~n25956 & n25962 ;
  assign n25964 = x644 | n25811 ;
  assign n25965 = n25811 ^ n16376 ^ 1'b0 ;
  assign n25966 = ( n25811 & n25838 ) | ( n25811 & ~n25965 ) | ( n25838 & ~n25965 ) ;
  assign n25967 = x644 & ~n25966 ;
  assign n25968 = ( x715 & n25964 ) | ( x715 & ~n25967 ) | ( n25964 & ~n25967 ) ;
  assign n25969 = ~x715 & n25968 ;
  assign n25970 = ( x1160 & n25963 ) | ( x1160 & ~n25969 ) | ( n25963 & ~n25969 ) ;
  assign n25971 = ~n25963 & n25970 ;
  assign n25972 = x644 & ~n25811 ;
  assign n25973 = x715 & ~n25972 ;
  assign n25974 = ( n25966 & n25967 ) | ( n25966 & n25973 ) | ( n25967 & n25973 ) ;
  assign n25975 = x644 & ~n25960 ;
  assign n25976 = x715 | n25975 ;
  assign n25977 = ( n25954 & n25956 ) | ( n25954 & ~n25976 ) | ( n25956 & ~n25976 ) ;
  assign n25978 = ( x1160 & ~n25974 ) | ( x1160 & n25977 ) | ( ~n25974 & n25977 ) ;
  assign n25979 = n25974 | n25978 ;
  assign n25980 = x790 & ~n25979 ;
  assign n25981 = ( x790 & n25971 ) | ( x790 & n25980 ) | ( n25971 & n25980 ) ;
  assign n25982 = x832 & ~n25981 ;
  assign n25983 = n25955 & n25982 ;
  assign n25984 = ~x183 & n7318 ;
  assign n25985 = x832 | n25984 ;
  assign n25986 = ~n25983 & n25985 ;
  assign n25987 = ( n25810 & n25983 ) | ( n25810 & ~n25986 ) | ( n25983 & ~n25986 ) ;
  assign n25988 = x184 | n15656 ;
  assign n25989 = x737 | n2069 ;
  assign n25990 = ~n25988 & n25989 ;
  assign n25991 = ( x38 & x184 ) | ( x38 & n16700 ) | ( x184 & n16700 ) ;
  assign n25992 = ~n2069 & n25991 ;
  assign n25993 = ( x184 & n16697 ) | ( x184 & ~n25992 ) | ( n16697 & ~n25992 ) ;
  assign n25994 = ~n25992 & n25993 ;
  assign n25995 = x184 | n15644 ;
  assign n25996 = n16185 & n25995 ;
  assign n25997 = x737 | n25996 ;
  assign n25998 = ( ~n25990 & n25994 ) | ( ~n25990 & n25997 ) | ( n25994 & n25997 ) ;
  assign n25999 = ~n25990 & n25998 ;
  assign n26000 = x625 & ~n25999 ;
  assign n26001 = x625 | n25988 ;
  assign n26002 = ( x1153 & n26000 ) | ( x1153 & n26001 ) | ( n26000 & n26001 ) ;
  assign n26003 = ~n26000 & n26002 ;
  assign n26004 = x625 & ~n25988 ;
  assign n26005 = x1153 | n26004 ;
  assign n26006 = ( x625 & n25999 ) | ( x625 & ~n26005 ) | ( n25999 & ~n26005 ) ;
  assign n26007 = ~n26005 & n26006 ;
  assign n26008 = n26003 | n26007 ;
  assign n26009 = n25999 ^ x778 ^ 1'b0 ;
  assign n26010 = ( n25999 & n26008 ) | ( n25999 & n26009 ) | ( n26008 & n26009 ) ;
  assign n26011 = n25988 ^ n16234 ^ 1'b0 ;
  assign n26012 = ( n25988 & n26010 ) | ( n25988 & ~n26011 ) | ( n26010 & ~n26011 ) ;
  assign n26013 = n25988 ^ n16254 ^ 1'b0 ;
  assign n26014 = ( n25988 & n26012 ) | ( n25988 & ~n26013 ) | ( n26012 & ~n26013 ) ;
  assign n26015 = n25988 ^ n16279 ^ 1'b0 ;
  assign n26016 = ( n25988 & n26014 ) | ( n25988 & ~n26015 ) | ( n26014 & ~n26015 ) ;
  assign n26017 = n25988 ^ n16318 ^ 1'b0 ;
  assign n26018 = ( n25988 & n26016 ) | ( n25988 & ~n26017 ) | ( n26016 & ~n26017 ) ;
  assign n26019 = x628 & ~n26018 ;
  assign n26020 = x628 | n25988 ;
  assign n26021 = ( x1156 & n26019 ) | ( x1156 & n26020 ) | ( n26019 & n26020 ) ;
  assign n26022 = ~n26019 & n26021 ;
  assign n26023 = x628 & ~n25988 ;
  assign n26024 = x1156 | n26023 ;
  assign n26025 = ( n26018 & n26019 ) | ( n26018 & ~n26024 ) | ( n26019 & ~n26024 ) ;
  assign n26026 = n26022 | n26025 ;
  assign n26027 = n26018 ^ x792 ^ 1'b0 ;
  assign n26028 = ( n26018 & n26026 ) | ( n26018 & n26027 ) | ( n26026 & n26027 ) ;
  assign n26029 = n25988 ^ x647 ^ 1'b0 ;
  assign n26030 = ( n25988 & n26028 ) | ( n25988 & ~n26029 ) | ( n26028 & ~n26029 ) ;
  assign n26031 = ( n25988 & n26028 ) | ( n25988 & n26029 ) | ( n26028 & n26029 ) ;
  assign n26032 = n26030 ^ x1157 ^ 1'b0 ;
  assign n26033 = ( n26030 & n26031 ) | ( n26030 & n26032 ) | ( n26031 & n26032 ) ;
  assign n26034 = n26028 ^ x787 ^ 1'b0 ;
  assign n26035 = ( n26028 & n26033 ) | ( n26028 & n26034 ) | ( n26033 & n26034 ) ;
  assign n26036 = x644 & ~n26035 ;
  assign n26037 = x715 | n26036 ;
  assign n26038 = x644 & ~n25988 ;
  assign n26039 = x715 & ~n26038 ;
  assign n26040 = n26039 ^ x1160 ^ 1'b0 ;
  assign n26041 = ~x777 & n15646 ;
  assign n26042 = n25995 & ~n26041 ;
  assign n26043 = ~x184 & x777 ;
  assign n26044 = ~n15488 & n26043 ;
  assign n26045 = ~x184 & n15587 ;
  assign n26046 = x184 & ~n15640 ;
  assign n26047 = x777 | n26046 ;
  assign n26048 = ( ~n26044 & n26045 ) | ( ~n26044 & n26047 ) | ( n26045 & n26047 ) ;
  assign n26049 = ~n26044 & n26048 ;
  assign n26050 = n26042 ^ x38 ^ 1'b0 ;
  assign n26051 = ( n26042 & n26049 ) | ( n26042 & ~n26050 ) | ( n26049 & ~n26050 ) ;
  assign n26052 = ~n2069 & n26051 ;
  assign n26053 = x184 & n2069 ;
  assign n26054 = n26052 | n26053 ;
  assign n26055 = n25988 ^ n15659 ^ 1'b0 ;
  assign n26056 = ( n25988 & n26054 ) | ( n25988 & ~n26055 ) | ( n26054 & ~n26055 ) ;
  assign n26057 = n15662 & n25988 ;
  assign n26058 = ( ~n15662 & n26052 ) | ( ~n15662 & n26053 ) | ( n26052 & n26053 ) ;
  assign n26059 = n26057 | n26058 ;
  assign n26060 = n26059 ^ n26056 ^ n25988 ;
  assign n26061 = n26060 ^ x1155 ^ 1'b0 ;
  assign n26062 = ( n26059 & n26060 ) | ( n26059 & ~n26061 ) | ( n26060 & ~n26061 ) ;
  assign n26063 = n26056 ^ x785 ^ 1'b0 ;
  assign n26064 = ( n26056 & n26062 ) | ( n26056 & n26063 ) | ( n26062 & n26063 ) ;
  assign n26065 = x618 & ~n26064 ;
  assign n26066 = x618 | n25988 ;
  assign n26067 = ( x1154 & n26065 ) | ( x1154 & n26066 ) | ( n26065 & n26066 ) ;
  assign n26068 = ~n26065 & n26067 ;
  assign n26069 = x618 & ~n25988 ;
  assign n26070 = x1154 | n26069 ;
  assign n26071 = ( n26064 & n26065 ) | ( n26064 & ~n26070 ) | ( n26065 & ~n26070 ) ;
  assign n26072 = n26068 | n26071 ;
  assign n26073 = n26064 ^ x781 ^ 1'b0 ;
  assign n26074 = ( n26064 & n26072 ) | ( n26064 & n26073 ) | ( n26072 & n26073 ) ;
  assign n26075 = x619 & ~n26074 ;
  assign n26076 = x619 | n25988 ;
  assign n26077 = ( x1159 & n26075 ) | ( x1159 & n26076 ) | ( n26075 & n26076 ) ;
  assign n26078 = ~n26075 & n26077 ;
  assign n26079 = x619 & ~n25988 ;
  assign n26080 = x1159 | n26079 ;
  assign n26081 = ( n26074 & n26075 ) | ( n26074 & ~n26080 ) | ( n26075 & ~n26080 ) ;
  assign n26082 = n26078 | n26081 ;
  assign n26083 = n26074 ^ x789 ^ 1'b0 ;
  assign n26084 = ( n26074 & n26082 ) | ( n26074 & n26083 ) | ( n26082 & n26083 ) ;
  assign n26085 = n25988 ^ n16518 ^ 1'b0 ;
  assign n26086 = ( n25988 & n26084 ) | ( n25988 & ~n26085 ) | ( n26084 & ~n26085 ) ;
  assign n26087 = n25988 ^ n16339 ^ 1'b0 ;
  assign n26088 = ( n25988 & n26086 ) | ( n25988 & ~n26087 ) | ( n26086 & ~n26087 ) ;
  assign n26089 = n25988 ^ n16376 ^ 1'b0 ;
  assign n26090 = ( n25988 & n26088 ) | ( n25988 & ~n26089 ) | ( n26088 & ~n26089 ) ;
  assign n26091 = x644 | n26090 ;
  assign n26092 = ( n26039 & ~n26040 ) | ( n26039 & n26091 ) | ( ~n26040 & n26091 ) ;
  assign n26093 = ( x1160 & n26040 ) | ( x1160 & n26092 ) | ( n26040 & n26092 ) ;
  assign n26094 = n26037 & ~n26093 ;
  assign n26095 = x644 & ~n26090 ;
  assign n26096 = ( ~x715 & n25988 ) | ( ~x715 & n26038 ) | ( n25988 & n26038 ) ;
  assign n26097 = x1160 & ~n26096 ;
  assign n26098 = ( x1160 & n26095 ) | ( x1160 & n26097 ) | ( n26095 & n26097 ) ;
  assign n26099 = ( x715 & n26035 ) | ( x715 & n26036 ) | ( n26035 & n26036 ) ;
  assign n26100 = n26098 & ~n26099 ;
  assign n26101 = ( x790 & n26094 ) | ( x790 & n26100 ) | ( n26094 & n26100 ) ;
  assign n26102 = n26100 ^ n26094 ^ 1'b0 ;
  assign n26103 = ( x790 & n26101 ) | ( x790 & n26102 ) | ( n26101 & n26102 ) ;
  assign n26104 = n19055 & n26088 ;
  assign n26105 = n16374 & n26030 ;
  assign n26106 = n16373 & n26031 ;
  assign n26107 = n26105 | n26106 ;
  assign n26108 = ( x787 & n26104 ) | ( x787 & n26107 ) | ( n26104 & n26107 ) ;
  assign n26109 = n26107 ^ n26104 ^ 1'b0 ;
  assign n26110 = ( x787 & n26108 ) | ( x787 & n26109 ) | ( n26108 & n26109 ) ;
  assign n26111 = x737 & ~n26051 ;
  assign n26112 = x184 & ~n16054 ;
  assign n26113 = ~x184 & n16048 ;
  assign n26114 = ( x777 & ~n26112 ) | ( x777 & n26113 ) | ( ~n26112 & n26113 ) ;
  assign n26115 = n26112 | n26114 ;
  assign n26116 = ~x184 & n16044 ;
  assign n26117 = x184 & ~n16029 ;
  assign n26118 = ( x777 & n26116 ) | ( x777 & ~n26117 ) | ( n26116 & ~n26117 ) ;
  assign n26119 = ~n26116 & n26118 ;
  assign n26120 = ( x39 & n26115 ) | ( x39 & ~n26119 ) | ( n26115 & ~n26119 ) ;
  assign n26121 = n26120 ^ n26115 ^ 1'b0 ;
  assign n26122 = ( x39 & n26120 ) | ( x39 & ~n26121 ) | ( n26120 & ~n26121 ) ;
  assign n26123 = x184 & n15795 ;
  assign n26124 = x777 & ~n26123 ;
  assign n26125 = x184 | n15876 ;
  assign n26126 = n26124 & n26125 ;
  assign n26127 = x184 & n15943 ;
  assign n26128 = x184 | n16003 ;
  assign n26129 = ( x777 & ~n26127 ) | ( x777 & n26128 ) | ( ~n26127 & n26128 ) ;
  assign n26130 = ~x777 & n26129 ;
  assign n26131 = ( x39 & n26126 ) | ( x39 & ~n26130 ) | ( n26126 & ~n26130 ) ;
  assign n26132 = ~n26126 & n26131 ;
  assign n26133 = ( x38 & n26122 ) | ( x38 & ~n26132 ) | ( n26122 & ~n26132 ) ;
  assign n26134 = ~x38 & n26133 ;
  assign n26135 = ~x777 & n15591 ;
  assign n26136 = n17156 | n26135 ;
  assign n26137 = x184 & ~n5017 ;
  assign n26138 = n26136 & n26137 ;
  assign n26139 = x38 & ~n26138 ;
  assign n26140 = n26139 ^ x737 ^ 1'b0 ;
  assign n26141 = x777 | n15968 ;
  assign n26142 = n17889 & n26141 ;
  assign n26143 = x184 | n26142 ;
  assign n26144 = ( n26139 & ~n26140 ) | ( n26139 & n26143 ) | ( ~n26140 & n26143 ) ;
  assign n26145 = ( x737 & n26140 ) | ( x737 & n26144 ) | ( n26140 & n26144 ) ;
  assign n26146 = ( ~n2069 & n26134 ) | ( ~n2069 & n26145 ) | ( n26134 & n26145 ) ;
  assign n26147 = ~n2069 & n26146 ;
  assign n26148 = n26147 ^ n26111 ^ 1'b0 ;
  assign n26149 = ( n26111 & n26147 ) | ( n26111 & n26148 ) | ( n26147 & n26148 ) ;
  assign n26150 = ( n26053 & ~n26111 ) | ( n26053 & n26149 ) | ( ~n26111 & n26149 ) ;
  assign n26151 = x625 & ~n26150 ;
  assign n26152 = x625 | n26054 ;
  assign n26153 = ( x1153 & n26151 ) | ( x1153 & n26152 ) | ( n26151 & n26152 ) ;
  assign n26154 = ~n26151 & n26153 ;
  assign n26155 = ( x608 & n26007 ) | ( x608 & ~n26154 ) | ( n26007 & ~n26154 ) ;
  assign n26156 = ~n26007 & n26155 ;
  assign n26157 = x608 | n26003 ;
  assign n26158 = x625 & ~n26054 ;
  assign n26159 = x1153 | n26158 ;
  assign n26160 = ( n26150 & n26151 ) | ( n26150 & ~n26159 ) | ( n26151 & ~n26159 ) ;
  assign n26161 = ( ~n26156 & n26157 ) | ( ~n26156 & n26160 ) | ( n26157 & n26160 ) ;
  assign n26162 = ~n26156 & n26161 ;
  assign n26163 = n26150 ^ x778 ^ 1'b0 ;
  assign n26164 = ( n26150 & n26162 ) | ( n26150 & n26163 ) | ( n26162 & n26163 ) ;
  assign n26165 = x609 & ~n26164 ;
  assign n26166 = x609 | n26010 ;
  assign n26167 = ( x1155 & n26165 ) | ( x1155 & n26166 ) | ( n26165 & n26166 ) ;
  assign n26168 = ~n26165 & n26167 ;
  assign n26169 = ~x1155 & n26059 ;
  assign n26170 = ( x660 & n26168 ) | ( x660 & ~n26169 ) | ( n26168 & ~n26169 ) ;
  assign n26171 = ~n26168 & n26170 ;
  assign n26172 = x1155 & n26060 ;
  assign n26173 = x660 | n26172 ;
  assign n26174 = x609 & ~n26010 ;
  assign n26175 = x1155 | n26174 ;
  assign n26176 = ( n26164 & n26165 ) | ( n26164 & ~n26175 ) | ( n26165 & ~n26175 ) ;
  assign n26177 = ( ~n26171 & n26173 ) | ( ~n26171 & n26176 ) | ( n26173 & n26176 ) ;
  assign n26178 = ~n26171 & n26177 ;
  assign n26179 = n26164 ^ x785 ^ 1'b0 ;
  assign n26180 = ( n26164 & n26178 ) | ( n26164 & n26179 ) | ( n26178 & n26179 ) ;
  assign n26181 = x618 & ~n26180 ;
  assign n26182 = x618 | n26012 ;
  assign n26183 = ( x1154 & n26181 ) | ( x1154 & n26182 ) | ( n26181 & n26182 ) ;
  assign n26184 = ~n26181 & n26183 ;
  assign n26185 = ( x627 & n26071 ) | ( x627 & ~n26184 ) | ( n26071 & ~n26184 ) ;
  assign n26186 = ~n26071 & n26185 ;
  assign n26187 = x627 | n26068 ;
  assign n26188 = x618 & ~n26012 ;
  assign n26189 = x1154 | n26188 ;
  assign n26190 = ( n26180 & n26181 ) | ( n26180 & ~n26189 ) | ( n26181 & ~n26189 ) ;
  assign n26191 = ( ~n26186 & n26187 ) | ( ~n26186 & n26190 ) | ( n26187 & n26190 ) ;
  assign n26192 = ~n26186 & n26191 ;
  assign n26193 = n26180 ^ x781 ^ 1'b0 ;
  assign n26194 = ( n26180 & n26192 ) | ( n26180 & n26193 ) | ( n26192 & n26193 ) ;
  assign n26195 = x619 | n26194 ;
  assign n26196 = x619 & ~n26014 ;
  assign n26197 = ( x1159 & n26195 ) | ( x1159 & ~n26196 ) | ( n26195 & ~n26196 ) ;
  assign n26198 = ~x1159 & n26197 ;
  assign n26199 = ( x648 & n26078 ) | ( x648 & ~n26198 ) | ( n26078 & ~n26198 ) ;
  assign n26200 = n26198 | n26199 ;
  assign n26201 = x619 & ~n26194 ;
  assign n26202 = x619 | n26014 ;
  assign n26203 = ( x1159 & n26201 ) | ( x1159 & n26202 ) | ( n26201 & n26202 ) ;
  assign n26204 = ~n26201 & n26203 ;
  assign n26205 = ( x648 & n26081 ) | ( x648 & ~n26204 ) | ( n26081 & ~n26204 ) ;
  assign n26206 = ~n26081 & n26205 ;
  assign n26207 = x789 & ~n26206 ;
  assign n26208 = n26200 & n26207 ;
  assign n26209 = ~x789 & n26194 ;
  assign n26210 = ( n16519 & ~n26208 ) | ( n16519 & n26209 ) | ( ~n26208 & n26209 ) ;
  assign n26211 = n26208 | n26210 ;
  assign n26212 = n26022 ^ x629 ^ 1'b0 ;
  assign n26213 = ( n26022 & n26025 ) | ( n26022 & n26212 ) | ( n26025 & n26212 ) ;
  assign n26214 = n19046 & n26086 ;
  assign n26215 = ( x792 & n26213 ) | ( x792 & n26214 ) | ( n26213 & n26214 ) ;
  assign n26216 = n26214 ^ n26213 ^ 1'b0 ;
  assign n26217 = ( x792 & n26215 ) | ( x792 & n26216 ) | ( n26215 & n26216 ) ;
  assign n26218 = n16459 & ~n26016 ;
  assign n26219 = ~x626 & n25988 ;
  assign n26220 = x626 & n26084 ;
  assign n26221 = ( n22317 & n26219 ) | ( n22317 & ~n26220 ) | ( n26219 & ~n26220 ) ;
  assign n26222 = ~n26219 & n26221 ;
  assign n26223 = ~x626 & n26084 ;
  assign n26224 = x626 & n25988 ;
  assign n26225 = ( n22322 & n26223 ) | ( n22322 & ~n26224 ) | ( n26223 & ~n26224 ) ;
  assign n26226 = ~n26223 & n26225 ;
  assign n26227 = ( ~n26218 & n26222 ) | ( ~n26218 & n26226 ) | ( n26222 & n26226 ) ;
  assign n26228 = n26218 | n26227 ;
  assign n26229 = ( x788 & ~n22314 ) | ( x788 & n26228 ) | ( ~n22314 & n26228 ) ;
  assign n26230 = ( n18482 & n22314 ) | ( n18482 & n26229 ) | ( n22314 & n26229 ) ;
  assign n26231 = ~n26217 & n26230 ;
  assign n26232 = ( n26211 & n26217 ) | ( n26211 & ~n26231 ) | ( n26217 & ~n26231 ) ;
  assign n26233 = ( ~n18484 & n26110 ) | ( ~n18484 & n26232 ) | ( n26110 & n26232 ) ;
  assign n26234 = n26110 ^ n18484 ^ 1'b0 ;
  assign n26235 = ( n26110 & n26233 ) | ( n26110 & ~n26234 ) | ( n26233 & ~n26234 ) ;
  assign n26236 = x644 | n26093 ;
  assign n26237 = x644 & n26098 ;
  assign n26238 = x790 & ~n26237 ;
  assign n26239 = n26236 & n26238 ;
  assign n26240 = ( ~n26103 & n26235 ) | ( ~n26103 & n26239 ) | ( n26235 & n26239 ) ;
  assign n26241 = ~n26103 & n26240 ;
  assign n26242 = ( x57 & n5193 ) | ( x57 & ~n26241 ) | ( n5193 & ~n26241 ) ;
  assign n26243 = n26241 | n26242 ;
  assign n26244 = x184 | n1611 ;
  assign n26245 = ~n26135 & n26244 ;
  assign n26246 = n16397 | n26245 ;
  assign n26247 = ~n15662 & n26135 ;
  assign n26248 = ~x1155 & n26244 ;
  assign n26249 = ~n26247 & n26248 ;
  assign n26250 = ( x1155 & n26246 ) | ( x1155 & n26247 ) | ( n26246 & n26247 ) ;
  assign n26251 = n26249 | n26250 ;
  assign n26252 = n26246 ^ x785 ^ 1'b0 ;
  assign n26253 = ( n26246 & n26251 ) | ( n26246 & n26252 ) | ( n26251 & n26252 ) ;
  assign n26254 = n16411 | n26253 ;
  assign n26255 = x1154 & n26254 ;
  assign n26256 = n16414 | n26253 ;
  assign n26257 = ~x1154 & n26256 ;
  assign n26258 = n26255 | n26257 ;
  assign n26259 = n26253 ^ x781 ^ 1'b0 ;
  assign n26260 = ( n26253 & n26258 ) | ( n26253 & n26259 ) | ( n26258 & n26259 ) ;
  assign n26261 = n21437 | n26260 ;
  assign n26262 = x1159 & n26261 ;
  assign n26263 = n21440 | n26260 ;
  assign n26264 = ~x1159 & n26263 ;
  assign n26265 = n26262 | n26264 ;
  assign n26266 = n26260 ^ x789 ^ 1'b0 ;
  assign n26267 = ( n26260 & n26265 ) | ( n26260 & n26266 ) | ( n26265 & n26266 ) ;
  assign n26268 = n26244 ^ n16518 ^ 1'b0 ;
  assign n26269 = ( n26244 & n26267 ) | ( n26244 & ~n26268 ) | ( n26267 & ~n26268 ) ;
  assign n26270 = n26244 ^ n16339 ^ 1'b0 ;
  assign n26271 = ( n26244 & n26269 ) | ( n26244 & ~n26270 ) | ( n26269 & ~n26270 ) ;
  assign n26272 = n19055 & n26271 ;
  assign n26273 = x647 & ~n26244 ;
  assign n26274 = x1157 | n26273 ;
  assign n26275 = ~x737 & n15778 ;
  assign n26276 = ~x625 & n26275 ;
  assign n26277 = ~x1153 & n26244 ;
  assign n26278 = ~n26276 & n26277 ;
  assign n26279 = x778 & ~n26278 ;
  assign n26280 = n26244 & ~n26275 ;
  assign n26281 = ( x1153 & n26276 ) | ( x1153 & n26280 ) | ( n26276 & n26280 ) ;
  assign n26282 = n26279 & ~n26281 ;
  assign n26283 = ( x778 & n26280 ) | ( x778 & ~n26282 ) | ( n26280 & ~n26282 ) ;
  assign n26284 = ~n26282 & n26283 ;
  assign n26285 = n16447 | n26284 ;
  assign n26286 = n16449 | n26285 ;
  assign n26287 = n16451 | n26286 ;
  assign n26288 = n16530 | n26287 ;
  assign n26289 = n16560 | n26288 ;
  assign n26290 = ( x647 & ~n26274 ) | ( x647 & n26289 ) | ( ~n26274 & n26289 ) ;
  assign n26291 = ~n26274 & n26290 ;
  assign n26292 = n26244 ^ x647 ^ 1'b0 ;
  assign n26293 = ( n26244 & n26289 ) | ( n26244 & n26292 ) | ( n26289 & n26292 ) ;
  assign n26294 = x1157 & n26293 ;
  assign n26295 = ( n16375 & n26291 ) | ( n16375 & n26294 ) | ( n26291 & n26294 ) ;
  assign n26296 = ( x787 & n26272 ) | ( x787 & n26295 ) | ( n26272 & n26295 ) ;
  assign n26297 = n26295 ^ n26272 ^ 1'b0 ;
  assign n26298 = ( x787 & n26296 ) | ( x787 & n26297 ) | ( n26296 & n26297 ) ;
  assign n26299 = ~x626 & n26244 ;
  assign n26300 = x626 & n26267 ;
  assign n26301 = ( n22317 & n26299 ) | ( n22317 & ~n26300 ) | ( n26299 & ~n26300 ) ;
  assign n26302 = ~n26299 & n26301 ;
  assign n26303 = ~x626 & n26267 ;
  assign n26304 = x626 & n26244 ;
  assign n26305 = ( n22322 & n26303 ) | ( n22322 & ~n26304 ) | ( n26303 & ~n26304 ) ;
  assign n26306 = ~n26303 & n26305 ;
  assign n26307 = n26287 & ~n26306 ;
  assign n26308 = ( n16459 & n26306 ) | ( n16459 & ~n26307 ) | ( n26306 & ~n26307 ) ;
  assign n26309 = ( x788 & n26302 ) | ( x788 & n26308 ) | ( n26302 & n26308 ) ;
  assign n26310 = n26308 ^ n26302 ^ 1'b0 ;
  assign n26311 = ( x788 & n26309 ) | ( x788 & n26310 ) | ( n26309 & n26310 ) ;
  assign n26312 = n15524 | n26280 ;
  assign n26313 = n26245 & n26312 ;
  assign n26314 = x625 & ~n26312 ;
  assign n26315 = ( n26277 & n26313 ) | ( n26277 & n26314 ) | ( n26313 & n26314 ) ;
  assign n26316 = ( x608 & n26281 ) | ( x608 & ~n26315 ) | ( n26281 & ~n26315 ) ;
  assign n26317 = n26315 | n26316 ;
  assign n26318 = x1153 & n26245 ;
  assign n26319 = ~n26314 & n26318 ;
  assign n26320 = x608 & ~n26278 ;
  assign n26321 = n26317 & ~n26320 ;
  assign n26322 = ( n26317 & n26319 ) | ( n26317 & n26321 ) | ( n26319 & n26321 ) ;
  assign n26323 = n26313 ^ x778 ^ 1'b0 ;
  assign n26324 = ( n26313 & n26322 ) | ( n26313 & n26323 ) | ( n26322 & n26323 ) ;
  assign n26325 = x609 & ~n26324 ;
  assign n26331 = x609 | n26284 ;
  assign n26332 = ( x1155 & n26325 ) | ( x1155 & n26331 ) | ( n26325 & n26331 ) ;
  assign n26333 = ~n26325 & n26332 ;
  assign n26334 = ( x660 & n26249 ) | ( x660 & ~n26333 ) | ( n26249 & ~n26333 ) ;
  assign n26335 = ~n26249 & n26334 ;
  assign n26326 = x609 & ~n26284 ;
  assign n26327 = x1155 | n26326 ;
  assign n26328 = ( n26324 & n26325 ) | ( n26324 & ~n26327 ) | ( n26325 & ~n26327 ) ;
  assign n26329 = ( x660 & n26250 ) | ( x660 & ~n26328 ) | ( n26250 & ~n26328 ) ;
  assign n26330 = n26328 | n26329 ;
  assign n26336 = n26335 ^ n26330 ^ 1'b0 ;
  assign n26337 = ( x785 & ~n26330 ) | ( x785 & n26335 ) | ( ~n26330 & n26335 ) ;
  assign n26338 = ( x785 & ~n26336 ) | ( x785 & n26337 ) | ( ~n26336 & n26337 ) ;
  assign n26339 = ( x785 & n26324 ) | ( x785 & ~n26338 ) | ( n26324 & ~n26338 ) ;
  assign n26340 = ~n26338 & n26339 ;
  assign n26341 = x618 & ~n26340 ;
  assign n26342 = x618 | n26285 ;
  assign n26343 = ( x1154 & n26341 ) | ( x1154 & n26342 ) | ( n26341 & n26342 ) ;
  assign n26344 = ~n26341 & n26343 ;
  assign n26345 = ( x627 & n26257 ) | ( x627 & ~n26344 ) | ( n26257 & ~n26344 ) ;
  assign n26346 = ~n26257 & n26345 ;
  assign n26347 = x627 | n26255 ;
  assign n26348 = x618 & ~n26285 ;
  assign n26349 = x1154 | n26348 ;
  assign n26350 = ( n26340 & n26341 ) | ( n26340 & ~n26349 ) | ( n26341 & ~n26349 ) ;
  assign n26351 = ( ~n26346 & n26347 ) | ( ~n26346 & n26350 ) | ( n26347 & n26350 ) ;
  assign n26352 = ~n26346 & n26351 ;
  assign n26353 = n26340 ^ x781 ^ 1'b0 ;
  assign n26354 = ( n26340 & n26352 ) | ( n26340 & n26353 ) | ( n26352 & n26353 ) ;
  assign n26355 = ~x789 & n26354 ;
  assign n26356 = x619 & ~n26286 ;
  assign n26357 = x1159 | n26356 ;
  assign n26358 = x619 & ~n26354 ;
  assign n26359 = ( n26354 & ~n26357 ) | ( n26354 & n26358 ) | ( ~n26357 & n26358 ) ;
  assign n26360 = ( x648 & n26262 ) | ( x648 & ~n26359 ) | ( n26262 & ~n26359 ) ;
  assign n26361 = n26359 | n26360 ;
  assign n26362 = x619 | n26286 ;
  assign n26363 = x1159 & ~n26358 ;
  assign n26364 = n26362 & n26363 ;
  assign n26365 = ( x648 & n26264 ) | ( x648 & ~n26364 ) | ( n26264 & ~n26364 ) ;
  assign n26366 = ~n26264 & n26365 ;
  assign n26367 = x789 & ~n26366 ;
  assign n26368 = n26361 & n26367 ;
  assign n26369 = ( n16519 & ~n26355 ) | ( n16519 & n26368 ) | ( ~n26355 & n26368 ) ;
  assign n26370 = n26355 | n26369 ;
  assign n26371 = n26370 ^ n26311 ^ 1'b0 ;
  assign n26372 = ( n26311 & n26370 ) | ( n26311 & n26371 ) | ( n26370 & n26371 ) ;
  assign n26373 = ( n18482 & ~n26311 ) | ( n18482 & n26372 ) | ( ~n26311 & n26372 ) ;
  assign n26374 = n19208 | n26288 ;
  assign n26375 = n16556 & ~n26269 ;
  assign n26376 = x629 & ~n26375 ;
  assign n26377 = n26374 & n26376 ;
  assign n26378 = n16557 & ~n26269 ;
  assign n26379 = n19212 & ~n26288 ;
  assign n26380 = n26378 | n26379 ;
  assign n26381 = ( x629 & ~n26377 ) | ( x629 & n26380 ) | ( ~n26377 & n26380 ) ;
  assign n26382 = ~n26377 & n26381 ;
  assign n26383 = ( x792 & ~n19206 ) | ( x792 & n26382 ) | ( ~n19206 & n26382 ) ;
  assign n26384 = ( n18484 & n19206 ) | ( n18484 & n26383 ) | ( n19206 & n26383 ) ;
  assign n26385 = ( n26298 & n26373 ) | ( n26298 & ~n26384 ) | ( n26373 & ~n26384 ) ;
  assign n26386 = n26385 ^ n26373 ^ 1'b0 ;
  assign n26387 = ( n26298 & n26385 ) | ( n26298 & ~n26386 ) | ( n26385 & ~n26386 ) ;
  assign n26388 = x790 | n26387 ;
  assign n26389 = x644 & ~n26387 ;
  assign n26390 = ( x787 & n26291 ) | ( x787 & ~n26294 ) | ( n26291 & ~n26294 ) ;
  assign n26391 = ~n26291 & n26390 ;
  assign n26392 = ( x787 & n26289 ) | ( x787 & ~n26391 ) | ( n26289 & ~n26391 ) ;
  assign n26393 = ~n26391 & n26392 ;
  assign n26394 = x644 | n26393 ;
  assign n26395 = ( x715 & n26389 ) | ( x715 & n26394 ) | ( n26389 & n26394 ) ;
  assign n26396 = ~n26389 & n26395 ;
  assign n26397 = x644 | n26244 ;
  assign n26398 = n26244 ^ n16376 ^ 1'b0 ;
  assign n26399 = ( n26244 & n26271 ) | ( n26244 & ~n26398 ) | ( n26271 & ~n26398 ) ;
  assign n26400 = x644 & ~n26399 ;
  assign n26401 = ( x715 & n26397 ) | ( x715 & ~n26400 ) | ( n26397 & ~n26400 ) ;
  assign n26402 = ~x715 & n26401 ;
  assign n26403 = ( x1160 & n26396 ) | ( x1160 & ~n26402 ) | ( n26396 & ~n26402 ) ;
  assign n26404 = ~n26396 & n26403 ;
  assign n26405 = x644 & ~n26244 ;
  assign n26406 = x715 & ~n26405 ;
  assign n26407 = ( n26399 & n26400 ) | ( n26399 & n26406 ) | ( n26400 & n26406 ) ;
  assign n26408 = x644 & ~n26393 ;
  assign n26409 = x715 | n26408 ;
  assign n26410 = ( n26387 & n26389 ) | ( n26387 & ~n26409 ) | ( n26389 & ~n26409 ) ;
  assign n26411 = ( x1160 & ~n26407 ) | ( x1160 & n26410 ) | ( ~n26407 & n26410 ) ;
  assign n26412 = n26407 | n26411 ;
  assign n26413 = x790 & ~n26412 ;
  assign n26414 = ( x790 & n26404 ) | ( x790 & n26413 ) | ( n26404 & n26413 ) ;
  assign n26415 = x832 & ~n26414 ;
  assign n26416 = n26388 & n26415 ;
  assign n26417 = ~x184 & n7318 ;
  assign n26418 = x832 | n26417 ;
  assign n26419 = ~n26416 & n26418 ;
  assign n26420 = ( n26243 & n26416 ) | ( n26243 & ~n26419 ) | ( n26416 & ~n26419 ) ;
  assign n26421 = x185 | n15656 ;
  assign n26422 = x701 | n2069 ;
  assign n26423 = ~n26421 & n26422 ;
  assign n26424 = ( x38 & x185 ) | ( x38 & n16700 ) | ( x185 & n16700 ) ;
  assign n26425 = ~n2069 & n26424 ;
  assign n26426 = ( x185 & n16697 ) | ( x185 & ~n26425 ) | ( n16697 & ~n26425 ) ;
  assign n26427 = ~n26425 & n26426 ;
  assign n26428 = x185 | n15644 ;
  assign n26429 = n16185 & n26428 ;
  assign n26430 = x701 | n26429 ;
  assign n26431 = ( ~n26423 & n26427 ) | ( ~n26423 & n26430 ) | ( n26427 & n26430 ) ;
  assign n26432 = ~n26423 & n26431 ;
  assign n26433 = x625 & ~n26432 ;
  assign n26434 = x625 | n26421 ;
  assign n26435 = ( x1153 & n26433 ) | ( x1153 & n26434 ) | ( n26433 & n26434 ) ;
  assign n26436 = ~n26433 & n26435 ;
  assign n26437 = x625 & ~n26421 ;
  assign n26438 = x1153 | n26437 ;
  assign n26439 = ( x625 & n26432 ) | ( x625 & ~n26438 ) | ( n26432 & ~n26438 ) ;
  assign n26440 = ~n26438 & n26439 ;
  assign n26441 = n26436 | n26440 ;
  assign n26442 = n26432 ^ x778 ^ 1'b0 ;
  assign n26443 = ( n26432 & n26441 ) | ( n26432 & n26442 ) | ( n26441 & n26442 ) ;
  assign n26444 = n26421 ^ n16234 ^ 1'b0 ;
  assign n26445 = ( n26421 & n26443 ) | ( n26421 & ~n26444 ) | ( n26443 & ~n26444 ) ;
  assign n26446 = n26421 ^ n16254 ^ 1'b0 ;
  assign n26447 = ( n26421 & n26445 ) | ( n26421 & ~n26446 ) | ( n26445 & ~n26446 ) ;
  assign n26448 = n26421 ^ n16279 ^ 1'b0 ;
  assign n26449 = ( n26421 & n26447 ) | ( n26421 & ~n26448 ) | ( n26447 & ~n26448 ) ;
  assign n26450 = n26421 ^ n16318 ^ 1'b0 ;
  assign n26451 = ( n26421 & n26449 ) | ( n26421 & ~n26450 ) | ( n26449 & ~n26450 ) ;
  assign n26452 = x628 & ~n26451 ;
  assign n26453 = x628 | n26421 ;
  assign n26454 = ( x1156 & n26452 ) | ( x1156 & n26453 ) | ( n26452 & n26453 ) ;
  assign n26455 = ~n26452 & n26454 ;
  assign n26456 = x628 & ~n26421 ;
  assign n26457 = x1156 | n26456 ;
  assign n26458 = ( n26451 & n26452 ) | ( n26451 & ~n26457 ) | ( n26452 & ~n26457 ) ;
  assign n26459 = n26455 | n26458 ;
  assign n26460 = n26451 ^ x792 ^ 1'b0 ;
  assign n26461 = ( n26451 & n26459 ) | ( n26451 & n26460 ) | ( n26459 & n26460 ) ;
  assign n26462 = n26421 ^ x647 ^ 1'b0 ;
  assign n26463 = ( n26421 & n26461 ) | ( n26421 & ~n26462 ) | ( n26461 & ~n26462 ) ;
  assign n26464 = ( n26421 & n26461 ) | ( n26421 & n26462 ) | ( n26461 & n26462 ) ;
  assign n26465 = n26463 ^ x1157 ^ 1'b0 ;
  assign n26466 = ( n26463 & n26464 ) | ( n26463 & n26465 ) | ( n26464 & n26465 ) ;
  assign n26467 = n26461 ^ x787 ^ 1'b0 ;
  assign n26468 = ( n26461 & n26466 ) | ( n26461 & n26467 ) | ( n26466 & n26467 ) ;
  assign n26469 = x644 & ~n26468 ;
  assign n26470 = x715 | n26469 ;
  assign n26471 = x644 & ~n26421 ;
  assign n26472 = x715 & ~n26471 ;
  assign n26473 = n26472 ^ x1160 ^ 1'b0 ;
  assign n26474 = x38 & n26428 ;
  assign n26475 = x751 & n15332 ;
  assign n26476 = x185 & ~n15638 ;
  assign n26477 = ( ~x39 & n26475 ) | ( ~x39 & n26476 ) | ( n26475 & n26476 ) ;
  assign n26478 = ~x39 & n26477 ;
  assign n26479 = n26478 ^ x185 ^ 1'b0 ;
  assign n26480 = ( ~x185 & x751 ) | ( ~x185 & n26479 ) | ( x751 & n26479 ) ;
  assign n26481 = ( x185 & n26478 ) | ( x185 & n26480 ) | ( n26478 & n26480 ) ;
  assign n26482 = n26480 ^ n26478 ^ x185 ;
  assign n26483 = ( n15587 & n26481 ) | ( n15587 & ~n26482 ) | ( n26481 & ~n26482 ) ;
  assign n26484 = x185 & ~n15631 ;
  assign n26485 = x751 & n15486 ;
  assign n26486 = ( x39 & n26484 ) | ( x39 & n26485 ) | ( n26484 & n26485 ) ;
  assign n26487 = n26485 ^ n26484 ^ 1'b0 ;
  assign n26488 = ( x39 & n26486 ) | ( x39 & n26487 ) | ( n26486 & n26487 ) ;
  assign n26489 = ( ~x38 & n26483 ) | ( ~x38 & n26488 ) | ( n26483 & n26488 ) ;
  assign n26490 = ~x38 & n26489 ;
  assign n26491 = ~x751 & n15646 ;
  assign n26492 = ~n26490 & n26491 ;
  assign n26493 = ( n26474 & n26490 ) | ( n26474 & ~n26492 ) | ( n26490 & ~n26492 ) ;
  assign n26494 = ~n2069 & n26493 ;
  assign n26495 = x185 & n2069 ;
  assign n26496 = n26494 | n26495 ;
  assign n26497 = n26421 ^ n15659 ^ 1'b0 ;
  assign n26498 = ( n26421 & n26496 ) | ( n26421 & ~n26497 ) | ( n26496 & ~n26497 ) ;
  assign n26499 = n15662 & n26421 ;
  assign n26500 = ( ~n15662 & n26494 ) | ( ~n15662 & n26495 ) | ( n26494 & n26495 ) ;
  assign n26501 = n26499 | n26500 ;
  assign n26502 = n26501 ^ n26498 ^ n26421 ;
  assign n26503 = n26502 ^ x1155 ^ 1'b0 ;
  assign n26504 = ( n26501 & n26502 ) | ( n26501 & ~n26503 ) | ( n26502 & ~n26503 ) ;
  assign n26505 = n26498 ^ x785 ^ 1'b0 ;
  assign n26506 = ( n26498 & n26504 ) | ( n26498 & n26505 ) | ( n26504 & n26505 ) ;
  assign n26507 = x618 & ~n26506 ;
  assign n26508 = x618 | n26421 ;
  assign n26509 = ( x1154 & n26507 ) | ( x1154 & n26508 ) | ( n26507 & n26508 ) ;
  assign n26510 = ~n26507 & n26509 ;
  assign n26511 = x618 & ~n26421 ;
  assign n26512 = x1154 | n26511 ;
  assign n26513 = ( n26506 & n26507 ) | ( n26506 & ~n26512 ) | ( n26507 & ~n26512 ) ;
  assign n26514 = n26510 | n26513 ;
  assign n26515 = n26506 ^ x781 ^ 1'b0 ;
  assign n26516 = ( n26506 & n26514 ) | ( n26506 & n26515 ) | ( n26514 & n26515 ) ;
  assign n26517 = x619 & ~n26516 ;
  assign n26518 = x619 | n26421 ;
  assign n26519 = ( x1159 & n26517 ) | ( x1159 & n26518 ) | ( n26517 & n26518 ) ;
  assign n26520 = ~n26517 & n26519 ;
  assign n26521 = x619 & ~n26421 ;
  assign n26522 = x1159 | n26521 ;
  assign n26523 = ( n26516 & n26517 ) | ( n26516 & ~n26522 ) | ( n26517 & ~n26522 ) ;
  assign n26524 = n26520 | n26523 ;
  assign n26525 = n26516 ^ x789 ^ 1'b0 ;
  assign n26526 = ( n26516 & n26524 ) | ( n26516 & n26525 ) | ( n26524 & n26525 ) ;
  assign n26527 = n26421 ^ n16518 ^ 1'b0 ;
  assign n26528 = ( n26421 & n26526 ) | ( n26421 & ~n26527 ) | ( n26526 & ~n26527 ) ;
  assign n26529 = n26421 ^ n16339 ^ 1'b0 ;
  assign n26530 = ( n26421 & n26528 ) | ( n26421 & ~n26529 ) | ( n26528 & ~n26529 ) ;
  assign n26531 = n26421 ^ n16376 ^ 1'b0 ;
  assign n26532 = ( n26421 & n26530 ) | ( n26421 & ~n26531 ) | ( n26530 & ~n26531 ) ;
  assign n26533 = x644 | n26532 ;
  assign n26534 = ( n26472 & ~n26473 ) | ( n26472 & n26533 ) | ( ~n26473 & n26533 ) ;
  assign n26535 = ( x1160 & n26473 ) | ( x1160 & n26534 ) | ( n26473 & n26534 ) ;
  assign n26536 = n26470 & ~n26535 ;
  assign n26537 = x644 & ~n26532 ;
  assign n26538 = ( ~x715 & n26421 ) | ( ~x715 & n26471 ) | ( n26421 & n26471 ) ;
  assign n26539 = x1160 & ~n26538 ;
  assign n26540 = ( x1160 & n26537 ) | ( x1160 & n26539 ) | ( n26537 & n26539 ) ;
  assign n26541 = ( x715 & n26468 ) | ( x715 & n26469 ) | ( n26468 & n26469 ) ;
  assign n26542 = n26540 & ~n26541 ;
  assign n26543 = ( x790 & n26536 ) | ( x790 & n26542 ) | ( n26536 & n26542 ) ;
  assign n26544 = n26542 ^ n26536 ^ 1'b0 ;
  assign n26545 = ( x790 & n26543 ) | ( x790 & n26544 ) | ( n26543 & n26544 ) ;
  assign n26546 = n19055 & n26530 ;
  assign n26547 = n16374 & n26463 ;
  assign n26548 = n16373 & n26464 ;
  assign n26549 = n26547 | n26548 ;
  assign n26550 = ( x787 & n26546 ) | ( x787 & n26549 ) | ( n26546 & n26549 ) ;
  assign n26551 = n26549 ^ n26546 ^ 1'b0 ;
  assign n26552 = ( x787 & n26550 ) | ( x787 & n26551 ) | ( n26550 & n26551 ) ;
  assign n26553 = x701 & ~n26493 ;
  assign n26554 = x185 & ~n16054 ;
  assign n26555 = ~x185 & n16048 ;
  assign n26556 = ( x751 & ~n26554 ) | ( x751 & n26555 ) | ( ~n26554 & n26555 ) ;
  assign n26557 = n26554 | n26556 ;
  assign n26558 = ~x185 & n16044 ;
  assign n26559 = x185 & ~n16029 ;
  assign n26560 = ( x751 & n26558 ) | ( x751 & ~n26559 ) | ( n26558 & ~n26559 ) ;
  assign n26561 = ~n26558 & n26560 ;
  assign n26562 = ( x39 & n26557 ) | ( x39 & ~n26561 ) | ( n26557 & ~n26561 ) ;
  assign n26563 = n26562 ^ n26557 ^ 1'b0 ;
  assign n26564 = ( x39 & n26562 ) | ( x39 & ~n26563 ) | ( n26562 & ~n26563 ) ;
  assign n26565 = x185 & n15795 ;
  assign n26566 = x751 & ~n26565 ;
  assign n26567 = x185 | n15876 ;
  assign n26568 = n26566 & n26567 ;
  assign n26569 = x185 & n15943 ;
  assign n26570 = x185 | n16003 ;
  assign n26571 = ( x751 & ~n26569 ) | ( x751 & n26570 ) | ( ~n26569 & n26570 ) ;
  assign n26572 = ~x751 & n26571 ;
  assign n26573 = ( x39 & n26568 ) | ( x39 & ~n26572 ) | ( n26568 & ~n26572 ) ;
  assign n26574 = ~n26568 & n26573 ;
  assign n26575 = ( x38 & n26564 ) | ( x38 & ~n26574 ) | ( n26564 & ~n26574 ) ;
  assign n26576 = ~x38 & n26575 ;
  assign n26577 = ~x751 & n15591 ;
  assign n26578 = n17156 | n26577 ;
  assign n26579 = x185 & ~n5017 ;
  assign n26580 = n26578 & n26579 ;
  assign n26581 = x38 & ~n26580 ;
  assign n26582 = n26581 ^ x701 ^ 1'b0 ;
  assign n26583 = x751 | n15968 ;
  assign n26584 = n17889 & n26583 ;
  assign n26585 = x185 | n26584 ;
  assign n26586 = ( n26581 & ~n26582 ) | ( n26581 & n26585 ) | ( ~n26582 & n26585 ) ;
  assign n26587 = ( x701 & n26582 ) | ( x701 & n26586 ) | ( n26582 & n26586 ) ;
  assign n26588 = ( ~n2069 & n26576 ) | ( ~n2069 & n26587 ) | ( n26576 & n26587 ) ;
  assign n26589 = ~n2069 & n26588 ;
  assign n26590 = n26589 ^ n26553 ^ 1'b0 ;
  assign n26591 = ( n26553 & n26589 ) | ( n26553 & n26590 ) | ( n26589 & n26590 ) ;
  assign n26592 = ( n26495 & ~n26553 ) | ( n26495 & n26591 ) | ( ~n26553 & n26591 ) ;
  assign n26593 = x625 & ~n26592 ;
  assign n26594 = x625 | n26496 ;
  assign n26595 = ( x1153 & n26593 ) | ( x1153 & n26594 ) | ( n26593 & n26594 ) ;
  assign n26596 = ~n26593 & n26595 ;
  assign n26597 = ( x608 & n26440 ) | ( x608 & ~n26596 ) | ( n26440 & ~n26596 ) ;
  assign n26598 = ~n26440 & n26597 ;
  assign n26599 = x608 | n26436 ;
  assign n26600 = x625 & ~n26496 ;
  assign n26601 = x1153 | n26600 ;
  assign n26602 = ( n26592 & n26593 ) | ( n26592 & ~n26601 ) | ( n26593 & ~n26601 ) ;
  assign n26603 = ( ~n26598 & n26599 ) | ( ~n26598 & n26602 ) | ( n26599 & n26602 ) ;
  assign n26604 = ~n26598 & n26603 ;
  assign n26605 = n26592 ^ x778 ^ 1'b0 ;
  assign n26606 = ( n26592 & n26604 ) | ( n26592 & n26605 ) | ( n26604 & n26605 ) ;
  assign n26607 = x609 & ~n26606 ;
  assign n26608 = x609 | n26443 ;
  assign n26609 = ( x1155 & n26607 ) | ( x1155 & n26608 ) | ( n26607 & n26608 ) ;
  assign n26610 = ~n26607 & n26609 ;
  assign n26611 = ~x1155 & n26501 ;
  assign n26612 = ( x660 & n26610 ) | ( x660 & ~n26611 ) | ( n26610 & ~n26611 ) ;
  assign n26613 = ~n26610 & n26612 ;
  assign n26614 = x1155 & n26502 ;
  assign n26615 = x660 | n26614 ;
  assign n26616 = x609 & ~n26443 ;
  assign n26617 = x1155 | n26616 ;
  assign n26618 = ( n26606 & n26607 ) | ( n26606 & ~n26617 ) | ( n26607 & ~n26617 ) ;
  assign n26619 = ( ~n26613 & n26615 ) | ( ~n26613 & n26618 ) | ( n26615 & n26618 ) ;
  assign n26620 = ~n26613 & n26619 ;
  assign n26621 = n26606 ^ x785 ^ 1'b0 ;
  assign n26622 = ( n26606 & n26620 ) | ( n26606 & n26621 ) | ( n26620 & n26621 ) ;
  assign n26623 = x618 & ~n26622 ;
  assign n26624 = x618 | n26445 ;
  assign n26625 = ( x1154 & n26623 ) | ( x1154 & n26624 ) | ( n26623 & n26624 ) ;
  assign n26626 = ~n26623 & n26625 ;
  assign n26627 = ( x627 & n26513 ) | ( x627 & ~n26626 ) | ( n26513 & ~n26626 ) ;
  assign n26628 = ~n26513 & n26627 ;
  assign n26629 = x627 | n26510 ;
  assign n26630 = x618 & ~n26445 ;
  assign n26631 = x1154 | n26630 ;
  assign n26632 = ( n26622 & n26623 ) | ( n26622 & ~n26631 ) | ( n26623 & ~n26631 ) ;
  assign n26633 = ( ~n26628 & n26629 ) | ( ~n26628 & n26632 ) | ( n26629 & n26632 ) ;
  assign n26634 = ~n26628 & n26633 ;
  assign n26635 = n26622 ^ x781 ^ 1'b0 ;
  assign n26636 = ( n26622 & n26634 ) | ( n26622 & n26635 ) | ( n26634 & n26635 ) ;
  assign n26637 = x619 | n26636 ;
  assign n26638 = x619 & ~n26447 ;
  assign n26639 = ( x1159 & n26637 ) | ( x1159 & ~n26638 ) | ( n26637 & ~n26638 ) ;
  assign n26640 = ~x1159 & n26639 ;
  assign n26641 = ( x648 & n26520 ) | ( x648 & ~n26640 ) | ( n26520 & ~n26640 ) ;
  assign n26642 = n26640 | n26641 ;
  assign n26643 = x619 & ~n26636 ;
  assign n26644 = x619 | n26447 ;
  assign n26645 = ( x1159 & n26643 ) | ( x1159 & n26644 ) | ( n26643 & n26644 ) ;
  assign n26646 = ~n26643 & n26645 ;
  assign n26647 = ( x648 & n26523 ) | ( x648 & ~n26646 ) | ( n26523 & ~n26646 ) ;
  assign n26648 = ~n26523 & n26647 ;
  assign n26649 = x789 & ~n26648 ;
  assign n26650 = n26642 & n26649 ;
  assign n26651 = ~x789 & n26636 ;
  assign n26652 = ( n16519 & ~n26650 ) | ( n16519 & n26651 ) | ( ~n26650 & n26651 ) ;
  assign n26653 = n26650 | n26652 ;
  assign n26654 = n26455 ^ x629 ^ 1'b0 ;
  assign n26655 = ( n26455 & n26458 ) | ( n26455 & n26654 ) | ( n26458 & n26654 ) ;
  assign n26656 = n19046 & n26528 ;
  assign n26657 = ( x792 & n26655 ) | ( x792 & n26656 ) | ( n26655 & n26656 ) ;
  assign n26658 = n26656 ^ n26655 ^ 1'b0 ;
  assign n26659 = ( x792 & n26657 ) | ( x792 & n26658 ) | ( n26657 & n26658 ) ;
  assign n26660 = n16459 & ~n26449 ;
  assign n26661 = ~x626 & n26421 ;
  assign n26662 = x626 & n26526 ;
  assign n26663 = ( n22317 & n26661 ) | ( n22317 & ~n26662 ) | ( n26661 & ~n26662 ) ;
  assign n26664 = ~n26661 & n26663 ;
  assign n26665 = ~x626 & n26526 ;
  assign n26666 = x626 & n26421 ;
  assign n26667 = ( n22322 & n26665 ) | ( n22322 & ~n26666 ) | ( n26665 & ~n26666 ) ;
  assign n26668 = ~n26665 & n26667 ;
  assign n26669 = ( ~n26660 & n26664 ) | ( ~n26660 & n26668 ) | ( n26664 & n26668 ) ;
  assign n26670 = n26660 | n26669 ;
  assign n26671 = ( x788 & ~n22314 ) | ( x788 & n26670 ) | ( ~n22314 & n26670 ) ;
  assign n26672 = ( n18482 & n22314 ) | ( n18482 & n26671 ) | ( n22314 & n26671 ) ;
  assign n26673 = ~n26659 & n26672 ;
  assign n26674 = ( n26653 & n26659 ) | ( n26653 & ~n26673 ) | ( n26659 & ~n26673 ) ;
  assign n26675 = ( ~n18484 & n26552 ) | ( ~n18484 & n26674 ) | ( n26552 & n26674 ) ;
  assign n26676 = n26552 ^ n18484 ^ 1'b0 ;
  assign n26677 = ( n26552 & n26675 ) | ( n26552 & ~n26676 ) | ( n26675 & ~n26676 ) ;
  assign n26678 = x644 | n26535 ;
  assign n26679 = x644 & n26540 ;
  assign n26680 = x790 & ~n26679 ;
  assign n26681 = n26678 & n26680 ;
  assign n26682 = ( ~n26545 & n26677 ) | ( ~n26545 & n26681 ) | ( n26677 & n26681 ) ;
  assign n26683 = ~n26545 & n26682 ;
  assign n26684 = ( x57 & n5193 ) | ( x57 & ~n26683 ) | ( n5193 & ~n26683 ) ;
  assign n26685 = n26683 | n26684 ;
  assign n26686 = x185 | n1611 ;
  assign n26687 = ~n26577 & n26686 ;
  assign n26688 = n16397 | n26687 ;
  assign n26689 = ~n15662 & n26577 ;
  assign n26690 = ~x1155 & n26686 ;
  assign n26691 = ~n26689 & n26690 ;
  assign n26692 = ( x1155 & n26688 ) | ( x1155 & n26689 ) | ( n26688 & n26689 ) ;
  assign n26693 = n26691 | n26692 ;
  assign n26694 = n26688 ^ x785 ^ 1'b0 ;
  assign n26695 = ( n26688 & n26693 ) | ( n26688 & n26694 ) | ( n26693 & n26694 ) ;
  assign n26696 = n16411 | n26695 ;
  assign n26697 = x1154 & n26696 ;
  assign n26698 = n16414 | n26695 ;
  assign n26699 = ~x1154 & n26698 ;
  assign n26700 = n26697 | n26699 ;
  assign n26701 = n26695 ^ x781 ^ 1'b0 ;
  assign n26702 = ( n26695 & n26700 ) | ( n26695 & n26701 ) | ( n26700 & n26701 ) ;
  assign n26703 = n21437 | n26702 ;
  assign n26704 = x1159 & n26703 ;
  assign n26705 = n21440 | n26702 ;
  assign n26706 = ~x1159 & n26705 ;
  assign n26707 = n26704 | n26706 ;
  assign n26708 = n26702 ^ x789 ^ 1'b0 ;
  assign n26709 = ( n26702 & n26707 ) | ( n26702 & n26708 ) | ( n26707 & n26708 ) ;
  assign n26710 = n26686 ^ n16518 ^ 1'b0 ;
  assign n26711 = ( n26686 & n26709 ) | ( n26686 & ~n26710 ) | ( n26709 & ~n26710 ) ;
  assign n26712 = n26686 ^ n16339 ^ 1'b0 ;
  assign n26713 = ( n26686 & n26711 ) | ( n26686 & ~n26712 ) | ( n26711 & ~n26712 ) ;
  assign n26714 = n19055 & n26713 ;
  assign n26715 = x647 & ~n26686 ;
  assign n26716 = x1157 | n26715 ;
  assign n26717 = ~x701 & n15778 ;
  assign n26718 = ~x625 & n26717 ;
  assign n26719 = ~x1153 & n26686 ;
  assign n26720 = ~n26718 & n26719 ;
  assign n26721 = x778 & ~n26720 ;
  assign n26722 = n26686 & ~n26717 ;
  assign n26723 = ( x1153 & n26718 ) | ( x1153 & n26722 ) | ( n26718 & n26722 ) ;
  assign n26724 = n26721 & ~n26723 ;
  assign n26725 = ( x778 & n26722 ) | ( x778 & ~n26724 ) | ( n26722 & ~n26724 ) ;
  assign n26726 = ~n26724 & n26725 ;
  assign n26727 = n16447 | n26726 ;
  assign n26728 = n16449 | n26727 ;
  assign n26729 = n16451 | n26728 ;
  assign n26730 = n16530 | n26729 ;
  assign n26731 = n16560 | n26730 ;
  assign n26732 = ( x647 & ~n26716 ) | ( x647 & n26731 ) | ( ~n26716 & n26731 ) ;
  assign n26733 = ~n26716 & n26732 ;
  assign n26734 = n26686 ^ x647 ^ 1'b0 ;
  assign n26735 = ( n26686 & n26731 ) | ( n26686 & n26734 ) | ( n26731 & n26734 ) ;
  assign n26736 = x1157 & n26735 ;
  assign n26737 = ( n16375 & n26733 ) | ( n16375 & n26736 ) | ( n26733 & n26736 ) ;
  assign n26738 = ( x787 & n26714 ) | ( x787 & n26737 ) | ( n26714 & n26737 ) ;
  assign n26739 = n26737 ^ n26714 ^ 1'b0 ;
  assign n26740 = ( x787 & n26738 ) | ( x787 & n26739 ) | ( n26738 & n26739 ) ;
  assign n26741 = ~x626 & n26686 ;
  assign n26742 = x626 & n26709 ;
  assign n26743 = ( n22317 & n26741 ) | ( n22317 & ~n26742 ) | ( n26741 & ~n26742 ) ;
  assign n26744 = ~n26741 & n26743 ;
  assign n26745 = ~x626 & n26709 ;
  assign n26746 = x626 & n26686 ;
  assign n26747 = ( n22322 & n26745 ) | ( n22322 & ~n26746 ) | ( n26745 & ~n26746 ) ;
  assign n26748 = ~n26745 & n26747 ;
  assign n26749 = n26729 & ~n26748 ;
  assign n26750 = ( n16459 & n26748 ) | ( n16459 & ~n26749 ) | ( n26748 & ~n26749 ) ;
  assign n26751 = ( x788 & n26744 ) | ( x788 & n26750 ) | ( n26744 & n26750 ) ;
  assign n26752 = n26750 ^ n26744 ^ 1'b0 ;
  assign n26753 = ( x788 & n26751 ) | ( x788 & n26752 ) | ( n26751 & n26752 ) ;
  assign n26754 = n15524 | n26722 ;
  assign n26755 = n26687 & n26754 ;
  assign n26756 = x625 & ~n26754 ;
  assign n26757 = ( n26719 & n26755 ) | ( n26719 & n26756 ) | ( n26755 & n26756 ) ;
  assign n26758 = ( x608 & n26723 ) | ( x608 & ~n26757 ) | ( n26723 & ~n26757 ) ;
  assign n26759 = n26757 | n26758 ;
  assign n26760 = x1153 & n26687 ;
  assign n26761 = ~n26756 & n26760 ;
  assign n26762 = x608 & ~n26720 ;
  assign n26763 = n26759 & ~n26762 ;
  assign n26764 = ( n26759 & n26761 ) | ( n26759 & n26763 ) | ( n26761 & n26763 ) ;
  assign n26765 = n26755 ^ x778 ^ 1'b0 ;
  assign n26766 = ( n26755 & n26764 ) | ( n26755 & n26765 ) | ( n26764 & n26765 ) ;
  assign n26767 = x609 & ~n26766 ;
  assign n26773 = x609 | n26726 ;
  assign n26774 = ( x1155 & n26767 ) | ( x1155 & n26773 ) | ( n26767 & n26773 ) ;
  assign n26775 = ~n26767 & n26774 ;
  assign n26776 = ( x660 & n26691 ) | ( x660 & ~n26775 ) | ( n26691 & ~n26775 ) ;
  assign n26777 = ~n26691 & n26776 ;
  assign n26768 = x609 & ~n26726 ;
  assign n26769 = x1155 | n26768 ;
  assign n26770 = ( n26766 & n26767 ) | ( n26766 & ~n26769 ) | ( n26767 & ~n26769 ) ;
  assign n26771 = ( x660 & n26692 ) | ( x660 & ~n26770 ) | ( n26692 & ~n26770 ) ;
  assign n26772 = n26770 | n26771 ;
  assign n26778 = n26777 ^ n26772 ^ 1'b0 ;
  assign n26779 = ( x785 & ~n26772 ) | ( x785 & n26777 ) | ( ~n26772 & n26777 ) ;
  assign n26780 = ( x785 & ~n26778 ) | ( x785 & n26779 ) | ( ~n26778 & n26779 ) ;
  assign n26781 = ( x785 & n26766 ) | ( x785 & ~n26780 ) | ( n26766 & ~n26780 ) ;
  assign n26782 = ~n26780 & n26781 ;
  assign n26783 = x618 & ~n26782 ;
  assign n26784 = x618 | n26727 ;
  assign n26785 = ( x1154 & n26783 ) | ( x1154 & n26784 ) | ( n26783 & n26784 ) ;
  assign n26786 = ~n26783 & n26785 ;
  assign n26787 = ( x627 & n26699 ) | ( x627 & ~n26786 ) | ( n26699 & ~n26786 ) ;
  assign n26788 = ~n26699 & n26787 ;
  assign n26789 = x627 | n26697 ;
  assign n26790 = x618 & ~n26727 ;
  assign n26791 = x1154 | n26790 ;
  assign n26792 = ( n26782 & n26783 ) | ( n26782 & ~n26791 ) | ( n26783 & ~n26791 ) ;
  assign n26793 = ( ~n26788 & n26789 ) | ( ~n26788 & n26792 ) | ( n26789 & n26792 ) ;
  assign n26794 = ~n26788 & n26793 ;
  assign n26795 = n26782 ^ x781 ^ 1'b0 ;
  assign n26796 = ( n26782 & n26794 ) | ( n26782 & n26795 ) | ( n26794 & n26795 ) ;
  assign n26797 = ~x789 & n26796 ;
  assign n26798 = x619 & ~n26728 ;
  assign n26799 = x1159 | n26798 ;
  assign n26800 = x619 & ~n26796 ;
  assign n26801 = ( n26796 & ~n26799 ) | ( n26796 & n26800 ) | ( ~n26799 & n26800 ) ;
  assign n26802 = ( x648 & n26704 ) | ( x648 & ~n26801 ) | ( n26704 & ~n26801 ) ;
  assign n26803 = n26801 | n26802 ;
  assign n26804 = x619 | n26728 ;
  assign n26805 = x1159 & ~n26800 ;
  assign n26806 = n26804 & n26805 ;
  assign n26807 = ( x648 & n26706 ) | ( x648 & ~n26806 ) | ( n26706 & ~n26806 ) ;
  assign n26808 = ~n26706 & n26807 ;
  assign n26809 = x789 & ~n26808 ;
  assign n26810 = n26803 & n26809 ;
  assign n26811 = ( n16519 & ~n26797 ) | ( n16519 & n26810 ) | ( ~n26797 & n26810 ) ;
  assign n26812 = n26797 | n26811 ;
  assign n26813 = n26812 ^ n26753 ^ 1'b0 ;
  assign n26814 = ( n26753 & n26812 ) | ( n26753 & n26813 ) | ( n26812 & n26813 ) ;
  assign n26815 = ( n18482 & ~n26753 ) | ( n18482 & n26814 ) | ( ~n26753 & n26814 ) ;
  assign n26816 = n19208 | n26730 ;
  assign n26817 = n16556 & ~n26711 ;
  assign n26818 = x629 & ~n26817 ;
  assign n26819 = n26816 & n26818 ;
  assign n26820 = n16557 & ~n26711 ;
  assign n26821 = n19212 & ~n26730 ;
  assign n26822 = n26820 | n26821 ;
  assign n26823 = ( x629 & ~n26819 ) | ( x629 & n26822 ) | ( ~n26819 & n26822 ) ;
  assign n26824 = ~n26819 & n26823 ;
  assign n26825 = ( x792 & ~n19206 ) | ( x792 & n26824 ) | ( ~n19206 & n26824 ) ;
  assign n26826 = ( n18484 & n19206 ) | ( n18484 & n26825 ) | ( n19206 & n26825 ) ;
  assign n26827 = ( n26740 & n26815 ) | ( n26740 & ~n26826 ) | ( n26815 & ~n26826 ) ;
  assign n26828 = n26827 ^ n26815 ^ 1'b0 ;
  assign n26829 = ( n26740 & n26827 ) | ( n26740 & ~n26828 ) | ( n26827 & ~n26828 ) ;
  assign n26830 = x790 | n26829 ;
  assign n26831 = x644 & ~n26829 ;
  assign n26832 = ( x787 & n26733 ) | ( x787 & ~n26736 ) | ( n26733 & ~n26736 ) ;
  assign n26833 = ~n26733 & n26832 ;
  assign n26834 = ( x787 & n26731 ) | ( x787 & ~n26833 ) | ( n26731 & ~n26833 ) ;
  assign n26835 = ~n26833 & n26834 ;
  assign n26836 = x644 | n26835 ;
  assign n26837 = ( x715 & n26831 ) | ( x715 & n26836 ) | ( n26831 & n26836 ) ;
  assign n26838 = ~n26831 & n26837 ;
  assign n26839 = x644 | n26686 ;
  assign n26840 = n26686 ^ n16376 ^ 1'b0 ;
  assign n26841 = ( n26686 & n26713 ) | ( n26686 & ~n26840 ) | ( n26713 & ~n26840 ) ;
  assign n26842 = x644 & ~n26841 ;
  assign n26843 = ( x715 & n26839 ) | ( x715 & ~n26842 ) | ( n26839 & ~n26842 ) ;
  assign n26844 = ~x715 & n26843 ;
  assign n26845 = ( x1160 & n26838 ) | ( x1160 & ~n26844 ) | ( n26838 & ~n26844 ) ;
  assign n26846 = ~n26838 & n26845 ;
  assign n26847 = x644 & ~n26686 ;
  assign n26848 = x715 & ~n26847 ;
  assign n26849 = ( n26841 & n26842 ) | ( n26841 & n26848 ) | ( n26842 & n26848 ) ;
  assign n26850 = x644 & ~n26835 ;
  assign n26851 = x715 | n26850 ;
  assign n26852 = ( n26829 & n26831 ) | ( n26829 & ~n26851 ) | ( n26831 & ~n26851 ) ;
  assign n26853 = ( x1160 & ~n26849 ) | ( x1160 & n26852 ) | ( ~n26849 & n26852 ) ;
  assign n26854 = n26849 | n26853 ;
  assign n26855 = x790 & ~n26854 ;
  assign n26856 = ( x790 & n26846 ) | ( x790 & n26855 ) | ( n26846 & n26855 ) ;
  assign n26857 = x832 & ~n26856 ;
  assign n26858 = n26830 & n26857 ;
  assign n26859 = ~x185 & n7318 ;
  assign n26860 = x832 | n26859 ;
  assign n26861 = ~n26858 & n26860 ;
  assign n26862 = ( n26685 & n26858 ) | ( n26685 & ~n26861 ) | ( n26858 & ~n26861 ) ;
  assign n26864 = x186 | x752 ;
  assign n26865 = n17843 & ~n26864 ;
  assign n26866 = x186 & ~n17846 ;
  assign n26867 = ( ~n17839 & n26865 ) | ( ~n17839 & n26866 ) | ( n26865 & n26866 ) ;
  assign n26868 = ~n17839 & n26867 ;
  assign n26869 = x186 | n15655 ;
  assign n26870 = n26868 ^ x752 ^ 1'b0 ;
  assign n26871 = ( ~x752 & n26869 ) | ( ~x752 & n26870 ) | ( n26869 & n26870 ) ;
  assign n26872 = ( x752 & n26868 ) | ( x752 & n26871 ) | ( n26868 & n26871 ) ;
  assign n26900 = x703 | n26872 ;
  assign n26901 = x752 & ~n17882 ;
  assign n26902 = x186 & n17886 ;
  assign n26903 = n26901 & ~n26902 ;
  assign n26904 = x186 | n17893 ;
  assign n26905 = n26903 & n26904 ;
  assign n26906 = x186 | n17902 ;
  assign n26907 = x186 & n17910 ;
  assign n26908 = ( x752 & n26906 ) | ( x752 & ~n26907 ) | ( n26906 & ~n26907 ) ;
  assign n26909 = ~x752 & n26908 ;
  assign n26910 = ( x703 & n26905 ) | ( x703 & ~n26909 ) | ( n26905 & ~n26909 ) ;
  assign n26911 = ~n26905 & n26910 ;
  assign n26912 = ( n2069 & n26900 ) | ( n2069 & ~n26911 ) | ( n26900 & ~n26911 ) ;
  assign n26913 = ~n2069 & n26912 ;
  assign n26914 = n26913 ^ x186 ^ 1'b0 ;
  assign n26915 = ( ~x186 & n2069 ) | ( ~x186 & n26914 ) | ( n2069 & n26914 ) ;
  assign n26916 = ( x186 & n26913 ) | ( x186 & n26915 ) | ( n26913 & n26915 ) ;
  assign n26917 = x625 & ~n26916 ;
  assign n26863 = x186 & n2069 ;
  assign n26873 = ~n2069 & n26872 ;
  assign n26874 = n26863 | n26873 ;
  assign n26918 = x625 | n26874 ;
  assign n26919 = ( x1153 & n26917 ) | ( x1153 & n26918 ) | ( n26917 & n26918 ) ;
  assign n26920 = ~n26917 & n26919 ;
  assign n26875 = x186 | n15656 ;
  assign n26921 = x625 & ~n26875 ;
  assign n26922 = x1153 | n26921 ;
  assign n26923 = ( x38 & x186 ) | ( x38 & n16700 ) | ( x186 & n16700 ) ;
  assign n26924 = ( x186 & n16697 ) | ( x186 & ~n26923 ) | ( n16697 & ~n26923 ) ;
  assign n26925 = ~n26923 & n26924 ;
  assign n26926 = x186 | n15644 ;
  assign n26927 = n16185 & n26926 ;
  assign n26928 = ( x703 & n26925 ) | ( x703 & ~n26927 ) | ( n26925 & ~n26927 ) ;
  assign n26929 = ~n26925 & n26928 ;
  assign n26930 = x703 | n26869 ;
  assign n26931 = ~n2069 & n26930 ;
  assign n26932 = n26931 ^ n26929 ^ 1'b0 ;
  assign n26933 = ( n26929 & n26931 ) | ( n26929 & n26932 ) | ( n26931 & n26932 ) ;
  assign n26934 = ( n26863 & ~n26929 ) | ( n26863 & n26933 ) | ( ~n26929 & n26933 ) ;
  assign n26935 = ( x625 & ~n26922 ) | ( x625 & n26934 ) | ( ~n26922 & n26934 ) ;
  assign n26936 = ~n26922 & n26935 ;
  assign n26937 = ( x608 & n26920 ) | ( x608 & ~n26936 ) | ( n26920 & ~n26936 ) ;
  assign n26938 = ~n26920 & n26937 ;
  assign n26939 = x625 & ~n26934 ;
  assign n26940 = x625 | n26875 ;
  assign n26941 = ( x1153 & n26939 ) | ( x1153 & n26940 ) | ( n26939 & n26940 ) ;
  assign n26942 = ~n26939 & n26941 ;
  assign n26943 = x608 | n26942 ;
  assign n26944 = x625 & ~n26874 ;
  assign n26945 = x1153 | n26944 ;
  assign n26946 = ( n26916 & n26917 ) | ( n26916 & ~n26945 ) | ( n26917 & ~n26945 ) ;
  assign n26947 = ( ~n26938 & n26943 ) | ( ~n26938 & n26946 ) | ( n26943 & n26946 ) ;
  assign n26948 = ~n26938 & n26947 ;
  assign n26949 = n26916 ^ x778 ^ 1'b0 ;
  assign n26950 = ( n26916 & n26948 ) | ( n26916 & n26949 ) | ( n26948 & n26949 ) ;
  assign n26951 = x609 & ~n26950 ;
  assign n26952 = n26936 | n26942 ;
  assign n26953 = n26934 ^ x778 ^ 1'b0 ;
  assign n26954 = ( n26934 & n26952 ) | ( n26934 & n26953 ) | ( n26952 & n26953 ) ;
  assign n26955 = x609 | n26954 ;
  assign n26956 = ( x1155 & n26951 ) | ( x1155 & n26955 ) | ( n26951 & n26955 ) ;
  assign n26957 = ~n26951 & n26956 ;
  assign n26878 = ~n15668 & n26875 ;
  assign n26879 = ( n15668 & n26863 ) | ( n15668 & n26873 ) | ( n26863 & n26873 ) ;
  assign n26880 = n26878 | n26879 ;
  assign n26876 = n26874 ^ n15659 ^ 1'b0 ;
  assign n26877 = ( n26874 & n26875 ) | ( n26874 & n26876 ) | ( n26875 & n26876 ) ;
  assign n26882 = n26880 ^ n26877 ^ n26875 ;
  assign n26958 = ~x1155 & n26882 ;
  assign n26959 = ( x660 & n26957 ) | ( x660 & ~n26958 ) | ( n26957 & ~n26958 ) ;
  assign n26960 = ~n26957 & n26959 ;
  assign n26961 = x1155 & n26880 ;
  assign n26962 = x660 | n26961 ;
  assign n26963 = x609 & ~n26954 ;
  assign n26964 = x1155 | n26963 ;
  assign n26965 = ( n26950 & n26951 ) | ( n26950 & ~n26964 ) | ( n26951 & ~n26964 ) ;
  assign n26966 = ( ~n26960 & n26962 ) | ( ~n26960 & n26965 ) | ( n26962 & n26965 ) ;
  assign n26967 = ~n26960 & n26966 ;
  assign n26968 = n26950 ^ x785 ^ 1'b0 ;
  assign n26969 = ( n26950 & n26967 ) | ( n26950 & n26968 ) | ( n26967 & n26968 ) ;
  assign n26970 = x618 & ~n26969 ;
  assign n26971 = n26875 ^ n16234 ^ 1'b0 ;
  assign n26972 = ( n26875 & n26954 ) | ( n26875 & ~n26971 ) | ( n26954 & ~n26971 ) ;
  assign n26973 = x618 | n26972 ;
  assign n26974 = ( x1154 & n26970 ) | ( x1154 & n26973 ) | ( n26970 & n26973 ) ;
  assign n26975 = ~n26970 & n26974 ;
  assign n26881 = n26880 ^ x1155 ^ 1'b0 ;
  assign n26883 = ( n26880 & ~n26881 ) | ( n26880 & n26882 ) | ( ~n26881 & n26882 ) ;
  assign n26884 = n26877 ^ x785 ^ 1'b0 ;
  assign n26885 = ( n26877 & n26883 ) | ( n26877 & n26884 ) | ( n26883 & n26884 ) ;
  assign n26886 = x618 & ~n26885 ;
  assign n26890 = x618 & ~n26875 ;
  assign n26891 = x1154 | n26890 ;
  assign n26892 = ( n26885 & n26886 ) | ( n26885 & ~n26891 ) | ( n26886 & ~n26891 ) ;
  assign n26976 = ( x627 & ~n26892 ) | ( x627 & n26975 ) | ( ~n26892 & n26975 ) ;
  assign n26977 = ~n26975 & n26976 ;
  assign n26887 = x618 | n26875 ;
  assign n26888 = ( x1154 & n26886 ) | ( x1154 & n26887 ) | ( n26886 & n26887 ) ;
  assign n26889 = ~n26886 & n26888 ;
  assign n26978 = x627 | n26889 ;
  assign n26979 = x618 & ~n26972 ;
  assign n26980 = x1154 | n26979 ;
  assign n26981 = ( n26969 & n26970 ) | ( n26969 & ~n26980 ) | ( n26970 & ~n26980 ) ;
  assign n26982 = ( ~n26977 & n26978 ) | ( ~n26977 & n26981 ) | ( n26978 & n26981 ) ;
  assign n26983 = ~n26977 & n26982 ;
  assign n26984 = n26969 ^ x781 ^ 1'b0 ;
  assign n26985 = ( n26969 & n26983 ) | ( n26969 & n26984 ) | ( n26983 & n26984 ) ;
  assign n26986 = x619 & ~n26985 ;
  assign n26987 = n26875 ^ n16254 ^ 1'b0 ;
  assign n26988 = ( n26875 & n26972 ) | ( n26875 & ~n26987 ) | ( n26972 & ~n26987 ) ;
  assign n26994 = x619 | n26988 ;
  assign n26995 = ( x1159 & n26986 ) | ( x1159 & n26994 ) | ( n26986 & n26994 ) ;
  assign n26996 = ~n26986 & n26995 ;
  assign n26893 = n26889 | n26892 ;
  assign n26894 = n26885 ^ x781 ^ 1'b0 ;
  assign n26895 = ( n26885 & n26893 ) | ( n26885 & n26894 ) | ( n26893 & n26894 ) ;
  assign n26896 = x619 & ~n26895 ;
  assign n26997 = x619 & ~n26875 ;
  assign n26998 = x1159 | n26997 ;
  assign n26999 = ( n26895 & n26896 ) | ( n26895 & ~n26998 ) | ( n26896 & ~n26998 ) ;
  assign n27000 = ( x648 & n26996 ) | ( x648 & ~n26999 ) | ( n26996 & ~n26999 ) ;
  assign n27001 = ~n26996 & n27000 ;
  assign n26897 = x619 | n26875 ;
  assign n26898 = ( x1159 & n26896 ) | ( x1159 & n26897 ) | ( n26896 & n26897 ) ;
  assign n26899 = ~n26896 & n26898 ;
  assign n26989 = x619 & ~n26988 ;
  assign n26990 = x1159 | n26989 ;
  assign n26991 = ( n26985 & n26986 ) | ( n26985 & ~n26990 ) | ( n26986 & ~n26990 ) ;
  assign n26992 = ( x648 & ~n26899 ) | ( x648 & n26991 ) | ( ~n26899 & n26991 ) ;
  assign n26993 = n26899 | n26992 ;
  assign n27002 = n27001 ^ n26993 ^ 1'b0 ;
  assign n27003 = ( x789 & ~n26993 ) | ( x789 & n27001 ) | ( ~n26993 & n27001 ) ;
  assign n27004 = ( x789 & ~n27002 ) | ( x789 & n27003 ) | ( ~n27002 & n27003 ) ;
  assign n27005 = ( x789 & n26985 ) | ( x789 & ~n27004 ) | ( n26985 & ~n27004 ) ;
  assign n27006 = ~n27004 & n27005 ;
  assign n27007 = ~x626 & n27006 ;
  assign n27008 = n26875 ^ n16279 ^ 1'b0 ;
  assign n27009 = ( n26875 & n26988 ) | ( n26875 & ~n27008 ) | ( n26988 & ~n27008 ) ;
  assign n27010 = x626 & n27009 ;
  assign n27011 = ( x641 & ~n27007 ) | ( x641 & n27010 ) | ( ~n27007 & n27010 ) ;
  assign n27012 = n27007 | n27011 ;
  assign n27013 = ~x626 & n26875 ;
  assign n27014 = n26899 | n26999 ;
  assign n27015 = n26895 ^ x789 ^ 1'b0 ;
  assign n27016 = ( n26895 & n27014 ) | ( n26895 & n27015 ) | ( n27014 & n27015 ) ;
  assign n27017 = x626 & n27016 ;
  assign n27018 = ( x641 & ~n27013 ) | ( x641 & n27017 ) | ( ~n27013 & n27017 ) ;
  assign n27019 = n27013 | n27018 ;
  assign n27020 = ~x626 & n27009 ;
  assign n27021 = x626 & n27006 ;
  assign n27022 = ( x641 & n27020 ) | ( x641 & ~n27021 ) | ( n27020 & ~n27021 ) ;
  assign n27023 = ~n27020 & n27022 ;
  assign n27024 = x1158 & ~n27023 ;
  assign n27025 = n27019 & n27024 ;
  assign n27026 = ~x626 & n27016 ;
  assign n27027 = x626 & n26875 ;
  assign n27028 = x641 & ~n27027 ;
  assign n27029 = n27028 ^ n27026 ^ 1'b0 ;
  assign n27030 = ( n27026 & n27028 ) | ( n27026 & n27029 ) | ( n27028 & n27029 ) ;
  assign n27031 = ( x1158 & ~n27026 ) | ( x1158 & n27030 ) | ( ~n27026 & n27030 ) ;
  assign n27032 = ~n27025 & n27031 ;
  assign n27033 = ( n27012 & n27025 ) | ( n27012 & ~n27032 ) | ( n27025 & ~n27032 ) ;
  assign n27034 = n27006 ^ x788 ^ 1'b0 ;
  assign n27035 = ( n27006 & n27033 ) | ( n27006 & n27034 ) | ( n27033 & n27034 ) ;
  assign n27036 = x628 & ~n27035 ;
  assign n27037 = n26875 ^ n16518 ^ 1'b0 ;
  assign n27038 = ( n26875 & n27016 ) | ( n26875 & ~n27037 ) | ( n27016 & ~n27037 ) ;
  assign n27039 = x628 | n27038 ;
  assign n27040 = ( x1156 & n27036 ) | ( x1156 & n27039 ) | ( n27036 & n27039 ) ;
  assign n27041 = ~n27036 & n27040 ;
  assign n27042 = x628 & ~n26875 ;
  assign n27043 = x1156 | n27042 ;
  assign n27044 = n26875 ^ n16318 ^ 1'b0 ;
  assign n27045 = ( n26875 & n27009 ) | ( n26875 & ~n27044 ) | ( n27009 & ~n27044 ) ;
  assign n27046 = x628 & ~n27045 ;
  assign n27047 = ( ~n27043 & n27045 ) | ( ~n27043 & n27046 ) | ( n27045 & n27046 ) ;
  assign n27048 = ( x629 & n27041 ) | ( x629 & ~n27047 ) | ( n27041 & ~n27047 ) ;
  assign n27049 = ~n27041 & n27048 ;
  assign n27050 = x628 | n26875 ;
  assign n27051 = ( x1156 & n27046 ) | ( x1156 & n27050 ) | ( n27046 & n27050 ) ;
  assign n27052 = ~n27046 & n27051 ;
  assign n27053 = x629 | n27052 ;
  assign n27054 = x628 & ~n27038 ;
  assign n27055 = x1156 | n27054 ;
  assign n27056 = ( n27035 & n27036 ) | ( n27035 & ~n27055 ) | ( n27036 & ~n27055 ) ;
  assign n27057 = ( ~n27049 & n27053 ) | ( ~n27049 & n27056 ) | ( n27053 & n27056 ) ;
  assign n27058 = ~n27049 & n27057 ;
  assign n27059 = n27035 ^ x792 ^ 1'b0 ;
  assign n27060 = ( n27035 & n27058 ) | ( n27035 & n27059 ) | ( n27058 & n27059 ) ;
  assign n27061 = x647 & ~n27060 ;
  assign n27062 = n26875 ^ n16339 ^ 1'b0 ;
  assign n27063 = ( n26875 & n27038 ) | ( n26875 & ~n27062 ) | ( n27038 & ~n27062 ) ;
  assign n27064 = x647 | n27063 ;
  assign n27065 = ( x1157 & n27061 ) | ( x1157 & n27064 ) | ( n27061 & n27064 ) ;
  assign n27066 = ~n27061 & n27065 ;
  assign n27067 = x647 & ~n26875 ;
  assign n27068 = x1157 | n27067 ;
  assign n27069 = n27047 | n27052 ;
  assign n27070 = n27045 ^ x792 ^ 1'b0 ;
  assign n27071 = ( n27045 & n27069 ) | ( n27045 & n27070 ) | ( n27069 & n27070 ) ;
  assign n27072 = x647 & ~n27071 ;
  assign n27073 = ( ~n27068 & n27071 ) | ( ~n27068 & n27072 ) | ( n27071 & n27072 ) ;
  assign n27074 = ( x630 & n27066 ) | ( x630 & ~n27073 ) | ( n27066 & ~n27073 ) ;
  assign n27075 = ~n27066 & n27074 ;
  assign n27076 = x647 | n26875 ;
  assign n27077 = ( x1157 & n27072 ) | ( x1157 & n27076 ) | ( n27072 & n27076 ) ;
  assign n27078 = ~n27072 & n27077 ;
  assign n27079 = x630 | n27078 ;
  assign n27080 = x647 & ~n27063 ;
  assign n27081 = x1157 | n27080 ;
  assign n27082 = ( n27060 & n27061 ) | ( n27060 & ~n27081 ) | ( n27061 & ~n27081 ) ;
  assign n27083 = ( ~n27075 & n27079 ) | ( ~n27075 & n27082 ) | ( n27079 & n27082 ) ;
  assign n27084 = ~n27075 & n27083 ;
  assign n27085 = n27060 ^ x787 ^ 1'b0 ;
  assign n27086 = ( n27060 & n27084 ) | ( n27060 & n27085 ) | ( n27084 & n27085 ) ;
  assign n27087 = x644 & ~n27086 ;
  assign n27088 = n27073 | n27078 ;
  assign n27089 = n27071 ^ x787 ^ 1'b0 ;
  assign n27090 = ( n27071 & n27088 ) | ( n27071 & n27089 ) | ( n27088 & n27089 ) ;
  assign n27091 = x644 | n27090 ;
  assign n27092 = ( x715 & n27087 ) | ( x715 & n27091 ) | ( n27087 & n27091 ) ;
  assign n27093 = ~n27087 & n27092 ;
  assign n27094 = x644 | n26875 ;
  assign n27095 = n26875 ^ n16376 ^ 1'b0 ;
  assign n27096 = ( n26875 & n27063 ) | ( n26875 & ~n27095 ) | ( n27063 & ~n27095 ) ;
  assign n27097 = x644 & ~n27096 ;
  assign n27098 = ( x715 & n27094 ) | ( x715 & ~n27097 ) | ( n27094 & ~n27097 ) ;
  assign n27099 = ~x715 & n27098 ;
  assign n27100 = ( x1160 & n27093 ) | ( x1160 & ~n27099 ) | ( n27093 & ~n27099 ) ;
  assign n27101 = ~n27093 & n27100 ;
  assign n27102 = x644 & ~n26875 ;
  assign n27103 = x715 & ~n27102 ;
  assign n27104 = ( n27096 & n27097 ) | ( n27096 & n27103 ) | ( n27097 & n27103 ) ;
  assign n27105 = x644 & ~n27090 ;
  assign n27106 = x715 | n27105 ;
  assign n27107 = ( n27086 & n27087 ) | ( n27086 & ~n27106 ) | ( n27087 & ~n27106 ) ;
  assign n27108 = ( x1160 & ~n27104 ) | ( x1160 & n27107 ) | ( ~n27104 & n27107 ) ;
  assign n27109 = n27104 | n27108 ;
  assign n27110 = ( x790 & n27101 ) | ( x790 & n27109 ) | ( n27101 & n27109 ) ;
  assign n27111 = ~n27101 & n27110 ;
  assign n27112 = ~x790 & n27086 ;
  assign n27113 = ( n7318 & ~n27111 ) | ( n7318 & n27112 ) | ( ~n27111 & n27112 ) ;
  assign n27114 = n27111 | n27113 ;
  assign n27115 = x186 | n1611 ;
  assign n27116 = ~x752 & n15591 ;
  assign n27117 = n27115 & ~n27116 ;
  assign n27118 = n16397 | n27117 ;
  assign n27119 = n16402 | n27117 ;
  assign n27120 = x1155 & n27119 ;
  assign n27121 = n16405 | n27118 ;
  assign n27122 = ~x1155 & n27121 ;
  assign n27123 = n27120 | n27122 ;
  assign n27124 = n27118 ^ x785 ^ 1'b0 ;
  assign n27125 = ( n27118 & n27123 ) | ( n27118 & n27124 ) | ( n27123 & n27124 ) ;
  assign n27126 = n16411 | n27125 ;
  assign n27127 = x1154 & n27126 ;
  assign n27128 = n16414 | n27125 ;
  assign n27129 = ~x1154 & n27128 ;
  assign n27130 = n27127 | n27129 ;
  assign n27131 = n27125 ^ x781 ^ 1'b0 ;
  assign n27132 = ( n27125 & n27130 ) | ( n27125 & n27131 ) | ( n27130 & n27131 ) ;
  assign n27133 = x619 & ~n27132 ;
  assign n27134 = x619 | n27115 ;
  assign n27135 = ( x1159 & n27133 ) | ( x1159 & n27134 ) | ( n27133 & n27134 ) ;
  assign n27136 = ~n27133 & n27135 ;
  assign n27137 = x619 & ~n27115 ;
  assign n27138 = x1159 | n27137 ;
  assign n27139 = ( n27132 & n27133 ) | ( n27132 & ~n27138 ) | ( n27133 & ~n27138 ) ;
  assign n27140 = n27136 | n27139 ;
  assign n27141 = n27132 ^ x789 ^ 1'b0 ;
  assign n27142 = ( n27132 & n27140 ) | ( n27132 & n27141 ) | ( n27140 & n27141 ) ;
  assign n27143 = n27115 ^ n16518 ^ 1'b0 ;
  assign n27144 = ( n27115 & n27142 ) | ( n27115 & ~n27143 ) | ( n27142 & ~n27143 ) ;
  assign n27145 = n27115 ^ n16339 ^ 1'b0 ;
  assign n27146 = ( n27115 & n27144 ) | ( n27115 & ~n27145 ) | ( n27144 & ~n27145 ) ;
  assign n27147 = n19055 & n27146 ;
  assign n27148 = x647 & ~n27115 ;
  assign n27149 = x1157 | n27148 ;
  assign n27150 = x703 & n15778 ;
  assign n27151 = n27115 & ~n27150 ;
  assign n27152 = ~x1153 & n27115 ;
  assign n27153 = ~x625 & n27150 ;
  assign n27154 = n27152 & ~n27153 ;
  assign n27155 = ( x1153 & n27151 ) | ( x1153 & n27153 ) | ( n27151 & n27153 ) ;
  assign n27156 = n27154 | n27155 ;
  assign n27157 = n27151 ^ x778 ^ 1'b0 ;
  assign n27158 = ( n27151 & n27156 ) | ( n27151 & n27157 ) | ( n27156 & n27157 ) ;
  assign n27159 = n16447 | n27158 ;
  assign n27160 = n16449 | n27159 ;
  assign n27161 = n16451 | n27160 ;
  assign n27162 = n16530 | n27161 ;
  assign n27163 = n16560 | n27162 ;
  assign n27164 = ( x647 & ~n27149 ) | ( x647 & n27163 ) | ( ~n27149 & n27163 ) ;
  assign n27165 = ~n27149 & n27164 ;
  assign n27166 = n27115 ^ x647 ^ 1'b0 ;
  assign n27167 = ( n27115 & n27163 ) | ( n27115 & n27166 ) | ( n27163 & n27166 ) ;
  assign n27168 = x1157 & n27167 ;
  assign n27169 = ( n16375 & n27165 ) | ( n16375 & n27168 ) | ( n27165 & n27168 ) ;
  assign n27170 = ( x787 & n27147 ) | ( x787 & n27169 ) | ( n27147 & n27169 ) ;
  assign n27171 = n27169 ^ n27147 ^ 1'b0 ;
  assign n27172 = ( x787 & n27170 ) | ( x787 & n27171 ) | ( n27170 & n27171 ) ;
  assign n27173 = ~x626 & n27115 ;
  assign n27174 = x626 & n27142 ;
  assign n27175 = ( n22317 & n27173 ) | ( n22317 & ~n27174 ) | ( n27173 & ~n27174 ) ;
  assign n27176 = ~n27173 & n27175 ;
  assign n27177 = ~x626 & n27142 ;
  assign n27178 = x626 & n27115 ;
  assign n27179 = ( n22322 & n27177 ) | ( n22322 & ~n27178 ) | ( n27177 & ~n27178 ) ;
  assign n27180 = ~n27177 & n27179 ;
  assign n27181 = n27161 & ~n27180 ;
  assign n27182 = ( n16459 & n27180 ) | ( n16459 & ~n27181 ) | ( n27180 & ~n27181 ) ;
  assign n27183 = ( x788 & n27176 ) | ( x788 & n27182 ) | ( n27176 & n27182 ) ;
  assign n27184 = n27182 ^ n27176 ^ 1'b0 ;
  assign n27185 = ( x788 & n27183 ) | ( x788 & n27184 ) | ( n27183 & n27184 ) ;
  assign n27186 = n15524 | n27151 ;
  assign n27187 = n27117 & n27186 ;
  assign n27188 = x625 & ~n27186 ;
  assign n27189 = ( n27152 & n27187 ) | ( n27152 & n27188 ) | ( n27187 & n27188 ) ;
  assign n27190 = ( x608 & n27155 ) | ( x608 & ~n27189 ) | ( n27155 & ~n27189 ) ;
  assign n27191 = n27189 | n27190 ;
  assign n27192 = x1153 & n27117 ;
  assign n27193 = ~n27188 & n27192 ;
  assign n27194 = x608 & ~n27154 ;
  assign n27195 = n27191 & ~n27194 ;
  assign n27196 = ( n27191 & n27193 ) | ( n27191 & n27195 ) | ( n27193 & n27195 ) ;
  assign n27197 = n27187 ^ x778 ^ 1'b0 ;
  assign n27198 = ( n27187 & n27196 ) | ( n27187 & n27197 ) | ( n27196 & n27197 ) ;
  assign n27199 = x609 & ~n27198 ;
  assign n27200 = x609 | n27158 ;
  assign n27201 = ( x1155 & n27199 ) | ( x1155 & n27200 ) | ( n27199 & n27200 ) ;
  assign n27202 = ~n27199 & n27201 ;
  assign n27203 = ( x660 & n27122 ) | ( x660 & ~n27202 ) | ( n27122 & ~n27202 ) ;
  assign n27204 = ~n27122 & n27203 ;
  assign n27205 = x660 | n27120 ;
  assign n27206 = x609 & ~n27158 ;
  assign n27207 = x1155 | n27206 ;
  assign n27208 = ( n27198 & n27199 ) | ( n27198 & ~n27207 ) | ( n27199 & ~n27207 ) ;
  assign n27209 = ( ~n27204 & n27205 ) | ( ~n27204 & n27208 ) | ( n27205 & n27208 ) ;
  assign n27210 = ~n27204 & n27209 ;
  assign n27211 = n27198 ^ x785 ^ 1'b0 ;
  assign n27212 = ( n27198 & n27210 ) | ( n27198 & n27211 ) | ( n27210 & n27211 ) ;
  assign n27213 = x618 & ~n27212 ;
  assign n27214 = x618 | n27159 ;
  assign n27215 = ( x1154 & n27213 ) | ( x1154 & n27214 ) | ( n27213 & n27214 ) ;
  assign n27216 = ~n27213 & n27215 ;
  assign n27217 = ( x627 & n27129 ) | ( x627 & ~n27216 ) | ( n27129 & ~n27216 ) ;
  assign n27218 = ~n27129 & n27217 ;
  assign n27219 = x627 | n27127 ;
  assign n27220 = x618 & ~n27159 ;
  assign n27221 = x1154 | n27220 ;
  assign n27222 = ( n27212 & n27213 ) | ( n27212 & ~n27221 ) | ( n27213 & ~n27221 ) ;
  assign n27223 = ( ~n27218 & n27219 ) | ( ~n27218 & n27222 ) | ( n27219 & n27222 ) ;
  assign n27224 = ~n27218 & n27223 ;
  assign n27225 = n27212 ^ x781 ^ 1'b0 ;
  assign n27226 = ( n27212 & n27224 ) | ( n27212 & n27225 ) | ( n27224 & n27225 ) ;
  assign n27227 = ~x789 & n27226 ;
  assign n27228 = x619 & ~n27160 ;
  assign n27229 = x1159 | n27228 ;
  assign n27230 = x619 & ~n27226 ;
  assign n27231 = ( n27226 & ~n27229 ) | ( n27226 & n27230 ) | ( ~n27229 & n27230 ) ;
  assign n27232 = ( x648 & n27136 ) | ( x648 & ~n27231 ) | ( n27136 & ~n27231 ) ;
  assign n27233 = n27231 | n27232 ;
  assign n27234 = x619 | n27160 ;
  assign n27235 = x1159 & ~n27230 ;
  assign n27236 = n27234 & n27235 ;
  assign n27237 = ( x648 & n27139 ) | ( x648 & ~n27236 ) | ( n27139 & ~n27236 ) ;
  assign n27238 = ~n27139 & n27237 ;
  assign n27239 = x789 & ~n27238 ;
  assign n27240 = n27233 & n27239 ;
  assign n27241 = ( n16519 & ~n27227 ) | ( n16519 & n27240 ) | ( ~n27227 & n27240 ) ;
  assign n27242 = n27227 | n27241 ;
  assign n27243 = n27242 ^ n27185 ^ 1'b0 ;
  assign n27244 = ( n27185 & n27242 ) | ( n27185 & n27243 ) | ( n27242 & n27243 ) ;
  assign n27245 = ( n18482 & ~n27185 ) | ( n18482 & n27244 ) | ( ~n27185 & n27244 ) ;
  assign n27246 = n19208 | n27162 ;
  assign n27247 = n16556 & ~n27144 ;
  assign n27248 = x629 & ~n27247 ;
  assign n27249 = n27246 & n27248 ;
  assign n27250 = n16557 & ~n27144 ;
  assign n27251 = n19212 & ~n27162 ;
  assign n27252 = n27250 | n27251 ;
  assign n27253 = ( x629 & ~n27249 ) | ( x629 & n27252 ) | ( ~n27249 & n27252 ) ;
  assign n27254 = ~n27249 & n27253 ;
  assign n27255 = ( x792 & ~n19206 ) | ( x792 & n27254 ) | ( ~n19206 & n27254 ) ;
  assign n27256 = ( n18484 & n19206 ) | ( n18484 & n27255 ) | ( n19206 & n27255 ) ;
  assign n27257 = ( n27172 & n27245 ) | ( n27172 & ~n27256 ) | ( n27245 & ~n27256 ) ;
  assign n27258 = n27257 ^ n27245 ^ 1'b0 ;
  assign n27259 = ( n27172 & n27257 ) | ( n27172 & ~n27258 ) | ( n27257 & ~n27258 ) ;
  assign n27260 = x790 | n27259 ;
  assign n27261 = x644 & ~n27259 ;
  assign n27262 = ( x787 & n27165 ) | ( x787 & ~n27168 ) | ( n27165 & ~n27168 ) ;
  assign n27263 = ~n27165 & n27262 ;
  assign n27264 = ( x787 & n27163 ) | ( x787 & ~n27263 ) | ( n27163 & ~n27263 ) ;
  assign n27265 = ~n27263 & n27264 ;
  assign n27266 = x644 | n27265 ;
  assign n27267 = ( x715 & n27261 ) | ( x715 & n27266 ) | ( n27261 & n27266 ) ;
  assign n27268 = ~n27261 & n27267 ;
  assign n27269 = x644 | n27115 ;
  assign n27270 = n27115 ^ n16376 ^ 1'b0 ;
  assign n27271 = ( n27115 & n27146 ) | ( n27115 & ~n27270 ) | ( n27146 & ~n27270 ) ;
  assign n27272 = x644 & ~n27271 ;
  assign n27273 = ( x715 & n27269 ) | ( x715 & ~n27272 ) | ( n27269 & ~n27272 ) ;
  assign n27274 = ~x715 & n27273 ;
  assign n27275 = ( x1160 & n27268 ) | ( x1160 & ~n27274 ) | ( n27268 & ~n27274 ) ;
  assign n27276 = ~n27268 & n27275 ;
  assign n27277 = x644 & ~n27115 ;
  assign n27278 = x715 & ~n27277 ;
  assign n27279 = ( n27271 & n27272 ) | ( n27271 & n27278 ) | ( n27272 & n27278 ) ;
  assign n27280 = x644 & ~n27265 ;
  assign n27281 = x715 | n27280 ;
  assign n27282 = ( n27259 & n27261 ) | ( n27259 & ~n27281 ) | ( n27261 & ~n27281 ) ;
  assign n27283 = ( x1160 & ~n27279 ) | ( x1160 & n27282 ) | ( ~n27279 & n27282 ) ;
  assign n27284 = n27279 | n27283 ;
  assign n27285 = x790 & ~n27284 ;
  assign n27286 = ( x790 & n27276 ) | ( x790 & n27285 ) | ( n27276 & n27285 ) ;
  assign n27287 = x832 & ~n27286 ;
  assign n27288 = n27260 & n27287 ;
  assign n27289 = ~x186 & n7318 ;
  assign n27290 = x832 | n27289 ;
  assign n27291 = ~n27288 & n27290 ;
  assign n27292 = ( n27114 & n27288 ) | ( n27114 & ~n27291 ) | ( n27288 & ~n27291 ) ;
  assign n27293 = x187 | n17839 ;
  assign n27294 = ( x770 & n22572 ) | ( x770 & n27293 ) | ( n22572 & n27293 ) ;
  assign n27295 = ~x770 & n27294 ;
  assign n27296 = ~x770 & n17843 ;
  assign n27297 = n19461 | n27296 ;
  assign n27298 = ( x187 & ~n27295 ) | ( x187 & n27297 ) | ( ~n27295 & n27297 ) ;
  assign n27299 = ~n27295 & n27298 ;
  assign n27330 = x726 | n27299 ;
  assign n27331 = x770 & ~n17882 ;
  assign n27332 = x187 & n17886 ;
  assign n27333 = n27331 & ~n27332 ;
  assign n27334 = x187 | n17893 ;
  assign n27335 = n27333 & n27334 ;
  assign n27336 = x187 | n17902 ;
  assign n27337 = x187 & n17910 ;
  assign n27338 = ( x770 & n27336 ) | ( x770 & ~n27337 ) | ( n27336 & ~n27337 ) ;
  assign n27339 = ~x770 & n27338 ;
  assign n27340 = ( x726 & n27335 ) | ( x726 & ~n27339 ) | ( n27335 & ~n27339 ) ;
  assign n27341 = ~n27335 & n27340 ;
  assign n27342 = ( n2069 & n27330 ) | ( n2069 & ~n27341 ) | ( n27330 & ~n27341 ) ;
  assign n27343 = ~n2069 & n27342 ;
  assign n27344 = n27343 ^ x187 ^ 1'b0 ;
  assign n27345 = ( ~x187 & n2069 ) | ( ~x187 & n27344 ) | ( n2069 & n27344 ) ;
  assign n27346 = ( x187 & n27343 ) | ( x187 & n27345 ) | ( n27343 & n27345 ) ;
  assign n27347 = x625 & ~n27346 ;
  assign n27300 = n27299 ^ n2069 ^ 1'b0 ;
  assign n27301 = ( x187 & n27299 ) | ( x187 & n27300 ) | ( n27299 & n27300 ) ;
  assign n27348 = x625 | n27301 ;
  assign n27349 = ( x1153 & n27347 ) | ( x1153 & n27348 ) | ( n27347 & n27348 ) ;
  assign n27350 = ~n27347 & n27349 ;
  assign n27302 = x187 | n15656 ;
  assign n27351 = x625 & ~n27302 ;
  assign n27352 = x1153 | n27351 ;
  assign n27353 = ( x38 & x187 ) | ( x38 & n16700 ) | ( x187 & n16700 ) ;
  assign n27354 = ( x187 & n16697 ) | ( x187 & ~n27353 ) | ( n16697 & ~n27353 ) ;
  assign n27355 = ~n27353 & n27354 ;
  assign n27356 = x187 | n15644 ;
  assign n27357 = n16185 & n27356 ;
  assign n27358 = ( x726 & n27355 ) | ( x726 & ~n27357 ) | ( n27355 & ~n27357 ) ;
  assign n27359 = ~n27355 & n27358 ;
  assign n27360 = x187 | x726 ;
  assign n27361 = n15655 | n27360 ;
  assign n27362 = ( n2069 & ~n27359 ) | ( n2069 & n27361 ) | ( ~n27359 & n27361 ) ;
  assign n27363 = ~n2069 & n27362 ;
  assign n27364 = n27363 ^ x187 ^ 1'b0 ;
  assign n27365 = ( ~x187 & n2069 ) | ( ~x187 & n27364 ) | ( n2069 & n27364 ) ;
  assign n27366 = ( x187 & n27363 ) | ( x187 & n27365 ) | ( n27363 & n27365 ) ;
  assign n27367 = ( x625 & ~n27352 ) | ( x625 & n27366 ) | ( ~n27352 & n27366 ) ;
  assign n27368 = ~n27352 & n27367 ;
  assign n27369 = ( x608 & n27350 ) | ( x608 & ~n27368 ) | ( n27350 & ~n27368 ) ;
  assign n27370 = ~n27350 & n27369 ;
  assign n27371 = x625 & ~n27301 ;
  assign n27372 = x1153 | n27371 ;
  assign n27373 = ( x625 & n27346 ) | ( x625 & ~n27372 ) | ( n27346 & ~n27372 ) ;
  assign n27374 = ~n27372 & n27373 ;
  assign n27375 = x625 & ~n27366 ;
  assign n27376 = x625 | n27302 ;
  assign n27377 = ( x1153 & n27375 ) | ( x1153 & n27376 ) | ( n27375 & n27376 ) ;
  assign n27378 = ~n27375 & n27377 ;
  assign n27379 = x608 | n27378 ;
  assign n27380 = ( ~n27370 & n27374 ) | ( ~n27370 & n27379 ) | ( n27374 & n27379 ) ;
  assign n27381 = ~n27370 & n27380 ;
  assign n27382 = n27346 ^ x778 ^ 1'b0 ;
  assign n27383 = ( n27346 & n27381 ) | ( n27346 & n27382 ) | ( n27381 & n27382 ) ;
  assign n27384 = x609 & ~n27383 ;
  assign n27385 = n27368 | n27378 ;
  assign n27386 = n27366 ^ x778 ^ 1'b0 ;
  assign n27387 = ( n27366 & n27385 ) | ( n27366 & n27386 ) | ( n27385 & n27386 ) ;
  assign n27388 = x609 | n27387 ;
  assign n27389 = ( x1155 & n27384 ) | ( x1155 & n27388 ) | ( n27384 & n27388 ) ;
  assign n27390 = ~n27384 & n27389 ;
  assign n27305 = ~n15659 & n27301 ;
  assign n27306 = ~x609 & n27305 ;
  assign n27307 = n15662 & n27302 ;
  assign n27308 = n27306 | n27307 ;
  assign n27391 = ~x1155 & n27308 ;
  assign n27392 = ( x660 & n27390 ) | ( x660 & ~n27391 ) | ( n27390 & ~n27391 ) ;
  assign n27393 = ~n27390 & n27392 ;
  assign n27309 = x609 & n27305 ;
  assign n27310 = ~n15668 & n27302 ;
  assign n27311 = n27309 | n27310 ;
  assign n27394 = x1155 & n27311 ;
  assign n27395 = x660 | n27394 ;
  assign n27396 = x609 & ~n27387 ;
  assign n27397 = x1155 | n27396 ;
  assign n27398 = ( n27383 & n27384 ) | ( n27383 & ~n27397 ) | ( n27384 & ~n27397 ) ;
  assign n27399 = ( ~n27393 & n27395 ) | ( ~n27393 & n27398 ) | ( n27395 & n27398 ) ;
  assign n27400 = ~n27393 & n27399 ;
  assign n27401 = n27383 ^ x785 ^ 1'b0 ;
  assign n27402 = ( n27383 & n27400 ) | ( n27383 & n27401 ) | ( n27400 & n27401 ) ;
  assign n27403 = x618 & ~n27402 ;
  assign n27404 = n27302 ^ n16234 ^ 1'b0 ;
  assign n27405 = ( n27302 & n27387 ) | ( n27302 & ~n27404 ) | ( n27387 & ~n27404 ) ;
  assign n27406 = x618 | n27405 ;
  assign n27407 = ( x1154 & n27403 ) | ( x1154 & n27406 ) | ( n27403 & n27406 ) ;
  assign n27408 = ~n27403 & n27407 ;
  assign n27303 = n27301 ^ n15659 ^ 1'b0 ;
  assign n27304 = ( n27301 & n27302 ) | ( n27301 & n27303 ) | ( n27302 & n27303 ) ;
  assign n27312 = n27311 ^ x1155 ^ 1'b0 ;
  assign n27313 = ( n27308 & n27311 ) | ( n27308 & ~n27312 ) | ( n27311 & ~n27312 ) ;
  assign n27314 = n27304 ^ x785 ^ 1'b0 ;
  assign n27315 = ( n27304 & n27313 ) | ( n27304 & n27314 ) | ( n27313 & n27314 ) ;
  assign n27316 = x618 & ~n27315 ;
  assign n27320 = x618 & ~n27302 ;
  assign n27321 = x1154 | n27320 ;
  assign n27322 = ( n27315 & n27316 ) | ( n27315 & ~n27321 ) | ( n27316 & ~n27321 ) ;
  assign n27409 = ( x627 & ~n27322 ) | ( x627 & n27408 ) | ( ~n27322 & n27408 ) ;
  assign n27410 = ~n27408 & n27409 ;
  assign n27317 = x618 | n27302 ;
  assign n27318 = ( x1154 & n27316 ) | ( x1154 & n27317 ) | ( n27316 & n27317 ) ;
  assign n27319 = ~n27316 & n27318 ;
  assign n27411 = x627 | n27319 ;
  assign n27412 = x618 & ~n27405 ;
  assign n27413 = x1154 | n27412 ;
  assign n27414 = ( n27402 & n27403 ) | ( n27402 & ~n27413 ) | ( n27403 & ~n27413 ) ;
  assign n27415 = ( ~n27410 & n27411 ) | ( ~n27410 & n27414 ) | ( n27411 & n27414 ) ;
  assign n27416 = ~n27410 & n27415 ;
  assign n27417 = n27402 ^ x781 ^ 1'b0 ;
  assign n27418 = ( n27402 & n27416 ) | ( n27402 & n27417 ) | ( n27416 & n27417 ) ;
  assign n27419 = x619 & ~n27418 ;
  assign n27420 = n27302 ^ n16254 ^ 1'b0 ;
  assign n27421 = ( n27302 & n27405 ) | ( n27302 & ~n27420 ) | ( n27405 & ~n27420 ) ;
  assign n27427 = x619 | n27421 ;
  assign n27428 = ( x1159 & n27419 ) | ( x1159 & n27427 ) | ( n27419 & n27427 ) ;
  assign n27429 = ~n27419 & n27428 ;
  assign n27323 = n27319 | n27322 ;
  assign n27324 = n27315 ^ x781 ^ 1'b0 ;
  assign n27325 = ( n27315 & n27323 ) | ( n27315 & n27324 ) | ( n27323 & n27324 ) ;
  assign n27326 = x619 & ~n27325 ;
  assign n27430 = x619 & ~n27302 ;
  assign n27431 = x1159 | n27430 ;
  assign n27432 = ( n27325 & n27326 ) | ( n27325 & ~n27431 ) | ( n27326 & ~n27431 ) ;
  assign n27433 = ( x648 & n27429 ) | ( x648 & ~n27432 ) | ( n27429 & ~n27432 ) ;
  assign n27434 = ~n27429 & n27433 ;
  assign n27327 = x619 | n27302 ;
  assign n27328 = ( x1159 & n27326 ) | ( x1159 & n27327 ) | ( n27326 & n27327 ) ;
  assign n27329 = ~n27326 & n27328 ;
  assign n27422 = x619 & ~n27421 ;
  assign n27423 = x1159 | n27422 ;
  assign n27424 = ( n27418 & n27419 ) | ( n27418 & ~n27423 ) | ( n27419 & ~n27423 ) ;
  assign n27425 = ( x648 & ~n27329 ) | ( x648 & n27424 ) | ( ~n27329 & n27424 ) ;
  assign n27426 = n27329 | n27425 ;
  assign n27435 = n27434 ^ n27426 ^ 1'b0 ;
  assign n27436 = ( x789 & ~n27426 ) | ( x789 & n27434 ) | ( ~n27426 & n27434 ) ;
  assign n27437 = ( x789 & ~n27435 ) | ( x789 & n27436 ) | ( ~n27435 & n27436 ) ;
  assign n27438 = ( x789 & n27418 ) | ( x789 & ~n27437 ) | ( n27418 & ~n27437 ) ;
  assign n27439 = ~n27437 & n27438 ;
  assign n27440 = ~x626 & n27439 ;
  assign n27441 = n27302 ^ n16279 ^ 1'b0 ;
  assign n27442 = ( n27302 & n27421 ) | ( n27302 & ~n27441 ) | ( n27421 & ~n27441 ) ;
  assign n27443 = x626 & n27442 ;
  assign n27444 = ( x641 & ~n27440 ) | ( x641 & n27443 ) | ( ~n27440 & n27443 ) ;
  assign n27445 = n27440 | n27444 ;
  assign n27446 = ~x626 & n27302 ;
  assign n27447 = n27329 | n27432 ;
  assign n27448 = n27325 ^ x789 ^ 1'b0 ;
  assign n27449 = ( n27325 & n27447 ) | ( n27325 & n27448 ) | ( n27447 & n27448 ) ;
  assign n27450 = x626 & n27449 ;
  assign n27451 = ( x641 & ~n27446 ) | ( x641 & n27450 ) | ( ~n27446 & n27450 ) ;
  assign n27452 = n27446 | n27451 ;
  assign n27453 = ~x626 & n27442 ;
  assign n27454 = x626 & n27439 ;
  assign n27455 = ( x641 & n27453 ) | ( x641 & ~n27454 ) | ( n27453 & ~n27454 ) ;
  assign n27456 = ~n27453 & n27455 ;
  assign n27457 = x1158 & ~n27456 ;
  assign n27458 = n27452 & n27457 ;
  assign n27459 = ~x626 & n27449 ;
  assign n27460 = x626 & n27302 ;
  assign n27461 = x641 & ~n27460 ;
  assign n27462 = n27461 ^ n27459 ^ 1'b0 ;
  assign n27463 = ( n27459 & n27461 ) | ( n27459 & n27462 ) | ( n27461 & n27462 ) ;
  assign n27464 = ( x1158 & ~n27459 ) | ( x1158 & n27463 ) | ( ~n27459 & n27463 ) ;
  assign n27465 = ~n27458 & n27464 ;
  assign n27466 = ( n27445 & n27458 ) | ( n27445 & ~n27465 ) | ( n27458 & ~n27465 ) ;
  assign n27467 = n27439 ^ x788 ^ 1'b0 ;
  assign n27468 = ( n27439 & n27466 ) | ( n27439 & n27467 ) | ( n27466 & n27467 ) ;
  assign n27469 = x628 & ~n27468 ;
  assign n27470 = n27302 ^ n16518 ^ 1'b0 ;
  assign n27471 = ( n27302 & n27449 ) | ( n27302 & ~n27470 ) | ( n27449 & ~n27470 ) ;
  assign n27472 = x628 | n27471 ;
  assign n27473 = ( x1156 & n27469 ) | ( x1156 & n27472 ) | ( n27469 & n27472 ) ;
  assign n27474 = ~n27469 & n27473 ;
  assign n27475 = x628 & ~n27302 ;
  assign n27476 = x1156 | n27475 ;
  assign n27477 = n27302 ^ n16318 ^ 1'b0 ;
  assign n27478 = ( n27302 & n27442 ) | ( n27302 & ~n27477 ) | ( n27442 & ~n27477 ) ;
  assign n27479 = x628 & ~n27478 ;
  assign n27480 = ( ~n27476 & n27478 ) | ( ~n27476 & n27479 ) | ( n27478 & n27479 ) ;
  assign n27481 = ( x629 & n27474 ) | ( x629 & ~n27480 ) | ( n27474 & ~n27480 ) ;
  assign n27482 = ~n27474 & n27481 ;
  assign n27483 = x628 | n27302 ;
  assign n27484 = ( x1156 & n27479 ) | ( x1156 & n27483 ) | ( n27479 & n27483 ) ;
  assign n27485 = ~n27479 & n27484 ;
  assign n27486 = x629 | n27485 ;
  assign n27487 = x628 & ~n27471 ;
  assign n27488 = x1156 | n27487 ;
  assign n27489 = ( n27468 & n27469 ) | ( n27468 & ~n27488 ) | ( n27469 & ~n27488 ) ;
  assign n27490 = ( ~n27482 & n27486 ) | ( ~n27482 & n27489 ) | ( n27486 & n27489 ) ;
  assign n27491 = ~n27482 & n27490 ;
  assign n27492 = n27468 ^ x792 ^ 1'b0 ;
  assign n27493 = ( n27468 & n27491 ) | ( n27468 & n27492 ) | ( n27491 & n27492 ) ;
  assign n27494 = x647 & ~n27493 ;
  assign n27495 = n27302 ^ n16339 ^ 1'b0 ;
  assign n27496 = ( n27302 & n27471 ) | ( n27302 & ~n27495 ) | ( n27471 & ~n27495 ) ;
  assign n27497 = x647 | n27496 ;
  assign n27498 = ( x1157 & n27494 ) | ( x1157 & n27497 ) | ( n27494 & n27497 ) ;
  assign n27499 = ~n27494 & n27498 ;
  assign n27500 = x647 & ~n27302 ;
  assign n27501 = x1157 | n27500 ;
  assign n27502 = n27480 | n27485 ;
  assign n27503 = n27478 ^ x792 ^ 1'b0 ;
  assign n27504 = ( n27478 & n27502 ) | ( n27478 & n27503 ) | ( n27502 & n27503 ) ;
  assign n27505 = x647 & ~n27504 ;
  assign n27506 = ( ~n27501 & n27504 ) | ( ~n27501 & n27505 ) | ( n27504 & n27505 ) ;
  assign n27507 = ( x630 & n27499 ) | ( x630 & ~n27506 ) | ( n27499 & ~n27506 ) ;
  assign n27508 = ~n27499 & n27507 ;
  assign n27509 = x647 | n27302 ;
  assign n27510 = ( x1157 & n27505 ) | ( x1157 & n27509 ) | ( n27505 & n27509 ) ;
  assign n27511 = ~n27505 & n27510 ;
  assign n27512 = x630 | n27511 ;
  assign n27513 = x647 & ~n27496 ;
  assign n27514 = x1157 | n27513 ;
  assign n27515 = ( n27493 & n27494 ) | ( n27493 & ~n27514 ) | ( n27494 & ~n27514 ) ;
  assign n27516 = ( ~n27508 & n27512 ) | ( ~n27508 & n27515 ) | ( n27512 & n27515 ) ;
  assign n27517 = ~n27508 & n27516 ;
  assign n27518 = n27493 ^ x787 ^ 1'b0 ;
  assign n27519 = ( n27493 & n27517 ) | ( n27493 & n27518 ) | ( n27517 & n27518 ) ;
  assign n27520 = x644 & ~n27519 ;
  assign n27521 = n27506 | n27511 ;
  assign n27522 = n27504 ^ x787 ^ 1'b0 ;
  assign n27523 = ( n27504 & n27521 ) | ( n27504 & n27522 ) | ( n27521 & n27522 ) ;
  assign n27524 = x644 | n27523 ;
  assign n27525 = ( x715 & n27520 ) | ( x715 & n27524 ) | ( n27520 & n27524 ) ;
  assign n27526 = ~n27520 & n27525 ;
  assign n27527 = x644 | n27302 ;
  assign n27528 = n27302 ^ n16376 ^ 1'b0 ;
  assign n27529 = ( n27302 & n27496 ) | ( n27302 & ~n27528 ) | ( n27496 & ~n27528 ) ;
  assign n27530 = x644 & ~n27529 ;
  assign n27531 = ( x715 & n27527 ) | ( x715 & ~n27530 ) | ( n27527 & ~n27530 ) ;
  assign n27532 = ~x715 & n27531 ;
  assign n27533 = ( x1160 & n27526 ) | ( x1160 & ~n27532 ) | ( n27526 & ~n27532 ) ;
  assign n27534 = ~n27526 & n27533 ;
  assign n27535 = x644 & ~n27302 ;
  assign n27536 = x715 & ~n27535 ;
  assign n27537 = ( n27529 & n27530 ) | ( n27529 & n27536 ) | ( n27530 & n27536 ) ;
  assign n27538 = x644 & ~n27523 ;
  assign n27539 = x715 | n27538 ;
  assign n27540 = ( n27519 & n27520 ) | ( n27519 & ~n27539 ) | ( n27520 & ~n27539 ) ;
  assign n27541 = ( x1160 & ~n27537 ) | ( x1160 & n27540 ) | ( ~n27537 & n27540 ) ;
  assign n27542 = n27537 | n27541 ;
  assign n27543 = ( x790 & n27534 ) | ( x790 & n27542 ) | ( n27534 & n27542 ) ;
  assign n27544 = ~n27534 & n27543 ;
  assign n27545 = ~x790 & n27519 ;
  assign n27546 = ( n7318 & ~n27544 ) | ( n7318 & n27545 ) | ( ~n27544 & n27545 ) ;
  assign n27547 = n27544 | n27546 ;
  assign n27548 = x187 | n1611 ;
  assign n27549 = ~x770 & n15591 ;
  assign n27550 = n27548 & ~n27549 ;
  assign n27551 = n16397 | n27550 ;
  assign n27552 = n16402 | n27550 ;
  assign n27553 = x1155 & n27552 ;
  assign n27554 = n16405 | n27551 ;
  assign n27555 = ~x1155 & n27554 ;
  assign n27556 = n27553 | n27555 ;
  assign n27557 = n27551 ^ x785 ^ 1'b0 ;
  assign n27558 = ( n27551 & n27556 ) | ( n27551 & n27557 ) | ( n27556 & n27557 ) ;
  assign n27559 = n16411 | n27558 ;
  assign n27560 = x1154 & n27559 ;
  assign n27561 = n16414 | n27558 ;
  assign n27562 = ~x1154 & n27561 ;
  assign n27563 = n27560 | n27562 ;
  assign n27564 = n27558 ^ x781 ^ 1'b0 ;
  assign n27565 = ( n27558 & n27563 ) | ( n27558 & n27564 ) | ( n27563 & n27564 ) ;
  assign n27566 = x619 & ~n27565 ;
  assign n27567 = x619 | n27548 ;
  assign n27568 = ( x1159 & n27566 ) | ( x1159 & n27567 ) | ( n27566 & n27567 ) ;
  assign n27569 = ~n27566 & n27568 ;
  assign n27570 = x619 & ~n27548 ;
  assign n27571 = x1159 | n27570 ;
  assign n27572 = ( n27565 & n27566 ) | ( n27565 & ~n27571 ) | ( n27566 & ~n27571 ) ;
  assign n27573 = n27569 | n27572 ;
  assign n27574 = n27565 ^ x789 ^ 1'b0 ;
  assign n27575 = ( n27565 & n27573 ) | ( n27565 & n27574 ) | ( n27573 & n27574 ) ;
  assign n27576 = n27548 ^ n16518 ^ 1'b0 ;
  assign n27577 = ( n27548 & n27575 ) | ( n27548 & ~n27576 ) | ( n27575 & ~n27576 ) ;
  assign n27578 = n27548 ^ n16339 ^ 1'b0 ;
  assign n27579 = ( n27548 & n27577 ) | ( n27548 & ~n27578 ) | ( n27577 & ~n27578 ) ;
  assign n27580 = n19055 & n27579 ;
  assign n27581 = x647 & ~n27548 ;
  assign n27582 = x1157 | n27581 ;
  assign n27583 = x726 & n15778 ;
  assign n27584 = n27548 & ~n27583 ;
  assign n27585 = ~x1153 & n27548 ;
  assign n27586 = ~x625 & n27583 ;
  assign n27587 = n27585 & ~n27586 ;
  assign n27588 = ( x1153 & n27584 ) | ( x1153 & n27586 ) | ( n27584 & n27586 ) ;
  assign n27589 = n27587 | n27588 ;
  assign n27590 = n27584 ^ x778 ^ 1'b0 ;
  assign n27591 = ( n27584 & n27589 ) | ( n27584 & n27590 ) | ( n27589 & n27590 ) ;
  assign n27592 = n16447 | n27591 ;
  assign n27593 = n16449 | n27592 ;
  assign n27594 = n16451 | n27593 ;
  assign n27595 = n16530 | n27594 ;
  assign n27596 = n16560 | n27595 ;
  assign n27597 = ( x647 & ~n27582 ) | ( x647 & n27596 ) | ( ~n27582 & n27596 ) ;
  assign n27598 = ~n27582 & n27597 ;
  assign n27599 = n27548 ^ x647 ^ 1'b0 ;
  assign n27600 = ( n27548 & n27596 ) | ( n27548 & n27599 ) | ( n27596 & n27599 ) ;
  assign n27601 = x1157 & n27600 ;
  assign n27602 = ( n16375 & n27598 ) | ( n16375 & n27601 ) | ( n27598 & n27601 ) ;
  assign n27603 = ( x787 & n27580 ) | ( x787 & n27602 ) | ( n27580 & n27602 ) ;
  assign n27604 = n27602 ^ n27580 ^ 1'b0 ;
  assign n27605 = ( x787 & n27603 ) | ( x787 & n27604 ) | ( n27603 & n27604 ) ;
  assign n27606 = ~x626 & n27548 ;
  assign n27607 = x626 & n27575 ;
  assign n27608 = ( n22317 & n27606 ) | ( n22317 & ~n27607 ) | ( n27606 & ~n27607 ) ;
  assign n27609 = ~n27606 & n27608 ;
  assign n27610 = ~x626 & n27575 ;
  assign n27611 = x626 & n27548 ;
  assign n27612 = ( n22322 & n27610 ) | ( n22322 & ~n27611 ) | ( n27610 & ~n27611 ) ;
  assign n27613 = ~n27610 & n27612 ;
  assign n27614 = n27594 & ~n27613 ;
  assign n27615 = ( n16459 & n27613 ) | ( n16459 & ~n27614 ) | ( n27613 & ~n27614 ) ;
  assign n27616 = ( x788 & n27609 ) | ( x788 & n27615 ) | ( n27609 & n27615 ) ;
  assign n27617 = n27615 ^ n27609 ^ 1'b0 ;
  assign n27618 = ( x788 & n27616 ) | ( x788 & n27617 ) | ( n27616 & n27617 ) ;
  assign n27619 = n15524 | n27584 ;
  assign n27620 = n27550 & n27619 ;
  assign n27621 = x625 & ~n27619 ;
  assign n27622 = ( n27585 & n27620 ) | ( n27585 & n27621 ) | ( n27620 & n27621 ) ;
  assign n27623 = ( x608 & n27588 ) | ( x608 & ~n27622 ) | ( n27588 & ~n27622 ) ;
  assign n27624 = n27622 | n27623 ;
  assign n27625 = x1153 & n27550 ;
  assign n27626 = ~n27621 & n27625 ;
  assign n27627 = x608 & ~n27587 ;
  assign n27628 = n27624 & ~n27627 ;
  assign n27629 = ( n27624 & n27626 ) | ( n27624 & n27628 ) | ( n27626 & n27628 ) ;
  assign n27630 = n27620 ^ x778 ^ 1'b0 ;
  assign n27631 = ( n27620 & n27629 ) | ( n27620 & n27630 ) | ( n27629 & n27630 ) ;
  assign n27632 = x609 & ~n27631 ;
  assign n27633 = x609 | n27591 ;
  assign n27634 = ( x1155 & n27632 ) | ( x1155 & n27633 ) | ( n27632 & n27633 ) ;
  assign n27635 = ~n27632 & n27634 ;
  assign n27636 = ( x660 & n27555 ) | ( x660 & ~n27635 ) | ( n27555 & ~n27635 ) ;
  assign n27637 = ~n27555 & n27636 ;
  assign n27638 = x660 | n27553 ;
  assign n27639 = x609 & ~n27591 ;
  assign n27640 = x1155 | n27639 ;
  assign n27641 = ( n27631 & n27632 ) | ( n27631 & ~n27640 ) | ( n27632 & ~n27640 ) ;
  assign n27642 = ( ~n27637 & n27638 ) | ( ~n27637 & n27641 ) | ( n27638 & n27641 ) ;
  assign n27643 = ~n27637 & n27642 ;
  assign n27644 = n27631 ^ x785 ^ 1'b0 ;
  assign n27645 = ( n27631 & n27643 ) | ( n27631 & n27644 ) | ( n27643 & n27644 ) ;
  assign n27646 = x618 & ~n27645 ;
  assign n27647 = x618 | n27592 ;
  assign n27648 = ( x1154 & n27646 ) | ( x1154 & n27647 ) | ( n27646 & n27647 ) ;
  assign n27649 = ~n27646 & n27648 ;
  assign n27650 = ( x627 & n27562 ) | ( x627 & ~n27649 ) | ( n27562 & ~n27649 ) ;
  assign n27651 = ~n27562 & n27650 ;
  assign n27652 = x627 | n27560 ;
  assign n27653 = x618 & ~n27592 ;
  assign n27654 = x1154 | n27653 ;
  assign n27655 = ( n27645 & n27646 ) | ( n27645 & ~n27654 ) | ( n27646 & ~n27654 ) ;
  assign n27656 = ( ~n27651 & n27652 ) | ( ~n27651 & n27655 ) | ( n27652 & n27655 ) ;
  assign n27657 = ~n27651 & n27656 ;
  assign n27658 = n27645 ^ x781 ^ 1'b0 ;
  assign n27659 = ( n27645 & n27657 ) | ( n27645 & n27658 ) | ( n27657 & n27658 ) ;
  assign n27660 = ~x789 & n27659 ;
  assign n27661 = x619 & ~n27593 ;
  assign n27662 = x1159 | n27661 ;
  assign n27663 = x619 & ~n27659 ;
  assign n27664 = ( n27659 & ~n27662 ) | ( n27659 & n27663 ) | ( ~n27662 & n27663 ) ;
  assign n27665 = ( x648 & n27569 ) | ( x648 & ~n27664 ) | ( n27569 & ~n27664 ) ;
  assign n27666 = n27664 | n27665 ;
  assign n27667 = x619 | n27593 ;
  assign n27668 = x1159 & ~n27663 ;
  assign n27669 = n27667 & n27668 ;
  assign n27670 = ( x648 & n27572 ) | ( x648 & ~n27669 ) | ( n27572 & ~n27669 ) ;
  assign n27671 = ~n27572 & n27670 ;
  assign n27672 = x789 & ~n27671 ;
  assign n27673 = n27666 & n27672 ;
  assign n27674 = ( n16519 & ~n27660 ) | ( n16519 & n27673 ) | ( ~n27660 & n27673 ) ;
  assign n27675 = n27660 | n27674 ;
  assign n27676 = n27675 ^ n27618 ^ 1'b0 ;
  assign n27677 = ( n27618 & n27675 ) | ( n27618 & n27676 ) | ( n27675 & n27676 ) ;
  assign n27678 = ( n18482 & ~n27618 ) | ( n18482 & n27677 ) | ( ~n27618 & n27677 ) ;
  assign n27679 = n19208 | n27595 ;
  assign n27680 = n16556 & ~n27577 ;
  assign n27681 = x629 & ~n27680 ;
  assign n27682 = n27679 & n27681 ;
  assign n27683 = n16557 & ~n27577 ;
  assign n27684 = n19212 & ~n27595 ;
  assign n27685 = n27683 | n27684 ;
  assign n27686 = ( x629 & ~n27682 ) | ( x629 & n27685 ) | ( ~n27682 & n27685 ) ;
  assign n27687 = ~n27682 & n27686 ;
  assign n27688 = ( x792 & ~n19206 ) | ( x792 & n27687 ) | ( ~n19206 & n27687 ) ;
  assign n27689 = ( n18484 & n19206 ) | ( n18484 & n27688 ) | ( n19206 & n27688 ) ;
  assign n27690 = ( n27605 & n27678 ) | ( n27605 & ~n27689 ) | ( n27678 & ~n27689 ) ;
  assign n27691 = n27690 ^ n27678 ^ 1'b0 ;
  assign n27692 = ( n27605 & n27690 ) | ( n27605 & ~n27691 ) | ( n27690 & ~n27691 ) ;
  assign n27693 = x790 | n27692 ;
  assign n27694 = x644 & ~n27692 ;
  assign n27695 = ( x787 & n27598 ) | ( x787 & ~n27601 ) | ( n27598 & ~n27601 ) ;
  assign n27696 = ~n27598 & n27695 ;
  assign n27697 = ( x787 & n27596 ) | ( x787 & ~n27696 ) | ( n27596 & ~n27696 ) ;
  assign n27698 = ~n27696 & n27697 ;
  assign n27699 = x644 | n27698 ;
  assign n27700 = ( x715 & n27694 ) | ( x715 & n27699 ) | ( n27694 & n27699 ) ;
  assign n27701 = ~n27694 & n27700 ;
  assign n27702 = x644 | n27548 ;
  assign n27703 = n27548 ^ n16376 ^ 1'b0 ;
  assign n27704 = ( n27548 & n27579 ) | ( n27548 & ~n27703 ) | ( n27579 & ~n27703 ) ;
  assign n27705 = x644 & ~n27704 ;
  assign n27706 = ( x715 & n27702 ) | ( x715 & ~n27705 ) | ( n27702 & ~n27705 ) ;
  assign n27707 = ~x715 & n27706 ;
  assign n27708 = ( x1160 & n27701 ) | ( x1160 & ~n27707 ) | ( n27701 & ~n27707 ) ;
  assign n27709 = ~n27701 & n27708 ;
  assign n27710 = x644 & ~n27548 ;
  assign n27711 = x715 & ~n27710 ;
  assign n27712 = ( n27704 & n27705 ) | ( n27704 & n27711 ) | ( n27705 & n27711 ) ;
  assign n27713 = x644 & ~n27698 ;
  assign n27714 = x715 | n27713 ;
  assign n27715 = ( n27692 & n27694 ) | ( n27692 & ~n27714 ) | ( n27694 & ~n27714 ) ;
  assign n27716 = ( x1160 & ~n27712 ) | ( x1160 & n27715 ) | ( ~n27712 & n27715 ) ;
  assign n27717 = n27712 | n27716 ;
  assign n27718 = x790 & ~n27717 ;
  assign n27719 = ( x790 & n27709 ) | ( x790 & n27718 ) | ( n27709 & n27718 ) ;
  assign n27720 = x832 & ~n27719 ;
  assign n27721 = n27693 & n27720 ;
  assign n27722 = ~x187 & n7318 ;
  assign n27723 = x832 | n27722 ;
  assign n27724 = ~n27721 & n27723 ;
  assign n27725 = ( n27547 & n27721 ) | ( n27547 & ~n27724 ) | ( n27721 & ~n27724 ) ;
  assign n27726 = x188 | n17839 ;
  assign n27727 = ( x768 & n22572 ) | ( x768 & n27726 ) | ( n22572 & n27726 ) ;
  assign n27728 = ~x768 & n27727 ;
  assign n27729 = n17843 ^ x768 ^ 1'b0 ;
  assign n27730 = ( n15655 & n17843 ) | ( n15655 & n27729 ) | ( n17843 & n27729 ) ;
  assign n27731 = ( x188 & ~n27728 ) | ( x188 & n27730 ) | ( ~n27728 & n27730 ) ;
  assign n27732 = ~n27728 & n27731 ;
  assign n27761 = x705 | n27732 ;
  assign n27762 = x768 & ~n17882 ;
  assign n27763 = x188 & n17886 ;
  assign n27764 = n27762 & ~n27763 ;
  assign n27765 = x188 | n17893 ;
  assign n27766 = n27764 & n27765 ;
  assign n27767 = x188 | n17902 ;
  assign n27768 = x188 & n17910 ;
  assign n27769 = ( x768 & n27767 ) | ( x768 & ~n27768 ) | ( n27767 & ~n27768 ) ;
  assign n27770 = ~x768 & n27769 ;
  assign n27771 = ( x705 & n27766 ) | ( x705 & ~n27770 ) | ( n27766 & ~n27770 ) ;
  assign n27772 = ~n27766 & n27771 ;
  assign n27773 = ( n2069 & n27761 ) | ( n2069 & ~n27772 ) | ( n27761 & ~n27772 ) ;
  assign n27774 = ~n2069 & n27773 ;
  assign n27775 = n27774 ^ x188 ^ 1'b0 ;
  assign n27776 = ( ~x188 & n2069 ) | ( ~x188 & n27775 ) | ( n2069 & n27775 ) ;
  assign n27777 = ( x188 & n27774 ) | ( x188 & n27776 ) | ( n27774 & n27776 ) ;
  assign n27778 = x625 & ~n27777 ;
  assign n27733 = n27732 ^ n2069 ^ 1'b0 ;
  assign n27734 = ( x188 & n27732 ) | ( x188 & n27733 ) | ( n27732 & n27733 ) ;
  assign n27779 = x625 | n27734 ;
  assign n27780 = ( x1153 & n27778 ) | ( x1153 & n27779 ) | ( n27778 & n27779 ) ;
  assign n27781 = ~n27778 & n27780 ;
  assign n27735 = x188 | n15656 ;
  assign n27782 = x625 & ~n27735 ;
  assign n27783 = x1153 | n27782 ;
  assign n27784 = ( x38 & x188 ) | ( x38 & n16700 ) | ( x188 & n16700 ) ;
  assign n27785 = ( x188 & n16697 ) | ( x188 & ~n27784 ) | ( n16697 & ~n27784 ) ;
  assign n27786 = ~n27784 & n27785 ;
  assign n27787 = x188 | n15644 ;
  assign n27788 = n16185 & n27787 ;
  assign n27789 = ( x705 & n27786 ) | ( x705 & ~n27788 ) | ( n27786 & ~n27788 ) ;
  assign n27790 = ~n27786 & n27789 ;
  assign n27791 = x188 | x705 ;
  assign n27792 = n15655 | n27791 ;
  assign n27793 = ( n2069 & ~n27790 ) | ( n2069 & n27792 ) | ( ~n27790 & n27792 ) ;
  assign n27794 = ~n2069 & n27793 ;
  assign n27795 = n27794 ^ x188 ^ 1'b0 ;
  assign n27796 = ( ~x188 & n2069 ) | ( ~x188 & n27795 ) | ( n2069 & n27795 ) ;
  assign n27797 = ( x188 & n27794 ) | ( x188 & n27796 ) | ( n27794 & n27796 ) ;
  assign n27798 = ( x625 & ~n27783 ) | ( x625 & n27797 ) | ( ~n27783 & n27797 ) ;
  assign n27799 = ~n27783 & n27798 ;
  assign n27800 = ( x608 & n27781 ) | ( x608 & ~n27799 ) | ( n27781 & ~n27799 ) ;
  assign n27801 = ~n27781 & n27800 ;
  assign n27802 = x625 & ~n27797 ;
  assign n27803 = x625 | n27735 ;
  assign n27804 = ( x1153 & n27802 ) | ( x1153 & n27803 ) | ( n27802 & n27803 ) ;
  assign n27805 = ~n27802 & n27804 ;
  assign n27806 = x608 | n27805 ;
  assign n27807 = x625 & ~n27734 ;
  assign n27808 = x1153 | n27807 ;
  assign n27809 = ( n27777 & n27778 ) | ( n27777 & ~n27808 ) | ( n27778 & ~n27808 ) ;
  assign n27810 = ( ~n27801 & n27806 ) | ( ~n27801 & n27809 ) | ( n27806 & n27809 ) ;
  assign n27811 = ~n27801 & n27810 ;
  assign n27812 = n27777 ^ x778 ^ 1'b0 ;
  assign n27813 = ( n27777 & n27811 ) | ( n27777 & n27812 ) | ( n27811 & n27812 ) ;
  assign n27814 = x609 & ~n27813 ;
  assign n27815 = n27799 | n27805 ;
  assign n27816 = n27797 ^ x778 ^ 1'b0 ;
  assign n27817 = ( n27797 & n27815 ) | ( n27797 & n27816 ) | ( n27815 & n27816 ) ;
  assign n27818 = x609 | n27817 ;
  assign n27819 = ( x1155 & n27814 ) | ( x1155 & n27818 ) | ( n27814 & n27818 ) ;
  assign n27820 = ~n27814 & n27819 ;
  assign n27738 = ~n15659 & n27734 ;
  assign n27739 = x609 & n27738 ;
  assign n27740 = ~n15668 & n27735 ;
  assign n27741 = n27739 | n27740 ;
  assign n27736 = n27734 ^ n15659 ^ 1'b0 ;
  assign n27737 = ( n27734 & n27735 ) | ( n27734 & n27736 ) | ( n27735 & n27736 ) ;
  assign n27743 = n27741 ^ n27737 ^ n27735 ;
  assign n27821 = ~x1155 & n27743 ;
  assign n27822 = ( x660 & n27820 ) | ( x660 & ~n27821 ) | ( n27820 & ~n27821 ) ;
  assign n27823 = ~n27820 & n27822 ;
  assign n27824 = x1155 & n27741 ;
  assign n27825 = x660 | n27824 ;
  assign n27826 = x609 & ~n27817 ;
  assign n27827 = x1155 | n27826 ;
  assign n27828 = ( n27813 & n27814 ) | ( n27813 & ~n27827 ) | ( n27814 & ~n27827 ) ;
  assign n27829 = ( ~n27823 & n27825 ) | ( ~n27823 & n27828 ) | ( n27825 & n27828 ) ;
  assign n27830 = ~n27823 & n27829 ;
  assign n27831 = n27813 ^ x785 ^ 1'b0 ;
  assign n27832 = ( n27813 & n27830 ) | ( n27813 & n27831 ) | ( n27830 & n27831 ) ;
  assign n27833 = x618 & ~n27832 ;
  assign n27834 = n27735 ^ n16234 ^ 1'b0 ;
  assign n27835 = ( n27735 & n27817 ) | ( n27735 & ~n27834 ) | ( n27817 & ~n27834 ) ;
  assign n27836 = x618 | n27835 ;
  assign n27837 = ( x1154 & n27833 ) | ( x1154 & n27836 ) | ( n27833 & n27836 ) ;
  assign n27838 = ~n27833 & n27837 ;
  assign n27742 = n27741 ^ x1155 ^ 1'b0 ;
  assign n27744 = ( n27741 & ~n27742 ) | ( n27741 & n27743 ) | ( ~n27742 & n27743 ) ;
  assign n27745 = n27737 ^ x785 ^ 1'b0 ;
  assign n27746 = ( n27737 & n27744 ) | ( n27737 & n27745 ) | ( n27744 & n27745 ) ;
  assign n27747 = x618 & ~n27746 ;
  assign n27751 = x618 & ~n27735 ;
  assign n27752 = x1154 | n27751 ;
  assign n27753 = ( n27746 & n27747 ) | ( n27746 & ~n27752 ) | ( n27747 & ~n27752 ) ;
  assign n27839 = ( x627 & ~n27753 ) | ( x627 & n27838 ) | ( ~n27753 & n27838 ) ;
  assign n27840 = ~n27838 & n27839 ;
  assign n27748 = x618 | n27735 ;
  assign n27749 = ( x1154 & n27747 ) | ( x1154 & n27748 ) | ( n27747 & n27748 ) ;
  assign n27750 = ~n27747 & n27749 ;
  assign n27841 = x627 | n27750 ;
  assign n27842 = x618 & ~n27835 ;
  assign n27843 = x1154 | n27842 ;
  assign n27844 = ( n27832 & n27833 ) | ( n27832 & ~n27843 ) | ( n27833 & ~n27843 ) ;
  assign n27845 = ( ~n27840 & n27841 ) | ( ~n27840 & n27844 ) | ( n27841 & n27844 ) ;
  assign n27846 = ~n27840 & n27845 ;
  assign n27847 = n27832 ^ x781 ^ 1'b0 ;
  assign n27848 = ( n27832 & n27846 ) | ( n27832 & n27847 ) | ( n27846 & n27847 ) ;
  assign n27849 = x619 & ~n27848 ;
  assign n27850 = n27735 ^ n16254 ^ 1'b0 ;
  assign n27851 = ( n27735 & n27835 ) | ( n27735 & ~n27850 ) | ( n27835 & ~n27850 ) ;
  assign n27857 = x619 | n27851 ;
  assign n27858 = ( x1159 & n27849 ) | ( x1159 & n27857 ) | ( n27849 & n27857 ) ;
  assign n27859 = ~n27849 & n27858 ;
  assign n27754 = n27750 | n27753 ;
  assign n27755 = n27746 ^ x781 ^ 1'b0 ;
  assign n27756 = ( n27746 & n27754 ) | ( n27746 & n27755 ) | ( n27754 & n27755 ) ;
  assign n27757 = x619 & ~n27756 ;
  assign n27860 = x619 & ~n27735 ;
  assign n27861 = x1159 | n27860 ;
  assign n27862 = ( n27756 & n27757 ) | ( n27756 & ~n27861 ) | ( n27757 & ~n27861 ) ;
  assign n27863 = ( x648 & n27859 ) | ( x648 & ~n27862 ) | ( n27859 & ~n27862 ) ;
  assign n27864 = ~n27859 & n27863 ;
  assign n27758 = x619 | n27735 ;
  assign n27759 = ( x1159 & n27757 ) | ( x1159 & n27758 ) | ( n27757 & n27758 ) ;
  assign n27760 = ~n27757 & n27759 ;
  assign n27852 = x619 & ~n27851 ;
  assign n27853 = x1159 | n27852 ;
  assign n27854 = ( n27848 & n27849 ) | ( n27848 & ~n27853 ) | ( n27849 & ~n27853 ) ;
  assign n27855 = ( x648 & ~n27760 ) | ( x648 & n27854 ) | ( ~n27760 & n27854 ) ;
  assign n27856 = n27760 | n27855 ;
  assign n27865 = n27864 ^ n27856 ^ 1'b0 ;
  assign n27866 = ( x789 & ~n27856 ) | ( x789 & n27864 ) | ( ~n27856 & n27864 ) ;
  assign n27867 = ( x789 & ~n27865 ) | ( x789 & n27866 ) | ( ~n27865 & n27866 ) ;
  assign n27868 = ( x789 & n27848 ) | ( x789 & ~n27867 ) | ( n27848 & ~n27867 ) ;
  assign n27869 = ~n27867 & n27868 ;
  assign n27870 = ~x626 & n27869 ;
  assign n27871 = n27735 ^ n16279 ^ 1'b0 ;
  assign n27872 = ( n27735 & n27851 ) | ( n27735 & ~n27871 ) | ( n27851 & ~n27871 ) ;
  assign n27873 = x626 & n27872 ;
  assign n27874 = ( x641 & ~n27870 ) | ( x641 & n27873 ) | ( ~n27870 & n27873 ) ;
  assign n27875 = n27870 | n27874 ;
  assign n27876 = ~x626 & n27735 ;
  assign n27877 = n27760 | n27862 ;
  assign n27878 = n27756 ^ x789 ^ 1'b0 ;
  assign n27879 = ( n27756 & n27877 ) | ( n27756 & n27878 ) | ( n27877 & n27878 ) ;
  assign n27880 = x626 & n27879 ;
  assign n27881 = ( x641 & ~n27876 ) | ( x641 & n27880 ) | ( ~n27876 & n27880 ) ;
  assign n27882 = n27876 | n27881 ;
  assign n27883 = ~x626 & n27872 ;
  assign n27884 = x626 & n27869 ;
  assign n27885 = ( x641 & n27883 ) | ( x641 & ~n27884 ) | ( n27883 & ~n27884 ) ;
  assign n27886 = ~n27883 & n27885 ;
  assign n27887 = x1158 & ~n27886 ;
  assign n27888 = n27882 & n27887 ;
  assign n27889 = ~x626 & n27879 ;
  assign n27890 = x626 & n27735 ;
  assign n27891 = x641 & ~n27890 ;
  assign n27892 = n27891 ^ n27889 ^ 1'b0 ;
  assign n27893 = ( n27889 & n27891 ) | ( n27889 & n27892 ) | ( n27891 & n27892 ) ;
  assign n27894 = ( x1158 & ~n27889 ) | ( x1158 & n27893 ) | ( ~n27889 & n27893 ) ;
  assign n27895 = ~n27888 & n27894 ;
  assign n27896 = ( n27875 & n27888 ) | ( n27875 & ~n27895 ) | ( n27888 & ~n27895 ) ;
  assign n27897 = n27869 ^ x788 ^ 1'b0 ;
  assign n27898 = ( n27869 & n27896 ) | ( n27869 & n27897 ) | ( n27896 & n27897 ) ;
  assign n27899 = x628 & ~n27898 ;
  assign n27900 = n27735 ^ n16518 ^ 1'b0 ;
  assign n27901 = ( n27735 & n27879 ) | ( n27735 & ~n27900 ) | ( n27879 & ~n27900 ) ;
  assign n27902 = x628 | n27901 ;
  assign n27903 = ( x1156 & n27899 ) | ( x1156 & n27902 ) | ( n27899 & n27902 ) ;
  assign n27904 = ~n27899 & n27903 ;
  assign n27905 = x628 & ~n27735 ;
  assign n27906 = x1156 | n27905 ;
  assign n27907 = n27735 ^ n16318 ^ 1'b0 ;
  assign n27908 = ( n27735 & n27872 ) | ( n27735 & ~n27907 ) | ( n27872 & ~n27907 ) ;
  assign n27909 = x628 & ~n27908 ;
  assign n27910 = ( ~n27906 & n27908 ) | ( ~n27906 & n27909 ) | ( n27908 & n27909 ) ;
  assign n27911 = ( x629 & n27904 ) | ( x629 & ~n27910 ) | ( n27904 & ~n27910 ) ;
  assign n27912 = ~n27904 & n27911 ;
  assign n27913 = x628 | n27735 ;
  assign n27914 = ( x1156 & n27909 ) | ( x1156 & n27913 ) | ( n27909 & n27913 ) ;
  assign n27915 = ~n27909 & n27914 ;
  assign n27916 = x629 | n27915 ;
  assign n27917 = x628 & ~n27901 ;
  assign n27918 = x1156 | n27917 ;
  assign n27919 = ( n27898 & n27899 ) | ( n27898 & ~n27918 ) | ( n27899 & ~n27918 ) ;
  assign n27920 = ( ~n27912 & n27916 ) | ( ~n27912 & n27919 ) | ( n27916 & n27919 ) ;
  assign n27921 = ~n27912 & n27920 ;
  assign n27922 = n27898 ^ x792 ^ 1'b0 ;
  assign n27923 = ( n27898 & n27921 ) | ( n27898 & n27922 ) | ( n27921 & n27922 ) ;
  assign n27924 = x647 & ~n27923 ;
  assign n27925 = n27735 ^ n16339 ^ 1'b0 ;
  assign n27926 = ( n27735 & n27901 ) | ( n27735 & ~n27925 ) | ( n27901 & ~n27925 ) ;
  assign n27927 = x647 | n27926 ;
  assign n27928 = ( x1157 & n27924 ) | ( x1157 & n27927 ) | ( n27924 & n27927 ) ;
  assign n27929 = ~n27924 & n27928 ;
  assign n27930 = x647 & ~n27735 ;
  assign n27931 = x1157 | n27930 ;
  assign n27932 = n27910 | n27915 ;
  assign n27933 = n27908 ^ x792 ^ 1'b0 ;
  assign n27934 = ( n27908 & n27932 ) | ( n27908 & n27933 ) | ( n27932 & n27933 ) ;
  assign n27935 = x647 & ~n27934 ;
  assign n27936 = ( ~n27931 & n27934 ) | ( ~n27931 & n27935 ) | ( n27934 & n27935 ) ;
  assign n27937 = ( x630 & n27929 ) | ( x630 & ~n27936 ) | ( n27929 & ~n27936 ) ;
  assign n27938 = ~n27929 & n27937 ;
  assign n27939 = x647 | n27735 ;
  assign n27940 = ( x1157 & n27935 ) | ( x1157 & n27939 ) | ( n27935 & n27939 ) ;
  assign n27941 = ~n27935 & n27940 ;
  assign n27942 = x630 | n27941 ;
  assign n27943 = x647 & ~n27926 ;
  assign n27944 = x1157 | n27943 ;
  assign n27945 = ( n27923 & n27924 ) | ( n27923 & ~n27944 ) | ( n27924 & ~n27944 ) ;
  assign n27946 = ( ~n27938 & n27942 ) | ( ~n27938 & n27945 ) | ( n27942 & n27945 ) ;
  assign n27947 = ~n27938 & n27946 ;
  assign n27948 = n27923 ^ x787 ^ 1'b0 ;
  assign n27949 = ( n27923 & n27947 ) | ( n27923 & n27948 ) | ( n27947 & n27948 ) ;
  assign n27950 = x644 & ~n27949 ;
  assign n27951 = n27936 | n27941 ;
  assign n27952 = n27934 ^ x787 ^ 1'b0 ;
  assign n27953 = ( n27934 & n27951 ) | ( n27934 & n27952 ) | ( n27951 & n27952 ) ;
  assign n27954 = x644 | n27953 ;
  assign n27955 = ( x715 & n27950 ) | ( x715 & n27954 ) | ( n27950 & n27954 ) ;
  assign n27956 = ~n27950 & n27955 ;
  assign n27957 = x644 | n27735 ;
  assign n27958 = n27735 ^ n16376 ^ 1'b0 ;
  assign n27959 = ( n27735 & n27926 ) | ( n27735 & ~n27958 ) | ( n27926 & ~n27958 ) ;
  assign n27960 = x644 & ~n27959 ;
  assign n27961 = ( x715 & n27957 ) | ( x715 & ~n27960 ) | ( n27957 & ~n27960 ) ;
  assign n27962 = ~x715 & n27961 ;
  assign n27963 = ( x1160 & n27956 ) | ( x1160 & ~n27962 ) | ( n27956 & ~n27962 ) ;
  assign n27964 = ~n27956 & n27963 ;
  assign n27965 = x644 & ~n27735 ;
  assign n27966 = x715 & ~n27965 ;
  assign n27967 = ( n27959 & n27960 ) | ( n27959 & n27966 ) | ( n27960 & n27966 ) ;
  assign n27968 = x644 & ~n27953 ;
  assign n27969 = x715 | n27968 ;
  assign n27970 = ( n27949 & n27950 ) | ( n27949 & ~n27969 ) | ( n27950 & ~n27969 ) ;
  assign n27971 = ( x1160 & ~n27967 ) | ( x1160 & n27970 ) | ( ~n27967 & n27970 ) ;
  assign n27972 = n27967 | n27971 ;
  assign n27973 = ( x790 & n27964 ) | ( x790 & n27972 ) | ( n27964 & n27972 ) ;
  assign n27974 = ~n27964 & n27973 ;
  assign n27975 = ~x790 & n27949 ;
  assign n27976 = ( n7318 & ~n27974 ) | ( n7318 & n27975 ) | ( ~n27974 & n27975 ) ;
  assign n27977 = n27974 | n27976 ;
  assign n27978 = x188 | n1611 ;
  assign n27979 = ~x768 & n15591 ;
  assign n27980 = n27978 & ~n27979 ;
  assign n27981 = n16397 | n27980 ;
  assign n27982 = n16402 | n27980 ;
  assign n27983 = x1155 & n27982 ;
  assign n27984 = n16405 | n27981 ;
  assign n27985 = ~x1155 & n27984 ;
  assign n27986 = n27983 | n27985 ;
  assign n27987 = n27981 ^ x785 ^ 1'b0 ;
  assign n27988 = ( n27981 & n27986 ) | ( n27981 & n27987 ) | ( n27986 & n27987 ) ;
  assign n27989 = n16411 | n27988 ;
  assign n27990 = x1154 & n27989 ;
  assign n27991 = n16414 | n27988 ;
  assign n27992 = ~x1154 & n27991 ;
  assign n27993 = n27990 | n27992 ;
  assign n27994 = n27988 ^ x781 ^ 1'b0 ;
  assign n27995 = ( n27988 & n27993 ) | ( n27988 & n27994 ) | ( n27993 & n27994 ) ;
  assign n27996 = x619 & ~n27995 ;
  assign n27997 = x619 | n27978 ;
  assign n27998 = ( x1159 & n27996 ) | ( x1159 & n27997 ) | ( n27996 & n27997 ) ;
  assign n27999 = ~n27996 & n27998 ;
  assign n28000 = x619 & ~n27978 ;
  assign n28001 = x1159 | n28000 ;
  assign n28002 = ( n27995 & n27996 ) | ( n27995 & ~n28001 ) | ( n27996 & ~n28001 ) ;
  assign n28003 = n27999 | n28002 ;
  assign n28004 = n27995 ^ x789 ^ 1'b0 ;
  assign n28005 = ( n27995 & n28003 ) | ( n27995 & n28004 ) | ( n28003 & n28004 ) ;
  assign n28006 = n27978 ^ n16518 ^ 1'b0 ;
  assign n28007 = ( n27978 & n28005 ) | ( n27978 & ~n28006 ) | ( n28005 & ~n28006 ) ;
  assign n28008 = n27978 ^ n16339 ^ 1'b0 ;
  assign n28009 = ( n27978 & n28007 ) | ( n27978 & ~n28008 ) | ( n28007 & ~n28008 ) ;
  assign n28010 = n19055 & n28009 ;
  assign n28011 = x647 & ~n27978 ;
  assign n28012 = x1157 | n28011 ;
  assign n28013 = x705 & n15778 ;
  assign n28014 = n27978 & ~n28013 ;
  assign n28015 = ~x1153 & n27978 ;
  assign n28016 = ~x625 & n28013 ;
  assign n28017 = n28015 & ~n28016 ;
  assign n28018 = ( x1153 & n28014 ) | ( x1153 & n28016 ) | ( n28014 & n28016 ) ;
  assign n28019 = n28017 | n28018 ;
  assign n28020 = n28014 ^ x778 ^ 1'b0 ;
  assign n28021 = ( n28014 & n28019 ) | ( n28014 & n28020 ) | ( n28019 & n28020 ) ;
  assign n28022 = n16447 | n28021 ;
  assign n28023 = n16449 | n28022 ;
  assign n28024 = n16451 | n28023 ;
  assign n28025 = n16530 | n28024 ;
  assign n28026 = n16560 | n28025 ;
  assign n28027 = ( x647 & ~n28012 ) | ( x647 & n28026 ) | ( ~n28012 & n28026 ) ;
  assign n28028 = ~n28012 & n28027 ;
  assign n28029 = n27978 ^ x647 ^ 1'b0 ;
  assign n28030 = ( n27978 & n28026 ) | ( n27978 & n28029 ) | ( n28026 & n28029 ) ;
  assign n28031 = x1157 & n28030 ;
  assign n28032 = ( n16375 & n28028 ) | ( n16375 & n28031 ) | ( n28028 & n28031 ) ;
  assign n28033 = ( x787 & n28010 ) | ( x787 & n28032 ) | ( n28010 & n28032 ) ;
  assign n28034 = n28032 ^ n28010 ^ 1'b0 ;
  assign n28035 = ( x787 & n28033 ) | ( x787 & n28034 ) | ( n28033 & n28034 ) ;
  assign n28036 = ~x626 & n27978 ;
  assign n28037 = x626 & n28005 ;
  assign n28038 = ( n22317 & n28036 ) | ( n22317 & ~n28037 ) | ( n28036 & ~n28037 ) ;
  assign n28039 = ~n28036 & n28038 ;
  assign n28040 = ~x626 & n28005 ;
  assign n28041 = x626 & n27978 ;
  assign n28042 = ( n22322 & n28040 ) | ( n22322 & ~n28041 ) | ( n28040 & ~n28041 ) ;
  assign n28043 = ~n28040 & n28042 ;
  assign n28044 = n28024 & ~n28043 ;
  assign n28045 = ( n16459 & n28043 ) | ( n16459 & ~n28044 ) | ( n28043 & ~n28044 ) ;
  assign n28046 = ( x788 & n28039 ) | ( x788 & n28045 ) | ( n28039 & n28045 ) ;
  assign n28047 = n28045 ^ n28039 ^ 1'b0 ;
  assign n28048 = ( x788 & n28046 ) | ( x788 & n28047 ) | ( n28046 & n28047 ) ;
  assign n28049 = n15524 | n28014 ;
  assign n28050 = n27980 & n28049 ;
  assign n28051 = x625 & ~n28049 ;
  assign n28052 = ( n28015 & n28050 ) | ( n28015 & n28051 ) | ( n28050 & n28051 ) ;
  assign n28053 = ( x608 & n28018 ) | ( x608 & ~n28052 ) | ( n28018 & ~n28052 ) ;
  assign n28054 = n28052 | n28053 ;
  assign n28055 = x1153 & n27980 ;
  assign n28056 = ~n28051 & n28055 ;
  assign n28057 = x608 & ~n28017 ;
  assign n28058 = n28054 & ~n28057 ;
  assign n28059 = ( n28054 & n28056 ) | ( n28054 & n28058 ) | ( n28056 & n28058 ) ;
  assign n28060 = n28050 ^ x778 ^ 1'b0 ;
  assign n28061 = ( n28050 & n28059 ) | ( n28050 & n28060 ) | ( n28059 & n28060 ) ;
  assign n28062 = x609 & ~n28061 ;
  assign n28063 = x609 | n28021 ;
  assign n28064 = ( x1155 & n28062 ) | ( x1155 & n28063 ) | ( n28062 & n28063 ) ;
  assign n28065 = ~n28062 & n28064 ;
  assign n28066 = ( x660 & n27985 ) | ( x660 & ~n28065 ) | ( n27985 & ~n28065 ) ;
  assign n28067 = ~n27985 & n28066 ;
  assign n28068 = x660 | n27983 ;
  assign n28069 = x609 & ~n28021 ;
  assign n28070 = x1155 | n28069 ;
  assign n28071 = ( n28061 & n28062 ) | ( n28061 & ~n28070 ) | ( n28062 & ~n28070 ) ;
  assign n28072 = ( ~n28067 & n28068 ) | ( ~n28067 & n28071 ) | ( n28068 & n28071 ) ;
  assign n28073 = ~n28067 & n28072 ;
  assign n28074 = n28061 ^ x785 ^ 1'b0 ;
  assign n28075 = ( n28061 & n28073 ) | ( n28061 & n28074 ) | ( n28073 & n28074 ) ;
  assign n28076 = x618 & ~n28075 ;
  assign n28077 = x618 | n28022 ;
  assign n28078 = ( x1154 & n28076 ) | ( x1154 & n28077 ) | ( n28076 & n28077 ) ;
  assign n28079 = ~n28076 & n28078 ;
  assign n28080 = ( x627 & n27992 ) | ( x627 & ~n28079 ) | ( n27992 & ~n28079 ) ;
  assign n28081 = ~n27992 & n28080 ;
  assign n28082 = x627 | n27990 ;
  assign n28083 = x618 & ~n28022 ;
  assign n28084 = x1154 | n28083 ;
  assign n28085 = ( n28075 & n28076 ) | ( n28075 & ~n28084 ) | ( n28076 & ~n28084 ) ;
  assign n28086 = ( ~n28081 & n28082 ) | ( ~n28081 & n28085 ) | ( n28082 & n28085 ) ;
  assign n28087 = ~n28081 & n28086 ;
  assign n28088 = n28075 ^ x781 ^ 1'b0 ;
  assign n28089 = ( n28075 & n28087 ) | ( n28075 & n28088 ) | ( n28087 & n28088 ) ;
  assign n28090 = ~x789 & n28089 ;
  assign n28091 = x619 & ~n28023 ;
  assign n28092 = x1159 | n28091 ;
  assign n28093 = x619 & ~n28089 ;
  assign n28094 = ( n28089 & ~n28092 ) | ( n28089 & n28093 ) | ( ~n28092 & n28093 ) ;
  assign n28095 = ( x648 & n27999 ) | ( x648 & ~n28094 ) | ( n27999 & ~n28094 ) ;
  assign n28096 = n28094 | n28095 ;
  assign n28097 = x619 | n28023 ;
  assign n28098 = x1159 & ~n28093 ;
  assign n28099 = n28097 & n28098 ;
  assign n28100 = ( x648 & n28002 ) | ( x648 & ~n28099 ) | ( n28002 & ~n28099 ) ;
  assign n28101 = ~n28002 & n28100 ;
  assign n28102 = x789 & ~n28101 ;
  assign n28103 = n28096 & n28102 ;
  assign n28104 = ( n16519 & ~n28090 ) | ( n16519 & n28103 ) | ( ~n28090 & n28103 ) ;
  assign n28105 = n28090 | n28104 ;
  assign n28106 = n28105 ^ n28048 ^ 1'b0 ;
  assign n28107 = ( n28048 & n28105 ) | ( n28048 & n28106 ) | ( n28105 & n28106 ) ;
  assign n28108 = ( n18482 & ~n28048 ) | ( n18482 & n28107 ) | ( ~n28048 & n28107 ) ;
  assign n28109 = n19208 | n28025 ;
  assign n28110 = n16556 & ~n28007 ;
  assign n28111 = x629 & ~n28110 ;
  assign n28112 = n28109 & n28111 ;
  assign n28113 = n16557 & ~n28007 ;
  assign n28114 = n19212 & ~n28025 ;
  assign n28115 = n28113 | n28114 ;
  assign n28116 = ( x629 & ~n28112 ) | ( x629 & n28115 ) | ( ~n28112 & n28115 ) ;
  assign n28117 = ~n28112 & n28116 ;
  assign n28118 = ( x792 & ~n19206 ) | ( x792 & n28117 ) | ( ~n19206 & n28117 ) ;
  assign n28119 = ( n18484 & n19206 ) | ( n18484 & n28118 ) | ( n19206 & n28118 ) ;
  assign n28120 = ( n28035 & n28108 ) | ( n28035 & ~n28119 ) | ( n28108 & ~n28119 ) ;
  assign n28121 = n28120 ^ n28108 ^ 1'b0 ;
  assign n28122 = ( n28035 & n28120 ) | ( n28035 & ~n28121 ) | ( n28120 & ~n28121 ) ;
  assign n28123 = x790 | n28122 ;
  assign n28124 = x644 & ~n28122 ;
  assign n28125 = ( x787 & n28028 ) | ( x787 & ~n28031 ) | ( n28028 & ~n28031 ) ;
  assign n28126 = ~n28028 & n28125 ;
  assign n28127 = ( x787 & n28026 ) | ( x787 & ~n28126 ) | ( n28026 & ~n28126 ) ;
  assign n28128 = ~n28126 & n28127 ;
  assign n28129 = x644 | n28128 ;
  assign n28130 = ( x715 & n28124 ) | ( x715 & n28129 ) | ( n28124 & n28129 ) ;
  assign n28131 = ~n28124 & n28130 ;
  assign n28132 = x644 | n27978 ;
  assign n28133 = n27978 ^ n16376 ^ 1'b0 ;
  assign n28134 = ( n27978 & n28009 ) | ( n27978 & ~n28133 ) | ( n28009 & ~n28133 ) ;
  assign n28135 = x644 & ~n28134 ;
  assign n28136 = ( x715 & n28132 ) | ( x715 & ~n28135 ) | ( n28132 & ~n28135 ) ;
  assign n28137 = ~x715 & n28136 ;
  assign n28138 = ( x1160 & n28131 ) | ( x1160 & ~n28137 ) | ( n28131 & ~n28137 ) ;
  assign n28139 = ~n28131 & n28138 ;
  assign n28140 = x644 & ~n27978 ;
  assign n28141 = x715 & ~n28140 ;
  assign n28142 = ( n28134 & n28135 ) | ( n28134 & n28141 ) | ( n28135 & n28141 ) ;
  assign n28143 = x644 & ~n28128 ;
  assign n28144 = x715 | n28143 ;
  assign n28145 = ( n28122 & n28124 ) | ( n28122 & ~n28144 ) | ( n28124 & ~n28144 ) ;
  assign n28146 = ( x1160 & ~n28142 ) | ( x1160 & n28145 ) | ( ~n28142 & n28145 ) ;
  assign n28147 = n28142 | n28146 ;
  assign n28148 = x790 & ~n28147 ;
  assign n28149 = ( x790 & n28139 ) | ( x790 & n28148 ) | ( n28139 & n28148 ) ;
  assign n28150 = x832 & ~n28149 ;
  assign n28151 = n28123 & n28150 ;
  assign n28152 = ~x188 & n7318 ;
  assign n28153 = x832 | n28152 ;
  assign n28154 = ~n28151 & n28153 ;
  assign n28155 = ( n27977 & n28151 ) | ( n27977 & ~n28154 ) | ( n28151 & ~n28154 ) ;
  assign n28156 = x189 & ~n1611 ;
  assign n28157 = x772 & n15591 ;
  assign n28158 = ~n18309 & n28157 ;
  assign n28159 = ~n18321 & n28158 ;
  assign n28160 = ~x626 & n28159 ;
  assign n28161 = n28156 | n28160 ;
  assign n28162 = ( x641 & x1158 ) | ( x641 & ~n28161 ) | ( x1158 & ~n28161 ) ;
  assign n28163 = ( x641 & ~n16317 ) | ( x641 & n28162 ) | ( ~n16317 & n28162 ) ;
  assign n28164 = x727 & n15778 ;
  assign n28165 = n28156 | n28164 ;
  assign n28166 = x1153 & ~n28156 ;
  assign n28167 = x625 & n28164 ;
  assign n28168 = n28166 & ~n28167 ;
  assign n28169 = n28167 ^ n28164 ^ n28156 ;
  assign n28170 = x1153 | n28169 ;
  assign n28171 = ~n28168 & n28170 ;
  assign n28172 = n28165 ^ x778 ^ 1'b0 ;
  assign n28173 = ( n28165 & n28171 ) | ( n28165 & n28172 ) | ( n28171 & n28172 ) ;
  assign n28174 = ~n17087 & n28173 ;
  assign n28175 = ~n16279 & n28174 ;
  assign n28176 = n28156 | n28175 ;
  assign n28177 = ( n16453 & ~n28163 ) | ( n16453 & n28176 ) | ( ~n28163 & n28176 ) ;
  assign n28178 = n28177 ^ n28163 ^ 1'b0 ;
  assign n28179 = ( n28163 & ~n28177 ) | ( n28163 & n28178 ) | ( ~n28177 & n28178 ) ;
  assign n28180 = x626 & n28159 ;
  assign n28181 = n28156 | n28180 ;
  assign n28182 = ( x1158 & ~n16317 ) | ( x1158 & n28181 ) | ( ~n16317 & n28181 ) ;
  assign n28183 = ( x641 & n16317 ) | ( x641 & n28182 ) | ( n16317 & n28182 ) ;
  assign n28184 = n28183 ^ n16454 ^ 1'b0 ;
  assign n28185 = ( ~n16454 & n28176 ) | ( ~n16454 & n28184 ) | ( n28176 & n28184 ) ;
  assign n28186 = ( n16454 & n28183 ) | ( n16454 & n28185 ) | ( n28183 & n28185 ) ;
  assign n28187 = ( x788 & n28179 ) | ( x788 & n28186 ) | ( n28179 & n28186 ) ;
  assign n28188 = ~n28179 & n28187 ;
  assign n28189 = ~n18315 & n28158 ;
  assign n28190 = n18451 & n28189 ;
  assign n28191 = n16276 & ~n28190 ;
  assign n28192 = ~n18374 & n28189 ;
  assign n28193 = ~n28191 & n28192 ;
  assign n28194 = ( n16277 & n28191 ) | ( n16277 & ~n28193 ) | ( n28191 & ~n28193 ) ;
  assign n28195 = n28174 & ~n28194 ;
  assign n28196 = ( n21630 & n28194 ) | ( n21630 & ~n28195 ) | ( n28194 & ~n28195 ) ;
  assign n28197 = n28196 ^ n16519 ^ 1'b0 ;
  assign n28198 = x789 & ~n28156 ;
  assign n28199 = ( n28196 & ~n28197 ) | ( n28196 & n28198 ) | ( ~n28197 & n28198 ) ;
  assign n28200 = ( n16519 & n28197 ) | ( n16519 & n28199 ) | ( n28197 & n28199 ) ;
  assign n28201 = x1154 | n28156 ;
  assign n28202 = ~n18378 & n28158 ;
  assign n28203 = n28201 | n28202 ;
  assign n28204 = ~n16234 & n28173 ;
  assign n28205 = n28156 | n28204 ;
  assign n28206 = ~x618 & n28205 ;
  assign n28207 = x608 | n28168 ;
  assign n28208 = n28156 | n28157 ;
  assign n28209 = x727 & n17156 ;
  assign n28210 = n28208 | n28209 ;
  assign n28211 = x625 & n28209 ;
  assign n28212 = n28210 & ~n28211 ;
  assign n28213 = ( x1153 & ~n28207 ) | ( x1153 & n28212 ) | ( ~n28207 & n28212 ) ;
  assign n28214 = ~n28207 & n28213 ;
  assign n28215 = x1153 & ~n28208 ;
  assign n28216 = ~n28211 & n28215 ;
  assign n28217 = ( x608 & n28170 ) | ( x608 & n28216 ) | ( n28170 & n28216 ) ;
  assign n28218 = ~n28216 & n28217 ;
  assign n28219 = ( x778 & n28214 ) | ( x778 & ~n28218 ) | ( n28214 & ~n28218 ) ;
  assign n28220 = ~n28214 & n28219 ;
  assign n28221 = ( x778 & n28210 ) | ( x778 & ~n28220 ) | ( n28210 & ~n28220 ) ;
  assign n28222 = ~n28220 & n28221 ;
  assign n28223 = ~x609 & n28222 ;
  assign n28224 = x609 & n28173 ;
  assign n28225 = ( x1155 & ~n28223 ) | ( x1155 & n28224 ) | ( ~n28223 & n28224 ) ;
  assign n28226 = n28223 | n28225 ;
  assign n28227 = x1155 | n28156 ;
  assign n28228 = ~n15662 & n28157 ;
  assign n28229 = n28227 | n28228 ;
  assign n28230 = ~x609 & n28173 ;
  assign n28231 = x609 & n28222 ;
  assign n28232 = ( x1155 & n28230 ) | ( x1155 & ~n28231 ) | ( n28230 & ~n28231 ) ;
  assign n28233 = ~n28230 & n28232 ;
  assign n28234 = x660 & ~n28233 ;
  assign n28235 = n28229 & n28234 ;
  assign n28236 = x1155 & ~n28156 ;
  assign n28237 = n15668 & n28157 ;
  assign n28238 = ( x660 & n28236 ) | ( x660 & ~n28237 ) | ( n28236 & ~n28237 ) ;
  assign n28239 = n28238 ^ n28236 ^ 1'b0 ;
  assign n28240 = ( x660 & n28238 ) | ( x660 & ~n28239 ) | ( n28238 & ~n28239 ) ;
  assign n28241 = ~n28235 & n28240 ;
  assign n28242 = ( n28226 & n28235 ) | ( n28226 & ~n28241 ) | ( n28235 & ~n28241 ) ;
  assign n28243 = n28222 ^ x785 ^ 1'b0 ;
  assign n28244 = ( n28222 & n28242 ) | ( n28222 & n28243 ) | ( n28242 & n28243 ) ;
  assign n28245 = x618 & n28244 ;
  assign n28246 = ( x1154 & n28206 ) | ( x1154 & ~n28245 ) | ( n28206 & ~n28245 ) ;
  assign n28247 = ~n28206 & n28246 ;
  assign n28248 = x627 & ~n28247 ;
  assign n28249 = n28203 & n28248 ;
  assign n28250 = ~x618 & n28244 ;
  assign n28251 = x618 & n28205 ;
  assign n28252 = ( x1154 & ~n28250 ) | ( x1154 & n28251 ) | ( ~n28250 & n28251 ) ;
  assign n28253 = n28250 | n28252 ;
  assign n28254 = x1154 & ~n28156 ;
  assign n28255 = n18431 & n28158 ;
  assign n28256 = n28254 & ~n28255 ;
  assign n28257 = ( x627 & n28253 ) | ( x627 & ~n28256 ) | ( n28253 & ~n28256 ) ;
  assign n28258 = ~x627 & n28257 ;
  assign n28259 = ( x781 & n28249 ) | ( x781 & n28258 ) | ( n28249 & n28258 ) ;
  assign n28260 = n28258 ^ n28249 ^ 1'b0 ;
  assign n28261 = ( x781 & n28259 ) | ( x781 & n28260 ) | ( n28259 & n28260 ) ;
  assign n28262 = ~x781 & n28244 ;
  assign n28263 = n21705 | n28262 ;
  assign n28264 = ( ~n28200 & n28261 ) | ( ~n28200 & n28263 ) | ( n28261 & n28263 ) ;
  assign n28265 = ~n28200 & n28264 ;
  assign n28266 = ( n18482 & ~n28188 ) | ( n18482 & n28265 ) | ( ~n28188 & n28265 ) ;
  assign n28267 = n28188 | n28266 ;
  assign n28268 = ~n17088 & n28173 ;
  assign n28269 = x628 & n28268 ;
  assign n28270 = ~n16518 & n28159 ;
  assign n28271 = x628 | n28270 ;
  assign n28272 = x629 & n28271 ;
  assign n28273 = ( x1156 & n28269 ) | ( x1156 & ~n28272 ) | ( n28269 & ~n28272 ) ;
  assign n28274 = ~n28269 & n28273 ;
  assign n28275 = x629 & ~n28268 ;
  assign n28276 = ~x629 & n28270 ;
  assign n28277 = ~n28275 & n28276 ;
  assign n28278 = ( x628 & n28275 ) | ( x628 & ~n28277 ) | ( n28275 & ~n28277 ) ;
  assign n28279 = ( ~x1156 & n28274 ) | ( ~x1156 & n28278 ) | ( n28274 & n28278 ) ;
  assign n28280 = n28274 ^ x1156 ^ 1'b0 ;
  assign n28281 = ( n28274 & n28279 ) | ( n28274 & ~n28280 ) | ( n28279 & ~n28280 ) ;
  assign n28282 = x792 & ~n28156 ;
  assign n28283 = n28281 & n28282 ;
  assign n28284 = ( n18484 & n28267 ) | ( n18484 & ~n28283 ) | ( n28267 & ~n28283 ) ;
  assign n28285 = n28284 ^ n28267 ^ 1'b0 ;
  assign n28286 = ( n18484 & n28284 ) | ( n18484 & ~n28285 ) | ( n28284 & ~n28285 ) ;
  assign n28289 = ~n17093 & n28268 ;
  assign n28290 = x630 & ~n28289 ;
  assign n28291 = ( x647 & n28289 ) | ( x647 & n28290 ) | ( n28289 & n28290 ) ;
  assign n28287 = ~n16339 & n28270 ;
  assign n28288 = x630 & n28287 ;
  assign n28292 = ( x1157 & ~n28288 ) | ( x1157 & n28291 ) | ( ~n28288 & n28291 ) ;
  assign n28293 = ~n28291 & n28292 ;
  assign n28294 = ~x630 & n28287 ;
  assign n28295 = ~n28290 & n28294 ;
  assign n28296 = ( x647 & n28290 ) | ( x647 & ~n28295 ) | ( n28290 & ~n28295 ) ;
  assign n28297 = ( ~x1157 & n28293 ) | ( ~x1157 & n28296 ) | ( n28293 & n28296 ) ;
  assign n28298 = n28293 ^ x1157 ^ 1'b0 ;
  assign n28299 = ( n28293 & n28297 ) | ( n28293 & ~n28298 ) | ( n28297 & ~n28298 ) ;
  assign n28300 = x787 & ~n28156 ;
  assign n28301 = n28286 & ~n28300 ;
  assign n28302 = ( n28286 & ~n28299 ) | ( n28286 & n28301 ) | ( ~n28299 & n28301 ) ;
  assign n28303 = ~x790 & n28302 ;
  assign n28304 = ~x644 & n28302 ;
  assign n28305 = ~n17273 & n28289 ;
  assign n28306 = n28156 | n28305 ;
  assign n28307 = x644 & n28306 ;
  assign n28308 = ( x715 & ~n28304 ) | ( x715 & n28307 ) | ( ~n28304 & n28307 ) ;
  assign n28309 = n28304 | n28308 ;
  assign n28310 = x715 & ~n28156 ;
  assign n28311 = n16518 | n21755 ;
  assign n28312 = n28159 & ~n28311 ;
  assign n28313 = ~x644 & n28312 ;
  assign n28314 = n28310 & ~n28313 ;
  assign n28315 = ( x1160 & n28309 ) | ( x1160 & ~n28314 ) | ( n28309 & ~n28314 ) ;
  assign n28316 = ~x1160 & n28315 ;
  assign n28317 = x715 | n28156 ;
  assign n28318 = x644 & n28312 ;
  assign n28319 = n28317 | n28318 ;
  assign n28320 = ~x644 & n28306 ;
  assign n28321 = x644 & n28302 ;
  assign n28322 = ( x715 & n28320 ) | ( x715 & ~n28321 ) | ( n28320 & ~n28321 ) ;
  assign n28323 = ~n28320 & n28322 ;
  assign n28324 = x1160 & ~n28323 ;
  assign n28325 = n28319 & n28324 ;
  assign n28326 = ( x790 & n28316 ) | ( x790 & n28325 ) | ( n28316 & n28325 ) ;
  assign n28327 = n28325 ^ n28316 ^ 1'b0 ;
  assign n28328 = ( x790 & n28326 ) | ( x790 & n28327 ) | ( n28326 & n28327 ) ;
  assign n28329 = ( x832 & n28303 ) | ( x832 & ~n28328 ) | ( n28303 & ~n28328 ) ;
  assign n28330 = ~n28303 & n28329 ;
  assign n28331 = ~x189 & n5193 ;
  assign n28332 = x189 & ~n15656 ;
  assign n28377 = ~x626 & n28332 ;
  assign n28378 = n28332 ^ n15659 ^ 1'b0 ;
  assign n28379 = x189 & n2069 ;
  assign n28338 = x189 | n15644 ;
  assign n28380 = x772 & n15524 ;
  assign n28381 = n15644 & ~n28380 ;
  assign n28382 = x38 & ~n28381 ;
  assign n28383 = n28338 & n28382 ;
  assign n28384 = ~x189 & x772 ;
  assign n28385 = n15640 & n28384 ;
  assign n28386 = x772 & ~n15585 ;
  assign n28387 = x39 & ~n20604 ;
  assign n28388 = ( x39 & n28386 ) | ( x39 & n28387 ) | ( n28386 & n28387 ) ;
  assign n28389 = x772 & n15509 ;
  assign n28390 = ~x772 & n15332 ;
  assign n28391 = x39 | n28390 ;
  assign n28392 = ( ~n28388 & n28389 ) | ( ~n28388 & n28391 ) | ( n28389 & n28391 ) ;
  assign n28393 = ~n28388 & n28392 ;
  assign n28394 = ~n28385 & n28393 ;
  assign n28395 = ( x189 & n28385 ) | ( x189 & ~n28394 ) | ( n28385 & ~n28394 ) ;
  assign n28396 = ( ~x38 & n28383 ) | ( ~x38 & n28395 ) | ( n28383 & n28395 ) ;
  assign n28397 = n28383 ^ x38 ^ 1'b0 ;
  assign n28398 = ( n28383 & n28396 ) | ( n28383 & ~n28397 ) | ( n28396 & ~n28397 ) ;
  assign n28399 = ~n2069 & n28398 ;
  assign n28400 = n28379 | n28399 ;
  assign n28401 = ( n28332 & ~n28378 ) | ( n28332 & n28400 ) | ( ~n28378 & n28400 ) ;
  assign n28402 = x609 & ~n28401 ;
  assign n28403 = x609 | n28332 ;
  assign n28404 = ( x1155 & n28402 ) | ( x1155 & n28403 ) | ( n28402 & n28403 ) ;
  assign n28405 = ~n28402 & n28404 ;
  assign n28406 = x609 & ~n28332 ;
  assign n28407 = x1155 | n28406 ;
  assign n28408 = ( n28401 & n28402 ) | ( n28401 & ~n28407 ) | ( n28402 & ~n28407 ) ;
  assign n28409 = n28405 | n28408 ;
  assign n28410 = n28401 ^ x785 ^ 1'b0 ;
  assign n28411 = ( n28401 & n28409 ) | ( n28401 & n28410 ) | ( n28409 & n28410 ) ;
  assign n28412 = x618 & ~n28411 ;
  assign n28413 = x618 | n28332 ;
  assign n28414 = ( x1154 & n28412 ) | ( x1154 & n28413 ) | ( n28412 & n28413 ) ;
  assign n28415 = ~n28412 & n28414 ;
  assign n28416 = x618 & ~n28332 ;
  assign n28417 = x1154 | n28416 ;
  assign n28418 = ( n28411 & n28412 ) | ( n28411 & ~n28417 ) | ( n28412 & ~n28417 ) ;
  assign n28419 = n28415 | n28418 ;
  assign n28420 = n28411 ^ x781 ^ 1'b0 ;
  assign n28421 = ( n28411 & n28419 ) | ( n28411 & n28420 ) | ( n28419 & n28420 ) ;
  assign n28422 = x619 & ~n28421 ;
  assign n28423 = x619 | n28332 ;
  assign n28424 = ( x1159 & n28422 ) | ( x1159 & n28423 ) | ( n28422 & n28423 ) ;
  assign n28425 = ~n28422 & n28424 ;
  assign n28426 = x619 & ~n28332 ;
  assign n28427 = x1159 | n28426 ;
  assign n28428 = ( n28421 & n28422 ) | ( n28421 & ~n28427 ) | ( n28422 & ~n28427 ) ;
  assign n28429 = n28425 | n28428 ;
  assign n28430 = n28421 ^ x789 ^ 1'b0 ;
  assign n28431 = ( n28421 & n28429 ) | ( n28421 & n28430 ) | ( n28429 & n28430 ) ;
  assign n28432 = x626 & n28431 ;
  assign n28433 = ( x641 & ~n28377 ) | ( x641 & n28432 ) | ( ~n28377 & n28432 ) ;
  assign n28434 = n28377 | n28433 ;
  assign n28333 = x189 | n16699 ;
  assign n28334 = x189 & n16697 ;
  assign n28335 = ( x38 & n28333 ) | ( x38 & ~n28334 ) | ( n28333 & ~n28334 ) ;
  assign n28336 = ~x38 & n28335 ;
  assign n28337 = x727 & ~n2069 ;
  assign n28339 = n18524 & n28338 ;
  assign n28340 = ( n28336 & n28337 ) | ( n28336 & ~n28339 ) | ( n28337 & ~n28339 ) ;
  assign n28341 = ~n28336 & n28340 ;
  assign n28342 = ( n28332 & n28337 ) | ( n28332 & ~n28341 ) | ( n28337 & ~n28341 ) ;
  assign n28343 = ~n28341 & n28342 ;
  assign n28344 = x625 & ~n28343 ;
  assign n28345 = x625 | n28332 ;
  assign n28346 = ( x1153 & n28344 ) | ( x1153 & n28345 ) | ( n28344 & n28345 ) ;
  assign n28347 = ~n28344 & n28346 ;
  assign n28348 = x625 & ~n28332 ;
  assign n28349 = x1153 | n28348 ;
  assign n28350 = ( x625 & n28343 ) | ( x625 & ~n28349 ) | ( n28343 & ~n28349 ) ;
  assign n28351 = ~n28349 & n28350 ;
  assign n28352 = n28347 | n28351 ;
  assign n28353 = n28343 ^ x778 ^ 1'b0 ;
  assign n28354 = ( n28343 & n28352 ) | ( n28343 & n28353 ) | ( n28352 & n28353 ) ;
  assign n28355 = n28332 ^ n16234 ^ 1'b0 ;
  assign n28356 = ( n28332 & n28354 ) | ( n28332 & ~n28355 ) | ( n28354 & ~n28355 ) ;
  assign n28357 = n28332 ^ n16254 ^ 1'b0 ;
  assign n28358 = ( n28332 & n28356 ) | ( n28332 & ~n28357 ) | ( n28356 & ~n28357 ) ;
  assign n28359 = n28332 ^ n16279 ^ 1'b0 ;
  assign n28360 = ( n28332 & n28358 ) | ( n28332 & ~n28359 ) | ( n28358 & ~n28359 ) ;
  assign n28435 = ~x626 & n28360 ;
  assign n28436 = x189 & n16048 ;
  assign n28437 = x189 | n16054 ;
  assign n28438 = ( x772 & n28436 ) | ( x772 & n28437 ) | ( n28436 & n28437 ) ;
  assign n28439 = ~n28436 & n28438 ;
  assign n28440 = x189 | n16029 ;
  assign n28441 = x189 & n16044 ;
  assign n28442 = ( x772 & n28440 ) | ( x772 & ~n28441 ) | ( n28440 & ~n28441 ) ;
  assign n28443 = ~x772 & n28442 ;
  assign n28444 = ( x39 & ~n28439 ) | ( x39 & n28443 ) | ( ~n28439 & n28443 ) ;
  assign n28445 = n28439 | n28444 ;
  assign n28446 = x189 | n15795 ;
  assign n28447 = x189 & n15876 ;
  assign n28448 = ( x772 & n28446 ) | ( x772 & ~n28447 ) | ( n28446 & ~n28447 ) ;
  assign n28449 = ~x772 & n28448 ;
  assign n28450 = x189 & n16003 ;
  assign n28451 = x189 | n15943 ;
  assign n28452 = ( x772 & n28450 ) | ( x772 & n28451 ) | ( n28450 & n28451 ) ;
  assign n28453 = ~n28450 & n28452 ;
  assign n28454 = ( x39 & n28449 ) | ( x39 & ~n28453 ) | ( n28449 & ~n28453 ) ;
  assign n28455 = ~n28449 & n28454 ;
  assign n28456 = ( x38 & n28445 ) | ( x38 & ~n28455 ) | ( n28445 & ~n28455 ) ;
  assign n28457 = ~x38 & n28456 ;
  assign n28458 = x727 & ~n17882 ;
  assign n28459 = ( n28383 & ~n28457 ) | ( n28383 & n28458 ) | ( ~n28457 & n28458 ) ;
  assign n28460 = ~n28383 & n28459 ;
  assign n28461 = ( n2051 & n2068 ) | ( n2051 & ~n28460 ) | ( n2068 & ~n28460 ) ;
  assign n28462 = n28460 | n28461 ;
  assign n28463 = ( x727 & n28398 ) | ( x727 & ~n28462 ) | ( n28398 & ~n28462 ) ;
  assign n28464 = ~n28462 & n28463 ;
  assign n28465 = n28464 ^ x189 ^ 1'b0 ;
  assign n28466 = ( ~x189 & n2069 ) | ( ~x189 & n28465 ) | ( n2069 & n28465 ) ;
  assign n28467 = ( x189 & n28464 ) | ( x189 & n28466 ) | ( n28464 & n28466 ) ;
  assign n28468 = x625 & ~n28467 ;
  assign n28474 = x625 | n28400 ;
  assign n28475 = ( x1153 & n28468 ) | ( x1153 & n28474 ) | ( n28468 & n28474 ) ;
  assign n28476 = ~n28468 & n28475 ;
  assign n28477 = ( x608 & ~n28351 ) | ( x608 & n28476 ) | ( ~n28351 & n28476 ) ;
  assign n28478 = ~n28476 & n28477 ;
  assign n28469 = x625 & ~n28400 ;
  assign n28470 = x1153 | n28469 ;
  assign n28471 = ( n28467 & n28468 ) | ( n28467 & ~n28470 ) | ( n28468 & ~n28470 ) ;
  assign n28472 = ( x608 & ~n28347 ) | ( x608 & n28471 ) | ( ~n28347 & n28471 ) ;
  assign n28473 = n28347 | n28472 ;
  assign n28479 = n28478 ^ n28473 ^ 1'b0 ;
  assign n28480 = ( x778 & ~n28473 ) | ( x778 & n28478 ) | ( ~n28473 & n28478 ) ;
  assign n28481 = ( x778 & ~n28479 ) | ( x778 & n28480 ) | ( ~n28479 & n28480 ) ;
  assign n28482 = ( x778 & n28467 ) | ( x778 & ~n28481 ) | ( n28467 & ~n28481 ) ;
  assign n28483 = ~n28481 & n28482 ;
  assign n28484 = x609 & ~n28483 ;
  assign n28490 = x609 | n28354 ;
  assign n28491 = ( x1155 & n28484 ) | ( x1155 & n28490 ) | ( n28484 & n28490 ) ;
  assign n28492 = ~n28484 & n28491 ;
  assign n28493 = ( x660 & ~n28408 ) | ( x660 & n28492 ) | ( ~n28408 & n28492 ) ;
  assign n28494 = ~n28492 & n28493 ;
  assign n28485 = x609 & ~n28354 ;
  assign n28486 = x1155 | n28485 ;
  assign n28487 = ( n28483 & n28484 ) | ( n28483 & ~n28486 ) | ( n28484 & ~n28486 ) ;
  assign n28488 = ( x660 & ~n28405 ) | ( x660 & n28487 ) | ( ~n28405 & n28487 ) ;
  assign n28489 = n28405 | n28488 ;
  assign n28495 = n28494 ^ n28489 ^ 1'b0 ;
  assign n28496 = ( x785 & ~n28489 ) | ( x785 & n28494 ) | ( ~n28489 & n28494 ) ;
  assign n28497 = ( x785 & ~n28495 ) | ( x785 & n28496 ) | ( ~n28495 & n28496 ) ;
  assign n28498 = ( x785 & n28483 ) | ( x785 & ~n28497 ) | ( n28483 & ~n28497 ) ;
  assign n28499 = ~n28497 & n28498 ;
  assign n28500 = x618 & ~n28499 ;
  assign n28506 = x618 | n28356 ;
  assign n28507 = ( x1154 & n28500 ) | ( x1154 & n28506 ) | ( n28500 & n28506 ) ;
  assign n28508 = ~n28500 & n28507 ;
  assign n28509 = ( x627 & ~n28418 ) | ( x627 & n28508 ) | ( ~n28418 & n28508 ) ;
  assign n28510 = ~n28508 & n28509 ;
  assign n28501 = x618 & ~n28356 ;
  assign n28502 = x1154 | n28501 ;
  assign n28503 = ( n28499 & n28500 ) | ( n28499 & ~n28502 ) | ( n28500 & ~n28502 ) ;
  assign n28504 = ( x627 & ~n28415 ) | ( x627 & n28503 ) | ( ~n28415 & n28503 ) ;
  assign n28505 = n28415 | n28504 ;
  assign n28511 = n28510 ^ n28505 ^ 1'b0 ;
  assign n28512 = ( x781 & ~n28505 ) | ( x781 & n28510 ) | ( ~n28505 & n28510 ) ;
  assign n28513 = ( x781 & ~n28511 ) | ( x781 & n28512 ) | ( ~n28511 & n28512 ) ;
  assign n28514 = ( x781 & n28499 ) | ( x781 & ~n28513 ) | ( n28499 & ~n28513 ) ;
  assign n28515 = ~n28513 & n28514 ;
  assign n28516 = x619 & ~n28515 ;
  assign n28522 = x619 | n28358 ;
  assign n28523 = ( x1159 & n28516 ) | ( x1159 & n28522 ) | ( n28516 & n28522 ) ;
  assign n28524 = ~n28516 & n28523 ;
  assign n28525 = ( x648 & ~n28428 ) | ( x648 & n28524 ) | ( ~n28428 & n28524 ) ;
  assign n28526 = ~n28524 & n28525 ;
  assign n28517 = x619 & ~n28358 ;
  assign n28518 = x1159 | n28517 ;
  assign n28519 = ( n28515 & n28516 ) | ( n28515 & ~n28518 ) | ( n28516 & ~n28518 ) ;
  assign n28520 = ( x648 & ~n28425 ) | ( x648 & n28519 ) | ( ~n28425 & n28519 ) ;
  assign n28521 = n28425 | n28520 ;
  assign n28527 = n28526 ^ n28521 ^ 1'b0 ;
  assign n28528 = ( x789 & ~n28521 ) | ( x789 & n28526 ) | ( ~n28521 & n28526 ) ;
  assign n28529 = ( x789 & ~n28527 ) | ( x789 & n28528 ) | ( ~n28527 & n28528 ) ;
  assign n28530 = ( x789 & n28515 ) | ( x789 & ~n28529 ) | ( n28515 & ~n28529 ) ;
  assign n28531 = ~n28529 & n28530 ;
  assign n28532 = x626 & n28531 ;
  assign n28533 = ( x641 & n28435 ) | ( x641 & ~n28532 ) | ( n28435 & ~n28532 ) ;
  assign n28534 = ~n28435 & n28533 ;
  assign n28535 = x1158 & ~n28534 ;
  assign n28536 = n28434 & n28535 ;
  assign n28537 = ~x626 & n28531 ;
  assign n28538 = x626 & n28360 ;
  assign n28539 = ( x641 & ~n28537 ) | ( x641 & n28538 ) | ( ~n28537 & n28538 ) ;
  assign n28540 = n28537 | n28539 ;
  assign n28541 = ~x626 & n28431 ;
  assign n28542 = x626 & n28332 ;
  assign n28543 = ( x641 & n28541 ) | ( x641 & ~n28542 ) | ( n28541 & ~n28542 ) ;
  assign n28544 = ~n28541 & n28543 ;
  assign n28545 = ( x1158 & n28540 ) | ( x1158 & ~n28544 ) | ( n28540 & ~n28544 ) ;
  assign n28546 = ~x1158 & n28545 ;
  assign n28547 = ( x788 & n28536 ) | ( x788 & ~n28546 ) | ( n28536 & ~n28546 ) ;
  assign n28548 = ~n28536 & n28547 ;
  assign n28549 = ( x788 & n28531 ) | ( x788 & ~n28548 ) | ( n28531 & ~n28548 ) ;
  assign n28550 = ~n28548 & n28549 ;
  assign n28551 = x628 & ~n28550 ;
  assign n28552 = n28332 ^ n16518 ^ 1'b0 ;
  assign n28553 = ( n28332 & n28431 ) | ( n28332 & ~n28552 ) | ( n28431 & ~n28552 ) ;
  assign n28559 = x628 | n28553 ;
  assign n28560 = ( x1156 & n28551 ) | ( x1156 & n28559 ) | ( n28551 & n28559 ) ;
  assign n28561 = ~n28551 & n28560 ;
  assign n28361 = n28332 ^ n16318 ^ 1'b0 ;
  assign n28362 = ( n28332 & n28360 ) | ( n28332 & ~n28361 ) | ( n28360 & ~n28361 ) ;
  assign n28363 = x628 & ~n28362 ;
  assign n28367 = x628 & ~n28332 ;
  assign n28368 = x1156 | n28367 ;
  assign n28369 = ( n28362 & n28363 ) | ( n28362 & ~n28368 ) | ( n28363 & ~n28368 ) ;
  assign n28562 = ( x629 & ~n28369 ) | ( x629 & n28561 ) | ( ~n28369 & n28561 ) ;
  assign n28563 = ~n28561 & n28562 ;
  assign n28364 = x628 | n28332 ;
  assign n28365 = ( x1156 & n28363 ) | ( x1156 & n28364 ) | ( n28363 & n28364 ) ;
  assign n28366 = ~n28363 & n28365 ;
  assign n28554 = x628 & ~n28553 ;
  assign n28555 = x1156 | n28554 ;
  assign n28556 = ( n28550 & n28551 ) | ( n28550 & ~n28555 ) | ( n28551 & ~n28555 ) ;
  assign n28557 = ( x629 & ~n28366 ) | ( x629 & n28556 ) | ( ~n28366 & n28556 ) ;
  assign n28558 = n28366 | n28557 ;
  assign n28564 = n28563 ^ n28558 ^ 1'b0 ;
  assign n28565 = ( x792 & ~n28558 ) | ( x792 & n28563 ) | ( ~n28558 & n28563 ) ;
  assign n28566 = ( x792 & ~n28564 ) | ( x792 & n28565 ) | ( ~n28564 & n28565 ) ;
  assign n28567 = ( x792 & n28550 ) | ( x792 & ~n28566 ) | ( n28550 & ~n28566 ) ;
  assign n28568 = ~n28566 & n28567 ;
  assign n28569 = x647 & ~n28568 ;
  assign n28570 = n28332 ^ n16339 ^ 1'b0 ;
  assign n28571 = ( n28332 & n28553 ) | ( n28332 & ~n28570 ) | ( n28553 & ~n28570 ) ;
  assign n28577 = x647 | n28571 ;
  assign n28578 = ( x1157 & n28569 ) | ( x1157 & n28577 ) | ( n28569 & n28577 ) ;
  assign n28579 = ~n28569 & n28578 ;
  assign n28370 = n28366 | n28369 ;
  assign n28371 = n28362 ^ x792 ^ 1'b0 ;
  assign n28372 = ( n28362 & n28370 ) | ( n28362 & n28371 ) | ( n28370 & n28371 ) ;
  assign n28373 = x647 & ~n28372 ;
  assign n28580 = x647 & ~n28332 ;
  assign n28581 = x1157 | n28580 ;
  assign n28582 = ( n28372 & n28373 ) | ( n28372 & ~n28581 ) | ( n28373 & ~n28581 ) ;
  assign n28583 = ( x630 & n28579 ) | ( x630 & ~n28582 ) | ( n28579 & ~n28582 ) ;
  assign n28584 = ~n28579 & n28583 ;
  assign n28374 = x647 | n28332 ;
  assign n28375 = ( x1157 & n28373 ) | ( x1157 & n28374 ) | ( n28373 & n28374 ) ;
  assign n28376 = ~n28373 & n28375 ;
  assign n28572 = x647 & ~n28571 ;
  assign n28573 = x1157 | n28572 ;
  assign n28574 = ( n28568 & n28569 ) | ( n28568 & ~n28573 ) | ( n28569 & ~n28573 ) ;
  assign n28575 = ( x630 & ~n28376 ) | ( x630 & n28574 ) | ( ~n28376 & n28574 ) ;
  assign n28576 = n28376 | n28575 ;
  assign n28585 = n28584 ^ n28576 ^ 1'b0 ;
  assign n28586 = ( x787 & ~n28576 ) | ( x787 & n28584 ) | ( ~n28576 & n28584 ) ;
  assign n28587 = ( x787 & ~n28585 ) | ( x787 & n28586 ) | ( ~n28585 & n28586 ) ;
  assign n28588 = ( x787 & n28568 ) | ( x787 & ~n28587 ) | ( n28568 & ~n28587 ) ;
  assign n28589 = ~n28587 & n28588 ;
  assign n28590 = ~x790 & n28589 ;
  assign n28598 = x644 & ~n28332 ;
  assign n28599 = x715 & ~n28598 ;
  assign n28600 = n28332 ^ n16376 ^ 1'b0 ;
  assign n28601 = ( n28332 & n28571 ) | ( n28332 & ~n28600 ) | ( n28571 & ~n28600 ) ;
  assign n28602 = x644 & ~n28601 ;
  assign n28603 = ( n28599 & n28601 ) | ( n28599 & n28602 ) | ( n28601 & n28602 ) ;
  assign n28591 = x644 | n28589 ;
  assign n28592 = n28376 | n28582 ;
  assign n28593 = n28372 ^ x787 ^ 1'b0 ;
  assign n28594 = ( n28372 & n28592 ) | ( n28372 & n28593 ) | ( n28592 & n28593 ) ;
  assign n28595 = x644 & ~n28594 ;
  assign n28596 = ( x715 & n28591 ) | ( x715 & ~n28595 ) | ( n28591 & ~n28595 ) ;
  assign n28597 = ~x715 & n28596 ;
  assign n28604 = ( x1160 & n28597 ) | ( x1160 & ~n28603 ) | ( n28597 & ~n28603 ) ;
  assign n28605 = n28603 | n28604 ;
  assign n28606 = x644 & ~n28589 ;
  assign n28607 = x644 | n28594 ;
  assign n28608 = ( x715 & n28606 ) | ( x715 & n28607 ) | ( n28606 & n28607 ) ;
  assign n28609 = ~n28606 & n28608 ;
  assign n28610 = x644 | n28332 ;
  assign n28611 = ( x715 & ~n28602 ) | ( x715 & n28610 ) | ( ~n28602 & n28610 ) ;
  assign n28612 = ~x715 & n28611 ;
  assign n28613 = ( x1160 & n28609 ) | ( x1160 & ~n28612 ) | ( n28609 & ~n28612 ) ;
  assign n28614 = ~n28609 & n28613 ;
  assign n28615 = x790 & ~n28614 ;
  assign n28616 = n28605 & n28615 ;
  assign n28617 = ( n5193 & ~n28590 ) | ( n5193 & n28616 ) | ( ~n28590 & n28616 ) ;
  assign n28618 = n28590 | n28617 ;
  assign n28619 = ( x57 & ~n28331 ) | ( x57 & n28618 ) | ( ~n28331 & n28618 ) ;
  assign n28620 = ~x57 & n28619 ;
  assign n28621 = x57 & x189 ;
  assign n28622 = x832 | n28621 ;
  assign n28623 = ( ~n28330 & n28620 ) | ( ~n28330 & n28622 ) | ( n28620 & n28622 ) ;
  assign n28624 = ~n28330 & n28623 ;
  assign n28625 = x190 | n15656 ;
  assign n28626 = x190 | n15644 ;
  assign n28627 = n16185 & n28626 ;
  assign n28628 = x190 | n16697 ;
  assign n28629 = x190 & n16699 ;
  assign n28630 = ( x38 & n28628 ) | ( x38 & ~n28629 ) | ( n28628 & ~n28629 ) ;
  assign n28631 = ~x38 & n28630 ;
  assign n28632 = ( x699 & n28627 ) | ( x699 & ~n28631 ) | ( n28627 & ~n28631 ) ;
  assign n28633 = ~n28627 & n28632 ;
  assign n28634 = x190 | x699 ;
  assign n28635 = n15655 | n28634 ;
  assign n28636 = ( n2069 & ~n28633 ) | ( n2069 & n28635 ) | ( ~n28633 & n28635 ) ;
  assign n28637 = ~n2069 & n28636 ;
  assign n28638 = n28637 ^ x190 ^ 1'b0 ;
  assign n28639 = ( ~x190 & n2069 ) | ( ~x190 & n28638 ) | ( n2069 & n28638 ) ;
  assign n28640 = ( x190 & n28637 ) | ( x190 & n28639 ) | ( n28637 & n28639 ) ;
  assign n28641 = x625 & ~n28640 ;
  assign n28642 = x625 | n28625 ;
  assign n28643 = ( x1153 & n28641 ) | ( x1153 & n28642 ) | ( n28641 & n28642 ) ;
  assign n28644 = ~n28641 & n28643 ;
  assign n28645 = x625 & ~n28625 ;
  assign n28646 = x1153 | n28645 ;
  assign n28647 = ( x625 & n28640 ) | ( x625 & ~n28646 ) | ( n28640 & ~n28646 ) ;
  assign n28648 = ~n28646 & n28647 ;
  assign n28649 = n28644 | n28648 ;
  assign n28650 = n28640 ^ x778 ^ 1'b0 ;
  assign n28651 = ( n28640 & n28649 ) | ( n28640 & n28650 ) | ( n28649 & n28650 ) ;
  assign n28652 = n28625 ^ n16234 ^ 1'b0 ;
  assign n28653 = ( n28625 & n28651 ) | ( n28625 & ~n28652 ) | ( n28651 & ~n28652 ) ;
  assign n28654 = n28625 ^ n16254 ^ 1'b0 ;
  assign n28655 = ( n28625 & n28653 ) | ( n28625 & ~n28654 ) | ( n28653 & ~n28654 ) ;
  assign n28656 = n28625 ^ n16279 ^ 1'b0 ;
  assign n28657 = ( n28625 & n28655 ) | ( n28625 & ~n28656 ) | ( n28655 & ~n28656 ) ;
  assign n28658 = n28625 ^ n16318 ^ 1'b0 ;
  assign n28659 = ( n28625 & n28657 ) | ( n28625 & ~n28658 ) | ( n28657 & ~n28658 ) ;
  assign n28660 = n28625 ^ x628 ^ 1'b0 ;
  assign n28661 = ( n28625 & n28659 ) | ( n28625 & ~n28660 ) | ( n28659 & ~n28660 ) ;
  assign n28662 = ( n28625 & n28659 ) | ( n28625 & n28660 ) | ( n28659 & n28660 ) ;
  assign n28663 = n28661 ^ x1156 ^ 1'b0 ;
  assign n28664 = ( n28661 & n28662 ) | ( n28661 & n28663 ) | ( n28662 & n28663 ) ;
  assign n28665 = n28659 ^ x792 ^ 1'b0 ;
  assign n28666 = ( n28659 & n28664 ) | ( n28659 & n28665 ) | ( n28664 & n28665 ) ;
  assign n28667 = n28625 ^ x647 ^ 1'b0 ;
  assign n28668 = ( n28625 & n28666 ) | ( n28625 & ~n28667 ) | ( n28666 & ~n28667 ) ;
  assign n28669 = ( n28625 & n28666 ) | ( n28625 & n28667 ) | ( n28666 & n28667 ) ;
  assign n28670 = n28668 ^ x1157 ^ 1'b0 ;
  assign n28671 = ( n28668 & n28669 ) | ( n28668 & n28670 ) | ( n28669 & n28670 ) ;
  assign n28672 = n28666 ^ x787 ^ 1'b0 ;
  assign n28673 = ( n28666 & n28671 ) | ( n28666 & n28672 ) | ( n28671 & n28672 ) ;
  assign n28674 = x644 & ~n28673 ;
  assign n28675 = x715 | n28674 ;
  assign n28676 = x644 & ~n28625 ;
  assign n28677 = x715 & ~n28676 ;
  assign n28678 = n28677 ^ x1160 ^ 1'b0 ;
  assign n28679 = x190 & n2069 ;
  assign n28680 = x38 & n28626 ;
  assign n28681 = ~x190 & x763 ;
  assign n28682 = n15587 & n28681 ;
  assign n28683 = x763 & n15639 ;
  assign n28684 = x190 & ~n28683 ;
  assign n28685 = ( n20789 & ~n28682 ) | ( n20789 & n28684 ) | ( ~n28682 & n28684 ) ;
  assign n28686 = n28682 | n28685 ;
  assign n28687 = x190 & ~n15631 ;
  assign n28688 = ~x763 & n15486 ;
  assign n28689 = ( x39 & n28687 ) | ( x39 & n28688 ) | ( n28687 & n28688 ) ;
  assign n28690 = n28688 ^ n28687 ^ 1'b0 ;
  assign n28691 = ( x39 & n28689 ) | ( x39 & n28690 ) | ( n28689 & n28690 ) ;
  assign n28692 = ( ~x38 & n28686 ) | ( ~x38 & n28691 ) | ( n28686 & n28691 ) ;
  assign n28693 = ~x38 & n28692 ;
  assign n28694 = x763 & n15646 ;
  assign n28695 = ~n28693 & n28694 ;
  assign n28696 = ( n28680 & n28693 ) | ( n28680 & ~n28695 ) | ( n28693 & ~n28695 ) ;
  assign n28697 = ~n2069 & n28696 ;
  assign n28698 = n28679 | n28697 ;
  assign n28699 = n28625 ^ n15659 ^ 1'b0 ;
  assign n28700 = ( n28625 & n28698 ) | ( n28625 & ~n28699 ) | ( n28698 & ~n28699 ) ;
  assign n28701 = n15662 & n28625 ;
  assign n28702 = ( ~n15662 & n28679 ) | ( ~n15662 & n28697 ) | ( n28679 & n28697 ) ;
  assign n28703 = n28701 | n28702 ;
  assign n28704 = n28703 ^ n28700 ^ n28625 ;
  assign n28705 = n28704 ^ x1155 ^ 1'b0 ;
  assign n28706 = ( n28703 & n28704 ) | ( n28703 & ~n28705 ) | ( n28704 & ~n28705 ) ;
  assign n28707 = n28700 ^ x785 ^ 1'b0 ;
  assign n28708 = ( n28700 & n28706 ) | ( n28700 & n28707 ) | ( n28706 & n28707 ) ;
  assign n28709 = x618 & ~n28708 ;
  assign n28710 = x618 | n28625 ;
  assign n28711 = ( x1154 & n28709 ) | ( x1154 & n28710 ) | ( n28709 & n28710 ) ;
  assign n28712 = ~n28709 & n28711 ;
  assign n28713 = x618 & ~n28625 ;
  assign n28714 = x1154 | n28713 ;
  assign n28715 = ( n28708 & n28709 ) | ( n28708 & ~n28714 ) | ( n28709 & ~n28714 ) ;
  assign n28716 = n28712 | n28715 ;
  assign n28717 = n28708 ^ x781 ^ 1'b0 ;
  assign n28718 = ( n28708 & n28716 ) | ( n28708 & n28717 ) | ( n28716 & n28717 ) ;
  assign n28719 = x619 | n28625 ;
  assign n28720 = x619 & ~n28718 ;
  assign n28721 = x1159 & ~n28720 ;
  assign n28722 = n28719 & n28721 ;
  assign n28723 = x619 & ~n28625 ;
  assign n28724 = x1159 | n28723 ;
  assign n28725 = ( n28718 & n28720 ) | ( n28718 & ~n28724 ) | ( n28720 & ~n28724 ) ;
  assign n28726 = n28722 | n28725 ;
  assign n28727 = n28718 ^ x789 ^ 1'b0 ;
  assign n28728 = ( n28718 & n28726 ) | ( n28718 & n28727 ) | ( n28726 & n28727 ) ;
  assign n28729 = n28625 ^ n16518 ^ 1'b0 ;
  assign n28730 = ( n28625 & n28728 ) | ( n28625 & ~n28729 ) | ( n28728 & ~n28729 ) ;
  assign n28731 = n28625 ^ n16339 ^ 1'b0 ;
  assign n28732 = ( n28625 & n28730 ) | ( n28625 & ~n28731 ) | ( n28730 & ~n28731 ) ;
  assign n28733 = n28625 ^ n16376 ^ 1'b0 ;
  assign n28734 = ( n28625 & n28732 ) | ( n28625 & ~n28733 ) | ( n28732 & ~n28733 ) ;
  assign n28735 = x644 | n28734 ;
  assign n28736 = ( n28677 & ~n28678 ) | ( n28677 & n28735 ) | ( ~n28678 & n28735 ) ;
  assign n28737 = ( x1160 & n28678 ) | ( x1160 & n28736 ) | ( n28678 & n28736 ) ;
  assign n28738 = n28675 & ~n28737 ;
  assign n28739 = x644 & ~n28734 ;
  assign n28740 = ( ~x715 & n28625 ) | ( ~x715 & n28676 ) | ( n28625 & n28676 ) ;
  assign n28741 = x1160 & ~n28740 ;
  assign n28742 = ( x1160 & n28739 ) | ( x1160 & n28741 ) | ( n28739 & n28741 ) ;
  assign n28743 = ( x715 & n28673 ) | ( x715 & n28674 ) | ( n28673 & n28674 ) ;
  assign n28744 = n28742 & ~n28743 ;
  assign n28745 = ( x790 & n28738 ) | ( x790 & n28744 ) | ( n28738 & n28744 ) ;
  assign n28746 = n28744 ^ n28738 ^ 1'b0 ;
  assign n28747 = ( x790 & n28745 ) | ( x790 & n28746 ) | ( n28745 & n28746 ) ;
  assign n28748 = n16374 & n28668 ;
  assign n28749 = n19055 & n28732 ;
  assign n28750 = n28748 | n28749 ;
  assign n28751 = n16373 & n28669 ;
  assign n28752 = ( x787 & n28750 ) | ( x787 & n28751 ) | ( n28750 & n28751 ) ;
  assign n28753 = n28751 ^ n28750 ^ 1'b0 ;
  assign n28754 = ( x787 & n28752 ) | ( x787 & n28753 ) | ( n28752 & n28753 ) ;
  assign n28755 = x619 & ~n28655 ;
  assign n28756 = x1159 | n28755 ;
  assign n28804 = x625 | n28698 ;
  assign n28758 = x699 | n28696 ;
  assign n28759 = x763 & n15591 ;
  assign n28760 = n17156 | n28759 ;
  assign n28761 = x190 & ~n5017 ;
  assign n28762 = n28760 & n28761 ;
  assign n28763 = ~x763 & n22207 ;
  assign n28764 = n15968 | n28763 ;
  assign n28765 = x39 | n28764 ;
  assign n28766 = ( ~x39 & x190 ) | ( ~x39 & n28765 ) | ( x190 & n28765 ) ;
  assign n28767 = ( x38 & n28762 ) | ( x38 & n28766 ) | ( n28762 & n28766 ) ;
  assign n28768 = ~n28762 & n28767 ;
  assign n28769 = x190 & n15795 ;
  assign n28770 = x763 | n28769 ;
  assign n28771 = ( x190 & n15876 ) | ( x190 & ~n28770 ) | ( n15876 & ~n28770 ) ;
  assign n28772 = ~n28770 & n28771 ;
  assign n28773 = x190 | n16003 ;
  assign n28774 = x190 & n15943 ;
  assign n28775 = x763 & ~n28774 ;
  assign n28776 = n28773 & n28775 ;
  assign n28777 = ( x39 & n28772 ) | ( x39 & ~n28776 ) | ( n28772 & ~n28776 ) ;
  assign n28778 = ~n28772 & n28777 ;
  assign n28779 = x190 & n16054 ;
  assign n28780 = x190 | n16048 ;
  assign n28781 = ( x763 & n28779 ) | ( x763 & n28780 ) | ( n28779 & n28780 ) ;
  assign n28782 = ~n28779 & n28781 ;
  assign n28783 = x190 | n16044 ;
  assign n28784 = x190 & n16029 ;
  assign n28785 = ( x763 & n28783 ) | ( x763 & ~n28784 ) | ( n28783 & ~n28784 ) ;
  assign n28786 = ~x763 & n28785 ;
  assign n28787 = ( x39 & ~n28782 ) | ( x39 & n28786 ) | ( ~n28782 & n28786 ) ;
  assign n28788 = n28782 | n28787 ;
  assign n28789 = ( x38 & ~n28778 ) | ( x38 & n28788 ) | ( ~n28778 & n28788 ) ;
  assign n28790 = ~x38 & n28789 ;
  assign n28791 = ( x699 & n28768 ) | ( x699 & ~n28790 ) | ( n28768 & ~n28790 ) ;
  assign n28792 = ~n28768 & n28791 ;
  assign n28793 = ( n2051 & n2068 ) | ( n2051 & ~n28792 ) | ( n2068 & ~n28792 ) ;
  assign n28794 = n28792 | n28793 ;
  assign n28795 = ( n28679 & n28758 ) | ( n28679 & ~n28794 ) | ( n28758 & ~n28794 ) ;
  assign n28796 = n28795 ^ n28758 ^ 1'b0 ;
  assign n28797 = ( n28679 & n28795 ) | ( n28679 & ~n28796 ) | ( n28795 & ~n28796 ) ;
  assign n28805 = x625 & ~n28797 ;
  assign n28806 = x1153 & ~n28805 ;
  assign n28807 = n28804 & n28806 ;
  assign n28808 = ( x608 & n28648 ) | ( x608 & ~n28807 ) | ( n28648 & ~n28807 ) ;
  assign n28809 = ~n28648 & n28808 ;
  assign n28798 = x625 | n28797 ;
  assign n28799 = x625 & ~n28698 ;
  assign n28800 = ( x1153 & n28798 ) | ( x1153 & ~n28799 ) | ( n28798 & ~n28799 ) ;
  assign n28801 = ~x1153 & n28800 ;
  assign n28802 = ( x608 & n28644 ) | ( x608 & ~n28801 ) | ( n28644 & ~n28801 ) ;
  assign n28803 = n28801 | n28802 ;
  assign n28810 = n28809 ^ n28803 ^ 1'b0 ;
  assign n28811 = ( x778 & ~n28803 ) | ( x778 & n28809 ) | ( ~n28803 & n28809 ) ;
  assign n28812 = ( x778 & ~n28810 ) | ( x778 & n28811 ) | ( ~n28810 & n28811 ) ;
  assign n28813 = ( x778 & n28797 ) | ( x778 & ~n28812 ) | ( n28797 & ~n28812 ) ;
  assign n28814 = ~n28812 & n28813 ;
  assign n28815 = x609 & ~n28814 ;
  assign n28821 = x609 | n28651 ;
  assign n28822 = ( x1155 & n28815 ) | ( x1155 & n28821 ) | ( n28815 & n28821 ) ;
  assign n28823 = ~n28815 & n28822 ;
  assign n28824 = ~x1155 & n28703 ;
  assign n28825 = ( x660 & n28823 ) | ( x660 & ~n28824 ) | ( n28823 & ~n28824 ) ;
  assign n28826 = ~n28823 & n28825 ;
  assign n28757 = x1155 & n28704 ;
  assign n28816 = x609 & ~n28651 ;
  assign n28817 = x1155 | n28816 ;
  assign n28818 = ( n28814 & n28815 ) | ( n28814 & ~n28817 ) | ( n28815 & ~n28817 ) ;
  assign n28819 = ( x660 & ~n28757 ) | ( x660 & n28818 ) | ( ~n28757 & n28818 ) ;
  assign n28820 = n28757 | n28819 ;
  assign n28827 = n28826 ^ n28820 ^ 1'b0 ;
  assign n28828 = ( x785 & ~n28820 ) | ( x785 & n28826 ) | ( ~n28820 & n28826 ) ;
  assign n28829 = ( x785 & ~n28827 ) | ( x785 & n28828 ) | ( ~n28827 & n28828 ) ;
  assign n28830 = ( x785 & n28814 ) | ( x785 & ~n28829 ) | ( n28814 & ~n28829 ) ;
  assign n28831 = ~n28829 & n28830 ;
  assign n28832 = x618 & ~n28831 ;
  assign n28838 = x618 | n28653 ;
  assign n28839 = ( x1154 & n28832 ) | ( x1154 & n28838 ) | ( n28832 & n28838 ) ;
  assign n28840 = ~n28832 & n28839 ;
  assign n28841 = ( x627 & n28715 ) | ( x627 & ~n28840 ) | ( n28715 & ~n28840 ) ;
  assign n28842 = ~n28715 & n28841 ;
  assign n28833 = x618 & ~n28653 ;
  assign n28834 = x1154 | n28833 ;
  assign n28835 = ( n28831 & n28832 ) | ( n28831 & ~n28834 ) | ( n28832 & ~n28834 ) ;
  assign n28836 = ( x627 & n28712 ) | ( x627 & ~n28835 ) | ( n28712 & ~n28835 ) ;
  assign n28837 = n28835 | n28836 ;
  assign n28843 = n28842 ^ n28837 ^ 1'b0 ;
  assign n28844 = ( x781 & ~n28837 ) | ( x781 & n28842 ) | ( ~n28837 & n28842 ) ;
  assign n28845 = ( x781 & ~n28843 ) | ( x781 & n28844 ) | ( ~n28843 & n28844 ) ;
  assign n28846 = ( x781 & n28831 ) | ( x781 & ~n28845 ) | ( n28831 & ~n28845 ) ;
  assign n28847 = ~n28845 & n28846 ;
  assign n28848 = x619 & ~n28847 ;
  assign n28849 = ( ~n28756 & n28847 ) | ( ~n28756 & n28848 ) | ( n28847 & n28848 ) ;
  assign n28850 = ( x648 & n28722 ) | ( x648 & ~n28849 ) | ( n28722 & ~n28849 ) ;
  assign n28851 = n28849 | n28850 ;
  assign n28852 = x619 | n28655 ;
  assign n28853 = x1159 & ~n28848 ;
  assign n28854 = n28852 & n28853 ;
  assign n28855 = ( x648 & n28725 ) | ( x648 & ~n28854 ) | ( n28725 & ~n28854 ) ;
  assign n28856 = ~n28725 & n28855 ;
  assign n28857 = x789 & ~n28856 ;
  assign n28858 = n28851 & n28857 ;
  assign n28859 = ~x789 & n28847 ;
  assign n28860 = ( n16519 & ~n28858 ) | ( n16519 & n28859 ) | ( ~n28858 & n28859 ) ;
  assign n28861 = n28858 | n28860 ;
  assign n28862 = n16337 & n28662 ;
  assign n28863 = n16338 & n28661 ;
  assign n28864 = n28862 | n28863 ;
  assign n28865 = n19046 & n28730 ;
  assign n28866 = ( x792 & n28864 ) | ( x792 & n28865 ) | ( n28864 & n28865 ) ;
  assign n28867 = n28865 ^ n28864 ^ 1'b0 ;
  assign n28868 = ( x792 & n28866 ) | ( x792 & n28867 ) | ( n28866 & n28867 ) ;
  assign n28869 = n16459 & ~n28657 ;
  assign n28870 = ~x626 & n28625 ;
  assign n28871 = x626 & n28728 ;
  assign n28872 = ( n22317 & n28870 ) | ( n22317 & ~n28871 ) | ( n28870 & ~n28871 ) ;
  assign n28873 = ~n28870 & n28872 ;
  assign n28874 = ~x626 & n28728 ;
  assign n28875 = x626 & n28625 ;
  assign n28876 = ( n22322 & n28874 ) | ( n22322 & ~n28875 ) | ( n28874 & ~n28875 ) ;
  assign n28877 = ~n28874 & n28876 ;
  assign n28878 = ( ~n28869 & n28873 ) | ( ~n28869 & n28877 ) | ( n28873 & n28877 ) ;
  assign n28879 = n28869 | n28878 ;
  assign n28880 = ( x788 & ~n22314 ) | ( x788 & n28879 ) | ( ~n22314 & n28879 ) ;
  assign n28881 = ( n18482 & n22314 ) | ( n18482 & n28880 ) | ( n22314 & n28880 ) ;
  assign n28882 = ~n28868 & n28881 ;
  assign n28883 = ( n28861 & n28868 ) | ( n28861 & ~n28882 ) | ( n28868 & ~n28882 ) ;
  assign n28884 = ( ~n18484 & n28754 ) | ( ~n18484 & n28883 ) | ( n28754 & n28883 ) ;
  assign n28885 = n28754 ^ n18484 ^ 1'b0 ;
  assign n28886 = ( n28754 & n28884 ) | ( n28754 & ~n28885 ) | ( n28884 & ~n28885 ) ;
  assign n28887 = x644 | n28737 ;
  assign n28888 = x644 & n28742 ;
  assign n28889 = x790 & ~n28888 ;
  assign n28890 = n28887 & n28889 ;
  assign n28891 = ( ~n28747 & n28886 ) | ( ~n28747 & n28890 ) | ( n28886 & n28890 ) ;
  assign n28892 = ~n28747 & n28891 ;
  assign n28893 = ( x57 & n5193 ) | ( x57 & ~n28892 ) | ( n5193 & ~n28892 ) ;
  assign n28894 = n28892 | n28893 ;
  assign n28895 = x190 | n1611 ;
  assign n28896 = ~n28759 & n28895 ;
  assign n28897 = n16397 | n28896 ;
  assign n28898 = ~n15662 & n28759 ;
  assign n28899 = ~x1155 & n28895 ;
  assign n28900 = ~n28898 & n28899 ;
  assign n28901 = ( x1155 & n28897 ) | ( x1155 & n28898 ) | ( n28897 & n28898 ) ;
  assign n28902 = n28900 | n28901 ;
  assign n28903 = n28897 ^ x785 ^ 1'b0 ;
  assign n28904 = ( n28897 & n28902 ) | ( n28897 & n28903 ) | ( n28902 & n28903 ) ;
  assign n28905 = n16411 | n28904 ;
  assign n28906 = x1154 & n28905 ;
  assign n28907 = n16414 | n28904 ;
  assign n28908 = ~x1154 & n28907 ;
  assign n28909 = n28906 | n28908 ;
  assign n28910 = n28904 ^ x781 ^ 1'b0 ;
  assign n28911 = ( n28904 & n28909 ) | ( n28904 & n28910 ) | ( n28909 & n28910 ) ;
  assign n28912 = n21437 | n28911 ;
  assign n28913 = x1159 & n28912 ;
  assign n28914 = n21440 | n28911 ;
  assign n28915 = ~x1159 & n28914 ;
  assign n28916 = n28913 | n28915 ;
  assign n28917 = n28911 ^ x789 ^ 1'b0 ;
  assign n28918 = ( n28911 & n28916 ) | ( n28911 & n28917 ) | ( n28916 & n28917 ) ;
  assign n28919 = n28895 ^ n16518 ^ 1'b0 ;
  assign n28920 = ( n28895 & n28918 ) | ( n28895 & ~n28919 ) | ( n28918 & ~n28919 ) ;
  assign n28921 = n28895 ^ n16339 ^ 1'b0 ;
  assign n28922 = ( n28895 & n28920 ) | ( n28895 & ~n28921 ) | ( n28920 & ~n28921 ) ;
  assign n28923 = n19055 & n28922 ;
  assign n28924 = x647 & ~n28895 ;
  assign n28925 = x1157 | n28924 ;
  assign n28926 = x699 & n15778 ;
  assign n28927 = ~x625 & n28926 ;
  assign n28928 = ~x1153 & n28895 ;
  assign n28929 = ~n28927 & n28928 ;
  assign n28930 = x778 & ~n28929 ;
  assign n28931 = n28895 & ~n28926 ;
  assign n28932 = ( x1153 & n28927 ) | ( x1153 & n28931 ) | ( n28927 & n28931 ) ;
  assign n28933 = n28930 & ~n28932 ;
  assign n28934 = ( x778 & n28931 ) | ( x778 & ~n28933 ) | ( n28931 & ~n28933 ) ;
  assign n28935 = ~n28933 & n28934 ;
  assign n28936 = n16447 | n28935 ;
  assign n28937 = n16449 | n28936 ;
  assign n28938 = n16451 | n28937 ;
  assign n28939 = n16530 | n28938 ;
  assign n28940 = n16560 | n28939 ;
  assign n28941 = ( x647 & ~n28925 ) | ( x647 & n28940 ) | ( ~n28925 & n28940 ) ;
  assign n28942 = ~n28925 & n28941 ;
  assign n28943 = n28895 ^ x647 ^ 1'b0 ;
  assign n28944 = ( n28895 & n28940 ) | ( n28895 & n28943 ) | ( n28940 & n28943 ) ;
  assign n28945 = x1157 & n28944 ;
  assign n28946 = ( n16375 & n28942 ) | ( n16375 & n28945 ) | ( n28942 & n28945 ) ;
  assign n28947 = ( x787 & n28923 ) | ( x787 & n28946 ) | ( n28923 & n28946 ) ;
  assign n28948 = n28946 ^ n28923 ^ 1'b0 ;
  assign n28949 = ( x787 & n28947 ) | ( x787 & n28948 ) | ( n28947 & n28948 ) ;
  assign n28950 = ~x626 & n28895 ;
  assign n28951 = x626 & n28918 ;
  assign n28952 = ( n22317 & n28950 ) | ( n22317 & ~n28951 ) | ( n28950 & ~n28951 ) ;
  assign n28953 = ~n28950 & n28952 ;
  assign n28954 = ~x626 & n28918 ;
  assign n28955 = x626 & n28895 ;
  assign n28956 = ( n22322 & n28954 ) | ( n22322 & ~n28955 ) | ( n28954 & ~n28955 ) ;
  assign n28957 = ~n28954 & n28956 ;
  assign n28958 = n28938 & ~n28957 ;
  assign n28959 = ( n16459 & n28957 ) | ( n16459 & ~n28958 ) | ( n28957 & ~n28958 ) ;
  assign n28960 = ( x788 & n28953 ) | ( x788 & n28959 ) | ( n28953 & n28959 ) ;
  assign n28961 = n28959 ^ n28953 ^ 1'b0 ;
  assign n28962 = ( x788 & n28960 ) | ( x788 & n28961 ) | ( n28960 & n28961 ) ;
  assign n28963 = n15524 | n28931 ;
  assign n28964 = n28896 & n28963 ;
  assign n28965 = x625 & ~n28963 ;
  assign n28966 = ( n28928 & n28964 ) | ( n28928 & n28965 ) | ( n28964 & n28965 ) ;
  assign n28967 = ( x608 & n28932 ) | ( x608 & ~n28966 ) | ( n28932 & ~n28966 ) ;
  assign n28968 = n28966 | n28967 ;
  assign n28969 = x1153 & n28896 ;
  assign n28970 = ~n28965 & n28969 ;
  assign n28971 = x608 & ~n28929 ;
  assign n28972 = n28968 & ~n28971 ;
  assign n28973 = ( n28968 & n28970 ) | ( n28968 & n28972 ) | ( n28970 & n28972 ) ;
  assign n28974 = n28964 ^ x778 ^ 1'b0 ;
  assign n28975 = ( n28964 & n28973 ) | ( n28964 & n28974 ) | ( n28973 & n28974 ) ;
  assign n28976 = x609 & ~n28975 ;
  assign n28982 = x609 | n28935 ;
  assign n28983 = ( x1155 & n28976 ) | ( x1155 & n28982 ) | ( n28976 & n28982 ) ;
  assign n28984 = ~n28976 & n28983 ;
  assign n28985 = ( x660 & n28900 ) | ( x660 & ~n28984 ) | ( n28900 & ~n28984 ) ;
  assign n28986 = ~n28900 & n28985 ;
  assign n28977 = x609 & ~n28935 ;
  assign n28978 = x1155 | n28977 ;
  assign n28979 = ( n28975 & n28976 ) | ( n28975 & ~n28978 ) | ( n28976 & ~n28978 ) ;
  assign n28980 = ( x660 & n28901 ) | ( x660 & ~n28979 ) | ( n28901 & ~n28979 ) ;
  assign n28981 = n28979 | n28980 ;
  assign n28987 = n28986 ^ n28981 ^ 1'b0 ;
  assign n28988 = ( x785 & ~n28981 ) | ( x785 & n28986 ) | ( ~n28981 & n28986 ) ;
  assign n28989 = ( x785 & ~n28987 ) | ( x785 & n28988 ) | ( ~n28987 & n28988 ) ;
  assign n28990 = ( x785 & n28975 ) | ( x785 & ~n28989 ) | ( n28975 & ~n28989 ) ;
  assign n28991 = ~n28989 & n28990 ;
  assign n28992 = x618 & ~n28991 ;
  assign n28993 = x618 | n28936 ;
  assign n28994 = ( x1154 & n28992 ) | ( x1154 & n28993 ) | ( n28992 & n28993 ) ;
  assign n28995 = ~n28992 & n28994 ;
  assign n28996 = ( x627 & n28908 ) | ( x627 & ~n28995 ) | ( n28908 & ~n28995 ) ;
  assign n28997 = ~n28908 & n28996 ;
  assign n28998 = x627 | n28906 ;
  assign n28999 = x618 & ~n28936 ;
  assign n29000 = x1154 | n28999 ;
  assign n29001 = ( n28991 & n28992 ) | ( n28991 & ~n29000 ) | ( n28992 & ~n29000 ) ;
  assign n29002 = ( ~n28997 & n28998 ) | ( ~n28997 & n29001 ) | ( n28998 & n29001 ) ;
  assign n29003 = ~n28997 & n29002 ;
  assign n29004 = n28991 ^ x781 ^ 1'b0 ;
  assign n29005 = ( n28991 & n29003 ) | ( n28991 & n29004 ) | ( n29003 & n29004 ) ;
  assign n29006 = ~x789 & n29005 ;
  assign n29007 = x619 & ~n28937 ;
  assign n29008 = x1159 | n29007 ;
  assign n29009 = x619 & ~n29005 ;
  assign n29010 = ( n29005 & ~n29008 ) | ( n29005 & n29009 ) | ( ~n29008 & n29009 ) ;
  assign n29011 = ( x648 & n28913 ) | ( x648 & ~n29010 ) | ( n28913 & ~n29010 ) ;
  assign n29012 = n29010 | n29011 ;
  assign n29013 = x619 | n28937 ;
  assign n29014 = x1159 & ~n29009 ;
  assign n29015 = n29013 & n29014 ;
  assign n29016 = ( x648 & n28915 ) | ( x648 & ~n29015 ) | ( n28915 & ~n29015 ) ;
  assign n29017 = ~n28915 & n29016 ;
  assign n29018 = x789 & ~n29017 ;
  assign n29019 = n29012 & n29018 ;
  assign n29020 = ( n16519 & ~n29006 ) | ( n16519 & n29019 ) | ( ~n29006 & n29019 ) ;
  assign n29021 = n29006 | n29020 ;
  assign n29022 = n29021 ^ n28962 ^ 1'b0 ;
  assign n29023 = ( n28962 & n29021 ) | ( n28962 & n29022 ) | ( n29021 & n29022 ) ;
  assign n29024 = ( n18482 & ~n28962 ) | ( n18482 & n29023 ) | ( ~n28962 & n29023 ) ;
  assign n29025 = n19208 | n28939 ;
  assign n29026 = n16556 & ~n28920 ;
  assign n29027 = x629 & ~n29026 ;
  assign n29028 = n29025 & n29027 ;
  assign n29029 = n16557 & ~n28920 ;
  assign n29030 = n19212 & ~n28939 ;
  assign n29031 = n29029 | n29030 ;
  assign n29032 = ( x629 & ~n29028 ) | ( x629 & n29031 ) | ( ~n29028 & n29031 ) ;
  assign n29033 = ~n29028 & n29032 ;
  assign n29034 = ( x792 & ~n19206 ) | ( x792 & n29033 ) | ( ~n19206 & n29033 ) ;
  assign n29035 = ( n18484 & n19206 ) | ( n18484 & n29034 ) | ( n19206 & n29034 ) ;
  assign n29036 = ( n28949 & n29024 ) | ( n28949 & ~n29035 ) | ( n29024 & ~n29035 ) ;
  assign n29037 = n29036 ^ n29024 ^ 1'b0 ;
  assign n29038 = ( n28949 & n29036 ) | ( n28949 & ~n29037 ) | ( n29036 & ~n29037 ) ;
  assign n29039 = x790 | n29038 ;
  assign n29040 = x644 & ~n29038 ;
  assign n29041 = ( x787 & n28942 ) | ( x787 & ~n28945 ) | ( n28942 & ~n28945 ) ;
  assign n29042 = ~n28942 & n29041 ;
  assign n29043 = ( x787 & n28940 ) | ( x787 & ~n29042 ) | ( n28940 & ~n29042 ) ;
  assign n29044 = ~n29042 & n29043 ;
  assign n29045 = x644 | n29044 ;
  assign n29046 = ( x715 & n29040 ) | ( x715 & n29045 ) | ( n29040 & n29045 ) ;
  assign n29047 = ~n29040 & n29046 ;
  assign n29048 = x644 | n28895 ;
  assign n29049 = n28895 ^ n16376 ^ 1'b0 ;
  assign n29050 = ( n28895 & n28922 ) | ( n28895 & ~n29049 ) | ( n28922 & ~n29049 ) ;
  assign n29051 = x644 & ~n29050 ;
  assign n29052 = ( x715 & n29048 ) | ( x715 & ~n29051 ) | ( n29048 & ~n29051 ) ;
  assign n29053 = ~x715 & n29052 ;
  assign n29054 = ( x1160 & n29047 ) | ( x1160 & ~n29053 ) | ( n29047 & ~n29053 ) ;
  assign n29055 = ~n29047 & n29054 ;
  assign n29056 = x644 & ~n28895 ;
  assign n29057 = x715 & ~n29056 ;
  assign n29058 = ( n29050 & n29051 ) | ( n29050 & n29057 ) | ( n29051 & n29057 ) ;
  assign n29059 = x644 & ~n29044 ;
  assign n29060 = x715 | n29059 ;
  assign n29061 = ( n29038 & n29040 ) | ( n29038 & ~n29060 ) | ( n29040 & ~n29060 ) ;
  assign n29062 = ( x1160 & ~n29058 ) | ( x1160 & n29061 ) | ( ~n29058 & n29061 ) ;
  assign n29063 = n29058 | n29062 ;
  assign n29064 = x790 & ~n29063 ;
  assign n29065 = ( x790 & n29055 ) | ( x790 & n29064 ) | ( n29055 & n29064 ) ;
  assign n29066 = x832 & ~n29065 ;
  assign n29067 = n29039 & n29066 ;
  assign n29068 = ~x190 & n7318 ;
  assign n29069 = x832 | n29068 ;
  assign n29070 = ~n29067 & n29069 ;
  assign n29071 = ( n28894 & n29067 ) | ( n28894 & ~n29070 ) | ( n29067 & ~n29070 ) ;
  assign n29072 = x191 | n15656 ;
  assign n29073 = x191 | n15644 ;
  assign n29074 = n16185 & n29073 ;
  assign n29075 = x191 | n16697 ;
  assign n29076 = x191 & n16699 ;
  assign n29077 = ( x38 & n29075 ) | ( x38 & ~n29076 ) | ( n29075 & ~n29076 ) ;
  assign n29078 = ~x38 & n29077 ;
  assign n29079 = ( x729 & n29074 ) | ( x729 & ~n29078 ) | ( n29074 & ~n29078 ) ;
  assign n29080 = ~n29074 & n29079 ;
  assign n29081 = x191 | x729 ;
  assign n29082 = n15655 | n29081 ;
  assign n29083 = ( n2069 & ~n29080 ) | ( n2069 & n29082 ) | ( ~n29080 & n29082 ) ;
  assign n29084 = ~n2069 & n29083 ;
  assign n29085 = n29084 ^ x191 ^ 1'b0 ;
  assign n29086 = ( ~x191 & n2069 ) | ( ~x191 & n29085 ) | ( n2069 & n29085 ) ;
  assign n29087 = ( x191 & n29084 ) | ( x191 & n29086 ) | ( n29084 & n29086 ) ;
  assign n29088 = x625 & ~n29087 ;
  assign n29089 = x625 | n29072 ;
  assign n29090 = ( x1153 & n29088 ) | ( x1153 & n29089 ) | ( n29088 & n29089 ) ;
  assign n29091 = ~n29088 & n29090 ;
  assign n29092 = x625 & ~n29072 ;
  assign n29093 = x1153 | n29092 ;
  assign n29094 = ( x625 & n29087 ) | ( x625 & ~n29093 ) | ( n29087 & ~n29093 ) ;
  assign n29095 = ~n29093 & n29094 ;
  assign n29096 = n29091 | n29095 ;
  assign n29097 = n29087 ^ x778 ^ 1'b0 ;
  assign n29098 = ( n29087 & n29096 ) | ( n29087 & n29097 ) | ( n29096 & n29097 ) ;
  assign n29099 = n29072 ^ n16234 ^ 1'b0 ;
  assign n29100 = ( n29072 & n29098 ) | ( n29072 & ~n29099 ) | ( n29098 & ~n29099 ) ;
  assign n29101 = n29072 ^ n16254 ^ 1'b0 ;
  assign n29102 = ( n29072 & n29100 ) | ( n29072 & ~n29101 ) | ( n29100 & ~n29101 ) ;
  assign n29103 = n29072 ^ n16279 ^ 1'b0 ;
  assign n29104 = ( n29072 & n29102 ) | ( n29072 & ~n29103 ) | ( n29102 & ~n29103 ) ;
  assign n29105 = n29072 ^ n16318 ^ 1'b0 ;
  assign n29106 = ( n29072 & n29104 ) | ( n29072 & ~n29105 ) | ( n29104 & ~n29105 ) ;
  assign n29107 = n29072 ^ x628 ^ 1'b0 ;
  assign n29108 = ( n29072 & n29106 ) | ( n29072 & ~n29107 ) | ( n29106 & ~n29107 ) ;
  assign n29109 = ( n29072 & n29106 ) | ( n29072 & n29107 ) | ( n29106 & n29107 ) ;
  assign n29110 = n29108 ^ x1156 ^ 1'b0 ;
  assign n29111 = ( n29108 & n29109 ) | ( n29108 & n29110 ) | ( n29109 & n29110 ) ;
  assign n29112 = n29106 ^ x792 ^ 1'b0 ;
  assign n29113 = ( n29106 & n29111 ) | ( n29106 & n29112 ) | ( n29111 & n29112 ) ;
  assign n29114 = n29072 ^ x647 ^ 1'b0 ;
  assign n29115 = ( n29072 & n29113 ) | ( n29072 & ~n29114 ) | ( n29113 & ~n29114 ) ;
  assign n29116 = ( n29072 & n29113 ) | ( n29072 & n29114 ) | ( n29113 & n29114 ) ;
  assign n29117 = n29115 ^ x1157 ^ 1'b0 ;
  assign n29118 = ( n29115 & n29116 ) | ( n29115 & n29117 ) | ( n29116 & n29117 ) ;
  assign n29119 = n29113 ^ x787 ^ 1'b0 ;
  assign n29120 = ( n29113 & n29118 ) | ( n29113 & n29119 ) | ( n29118 & n29119 ) ;
  assign n29121 = x644 & ~n29120 ;
  assign n29122 = x715 | n29121 ;
  assign n29123 = x644 & ~n29072 ;
  assign n29124 = x715 & ~n29123 ;
  assign n29125 = n29124 ^ x1160 ^ 1'b0 ;
  assign n29126 = x191 & n2069 ;
  assign n29127 = x38 & n29073 ;
  assign n29128 = ~x191 & x746 ;
  assign n29129 = n15587 & n29128 ;
  assign n29130 = x746 & n15639 ;
  assign n29131 = x191 & ~n29130 ;
  assign n29132 = ( n20873 & ~n29129 ) | ( n20873 & n29131 ) | ( ~n29129 & n29131 ) ;
  assign n29133 = n29129 | n29132 ;
  assign n29134 = x191 & ~n15631 ;
  assign n29135 = ~x746 & n15486 ;
  assign n29136 = ( x39 & n29134 ) | ( x39 & n29135 ) | ( n29134 & n29135 ) ;
  assign n29137 = n29135 ^ n29134 ^ 1'b0 ;
  assign n29138 = ( x39 & n29136 ) | ( x39 & n29137 ) | ( n29136 & n29137 ) ;
  assign n29139 = ( ~x38 & n29133 ) | ( ~x38 & n29138 ) | ( n29133 & n29138 ) ;
  assign n29140 = ~x38 & n29139 ;
  assign n29141 = x746 & n15646 ;
  assign n29142 = ~n29140 & n29141 ;
  assign n29143 = ( n29127 & n29140 ) | ( n29127 & ~n29142 ) | ( n29140 & ~n29142 ) ;
  assign n29144 = ~n2069 & n29143 ;
  assign n29145 = n29126 | n29144 ;
  assign n29146 = n29072 ^ n15659 ^ 1'b0 ;
  assign n29147 = ( n29072 & n29145 ) | ( n29072 & ~n29146 ) | ( n29145 & ~n29146 ) ;
  assign n29148 = n15662 & n29072 ;
  assign n29149 = ( ~n15662 & n29126 ) | ( ~n15662 & n29144 ) | ( n29126 & n29144 ) ;
  assign n29150 = n29148 | n29149 ;
  assign n29151 = n29150 ^ n29147 ^ n29072 ;
  assign n29152 = n29151 ^ x1155 ^ 1'b0 ;
  assign n29153 = ( n29150 & n29151 ) | ( n29150 & ~n29152 ) | ( n29151 & ~n29152 ) ;
  assign n29154 = n29147 ^ x785 ^ 1'b0 ;
  assign n29155 = ( n29147 & n29153 ) | ( n29147 & n29154 ) | ( n29153 & n29154 ) ;
  assign n29156 = x618 & ~n29155 ;
  assign n29157 = x618 | n29072 ;
  assign n29158 = ( x1154 & n29156 ) | ( x1154 & n29157 ) | ( n29156 & n29157 ) ;
  assign n29159 = ~n29156 & n29158 ;
  assign n29160 = x618 & ~n29072 ;
  assign n29161 = x1154 | n29160 ;
  assign n29162 = ( n29155 & n29156 ) | ( n29155 & ~n29161 ) | ( n29156 & ~n29161 ) ;
  assign n29163 = n29159 | n29162 ;
  assign n29164 = n29155 ^ x781 ^ 1'b0 ;
  assign n29165 = ( n29155 & n29163 ) | ( n29155 & n29164 ) | ( n29163 & n29164 ) ;
  assign n29166 = x619 | n29072 ;
  assign n29167 = x619 & ~n29165 ;
  assign n29168 = x1159 & ~n29167 ;
  assign n29169 = n29166 & n29168 ;
  assign n29170 = x619 & ~n29072 ;
  assign n29171 = x1159 | n29170 ;
  assign n29172 = ( n29165 & n29167 ) | ( n29165 & ~n29171 ) | ( n29167 & ~n29171 ) ;
  assign n29173 = n29169 | n29172 ;
  assign n29174 = n29165 ^ x789 ^ 1'b0 ;
  assign n29175 = ( n29165 & n29173 ) | ( n29165 & n29174 ) | ( n29173 & n29174 ) ;
  assign n29176 = n29072 ^ n16518 ^ 1'b0 ;
  assign n29177 = ( n29072 & n29175 ) | ( n29072 & ~n29176 ) | ( n29175 & ~n29176 ) ;
  assign n29178 = n29072 ^ n16339 ^ 1'b0 ;
  assign n29179 = ( n29072 & n29177 ) | ( n29072 & ~n29178 ) | ( n29177 & ~n29178 ) ;
  assign n29180 = n29072 ^ n16376 ^ 1'b0 ;
  assign n29181 = ( n29072 & n29179 ) | ( n29072 & ~n29180 ) | ( n29179 & ~n29180 ) ;
  assign n29182 = x644 | n29181 ;
  assign n29183 = ( n29124 & ~n29125 ) | ( n29124 & n29182 ) | ( ~n29125 & n29182 ) ;
  assign n29184 = ( x1160 & n29125 ) | ( x1160 & n29183 ) | ( n29125 & n29183 ) ;
  assign n29185 = n29122 & ~n29184 ;
  assign n29186 = x644 & ~n29181 ;
  assign n29187 = ( ~x715 & n29072 ) | ( ~x715 & n29123 ) | ( n29072 & n29123 ) ;
  assign n29188 = x1160 & ~n29187 ;
  assign n29189 = ( x1160 & n29186 ) | ( x1160 & n29188 ) | ( n29186 & n29188 ) ;
  assign n29190 = ( x715 & n29120 ) | ( x715 & n29121 ) | ( n29120 & n29121 ) ;
  assign n29191 = n29189 & ~n29190 ;
  assign n29192 = ( x790 & n29185 ) | ( x790 & n29191 ) | ( n29185 & n29191 ) ;
  assign n29193 = n29191 ^ n29185 ^ 1'b0 ;
  assign n29194 = ( x790 & n29192 ) | ( x790 & n29193 ) | ( n29192 & n29193 ) ;
  assign n29195 = n16374 & n29115 ;
  assign n29196 = n19055 & n29179 ;
  assign n29197 = n29195 | n29196 ;
  assign n29198 = n16373 & n29116 ;
  assign n29199 = ( x787 & n29197 ) | ( x787 & n29198 ) | ( n29197 & n29198 ) ;
  assign n29200 = n29198 ^ n29197 ^ 1'b0 ;
  assign n29201 = ( x787 & n29199 ) | ( x787 & n29200 ) | ( n29199 & n29200 ) ;
  assign n29202 = x619 & ~n29102 ;
  assign n29203 = x1159 | n29202 ;
  assign n29251 = x625 | n29145 ;
  assign n29205 = x729 | n29143 ;
  assign n29206 = x746 & n15591 ;
  assign n29207 = n17156 | n29206 ;
  assign n29208 = x191 & ~n5017 ;
  assign n29209 = n29207 & n29208 ;
  assign n29210 = ~x746 & n22207 ;
  assign n29211 = n15968 | n29210 ;
  assign n29212 = x39 | n29211 ;
  assign n29213 = ( ~x39 & x191 ) | ( ~x39 & n29212 ) | ( x191 & n29212 ) ;
  assign n29214 = ( x38 & n29209 ) | ( x38 & n29213 ) | ( n29209 & n29213 ) ;
  assign n29215 = ~n29209 & n29214 ;
  assign n29216 = x191 & n15795 ;
  assign n29217 = x746 | n29216 ;
  assign n29218 = ( x191 & n15876 ) | ( x191 & ~n29217 ) | ( n15876 & ~n29217 ) ;
  assign n29219 = ~n29217 & n29218 ;
  assign n29220 = x191 | n16003 ;
  assign n29221 = x191 & n15943 ;
  assign n29222 = x746 & ~n29221 ;
  assign n29223 = n29220 & n29222 ;
  assign n29224 = ( x39 & n29219 ) | ( x39 & ~n29223 ) | ( n29219 & ~n29223 ) ;
  assign n29225 = ~n29219 & n29224 ;
  assign n29226 = x191 & n16054 ;
  assign n29227 = x191 | n16048 ;
  assign n29228 = ( x746 & n29226 ) | ( x746 & n29227 ) | ( n29226 & n29227 ) ;
  assign n29229 = ~n29226 & n29228 ;
  assign n29230 = x191 | n16044 ;
  assign n29231 = x191 & n16029 ;
  assign n29232 = ( x746 & n29230 ) | ( x746 & ~n29231 ) | ( n29230 & ~n29231 ) ;
  assign n29233 = ~x746 & n29232 ;
  assign n29234 = ( x39 & ~n29229 ) | ( x39 & n29233 ) | ( ~n29229 & n29233 ) ;
  assign n29235 = n29229 | n29234 ;
  assign n29236 = ( x38 & ~n29225 ) | ( x38 & n29235 ) | ( ~n29225 & n29235 ) ;
  assign n29237 = ~x38 & n29236 ;
  assign n29238 = ( x729 & n29215 ) | ( x729 & ~n29237 ) | ( n29215 & ~n29237 ) ;
  assign n29239 = ~n29215 & n29238 ;
  assign n29240 = ( n2051 & n2068 ) | ( n2051 & ~n29239 ) | ( n2068 & ~n29239 ) ;
  assign n29241 = n29239 | n29240 ;
  assign n29242 = ( n29126 & n29205 ) | ( n29126 & ~n29241 ) | ( n29205 & ~n29241 ) ;
  assign n29243 = n29242 ^ n29205 ^ 1'b0 ;
  assign n29244 = ( n29126 & n29242 ) | ( n29126 & ~n29243 ) | ( n29242 & ~n29243 ) ;
  assign n29252 = x625 & ~n29244 ;
  assign n29253 = x1153 & ~n29252 ;
  assign n29254 = n29251 & n29253 ;
  assign n29255 = ( x608 & n29095 ) | ( x608 & ~n29254 ) | ( n29095 & ~n29254 ) ;
  assign n29256 = ~n29095 & n29255 ;
  assign n29245 = x625 | n29244 ;
  assign n29246 = x625 & ~n29145 ;
  assign n29247 = ( x1153 & n29245 ) | ( x1153 & ~n29246 ) | ( n29245 & ~n29246 ) ;
  assign n29248 = ~x1153 & n29247 ;
  assign n29249 = ( x608 & n29091 ) | ( x608 & ~n29248 ) | ( n29091 & ~n29248 ) ;
  assign n29250 = n29248 | n29249 ;
  assign n29257 = n29256 ^ n29250 ^ 1'b0 ;
  assign n29258 = ( x778 & ~n29250 ) | ( x778 & n29256 ) | ( ~n29250 & n29256 ) ;
  assign n29259 = ( x778 & ~n29257 ) | ( x778 & n29258 ) | ( ~n29257 & n29258 ) ;
  assign n29260 = ( x778 & n29244 ) | ( x778 & ~n29259 ) | ( n29244 & ~n29259 ) ;
  assign n29261 = ~n29259 & n29260 ;
  assign n29262 = x609 & ~n29261 ;
  assign n29268 = x609 | n29098 ;
  assign n29269 = ( x1155 & n29262 ) | ( x1155 & n29268 ) | ( n29262 & n29268 ) ;
  assign n29270 = ~n29262 & n29269 ;
  assign n29271 = ~x1155 & n29150 ;
  assign n29272 = ( x660 & n29270 ) | ( x660 & ~n29271 ) | ( n29270 & ~n29271 ) ;
  assign n29273 = ~n29270 & n29272 ;
  assign n29204 = x1155 & n29151 ;
  assign n29263 = x609 & ~n29098 ;
  assign n29264 = x1155 | n29263 ;
  assign n29265 = ( n29261 & n29262 ) | ( n29261 & ~n29264 ) | ( n29262 & ~n29264 ) ;
  assign n29266 = ( x660 & ~n29204 ) | ( x660 & n29265 ) | ( ~n29204 & n29265 ) ;
  assign n29267 = n29204 | n29266 ;
  assign n29274 = n29273 ^ n29267 ^ 1'b0 ;
  assign n29275 = ( x785 & ~n29267 ) | ( x785 & n29273 ) | ( ~n29267 & n29273 ) ;
  assign n29276 = ( x785 & ~n29274 ) | ( x785 & n29275 ) | ( ~n29274 & n29275 ) ;
  assign n29277 = ( x785 & n29261 ) | ( x785 & ~n29276 ) | ( n29261 & ~n29276 ) ;
  assign n29278 = ~n29276 & n29277 ;
  assign n29279 = x618 & ~n29278 ;
  assign n29285 = x618 | n29100 ;
  assign n29286 = ( x1154 & n29279 ) | ( x1154 & n29285 ) | ( n29279 & n29285 ) ;
  assign n29287 = ~n29279 & n29286 ;
  assign n29288 = ( x627 & n29162 ) | ( x627 & ~n29287 ) | ( n29162 & ~n29287 ) ;
  assign n29289 = ~n29162 & n29288 ;
  assign n29280 = x618 & ~n29100 ;
  assign n29281 = x1154 | n29280 ;
  assign n29282 = ( n29278 & n29279 ) | ( n29278 & ~n29281 ) | ( n29279 & ~n29281 ) ;
  assign n29283 = ( x627 & n29159 ) | ( x627 & ~n29282 ) | ( n29159 & ~n29282 ) ;
  assign n29284 = n29282 | n29283 ;
  assign n29290 = n29289 ^ n29284 ^ 1'b0 ;
  assign n29291 = ( x781 & ~n29284 ) | ( x781 & n29289 ) | ( ~n29284 & n29289 ) ;
  assign n29292 = ( x781 & ~n29290 ) | ( x781 & n29291 ) | ( ~n29290 & n29291 ) ;
  assign n29293 = ( x781 & n29278 ) | ( x781 & ~n29292 ) | ( n29278 & ~n29292 ) ;
  assign n29294 = ~n29292 & n29293 ;
  assign n29295 = x619 & ~n29294 ;
  assign n29296 = ( ~n29203 & n29294 ) | ( ~n29203 & n29295 ) | ( n29294 & n29295 ) ;
  assign n29297 = ( x648 & n29169 ) | ( x648 & ~n29296 ) | ( n29169 & ~n29296 ) ;
  assign n29298 = n29296 | n29297 ;
  assign n29299 = x619 | n29102 ;
  assign n29300 = x1159 & ~n29295 ;
  assign n29301 = n29299 & n29300 ;
  assign n29302 = ( x648 & n29172 ) | ( x648 & ~n29301 ) | ( n29172 & ~n29301 ) ;
  assign n29303 = ~n29172 & n29302 ;
  assign n29304 = x789 & ~n29303 ;
  assign n29305 = n29298 & n29304 ;
  assign n29306 = ~x789 & n29294 ;
  assign n29307 = ( n16519 & ~n29305 ) | ( n16519 & n29306 ) | ( ~n29305 & n29306 ) ;
  assign n29308 = n29305 | n29307 ;
  assign n29309 = n16337 & n29109 ;
  assign n29310 = n16338 & n29108 ;
  assign n29311 = n29309 | n29310 ;
  assign n29312 = n19046 & n29177 ;
  assign n29313 = ( x792 & n29311 ) | ( x792 & n29312 ) | ( n29311 & n29312 ) ;
  assign n29314 = n29312 ^ n29311 ^ 1'b0 ;
  assign n29315 = ( x792 & n29313 ) | ( x792 & n29314 ) | ( n29313 & n29314 ) ;
  assign n29316 = n16459 & ~n29104 ;
  assign n29317 = ~x626 & n29072 ;
  assign n29318 = x626 & n29175 ;
  assign n29319 = ( n22317 & n29317 ) | ( n22317 & ~n29318 ) | ( n29317 & ~n29318 ) ;
  assign n29320 = ~n29317 & n29319 ;
  assign n29321 = ~x626 & n29175 ;
  assign n29322 = x626 & n29072 ;
  assign n29323 = ( n22322 & n29321 ) | ( n22322 & ~n29322 ) | ( n29321 & ~n29322 ) ;
  assign n29324 = ~n29321 & n29323 ;
  assign n29325 = ( ~n29316 & n29320 ) | ( ~n29316 & n29324 ) | ( n29320 & n29324 ) ;
  assign n29326 = n29316 | n29325 ;
  assign n29327 = ( x788 & ~n22314 ) | ( x788 & n29326 ) | ( ~n22314 & n29326 ) ;
  assign n29328 = ( n18482 & n22314 ) | ( n18482 & n29327 ) | ( n22314 & n29327 ) ;
  assign n29329 = ~n29315 & n29328 ;
  assign n29330 = ( n29308 & n29315 ) | ( n29308 & ~n29329 ) | ( n29315 & ~n29329 ) ;
  assign n29331 = ( ~n18484 & n29201 ) | ( ~n18484 & n29330 ) | ( n29201 & n29330 ) ;
  assign n29332 = n29201 ^ n18484 ^ 1'b0 ;
  assign n29333 = ( n29201 & n29331 ) | ( n29201 & ~n29332 ) | ( n29331 & ~n29332 ) ;
  assign n29334 = x644 | n29184 ;
  assign n29335 = x644 & n29189 ;
  assign n29336 = x790 & ~n29335 ;
  assign n29337 = n29334 & n29336 ;
  assign n29338 = ( ~n29194 & n29333 ) | ( ~n29194 & n29337 ) | ( n29333 & n29337 ) ;
  assign n29339 = ~n29194 & n29338 ;
  assign n29340 = ( x57 & n5193 ) | ( x57 & ~n29339 ) | ( n5193 & ~n29339 ) ;
  assign n29341 = n29339 | n29340 ;
  assign n29342 = x191 | n1611 ;
  assign n29343 = ~n29206 & n29342 ;
  assign n29344 = n16397 | n29343 ;
  assign n29345 = ~n15662 & n29206 ;
  assign n29346 = ~x1155 & n29342 ;
  assign n29347 = ~n29345 & n29346 ;
  assign n29348 = ( x1155 & n29344 ) | ( x1155 & n29345 ) | ( n29344 & n29345 ) ;
  assign n29349 = n29347 | n29348 ;
  assign n29350 = n29344 ^ x785 ^ 1'b0 ;
  assign n29351 = ( n29344 & n29349 ) | ( n29344 & n29350 ) | ( n29349 & n29350 ) ;
  assign n29352 = n16411 | n29351 ;
  assign n29353 = x1154 & n29352 ;
  assign n29354 = n16414 | n29351 ;
  assign n29355 = ~x1154 & n29354 ;
  assign n29356 = n29353 | n29355 ;
  assign n29357 = n29351 ^ x781 ^ 1'b0 ;
  assign n29358 = ( n29351 & n29356 ) | ( n29351 & n29357 ) | ( n29356 & n29357 ) ;
  assign n29359 = n21437 | n29358 ;
  assign n29360 = x1159 & n29359 ;
  assign n29361 = n21440 | n29358 ;
  assign n29362 = ~x1159 & n29361 ;
  assign n29363 = n29360 | n29362 ;
  assign n29364 = n29358 ^ x789 ^ 1'b0 ;
  assign n29365 = ( n29358 & n29363 ) | ( n29358 & n29364 ) | ( n29363 & n29364 ) ;
  assign n29366 = n29342 ^ n16518 ^ 1'b0 ;
  assign n29367 = ( n29342 & n29365 ) | ( n29342 & ~n29366 ) | ( n29365 & ~n29366 ) ;
  assign n29368 = n29342 ^ n16339 ^ 1'b0 ;
  assign n29369 = ( n29342 & n29367 ) | ( n29342 & ~n29368 ) | ( n29367 & ~n29368 ) ;
  assign n29370 = n19055 & n29369 ;
  assign n29371 = x647 & ~n29342 ;
  assign n29372 = x1157 | n29371 ;
  assign n29373 = x729 & n15778 ;
  assign n29374 = ~x625 & n29373 ;
  assign n29375 = ~x1153 & n29342 ;
  assign n29376 = ~n29374 & n29375 ;
  assign n29377 = x778 & ~n29376 ;
  assign n29378 = n29342 & ~n29373 ;
  assign n29379 = ( x1153 & n29374 ) | ( x1153 & n29378 ) | ( n29374 & n29378 ) ;
  assign n29380 = n29377 & ~n29379 ;
  assign n29381 = ( x778 & n29378 ) | ( x778 & ~n29380 ) | ( n29378 & ~n29380 ) ;
  assign n29382 = ~n29380 & n29381 ;
  assign n29383 = n16447 | n29382 ;
  assign n29384 = n16449 | n29383 ;
  assign n29385 = n16451 | n29384 ;
  assign n29386 = n16530 | n29385 ;
  assign n29387 = n16560 | n29386 ;
  assign n29388 = ( x647 & ~n29372 ) | ( x647 & n29387 ) | ( ~n29372 & n29387 ) ;
  assign n29389 = ~n29372 & n29388 ;
  assign n29390 = n29342 ^ x647 ^ 1'b0 ;
  assign n29391 = ( n29342 & n29387 ) | ( n29342 & n29390 ) | ( n29387 & n29390 ) ;
  assign n29392 = x1157 & n29391 ;
  assign n29393 = ( n16375 & n29389 ) | ( n16375 & n29392 ) | ( n29389 & n29392 ) ;
  assign n29394 = ( x787 & n29370 ) | ( x787 & n29393 ) | ( n29370 & n29393 ) ;
  assign n29395 = n29393 ^ n29370 ^ 1'b0 ;
  assign n29396 = ( x787 & n29394 ) | ( x787 & n29395 ) | ( n29394 & n29395 ) ;
  assign n29397 = ~x626 & n29342 ;
  assign n29398 = x626 & n29365 ;
  assign n29399 = ( n22317 & n29397 ) | ( n22317 & ~n29398 ) | ( n29397 & ~n29398 ) ;
  assign n29400 = ~n29397 & n29399 ;
  assign n29401 = ~x626 & n29365 ;
  assign n29402 = x626 & n29342 ;
  assign n29403 = ( n22322 & n29401 ) | ( n22322 & ~n29402 ) | ( n29401 & ~n29402 ) ;
  assign n29404 = ~n29401 & n29403 ;
  assign n29405 = n29385 & ~n29404 ;
  assign n29406 = ( n16459 & n29404 ) | ( n16459 & ~n29405 ) | ( n29404 & ~n29405 ) ;
  assign n29407 = ( x788 & n29400 ) | ( x788 & n29406 ) | ( n29400 & n29406 ) ;
  assign n29408 = n29406 ^ n29400 ^ 1'b0 ;
  assign n29409 = ( x788 & n29407 ) | ( x788 & n29408 ) | ( n29407 & n29408 ) ;
  assign n29410 = n15524 | n29378 ;
  assign n29411 = n29343 & n29410 ;
  assign n29412 = x625 & ~n29410 ;
  assign n29413 = ( n29375 & n29411 ) | ( n29375 & n29412 ) | ( n29411 & n29412 ) ;
  assign n29414 = ( x608 & n29379 ) | ( x608 & ~n29413 ) | ( n29379 & ~n29413 ) ;
  assign n29415 = n29413 | n29414 ;
  assign n29416 = x1153 & n29343 ;
  assign n29417 = ~n29412 & n29416 ;
  assign n29418 = x608 & ~n29376 ;
  assign n29419 = n29415 & ~n29418 ;
  assign n29420 = ( n29415 & n29417 ) | ( n29415 & n29419 ) | ( n29417 & n29419 ) ;
  assign n29421 = n29411 ^ x778 ^ 1'b0 ;
  assign n29422 = ( n29411 & n29420 ) | ( n29411 & n29421 ) | ( n29420 & n29421 ) ;
  assign n29423 = x609 & ~n29422 ;
  assign n29429 = x609 | n29382 ;
  assign n29430 = ( x1155 & n29423 ) | ( x1155 & n29429 ) | ( n29423 & n29429 ) ;
  assign n29431 = ~n29423 & n29430 ;
  assign n29432 = ( x660 & n29347 ) | ( x660 & ~n29431 ) | ( n29347 & ~n29431 ) ;
  assign n29433 = ~n29347 & n29432 ;
  assign n29424 = x609 & ~n29382 ;
  assign n29425 = x1155 | n29424 ;
  assign n29426 = ( n29422 & n29423 ) | ( n29422 & ~n29425 ) | ( n29423 & ~n29425 ) ;
  assign n29427 = ( x660 & n29348 ) | ( x660 & ~n29426 ) | ( n29348 & ~n29426 ) ;
  assign n29428 = n29426 | n29427 ;
  assign n29434 = n29433 ^ n29428 ^ 1'b0 ;
  assign n29435 = ( x785 & ~n29428 ) | ( x785 & n29433 ) | ( ~n29428 & n29433 ) ;
  assign n29436 = ( x785 & ~n29434 ) | ( x785 & n29435 ) | ( ~n29434 & n29435 ) ;
  assign n29437 = ( x785 & n29422 ) | ( x785 & ~n29436 ) | ( n29422 & ~n29436 ) ;
  assign n29438 = ~n29436 & n29437 ;
  assign n29439 = x618 & ~n29438 ;
  assign n29440 = x618 | n29383 ;
  assign n29441 = ( x1154 & n29439 ) | ( x1154 & n29440 ) | ( n29439 & n29440 ) ;
  assign n29442 = ~n29439 & n29441 ;
  assign n29443 = ( x627 & n29355 ) | ( x627 & ~n29442 ) | ( n29355 & ~n29442 ) ;
  assign n29444 = ~n29355 & n29443 ;
  assign n29445 = x627 | n29353 ;
  assign n29446 = x618 & ~n29383 ;
  assign n29447 = x1154 | n29446 ;
  assign n29448 = ( n29438 & n29439 ) | ( n29438 & ~n29447 ) | ( n29439 & ~n29447 ) ;
  assign n29449 = ( ~n29444 & n29445 ) | ( ~n29444 & n29448 ) | ( n29445 & n29448 ) ;
  assign n29450 = ~n29444 & n29449 ;
  assign n29451 = n29438 ^ x781 ^ 1'b0 ;
  assign n29452 = ( n29438 & n29450 ) | ( n29438 & n29451 ) | ( n29450 & n29451 ) ;
  assign n29453 = ~x789 & n29452 ;
  assign n29454 = x619 & ~n29384 ;
  assign n29455 = x1159 | n29454 ;
  assign n29456 = x619 & ~n29452 ;
  assign n29457 = ( n29452 & ~n29455 ) | ( n29452 & n29456 ) | ( ~n29455 & n29456 ) ;
  assign n29458 = ( x648 & n29360 ) | ( x648 & ~n29457 ) | ( n29360 & ~n29457 ) ;
  assign n29459 = n29457 | n29458 ;
  assign n29460 = x619 | n29384 ;
  assign n29461 = x1159 & ~n29456 ;
  assign n29462 = n29460 & n29461 ;
  assign n29463 = ( x648 & n29362 ) | ( x648 & ~n29462 ) | ( n29362 & ~n29462 ) ;
  assign n29464 = ~n29362 & n29463 ;
  assign n29465 = x789 & ~n29464 ;
  assign n29466 = n29459 & n29465 ;
  assign n29467 = ( n16519 & ~n29453 ) | ( n16519 & n29466 ) | ( ~n29453 & n29466 ) ;
  assign n29468 = n29453 | n29467 ;
  assign n29469 = n29468 ^ n29409 ^ 1'b0 ;
  assign n29470 = ( n29409 & n29468 ) | ( n29409 & n29469 ) | ( n29468 & n29469 ) ;
  assign n29471 = ( n18482 & ~n29409 ) | ( n18482 & n29470 ) | ( ~n29409 & n29470 ) ;
  assign n29472 = n19208 | n29386 ;
  assign n29473 = n16556 & ~n29367 ;
  assign n29474 = x629 & ~n29473 ;
  assign n29475 = n29472 & n29474 ;
  assign n29476 = n16557 & ~n29367 ;
  assign n29477 = n19212 & ~n29386 ;
  assign n29478 = n29476 | n29477 ;
  assign n29479 = ( x629 & ~n29475 ) | ( x629 & n29478 ) | ( ~n29475 & n29478 ) ;
  assign n29480 = ~n29475 & n29479 ;
  assign n29481 = ( x792 & ~n19206 ) | ( x792 & n29480 ) | ( ~n19206 & n29480 ) ;
  assign n29482 = ( n18484 & n19206 ) | ( n18484 & n29481 ) | ( n19206 & n29481 ) ;
  assign n29483 = ( n29396 & n29471 ) | ( n29396 & ~n29482 ) | ( n29471 & ~n29482 ) ;
  assign n29484 = n29483 ^ n29471 ^ 1'b0 ;
  assign n29485 = ( n29396 & n29483 ) | ( n29396 & ~n29484 ) | ( n29483 & ~n29484 ) ;
  assign n29486 = x790 | n29485 ;
  assign n29487 = x644 & ~n29485 ;
  assign n29488 = ( x787 & n29389 ) | ( x787 & ~n29392 ) | ( n29389 & ~n29392 ) ;
  assign n29489 = ~n29389 & n29488 ;
  assign n29490 = ( x787 & n29387 ) | ( x787 & ~n29489 ) | ( n29387 & ~n29489 ) ;
  assign n29491 = ~n29489 & n29490 ;
  assign n29492 = x644 | n29491 ;
  assign n29493 = ( x715 & n29487 ) | ( x715 & n29492 ) | ( n29487 & n29492 ) ;
  assign n29494 = ~n29487 & n29493 ;
  assign n29495 = x644 | n29342 ;
  assign n29496 = n29342 ^ n16376 ^ 1'b0 ;
  assign n29497 = ( n29342 & n29369 ) | ( n29342 & ~n29496 ) | ( n29369 & ~n29496 ) ;
  assign n29498 = x644 & ~n29497 ;
  assign n29499 = ( x715 & n29495 ) | ( x715 & ~n29498 ) | ( n29495 & ~n29498 ) ;
  assign n29500 = ~x715 & n29499 ;
  assign n29501 = ( x1160 & n29494 ) | ( x1160 & ~n29500 ) | ( n29494 & ~n29500 ) ;
  assign n29502 = ~n29494 & n29501 ;
  assign n29503 = x644 & ~n29342 ;
  assign n29504 = x715 & ~n29503 ;
  assign n29505 = ( n29497 & n29498 ) | ( n29497 & n29504 ) | ( n29498 & n29504 ) ;
  assign n29506 = x644 & ~n29491 ;
  assign n29507 = x715 | n29506 ;
  assign n29508 = ( n29485 & n29487 ) | ( n29485 & ~n29507 ) | ( n29487 & ~n29507 ) ;
  assign n29509 = ( x1160 & ~n29505 ) | ( x1160 & n29508 ) | ( ~n29505 & n29508 ) ;
  assign n29510 = n29505 | n29509 ;
  assign n29511 = x790 & ~n29510 ;
  assign n29512 = ( x790 & n29502 ) | ( x790 & n29511 ) | ( n29502 & n29511 ) ;
  assign n29513 = x832 & ~n29512 ;
  assign n29514 = n29486 & n29513 ;
  assign n29515 = ~x191 & n7318 ;
  assign n29516 = x832 | n29515 ;
  assign n29517 = ~n29514 & n29516 ;
  assign n29518 = ( n29341 & n29514 ) | ( n29341 & ~n29517 ) | ( n29514 & ~n29517 ) ;
  assign n29519 = x192 | n15656 ;
  assign n29520 = x192 | n15644 ;
  assign n29521 = n16185 & n29520 ;
  assign n29522 = x192 | n16697 ;
  assign n29523 = x192 & n16699 ;
  assign n29524 = ( x38 & n29522 ) | ( x38 & ~n29523 ) | ( n29522 & ~n29523 ) ;
  assign n29525 = ~x38 & n29524 ;
  assign n29526 = ( x691 & n29521 ) | ( x691 & ~n29525 ) | ( n29521 & ~n29525 ) ;
  assign n29527 = ~n29521 & n29526 ;
  assign n29528 = x192 | x691 ;
  assign n29529 = n15655 | n29528 ;
  assign n29530 = ( n2069 & ~n29527 ) | ( n2069 & n29529 ) | ( ~n29527 & n29529 ) ;
  assign n29531 = ~n2069 & n29530 ;
  assign n29532 = n29531 ^ x192 ^ 1'b0 ;
  assign n29533 = ( ~x192 & n2069 ) | ( ~x192 & n29532 ) | ( n2069 & n29532 ) ;
  assign n29534 = ( x192 & n29531 ) | ( x192 & n29533 ) | ( n29531 & n29533 ) ;
  assign n29535 = x625 & ~n29534 ;
  assign n29536 = x625 | n29519 ;
  assign n29537 = ( x1153 & n29535 ) | ( x1153 & n29536 ) | ( n29535 & n29536 ) ;
  assign n29538 = ~n29535 & n29537 ;
  assign n29539 = x625 & ~n29519 ;
  assign n29540 = x1153 | n29539 ;
  assign n29541 = ( x625 & n29534 ) | ( x625 & ~n29540 ) | ( n29534 & ~n29540 ) ;
  assign n29542 = ~n29540 & n29541 ;
  assign n29543 = n29538 | n29542 ;
  assign n29544 = n29534 ^ x778 ^ 1'b0 ;
  assign n29545 = ( n29534 & n29543 ) | ( n29534 & n29544 ) | ( n29543 & n29544 ) ;
  assign n29546 = n29519 ^ n16234 ^ 1'b0 ;
  assign n29547 = ( n29519 & n29545 ) | ( n29519 & ~n29546 ) | ( n29545 & ~n29546 ) ;
  assign n29548 = n29519 ^ n16254 ^ 1'b0 ;
  assign n29549 = ( n29519 & n29547 ) | ( n29519 & ~n29548 ) | ( n29547 & ~n29548 ) ;
  assign n29550 = n29519 ^ n16279 ^ 1'b0 ;
  assign n29551 = ( n29519 & n29549 ) | ( n29519 & ~n29550 ) | ( n29549 & ~n29550 ) ;
  assign n29552 = n29519 ^ n16318 ^ 1'b0 ;
  assign n29553 = ( n29519 & n29551 ) | ( n29519 & ~n29552 ) | ( n29551 & ~n29552 ) ;
  assign n29554 = n29519 ^ x628 ^ 1'b0 ;
  assign n29555 = ( n29519 & n29553 ) | ( n29519 & ~n29554 ) | ( n29553 & ~n29554 ) ;
  assign n29556 = ( n29519 & n29553 ) | ( n29519 & n29554 ) | ( n29553 & n29554 ) ;
  assign n29557 = n29555 ^ x1156 ^ 1'b0 ;
  assign n29558 = ( n29555 & n29556 ) | ( n29555 & n29557 ) | ( n29556 & n29557 ) ;
  assign n29559 = n29553 ^ x792 ^ 1'b0 ;
  assign n29560 = ( n29553 & n29558 ) | ( n29553 & n29559 ) | ( n29558 & n29559 ) ;
  assign n29561 = n29519 ^ x647 ^ 1'b0 ;
  assign n29562 = ( n29519 & n29560 ) | ( n29519 & ~n29561 ) | ( n29560 & ~n29561 ) ;
  assign n29563 = ( n29519 & n29560 ) | ( n29519 & n29561 ) | ( n29560 & n29561 ) ;
  assign n29564 = n29562 ^ x1157 ^ 1'b0 ;
  assign n29565 = ( n29562 & n29563 ) | ( n29562 & n29564 ) | ( n29563 & n29564 ) ;
  assign n29566 = n29560 ^ x787 ^ 1'b0 ;
  assign n29567 = ( n29560 & n29565 ) | ( n29560 & n29566 ) | ( n29565 & n29566 ) ;
  assign n29568 = x644 & ~n29567 ;
  assign n29569 = x715 | n29568 ;
  assign n29570 = x644 & ~n29519 ;
  assign n29571 = x715 & ~n29570 ;
  assign n29572 = n29571 ^ x1160 ^ 1'b0 ;
  assign n29573 = x192 & n2069 ;
  assign n29574 = x38 & n29520 ;
  assign n29575 = ~x192 & x764 ;
  assign n29576 = n15587 & n29575 ;
  assign n29577 = x764 & n15639 ;
  assign n29578 = x192 & ~n29577 ;
  assign n29579 = ( n21038 & ~n29576 ) | ( n21038 & n29578 ) | ( ~n29576 & n29578 ) ;
  assign n29580 = n29576 | n29579 ;
  assign n29581 = x192 & ~n15631 ;
  assign n29582 = ~x764 & n15486 ;
  assign n29583 = ( x39 & n29581 ) | ( x39 & n29582 ) | ( n29581 & n29582 ) ;
  assign n29584 = n29582 ^ n29581 ^ 1'b0 ;
  assign n29585 = ( x39 & n29583 ) | ( x39 & n29584 ) | ( n29583 & n29584 ) ;
  assign n29586 = ( ~x38 & n29580 ) | ( ~x38 & n29585 ) | ( n29580 & n29585 ) ;
  assign n29587 = ~x38 & n29586 ;
  assign n29588 = x764 & n15646 ;
  assign n29589 = ~n29587 & n29588 ;
  assign n29590 = ( n29574 & n29587 ) | ( n29574 & ~n29589 ) | ( n29587 & ~n29589 ) ;
  assign n29591 = ~n2069 & n29590 ;
  assign n29592 = n29573 | n29591 ;
  assign n29593 = n29519 ^ n15659 ^ 1'b0 ;
  assign n29594 = ( n29519 & n29592 ) | ( n29519 & ~n29593 ) | ( n29592 & ~n29593 ) ;
  assign n29595 = n15662 & n29519 ;
  assign n29596 = ( ~n15662 & n29573 ) | ( ~n15662 & n29591 ) | ( n29573 & n29591 ) ;
  assign n29597 = n29595 | n29596 ;
  assign n29598 = n29597 ^ n29594 ^ n29519 ;
  assign n29599 = n29598 ^ x1155 ^ 1'b0 ;
  assign n29600 = ( n29597 & n29598 ) | ( n29597 & ~n29599 ) | ( n29598 & ~n29599 ) ;
  assign n29601 = n29594 ^ x785 ^ 1'b0 ;
  assign n29602 = ( n29594 & n29600 ) | ( n29594 & n29601 ) | ( n29600 & n29601 ) ;
  assign n29603 = x618 & ~n29602 ;
  assign n29604 = x618 | n29519 ;
  assign n29605 = ( x1154 & n29603 ) | ( x1154 & n29604 ) | ( n29603 & n29604 ) ;
  assign n29606 = ~n29603 & n29605 ;
  assign n29607 = x618 & ~n29519 ;
  assign n29608 = x1154 | n29607 ;
  assign n29609 = ( n29602 & n29603 ) | ( n29602 & ~n29608 ) | ( n29603 & ~n29608 ) ;
  assign n29610 = n29606 | n29609 ;
  assign n29611 = n29602 ^ x781 ^ 1'b0 ;
  assign n29612 = ( n29602 & n29610 ) | ( n29602 & n29611 ) | ( n29610 & n29611 ) ;
  assign n29613 = x619 | n29519 ;
  assign n29614 = x619 & ~n29612 ;
  assign n29615 = x1159 & ~n29614 ;
  assign n29616 = n29613 & n29615 ;
  assign n29617 = x619 & ~n29519 ;
  assign n29618 = x1159 | n29617 ;
  assign n29619 = ( n29612 & n29614 ) | ( n29612 & ~n29618 ) | ( n29614 & ~n29618 ) ;
  assign n29620 = n29616 | n29619 ;
  assign n29621 = n29612 ^ x789 ^ 1'b0 ;
  assign n29622 = ( n29612 & n29620 ) | ( n29612 & n29621 ) | ( n29620 & n29621 ) ;
  assign n29623 = n29519 ^ n16518 ^ 1'b0 ;
  assign n29624 = ( n29519 & n29622 ) | ( n29519 & ~n29623 ) | ( n29622 & ~n29623 ) ;
  assign n29625 = n29519 ^ n16339 ^ 1'b0 ;
  assign n29626 = ( n29519 & n29624 ) | ( n29519 & ~n29625 ) | ( n29624 & ~n29625 ) ;
  assign n29627 = n29519 ^ n16376 ^ 1'b0 ;
  assign n29628 = ( n29519 & n29626 ) | ( n29519 & ~n29627 ) | ( n29626 & ~n29627 ) ;
  assign n29629 = x644 | n29628 ;
  assign n29630 = ( n29571 & ~n29572 ) | ( n29571 & n29629 ) | ( ~n29572 & n29629 ) ;
  assign n29631 = ( x1160 & n29572 ) | ( x1160 & n29630 ) | ( n29572 & n29630 ) ;
  assign n29632 = n29569 & ~n29631 ;
  assign n29633 = x644 & ~n29628 ;
  assign n29634 = ( ~x715 & n29519 ) | ( ~x715 & n29570 ) | ( n29519 & n29570 ) ;
  assign n29635 = x1160 & ~n29634 ;
  assign n29636 = ( x1160 & n29633 ) | ( x1160 & n29635 ) | ( n29633 & n29635 ) ;
  assign n29637 = ( x715 & n29567 ) | ( x715 & n29568 ) | ( n29567 & n29568 ) ;
  assign n29638 = n29636 & ~n29637 ;
  assign n29639 = ( x790 & n29632 ) | ( x790 & n29638 ) | ( n29632 & n29638 ) ;
  assign n29640 = n29638 ^ n29632 ^ 1'b0 ;
  assign n29641 = ( x790 & n29639 ) | ( x790 & n29640 ) | ( n29639 & n29640 ) ;
  assign n29642 = n16374 & n29562 ;
  assign n29643 = n19055 & n29626 ;
  assign n29644 = n29642 | n29643 ;
  assign n29645 = n16373 & n29563 ;
  assign n29646 = ( x787 & n29644 ) | ( x787 & n29645 ) | ( n29644 & n29645 ) ;
  assign n29647 = n29645 ^ n29644 ^ 1'b0 ;
  assign n29648 = ( x787 & n29646 ) | ( x787 & n29647 ) | ( n29646 & n29647 ) ;
  assign n29649 = x619 & ~n29549 ;
  assign n29650 = x1159 | n29649 ;
  assign n29698 = x625 | n29592 ;
  assign n29652 = x691 | n29590 ;
  assign n29653 = x764 & n15591 ;
  assign n29654 = n17156 | n29653 ;
  assign n29655 = x192 & ~n5017 ;
  assign n29656 = n29654 & n29655 ;
  assign n29657 = ~x764 & n22207 ;
  assign n29658 = n15968 | n29657 ;
  assign n29659 = x39 | n29658 ;
  assign n29660 = ( ~x39 & x192 ) | ( ~x39 & n29659 ) | ( x192 & n29659 ) ;
  assign n29661 = ( x38 & n29656 ) | ( x38 & n29660 ) | ( n29656 & n29660 ) ;
  assign n29662 = ~n29656 & n29661 ;
  assign n29663 = x192 & n15795 ;
  assign n29664 = x764 | n29663 ;
  assign n29665 = ( x192 & n15876 ) | ( x192 & ~n29664 ) | ( n15876 & ~n29664 ) ;
  assign n29666 = ~n29664 & n29665 ;
  assign n29667 = x192 | n16003 ;
  assign n29668 = x192 & n15943 ;
  assign n29669 = x764 & ~n29668 ;
  assign n29670 = n29667 & n29669 ;
  assign n29671 = ( x39 & n29666 ) | ( x39 & ~n29670 ) | ( n29666 & ~n29670 ) ;
  assign n29672 = ~n29666 & n29671 ;
  assign n29673 = x192 & n16054 ;
  assign n29674 = x192 | n16048 ;
  assign n29675 = ( x764 & n29673 ) | ( x764 & n29674 ) | ( n29673 & n29674 ) ;
  assign n29676 = ~n29673 & n29675 ;
  assign n29677 = x192 | n16044 ;
  assign n29678 = x192 & n16029 ;
  assign n29679 = ( x764 & n29677 ) | ( x764 & ~n29678 ) | ( n29677 & ~n29678 ) ;
  assign n29680 = ~x764 & n29679 ;
  assign n29681 = ( x39 & ~n29676 ) | ( x39 & n29680 ) | ( ~n29676 & n29680 ) ;
  assign n29682 = n29676 | n29681 ;
  assign n29683 = ( x38 & ~n29672 ) | ( x38 & n29682 ) | ( ~n29672 & n29682 ) ;
  assign n29684 = ~x38 & n29683 ;
  assign n29685 = ( x691 & n29662 ) | ( x691 & ~n29684 ) | ( n29662 & ~n29684 ) ;
  assign n29686 = ~n29662 & n29685 ;
  assign n29687 = ( n2051 & n2068 ) | ( n2051 & ~n29686 ) | ( n2068 & ~n29686 ) ;
  assign n29688 = n29686 | n29687 ;
  assign n29689 = ( n29573 & n29652 ) | ( n29573 & ~n29688 ) | ( n29652 & ~n29688 ) ;
  assign n29690 = n29689 ^ n29652 ^ 1'b0 ;
  assign n29691 = ( n29573 & n29689 ) | ( n29573 & ~n29690 ) | ( n29689 & ~n29690 ) ;
  assign n29699 = x625 & ~n29691 ;
  assign n29700 = x1153 & ~n29699 ;
  assign n29701 = n29698 & n29700 ;
  assign n29702 = ( x608 & n29542 ) | ( x608 & ~n29701 ) | ( n29542 & ~n29701 ) ;
  assign n29703 = ~n29542 & n29702 ;
  assign n29692 = x625 | n29691 ;
  assign n29693 = x625 & ~n29592 ;
  assign n29694 = ( x1153 & n29692 ) | ( x1153 & ~n29693 ) | ( n29692 & ~n29693 ) ;
  assign n29695 = ~x1153 & n29694 ;
  assign n29696 = ( x608 & n29538 ) | ( x608 & ~n29695 ) | ( n29538 & ~n29695 ) ;
  assign n29697 = n29695 | n29696 ;
  assign n29704 = n29703 ^ n29697 ^ 1'b0 ;
  assign n29705 = ( x778 & ~n29697 ) | ( x778 & n29703 ) | ( ~n29697 & n29703 ) ;
  assign n29706 = ( x778 & ~n29704 ) | ( x778 & n29705 ) | ( ~n29704 & n29705 ) ;
  assign n29707 = ( x778 & n29691 ) | ( x778 & ~n29706 ) | ( n29691 & ~n29706 ) ;
  assign n29708 = ~n29706 & n29707 ;
  assign n29709 = x609 & ~n29708 ;
  assign n29715 = x609 | n29545 ;
  assign n29716 = ( x1155 & n29709 ) | ( x1155 & n29715 ) | ( n29709 & n29715 ) ;
  assign n29717 = ~n29709 & n29716 ;
  assign n29718 = ~x1155 & n29597 ;
  assign n29719 = ( x660 & n29717 ) | ( x660 & ~n29718 ) | ( n29717 & ~n29718 ) ;
  assign n29720 = ~n29717 & n29719 ;
  assign n29651 = x1155 & n29598 ;
  assign n29710 = x609 & ~n29545 ;
  assign n29711 = x1155 | n29710 ;
  assign n29712 = ( n29708 & n29709 ) | ( n29708 & ~n29711 ) | ( n29709 & ~n29711 ) ;
  assign n29713 = ( x660 & ~n29651 ) | ( x660 & n29712 ) | ( ~n29651 & n29712 ) ;
  assign n29714 = n29651 | n29713 ;
  assign n29721 = n29720 ^ n29714 ^ 1'b0 ;
  assign n29722 = ( x785 & ~n29714 ) | ( x785 & n29720 ) | ( ~n29714 & n29720 ) ;
  assign n29723 = ( x785 & ~n29721 ) | ( x785 & n29722 ) | ( ~n29721 & n29722 ) ;
  assign n29724 = ( x785 & n29708 ) | ( x785 & ~n29723 ) | ( n29708 & ~n29723 ) ;
  assign n29725 = ~n29723 & n29724 ;
  assign n29726 = x618 & ~n29725 ;
  assign n29732 = x618 | n29547 ;
  assign n29733 = ( x1154 & n29726 ) | ( x1154 & n29732 ) | ( n29726 & n29732 ) ;
  assign n29734 = ~n29726 & n29733 ;
  assign n29735 = ( x627 & n29609 ) | ( x627 & ~n29734 ) | ( n29609 & ~n29734 ) ;
  assign n29736 = ~n29609 & n29735 ;
  assign n29727 = x618 & ~n29547 ;
  assign n29728 = x1154 | n29727 ;
  assign n29729 = ( n29725 & n29726 ) | ( n29725 & ~n29728 ) | ( n29726 & ~n29728 ) ;
  assign n29730 = ( x627 & n29606 ) | ( x627 & ~n29729 ) | ( n29606 & ~n29729 ) ;
  assign n29731 = n29729 | n29730 ;
  assign n29737 = n29736 ^ n29731 ^ 1'b0 ;
  assign n29738 = ( x781 & ~n29731 ) | ( x781 & n29736 ) | ( ~n29731 & n29736 ) ;
  assign n29739 = ( x781 & ~n29737 ) | ( x781 & n29738 ) | ( ~n29737 & n29738 ) ;
  assign n29740 = ( x781 & n29725 ) | ( x781 & ~n29739 ) | ( n29725 & ~n29739 ) ;
  assign n29741 = ~n29739 & n29740 ;
  assign n29742 = x619 & ~n29741 ;
  assign n29743 = ( ~n29650 & n29741 ) | ( ~n29650 & n29742 ) | ( n29741 & n29742 ) ;
  assign n29744 = ( x648 & n29616 ) | ( x648 & ~n29743 ) | ( n29616 & ~n29743 ) ;
  assign n29745 = n29743 | n29744 ;
  assign n29746 = x619 | n29549 ;
  assign n29747 = x1159 & ~n29742 ;
  assign n29748 = n29746 & n29747 ;
  assign n29749 = ( x648 & n29619 ) | ( x648 & ~n29748 ) | ( n29619 & ~n29748 ) ;
  assign n29750 = ~n29619 & n29749 ;
  assign n29751 = x789 & ~n29750 ;
  assign n29752 = n29745 & n29751 ;
  assign n29753 = ~x789 & n29741 ;
  assign n29754 = ( n16519 & ~n29752 ) | ( n16519 & n29753 ) | ( ~n29752 & n29753 ) ;
  assign n29755 = n29752 | n29754 ;
  assign n29756 = n16337 & n29556 ;
  assign n29757 = n16338 & n29555 ;
  assign n29758 = n29756 | n29757 ;
  assign n29759 = n19046 & n29624 ;
  assign n29760 = ( x792 & n29758 ) | ( x792 & n29759 ) | ( n29758 & n29759 ) ;
  assign n29761 = n29759 ^ n29758 ^ 1'b0 ;
  assign n29762 = ( x792 & n29760 ) | ( x792 & n29761 ) | ( n29760 & n29761 ) ;
  assign n29763 = n16459 & ~n29551 ;
  assign n29764 = ~x626 & n29519 ;
  assign n29765 = x626 & n29622 ;
  assign n29766 = ( n22317 & n29764 ) | ( n22317 & ~n29765 ) | ( n29764 & ~n29765 ) ;
  assign n29767 = ~n29764 & n29766 ;
  assign n29768 = ~x626 & n29622 ;
  assign n29769 = x626 & n29519 ;
  assign n29770 = ( n22322 & n29768 ) | ( n22322 & ~n29769 ) | ( n29768 & ~n29769 ) ;
  assign n29771 = ~n29768 & n29770 ;
  assign n29772 = ( ~n29763 & n29767 ) | ( ~n29763 & n29771 ) | ( n29767 & n29771 ) ;
  assign n29773 = n29763 | n29772 ;
  assign n29774 = ( x788 & ~n22314 ) | ( x788 & n29773 ) | ( ~n22314 & n29773 ) ;
  assign n29775 = ( n18482 & n22314 ) | ( n18482 & n29774 ) | ( n22314 & n29774 ) ;
  assign n29776 = ~n29762 & n29775 ;
  assign n29777 = ( n29755 & n29762 ) | ( n29755 & ~n29776 ) | ( n29762 & ~n29776 ) ;
  assign n29778 = ( ~n18484 & n29648 ) | ( ~n18484 & n29777 ) | ( n29648 & n29777 ) ;
  assign n29779 = n29648 ^ n18484 ^ 1'b0 ;
  assign n29780 = ( n29648 & n29778 ) | ( n29648 & ~n29779 ) | ( n29778 & ~n29779 ) ;
  assign n29781 = x644 | n29631 ;
  assign n29782 = x644 & n29636 ;
  assign n29783 = x790 & ~n29782 ;
  assign n29784 = n29781 & n29783 ;
  assign n29785 = ( ~n29641 & n29780 ) | ( ~n29641 & n29784 ) | ( n29780 & n29784 ) ;
  assign n29786 = ~n29641 & n29785 ;
  assign n29787 = ( x57 & n5193 ) | ( x57 & ~n29786 ) | ( n5193 & ~n29786 ) ;
  assign n29788 = n29786 | n29787 ;
  assign n29789 = x192 | n1611 ;
  assign n29790 = ~n29653 & n29789 ;
  assign n29791 = n16397 | n29790 ;
  assign n29792 = ~n15662 & n29653 ;
  assign n29793 = ~x1155 & n29789 ;
  assign n29794 = ~n29792 & n29793 ;
  assign n29795 = ( x1155 & n29791 ) | ( x1155 & n29792 ) | ( n29791 & n29792 ) ;
  assign n29796 = n29794 | n29795 ;
  assign n29797 = n29791 ^ x785 ^ 1'b0 ;
  assign n29798 = ( n29791 & n29796 ) | ( n29791 & n29797 ) | ( n29796 & n29797 ) ;
  assign n29799 = n16411 | n29798 ;
  assign n29800 = x1154 & n29799 ;
  assign n29801 = n16414 | n29798 ;
  assign n29802 = ~x1154 & n29801 ;
  assign n29803 = n29800 | n29802 ;
  assign n29804 = n29798 ^ x781 ^ 1'b0 ;
  assign n29805 = ( n29798 & n29803 ) | ( n29798 & n29804 ) | ( n29803 & n29804 ) ;
  assign n29806 = n21437 | n29805 ;
  assign n29807 = x1159 & n29806 ;
  assign n29808 = n21440 | n29805 ;
  assign n29809 = ~x1159 & n29808 ;
  assign n29810 = n29807 | n29809 ;
  assign n29811 = n29805 ^ x789 ^ 1'b0 ;
  assign n29812 = ( n29805 & n29810 ) | ( n29805 & n29811 ) | ( n29810 & n29811 ) ;
  assign n29813 = n29789 ^ n16518 ^ 1'b0 ;
  assign n29814 = ( n29789 & n29812 ) | ( n29789 & ~n29813 ) | ( n29812 & ~n29813 ) ;
  assign n29815 = n29789 ^ n16339 ^ 1'b0 ;
  assign n29816 = ( n29789 & n29814 ) | ( n29789 & ~n29815 ) | ( n29814 & ~n29815 ) ;
  assign n29817 = n19055 & n29816 ;
  assign n29818 = x647 & ~n29789 ;
  assign n29819 = x1157 | n29818 ;
  assign n29820 = x691 & n15778 ;
  assign n29821 = ~x625 & n29820 ;
  assign n29822 = ~x1153 & n29789 ;
  assign n29823 = ~n29821 & n29822 ;
  assign n29824 = x778 & ~n29823 ;
  assign n29825 = n29789 & ~n29820 ;
  assign n29826 = ( x1153 & n29821 ) | ( x1153 & n29825 ) | ( n29821 & n29825 ) ;
  assign n29827 = n29824 & ~n29826 ;
  assign n29828 = ( x778 & n29825 ) | ( x778 & ~n29827 ) | ( n29825 & ~n29827 ) ;
  assign n29829 = ~n29827 & n29828 ;
  assign n29830 = n16447 | n29829 ;
  assign n29831 = n16449 | n29830 ;
  assign n29832 = n16451 | n29831 ;
  assign n29833 = n16530 | n29832 ;
  assign n29834 = n16560 | n29833 ;
  assign n29835 = ( x647 & ~n29819 ) | ( x647 & n29834 ) | ( ~n29819 & n29834 ) ;
  assign n29836 = ~n29819 & n29835 ;
  assign n29837 = n29789 ^ x647 ^ 1'b0 ;
  assign n29838 = ( n29789 & n29834 ) | ( n29789 & n29837 ) | ( n29834 & n29837 ) ;
  assign n29839 = x1157 & n29838 ;
  assign n29840 = ( n16375 & n29836 ) | ( n16375 & n29839 ) | ( n29836 & n29839 ) ;
  assign n29841 = ( x787 & n29817 ) | ( x787 & n29840 ) | ( n29817 & n29840 ) ;
  assign n29842 = n29840 ^ n29817 ^ 1'b0 ;
  assign n29843 = ( x787 & n29841 ) | ( x787 & n29842 ) | ( n29841 & n29842 ) ;
  assign n29844 = ~x626 & n29789 ;
  assign n29845 = x626 & n29812 ;
  assign n29846 = ( n22317 & n29844 ) | ( n22317 & ~n29845 ) | ( n29844 & ~n29845 ) ;
  assign n29847 = ~n29844 & n29846 ;
  assign n29848 = ~x626 & n29812 ;
  assign n29849 = x626 & n29789 ;
  assign n29850 = ( n22322 & n29848 ) | ( n22322 & ~n29849 ) | ( n29848 & ~n29849 ) ;
  assign n29851 = ~n29848 & n29850 ;
  assign n29852 = n29832 & ~n29851 ;
  assign n29853 = ( n16459 & n29851 ) | ( n16459 & ~n29852 ) | ( n29851 & ~n29852 ) ;
  assign n29854 = ( x788 & n29847 ) | ( x788 & n29853 ) | ( n29847 & n29853 ) ;
  assign n29855 = n29853 ^ n29847 ^ 1'b0 ;
  assign n29856 = ( x788 & n29854 ) | ( x788 & n29855 ) | ( n29854 & n29855 ) ;
  assign n29857 = n15524 | n29825 ;
  assign n29858 = n29790 & n29857 ;
  assign n29859 = x625 & ~n29857 ;
  assign n29860 = ( n29822 & n29858 ) | ( n29822 & n29859 ) | ( n29858 & n29859 ) ;
  assign n29861 = ( x608 & n29826 ) | ( x608 & ~n29860 ) | ( n29826 & ~n29860 ) ;
  assign n29862 = n29860 | n29861 ;
  assign n29863 = x1153 & n29790 ;
  assign n29864 = ~n29859 & n29863 ;
  assign n29865 = x608 & ~n29823 ;
  assign n29866 = n29862 & ~n29865 ;
  assign n29867 = ( n29862 & n29864 ) | ( n29862 & n29866 ) | ( n29864 & n29866 ) ;
  assign n29868 = n29858 ^ x778 ^ 1'b0 ;
  assign n29869 = ( n29858 & n29867 ) | ( n29858 & n29868 ) | ( n29867 & n29868 ) ;
  assign n29870 = x609 & ~n29869 ;
  assign n29876 = x609 | n29829 ;
  assign n29877 = ( x1155 & n29870 ) | ( x1155 & n29876 ) | ( n29870 & n29876 ) ;
  assign n29878 = ~n29870 & n29877 ;
  assign n29879 = ( x660 & n29794 ) | ( x660 & ~n29878 ) | ( n29794 & ~n29878 ) ;
  assign n29880 = ~n29794 & n29879 ;
  assign n29871 = x609 & ~n29829 ;
  assign n29872 = x1155 | n29871 ;
  assign n29873 = ( n29869 & n29870 ) | ( n29869 & ~n29872 ) | ( n29870 & ~n29872 ) ;
  assign n29874 = ( x660 & n29795 ) | ( x660 & ~n29873 ) | ( n29795 & ~n29873 ) ;
  assign n29875 = n29873 | n29874 ;
  assign n29881 = n29880 ^ n29875 ^ 1'b0 ;
  assign n29882 = ( x785 & ~n29875 ) | ( x785 & n29880 ) | ( ~n29875 & n29880 ) ;
  assign n29883 = ( x785 & ~n29881 ) | ( x785 & n29882 ) | ( ~n29881 & n29882 ) ;
  assign n29884 = ( x785 & n29869 ) | ( x785 & ~n29883 ) | ( n29869 & ~n29883 ) ;
  assign n29885 = ~n29883 & n29884 ;
  assign n29886 = x618 & ~n29885 ;
  assign n29887 = x618 | n29830 ;
  assign n29888 = ( x1154 & n29886 ) | ( x1154 & n29887 ) | ( n29886 & n29887 ) ;
  assign n29889 = ~n29886 & n29888 ;
  assign n29890 = ( x627 & n29802 ) | ( x627 & ~n29889 ) | ( n29802 & ~n29889 ) ;
  assign n29891 = ~n29802 & n29890 ;
  assign n29892 = x627 | n29800 ;
  assign n29893 = x618 & ~n29830 ;
  assign n29894 = x1154 | n29893 ;
  assign n29895 = ( n29885 & n29886 ) | ( n29885 & ~n29894 ) | ( n29886 & ~n29894 ) ;
  assign n29896 = ( ~n29891 & n29892 ) | ( ~n29891 & n29895 ) | ( n29892 & n29895 ) ;
  assign n29897 = ~n29891 & n29896 ;
  assign n29898 = n29885 ^ x781 ^ 1'b0 ;
  assign n29899 = ( n29885 & n29897 ) | ( n29885 & n29898 ) | ( n29897 & n29898 ) ;
  assign n29900 = ~x789 & n29899 ;
  assign n29901 = x619 & ~n29831 ;
  assign n29902 = x1159 | n29901 ;
  assign n29903 = x619 & ~n29899 ;
  assign n29904 = ( n29899 & ~n29902 ) | ( n29899 & n29903 ) | ( ~n29902 & n29903 ) ;
  assign n29905 = ( x648 & n29807 ) | ( x648 & ~n29904 ) | ( n29807 & ~n29904 ) ;
  assign n29906 = n29904 | n29905 ;
  assign n29907 = x619 | n29831 ;
  assign n29908 = x1159 & ~n29903 ;
  assign n29909 = n29907 & n29908 ;
  assign n29910 = ( x648 & n29809 ) | ( x648 & ~n29909 ) | ( n29809 & ~n29909 ) ;
  assign n29911 = ~n29809 & n29910 ;
  assign n29912 = x789 & ~n29911 ;
  assign n29913 = n29906 & n29912 ;
  assign n29914 = ( n16519 & ~n29900 ) | ( n16519 & n29913 ) | ( ~n29900 & n29913 ) ;
  assign n29915 = n29900 | n29914 ;
  assign n29916 = n29915 ^ n29856 ^ 1'b0 ;
  assign n29917 = ( n29856 & n29915 ) | ( n29856 & n29916 ) | ( n29915 & n29916 ) ;
  assign n29918 = ( n18482 & ~n29856 ) | ( n18482 & n29917 ) | ( ~n29856 & n29917 ) ;
  assign n29919 = n19208 | n29833 ;
  assign n29920 = n16556 & ~n29814 ;
  assign n29921 = x629 & ~n29920 ;
  assign n29922 = n29919 & n29921 ;
  assign n29923 = n16557 & ~n29814 ;
  assign n29924 = n19212 & ~n29833 ;
  assign n29925 = n29923 | n29924 ;
  assign n29926 = ( x629 & ~n29922 ) | ( x629 & n29925 ) | ( ~n29922 & n29925 ) ;
  assign n29927 = ~n29922 & n29926 ;
  assign n29928 = ( x792 & ~n19206 ) | ( x792 & n29927 ) | ( ~n19206 & n29927 ) ;
  assign n29929 = ( n18484 & n19206 ) | ( n18484 & n29928 ) | ( n19206 & n29928 ) ;
  assign n29930 = ( n29843 & n29918 ) | ( n29843 & ~n29929 ) | ( n29918 & ~n29929 ) ;
  assign n29931 = n29930 ^ n29918 ^ 1'b0 ;
  assign n29932 = ( n29843 & n29930 ) | ( n29843 & ~n29931 ) | ( n29930 & ~n29931 ) ;
  assign n29933 = x790 | n29932 ;
  assign n29934 = x644 & ~n29932 ;
  assign n29935 = ( x787 & n29836 ) | ( x787 & ~n29839 ) | ( n29836 & ~n29839 ) ;
  assign n29936 = ~n29836 & n29935 ;
  assign n29937 = ( x787 & n29834 ) | ( x787 & ~n29936 ) | ( n29834 & ~n29936 ) ;
  assign n29938 = ~n29936 & n29937 ;
  assign n29939 = x644 | n29938 ;
  assign n29940 = ( x715 & n29934 ) | ( x715 & n29939 ) | ( n29934 & n29939 ) ;
  assign n29941 = ~n29934 & n29940 ;
  assign n29942 = x644 | n29789 ;
  assign n29943 = n29789 ^ n16376 ^ 1'b0 ;
  assign n29944 = ( n29789 & n29816 ) | ( n29789 & ~n29943 ) | ( n29816 & ~n29943 ) ;
  assign n29945 = x644 & ~n29944 ;
  assign n29946 = ( x715 & n29942 ) | ( x715 & ~n29945 ) | ( n29942 & ~n29945 ) ;
  assign n29947 = ~x715 & n29946 ;
  assign n29948 = ( x1160 & n29941 ) | ( x1160 & ~n29947 ) | ( n29941 & ~n29947 ) ;
  assign n29949 = ~n29941 & n29948 ;
  assign n29950 = x644 & ~n29789 ;
  assign n29951 = x715 & ~n29950 ;
  assign n29952 = ( n29944 & n29945 ) | ( n29944 & n29951 ) | ( n29945 & n29951 ) ;
  assign n29953 = x644 & ~n29938 ;
  assign n29954 = x715 | n29953 ;
  assign n29955 = ( n29932 & n29934 ) | ( n29932 & ~n29954 ) | ( n29934 & ~n29954 ) ;
  assign n29956 = ( x1160 & ~n29952 ) | ( x1160 & n29955 ) | ( ~n29952 & n29955 ) ;
  assign n29957 = n29952 | n29956 ;
  assign n29958 = x790 & ~n29957 ;
  assign n29959 = ( x790 & n29949 ) | ( x790 & n29958 ) | ( n29949 & n29958 ) ;
  assign n29960 = x832 & ~n29959 ;
  assign n29961 = n29933 & n29960 ;
  assign n29962 = ~x192 & n7318 ;
  assign n29963 = x832 | n29962 ;
  assign n29964 = ~n29961 & n29963 ;
  assign n29965 = ( n29788 & n29961 ) | ( n29788 & ~n29964 ) | ( n29961 & ~n29964 ) ;
  assign n29966 = x193 | n15656 ;
  assign n29967 = ( x38 & x193 ) | ( x38 & n16700 ) | ( x193 & n16700 ) ;
  assign n29968 = ~n2069 & n29967 ;
  assign n29969 = ( x193 & n16697 ) | ( x193 & ~n29968 ) | ( n16697 & ~n29968 ) ;
  assign n29970 = ~n29968 & n29969 ;
  assign n29971 = x193 | n15644 ;
  assign n29972 = n16185 & n29971 ;
  assign n29973 = ( x690 & n29970 ) | ( x690 & ~n29972 ) | ( n29970 & ~n29972 ) ;
  assign n29974 = ~n29970 & n29973 ;
  assign n29975 = x690 & ~n2069 ;
  assign n29976 = ( n29966 & ~n29974 ) | ( n29966 & n29975 ) | ( ~n29974 & n29975 ) ;
  assign n29977 = ~n29974 & n29976 ;
  assign n29978 = x625 & ~n29977 ;
  assign n29979 = x625 | n29966 ;
  assign n29980 = ( x1153 & n29978 ) | ( x1153 & n29979 ) | ( n29978 & n29979 ) ;
  assign n29981 = ~n29978 & n29980 ;
  assign n29982 = x625 & ~n29966 ;
  assign n29983 = x1153 | n29982 ;
  assign n29984 = ( x625 & n29977 ) | ( x625 & ~n29983 ) | ( n29977 & ~n29983 ) ;
  assign n29985 = ~n29983 & n29984 ;
  assign n29986 = n29981 | n29985 ;
  assign n29987 = n29977 ^ x778 ^ 1'b0 ;
  assign n29988 = ( n29977 & n29986 ) | ( n29977 & n29987 ) | ( n29986 & n29987 ) ;
  assign n29989 = n29966 ^ n16234 ^ 1'b0 ;
  assign n29990 = ( n29966 & n29988 ) | ( n29966 & ~n29989 ) | ( n29988 & ~n29989 ) ;
  assign n29991 = n29966 ^ n16254 ^ 1'b0 ;
  assign n29992 = ( n29966 & n29990 ) | ( n29966 & ~n29991 ) | ( n29990 & ~n29991 ) ;
  assign n29993 = n29966 ^ n16279 ^ 1'b0 ;
  assign n29994 = ( n29966 & n29992 ) | ( n29966 & ~n29993 ) | ( n29992 & ~n29993 ) ;
  assign n29995 = n29966 ^ n16318 ^ 1'b0 ;
  assign n29996 = ( n29966 & n29994 ) | ( n29966 & ~n29995 ) | ( n29994 & ~n29995 ) ;
  assign n29997 = x628 & ~n29996 ;
  assign n29998 = x628 | n29966 ;
  assign n29999 = ( x1156 & n29997 ) | ( x1156 & n29998 ) | ( n29997 & n29998 ) ;
  assign n30000 = ~n29997 & n29999 ;
  assign n30001 = x628 & ~n29966 ;
  assign n30002 = x1156 | n30001 ;
  assign n30003 = ( n29996 & n29997 ) | ( n29996 & ~n30002 ) | ( n29997 & ~n30002 ) ;
  assign n30004 = n30000 | n30003 ;
  assign n30005 = n29996 ^ x792 ^ 1'b0 ;
  assign n30006 = ( n29996 & n30004 ) | ( n29996 & n30005 ) | ( n30004 & n30005 ) ;
  assign n30007 = n29966 ^ x647 ^ 1'b0 ;
  assign n30008 = ( n29966 & n30006 ) | ( n29966 & ~n30007 ) | ( n30006 & ~n30007 ) ;
  assign n30009 = ( n29966 & n30006 ) | ( n29966 & n30007 ) | ( n30006 & n30007 ) ;
  assign n30010 = n30008 ^ x1157 ^ 1'b0 ;
  assign n30011 = ( n30008 & n30009 ) | ( n30008 & n30010 ) | ( n30009 & n30010 ) ;
  assign n30012 = n30006 ^ x787 ^ 1'b0 ;
  assign n30013 = ( n30006 & n30011 ) | ( n30006 & n30012 ) | ( n30011 & n30012 ) ;
  assign n30014 = x644 & ~n30013 ;
  assign n30015 = x715 | n30014 ;
  assign n30016 = x644 & ~n29966 ;
  assign n30017 = x715 & ~n30016 ;
  assign n30018 = n30017 ^ x1160 ^ 1'b0 ;
  assign n30019 = x739 & n15646 ;
  assign n30020 = n29971 & ~n30019 ;
  assign n30021 = ~x193 & n15587 ;
  assign n30022 = x193 & ~n15640 ;
  assign n30023 = ( x739 & n30021 ) | ( x739 & ~n30022 ) | ( n30021 & ~n30022 ) ;
  assign n30024 = ~n30021 & n30023 ;
  assign n30025 = x193 | x739 ;
  assign n30026 = ( n15488 & ~n30024 ) | ( n15488 & n30025 ) | ( ~n30024 & n30025 ) ;
  assign n30027 = ~n30024 & n30026 ;
  assign n30028 = n30020 ^ x38 ^ 1'b0 ;
  assign n30029 = ( n30020 & n30027 ) | ( n30020 & ~n30028 ) | ( n30027 & ~n30028 ) ;
  assign n30030 = ~n2069 & n30029 ;
  assign n30031 = x193 & n2069 ;
  assign n30032 = n30030 | n30031 ;
  assign n30033 = n29966 ^ n15659 ^ 1'b0 ;
  assign n30034 = ( n29966 & n30032 ) | ( n29966 & ~n30033 ) | ( n30032 & ~n30033 ) ;
  assign n30035 = n15662 & n29966 ;
  assign n30036 = ( ~n15662 & n30030 ) | ( ~n15662 & n30031 ) | ( n30030 & n30031 ) ;
  assign n30037 = n30035 | n30036 ;
  assign n30038 = n30037 ^ n30034 ^ n29966 ;
  assign n30039 = n30038 ^ x1155 ^ 1'b0 ;
  assign n30040 = ( n30037 & n30038 ) | ( n30037 & ~n30039 ) | ( n30038 & ~n30039 ) ;
  assign n30041 = n30034 ^ x785 ^ 1'b0 ;
  assign n30042 = ( n30034 & n30040 ) | ( n30034 & n30041 ) | ( n30040 & n30041 ) ;
  assign n30043 = x618 & ~n30042 ;
  assign n30044 = x618 | n29966 ;
  assign n30045 = ( x1154 & n30043 ) | ( x1154 & n30044 ) | ( n30043 & n30044 ) ;
  assign n30046 = ~n30043 & n30045 ;
  assign n30047 = x618 & ~n29966 ;
  assign n30048 = x1154 | n30047 ;
  assign n30049 = ( n30042 & n30043 ) | ( n30042 & ~n30048 ) | ( n30043 & ~n30048 ) ;
  assign n30050 = n30046 | n30049 ;
  assign n30051 = n30042 ^ x781 ^ 1'b0 ;
  assign n30052 = ( n30042 & n30050 ) | ( n30042 & n30051 ) | ( n30050 & n30051 ) ;
  assign n30053 = x619 & ~n30052 ;
  assign n30054 = x619 | n29966 ;
  assign n30055 = ( x1159 & n30053 ) | ( x1159 & n30054 ) | ( n30053 & n30054 ) ;
  assign n30056 = ~n30053 & n30055 ;
  assign n30057 = x619 & ~n29966 ;
  assign n30058 = x1159 | n30057 ;
  assign n30059 = ( n30052 & n30053 ) | ( n30052 & ~n30058 ) | ( n30053 & ~n30058 ) ;
  assign n30060 = n30056 | n30059 ;
  assign n30061 = n30052 ^ x789 ^ 1'b0 ;
  assign n30062 = ( n30052 & n30060 ) | ( n30052 & n30061 ) | ( n30060 & n30061 ) ;
  assign n30063 = n29966 ^ n16518 ^ 1'b0 ;
  assign n30064 = ( n29966 & n30062 ) | ( n29966 & ~n30063 ) | ( n30062 & ~n30063 ) ;
  assign n30065 = n29966 ^ n16339 ^ 1'b0 ;
  assign n30066 = ( n29966 & n30064 ) | ( n29966 & ~n30065 ) | ( n30064 & ~n30065 ) ;
  assign n30067 = n29966 ^ n16376 ^ 1'b0 ;
  assign n30068 = ( n29966 & n30066 ) | ( n29966 & ~n30067 ) | ( n30066 & ~n30067 ) ;
  assign n30069 = x644 | n30068 ;
  assign n30070 = ( n30017 & ~n30018 ) | ( n30017 & n30069 ) | ( ~n30018 & n30069 ) ;
  assign n30071 = ( x1160 & n30018 ) | ( x1160 & n30070 ) | ( n30018 & n30070 ) ;
  assign n30072 = n30015 & ~n30071 ;
  assign n30073 = x644 & ~n30068 ;
  assign n30074 = ( ~x715 & n29966 ) | ( ~x715 & n30016 ) | ( n29966 & n30016 ) ;
  assign n30075 = x1160 & ~n30074 ;
  assign n30076 = ( x1160 & n30073 ) | ( x1160 & n30075 ) | ( n30073 & n30075 ) ;
  assign n30077 = ( x715 & n30013 ) | ( x715 & n30014 ) | ( n30013 & n30014 ) ;
  assign n30078 = n30076 & ~n30077 ;
  assign n30079 = ( x790 & n30072 ) | ( x790 & n30078 ) | ( n30072 & n30078 ) ;
  assign n30080 = n30078 ^ n30072 ^ 1'b0 ;
  assign n30081 = ( x790 & n30079 ) | ( x790 & n30080 ) | ( n30079 & n30080 ) ;
  assign n30082 = n19055 & n30066 ;
  assign n30083 = n16374 & n30008 ;
  assign n30084 = n16373 & n30009 ;
  assign n30085 = n30083 | n30084 ;
  assign n30086 = ( x787 & n30082 ) | ( x787 & n30085 ) | ( n30082 & n30085 ) ;
  assign n30087 = n30085 ^ n30082 ^ 1'b0 ;
  assign n30088 = ( x787 & n30086 ) | ( x787 & n30087 ) | ( n30086 & n30087 ) ;
  assign n30089 = x690 | n30029 ;
  assign n30090 = x193 & ~n16029 ;
  assign n30091 = ~x193 & n16044 ;
  assign n30092 = ( x739 & ~n30090 ) | ( x739 & n30091 ) | ( ~n30090 & n30091 ) ;
  assign n30093 = n30090 | n30092 ;
  assign n30094 = ~x193 & n16048 ;
  assign n30095 = x193 & ~n16054 ;
  assign n30096 = ( x739 & n30094 ) | ( x739 & ~n30095 ) | ( n30094 & ~n30095 ) ;
  assign n30097 = ~n30094 & n30096 ;
  assign n30098 = ( x39 & n30093 ) | ( x39 & ~n30097 ) | ( n30093 & ~n30097 ) ;
  assign n30099 = n30098 ^ n30093 ^ 1'b0 ;
  assign n30100 = ( x39 & n30098 ) | ( x39 & ~n30099 ) | ( n30098 & ~n30099 ) ;
  assign n30101 = ( x739 & n15795 ) | ( x739 & n30025 ) | ( n15795 & n30025 ) ;
  assign n30102 = ( x193 & n15876 ) | ( x193 & ~n30101 ) | ( n15876 & ~n30101 ) ;
  assign n30103 = ~n30101 & n30102 ;
  assign n30104 = x193 | n16003 ;
  assign n30105 = x193 & n15943 ;
  assign n30106 = x739 & ~n30105 ;
  assign n30107 = n30104 & n30106 ;
  assign n30108 = ( x39 & n30103 ) | ( x39 & ~n30107 ) | ( n30103 & ~n30107 ) ;
  assign n30109 = ~n30103 & n30108 ;
  assign n30110 = ( x38 & n30100 ) | ( x38 & ~n30109 ) | ( n30100 & ~n30109 ) ;
  assign n30111 = ~x38 & n30110 ;
  assign n30112 = x739 & n15591 ;
  assign n30113 = n17156 | n30112 ;
  assign n30114 = x193 & ~n5017 ;
  assign n30115 = n30113 & n30114 ;
  assign n30116 = ~x739 & n22207 ;
  assign n30117 = n15968 | n30116 ;
  assign n30118 = x39 | n30117 ;
  assign n30119 = ( ~x39 & x193 ) | ( ~x39 & n30118 ) | ( x193 & n30118 ) ;
  assign n30120 = ( x38 & n30115 ) | ( x38 & n30119 ) | ( n30115 & n30119 ) ;
  assign n30121 = ~n30115 & n30120 ;
  assign n30122 = ( x690 & n30111 ) | ( x690 & ~n30121 ) | ( n30111 & ~n30121 ) ;
  assign n30123 = ~n30111 & n30122 ;
  assign n30124 = ( n2051 & n2068 ) | ( n2051 & ~n30123 ) | ( n2068 & ~n30123 ) ;
  assign n30125 = n30123 | n30124 ;
  assign n30126 = ( n30031 & n30089 ) | ( n30031 & ~n30125 ) | ( n30089 & ~n30125 ) ;
  assign n30127 = n30126 ^ n30089 ^ 1'b0 ;
  assign n30128 = ( n30031 & n30126 ) | ( n30031 & ~n30127 ) | ( n30126 & ~n30127 ) ;
  assign n30129 = x625 & ~n30128 ;
  assign n30130 = x625 | n30032 ;
  assign n30131 = ( x1153 & n30129 ) | ( x1153 & n30130 ) | ( n30129 & n30130 ) ;
  assign n30132 = ~n30129 & n30131 ;
  assign n30133 = ( x608 & n29985 ) | ( x608 & ~n30132 ) | ( n29985 & ~n30132 ) ;
  assign n30134 = ~n29985 & n30133 ;
  assign n30135 = x608 | n29981 ;
  assign n30136 = x625 & ~n30032 ;
  assign n30137 = x1153 | n30136 ;
  assign n30138 = ( n30128 & n30129 ) | ( n30128 & ~n30137 ) | ( n30129 & ~n30137 ) ;
  assign n30139 = ( ~n30134 & n30135 ) | ( ~n30134 & n30138 ) | ( n30135 & n30138 ) ;
  assign n30140 = ~n30134 & n30139 ;
  assign n30141 = n30128 ^ x778 ^ 1'b0 ;
  assign n30142 = ( n30128 & n30140 ) | ( n30128 & n30141 ) | ( n30140 & n30141 ) ;
  assign n30143 = x609 & ~n30142 ;
  assign n30144 = x609 | n29988 ;
  assign n30145 = ( x1155 & n30143 ) | ( x1155 & n30144 ) | ( n30143 & n30144 ) ;
  assign n30146 = ~n30143 & n30145 ;
  assign n30147 = ~x1155 & n30037 ;
  assign n30148 = ( x660 & n30146 ) | ( x660 & ~n30147 ) | ( n30146 & ~n30147 ) ;
  assign n30149 = ~n30146 & n30148 ;
  assign n30150 = x1155 & n30038 ;
  assign n30151 = x660 | n30150 ;
  assign n30152 = x609 & ~n29988 ;
  assign n30153 = x1155 | n30152 ;
  assign n30154 = ( n30142 & n30143 ) | ( n30142 & ~n30153 ) | ( n30143 & ~n30153 ) ;
  assign n30155 = ( ~n30149 & n30151 ) | ( ~n30149 & n30154 ) | ( n30151 & n30154 ) ;
  assign n30156 = ~n30149 & n30155 ;
  assign n30157 = n30142 ^ x785 ^ 1'b0 ;
  assign n30158 = ( n30142 & n30156 ) | ( n30142 & n30157 ) | ( n30156 & n30157 ) ;
  assign n30159 = x618 & ~n30158 ;
  assign n30160 = x618 | n29990 ;
  assign n30161 = ( x1154 & n30159 ) | ( x1154 & n30160 ) | ( n30159 & n30160 ) ;
  assign n30162 = ~n30159 & n30161 ;
  assign n30163 = ( x627 & n30049 ) | ( x627 & ~n30162 ) | ( n30049 & ~n30162 ) ;
  assign n30164 = ~n30049 & n30163 ;
  assign n30165 = x627 | n30046 ;
  assign n30166 = x618 & ~n29990 ;
  assign n30167 = x1154 | n30166 ;
  assign n30168 = ( n30158 & n30159 ) | ( n30158 & ~n30167 ) | ( n30159 & ~n30167 ) ;
  assign n30169 = ( ~n30164 & n30165 ) | ( ~n30164 & n30168 ) | ( n30165 & n30168 ) ;
  assign n30170 = ~n30164 & n30169 ;
  assign n30171 = n30158 ^ x781 ^ 1'b0 ;
  assign n30172 = ( n30158 & n30170 ) | ( n30158 & n30171 ) | ( n30170 & n30171 ) ;
  assign n30173 = x619 | n30172 ;
  assign n30174 = x619 & ~n29992 ;
  assign n30175 = ( x1159 & n30173 ) | ( x1159 & ~n30174 ) | ( n30173 & ~n30174 ) ;
  assign n30176 = ~x1159 & n30175 ;
  assign n30177 = ( x648 & n30056 ) | ( x648 & ~n30176 ) | ( n30056 & ~n30176 ) ;
  assign n30178 = n30176 | n30177 ;
  assign n30179 = x619 & ~n30172 ;
  assign n30180 = x619 | n29992 ;
  assign n30181 = ( x1159 & n30179 ) | ( x1159 & n30180 ) | ( n30179 & n30180 ) ;
  assign n30182 = ~n30179 & n30181 ;
  assign n30183 = ( x648 & n30059 ) | ( x648 & ~n30182 ) | ( n30059 & ~n30182 ) ;
  assign n30184 = ~n30059 & n30183 ;
  assign n30185 = x789 & ~n30184 ;
  assign n30186 = n30178 & n30185 ;
  assign n30187 = ~x789 & n30172 ;
  assign n30188 = ( n16519 & ~n30186 ) | ( n16519 & n30187 ) | ( ~n30186 & n30187 ) ;
  assign n30189 = n30186 | n30188 ;
  assign n30190 = n30000 ^ x629 ^ 1'b0 ;
  assign n30191 = ( n30000 & n30003 ) | ( n30000 & n30190 ) | ( n30003 & n30190 ) ;
  assign n30192 = n19046 & n30064 ;
  assign n30193 = ( x792 & n30191 ) | ( x792 & n30192 ) | ( n30191 & n30192 ) ;
  assign n30194 = n30192 ^ n30191 ^ 1'b0 ;
  assign n30195 = ( x792 & n30193 ) | ( x792 & n30194 ) | ( n30193 & n30194 ) ;
  assign n30196 = n16459 & ~n29994 ;
  assign n30197 = ~x626 & n29966 ;
  assign n30198 = x626 & n30062 ;
  assign n30199 = ( n22317 & n30197 ) | ( n22317 & ~n30198 ) | ( n30197 & ~n30198 ) ;
  assign n30200 = ~n30197 & n30199 ;
  assign n30201 = ~x626 & n30062 ;
  assign n30202 = x626 & n29966 ;
  assign n30203 = ( n22322 & n30201 ) | ( n22322 & ~n30202 ) | ( n30201 & ~n30202 ) ;
  assign n30204 = ~n30201 & n30203 ;
  assign n30205 = ( ~n30196 & n30200 ) | ( ~n30196 & n30204 ) | ( n30200 & n30204 ) ;
  assign n30206 = n30196 | n30205 ;
  assign n30207 = ( x788 & ~n22314 ) | ( x788 & n30206 ) | ( ~n22314 & n30206 ) ;
  assign n30208 = ( n18482 & n22314 ) | ( n18482 & n30207 ) | ( n22314 & n30207 ) ;
  assign n30209 = ~n30195 & n30208 ;
  assign n30210 = ( n30189 & n30195 ) | ( n30189 & ~n30209 ) | ( n30195 & ~n30209 ) ;
  assign n30211 = ( ~n18484 & n30088 ) | ( ~n18484 & n30210 ) | ( n30088 & n30210 ) ;
  assign n30212 = n30088 ^ n18484 ^ 1'b0 ;
  assign n30213 = ( n30088 & n30211 ) | ( n30088 & ~n30212 ) | ( n30211 & ~n30212 ) ;
  assign n30214 = x644 | n30071 ;
  assign n30215 = x644 & n30076 ;
  assign n30216 = x790 & ~n30215 ;
  assign n30217 = n30214 & n30216 ;
  assign n30218 = ( ~n30081 & n30213 ) | ( ~n30081 & n30217 ) | ( n30213 & n30217 ) ;
  assign n30219 = ~n30081 & n30218 ;
  assign n30220 = ( x57 & n5193 ) | ( x57 & ~n30219 ) | ( n5193 & ~n30219 ) ;
  assign n30221 = n30219 | n30220 ;
  assign n30222 = x193 | n1611 ;
  assign n30223 = ~n30112 & n30222 ;
  assign n30224 = n16397 | n30223 ;
  assign n30225 = ~n15662 & n30112 ;
  assign n30226 = ~x1155 & n30222 ;
  assign n30227 = ~n30225 & n30226 ;
  assign n30228 = ( x1155 & n30224 ) | ( x1155 & n30225 ) | ( n30224 & n30225 ) ;
  assign n30229 = n30227 | n30228 ;
  assign n30230 = n30224 ^ x785 ^ 1'b0 ;
  assign n30231 = ( n30224 & n30229 ) | ( n30224 & n30230 ) | ( n30229 & n30230 ) ;
  assign n30232 = n16411 | n30231 ;
  assign n30233 = x1154 & n30232 ;
  assign n30234 = n16414 | n30231 ;
  assign n30235 = ~x1154 & n30234 ;
  assign n30236 = n30233 | n30235 ;
  assign n30237 = n30231 ^ x781 ^ 1'b0 ;
  assign n30238 = ( n30231 & n30236 ) | ( n30231 & n30237 ) | ( n30236 & n30237 ) ;
  assign n30239 = n21437 | n30238 ;
  assign n30240 = x1159 & n30239 ;
  assign n30241 = n21440 | n30238 ;
  assign n30242 = ~x1159 & n30241 ;
  assign n30243 = n30240 | n30242 ;
  assign n30244 = n30238 ^ x789 ^ 1'b0 ;
  assign n30245 = ( n30238 & n30243 ) | ( n30238 & n30244 ) | ( n30243 & n30244 ) ;
  assign n30246 = n30222 ^ n16518 ^ 1'b0 ;
  assign n30247 = ( n30222 & n30245 ) | ( n30222 & ~n30246 ) | ( n30245 & ~n30246 ) ;
  assign n30248 = n30222 ^ n16339 ^ 1'b0 ;
  assign n30249 = ( n30222 & n30247 ) | ( n30222 & ~n30248 ) | ( n30247 & ~n30248 ) ;
  assign n30250 = n19055 & n30249 ;
  assign n30251 = x647 & ~n30222 ;
  assign n30252 = x1157 | n30251 ;
  assign n30253 = x690 & n15778 ;
  assign n30254 = ~x625 & n30253 ;
  assign n30255 = ~x1153 & n30222 ;
  assign n30256 = ~n30254 & n30255 ;
  assign n30257 = x778 & ~n30256 ;
  assign n30258 = n30222 & ~n30253 ;
  assign n30259 = ( x1153 & n30254 ) | ( x1153 & n30258 ) | ( n30254 & n30258 ) ;
  assign n30260 = n30257 & ~n30259 ;
  assign n30261 = ( x778 & n30258 ) | ( x778 & ~n30260 ) | ( n30258 & ~n30260 ) ;
  assign n30262 = ~n30260 & n30261 ;
  assign n30263 = n16447 | n30262 ;
  assign n30264 = n16449 | n30263 ;
  assign n30265 = n16451 | n30264 ;
  assign n30266 = n16530 | n30265 ;
  assign n30267 = n16560 | n30266 ;
  assign n30268 = ( x647 & ~n30252 ) | ( x647 & n30267 ) | ( ~n30252 & n30267 ) ;
  assign n30269 = ~n30252 & n30268 ;
  assign n30270 = n30222 ^ x647 ^ 1'b0 ;
  assign n30271 = ( n30222 & n30267 ) | ( n30222 & n30270 ) | ( n30267 & n30270 ) ;
  assign n30272 = x1157 & n30271 ;
  assign n30273 = ( n16375 & n30269 ) | ( n16375 & n30272 ) | ( n30269 & n30272 ) ;
  assign n30274 = ( x787 & n30250 ) | ( x787 & n30273 ) | ( n30250 & n30273 ) ;
  assign n30275 = n30273 ^ n30250 ^ 1'b0 ;
  assign n30276 = ( x787 & n30274 ) | ( x787 & n30275 ) | ( n30274 & n30275 ) ;
  assign n30277 = ~x626 & n30222 ;
  assign n30278 = x626 & n30245 ;
  assign n30279 = ( n22317 & n30277 ) | ( n22317 & ~n30278 ) | ( n30277 & ~n30278 ) ;
  assign n30280 = ~n30277 & n30279 ;
  assign n30281 = ~x626 & n30245 ;
  assign n30282 = x626 & n30222 ;
  assign n30283 = ( n22322 & n30281 ) | ( n22322 & ~n30282 ) | ( n30281 & ~n30282 ) ;
  assign n30284 = ~n30281 & n30283 ;
  assign n30285 = n30265 & ~n30284 ;
  assign n30286 = ( n16459 & n30284 ) | ( n16459 & ~n30285 ) | ( n30284 & ~n30285 ) ;
  assign n30287 = ( x788 & n30280 ) | ( x788 & n30286 ) | ( n30280 & n30286 ) ;
  assign n30288 = n30286 ^ n30280 ^ 1'b0 ;
  assign n30289 = ( x788 & n30287 ) | ( x788 & n30288 ) | ( n30287 & n30288 ) ;
  assign n30290 = n15524 | n30258 ;
  assign n30291 = n30223 & n30290 ;
  assign n30292 = x625 & ~n30290 ;
  assign n30293 = ( n30255 & n30291 ) | ( n30255 & n30292 ) | ( n30291 & n30292 ) ;
  assign n30294 = ( x608 & n30259 ) | ( x608 & ~n30293 ) | ( n30259 & ~n30293 ) ;
  assign n30295 = n30293 | n30294 ;
  assign n30296 = x1153 & n30223 ;
  assign n30297 = ~n30292 & n30296 ;
  assign n30298 = x608 & ~n30256 ;
  assign n30299 = n30295 & ~n30298 ;
  assign n30300 = ( n30295 & n30297 ) | ( n30295 & n30299 ) | ( n30297 & n30299 ) ;
  assign n30301 = n30291 ^ x778 ^ 1'b0 ;
  assign n30302 = ( n30291 & n30300 ) | ( n30291 & n30301 ) | ( n30300 & n30301 ) ;
  assign n30303 = x609 & ~n30302 ;
  assign n30309 = x609 | n30262 ;
  assign n30310 = ( x1155 & n30303 ) | ( x1155 & n30309 ) | ( n30303 & n30309 ) ;
  assign n30311 = ~n30303 & n30310 ;
  assign n30312 = ( x660 & n30227 ) | ( x660 & ~n30311 ) | ( n30227 & ~n30311 ) ;
  assign n30313 = ~n30227 & n30312 ;
  assign n30304 = x609 & ~n30262 ;
  assign n30305 = x1155 | n30304 ;
  assign n30306 = ( n30302 & n30303 ) | ( n30302 & ~n30305 ) | ( n30303 & ~n30305 ) ;
  assign n30307 = ( x660 & n30228 ) | ( x660 & ~n30306 ) | ( n30228 & ~n30306 ) ;
  assign n30308 = n30306 | n30307 ;
  assign n30314 = n30313 ^ n30308 ^ 1'b0 ;
  assign n30315 = ( x785 & ~n30308 ) | ( x785 & n30313 ) | ( ~n30308 & n30313 ) ;
  assign n30316 = ( x785 & ~n30314 ) | ( x785 & n30315 ) | ( ~n30314 & n30315 ) ;
  assign n30317 = ( x785 & n30302 ) | ( x785 & ~n30316 ) | ( n30302 & ~n30316 ) ;
  assign n30318 = ~n30316 & n30317 ;
  assign n30319 = x618 & ~n30318 ;
  assign n30320 = x618 | n30263 ;
  assign n30321 = ( x1154 & n30319 ) | ( x1154 & n30320 ) | ( n30319 & n30320 ) ;
  assign n30322 = ~n30319 & n30321 ;
  assign n30323 = ( x627 & n30235 ) | ( x627 & ~n30322 ) | ( n30235 & ~n30322 ) ;
  assign n30324 = ~n30235 & n30323 ;
  assign n30325 = x627 | n30233 ;
  assign n30326 = x618 & ~n30263 ;
  assign n30327 = x1154 | n30326 ;
  assign n30328 = ( n30318 & n30319 ) | ( n30318 & ~n30327 ) | ( n30319 & ~n30327 ) ;
  assign n30329 = ( ~n30324 & n30325 ) | ( ~n30324 & n30328 ) | ( n30325 & n30328 ) ;
  assign n30330 = ~n30324 & n30329 ;
  assign n30331 = n30318 ^ x781 ^ 1'b0 ;
  assign n30332 = ( n30318 & n30330 ) | ( n30318 & n30331 ) | ( n30330 & n30331 ) ;
  assign n30333 = ~x789 & n30332 ;
  assign n30334 = x619 & ~n30264 ;
  assign n30335 = x1159 | n30334 ;
  assign n30336 = x619 & ~n30332 ;
  assign n30337 = ( n30332 & ~n30335 ) | ( n30332 & n30336 ) | ( ~n30335 & n30336 ) ;
  assign n30338 = ( x648 & n30240 ) | ( x648 & ~n30337 ) | ( n30240 & ~n30337 ) ;
  assign n30339 = n30337 | n30338 ;
  assign n30340 = x619 | n30264 ;
  assign n30341 = x1159 & ~n30336 ;
  assign n30342 = n30340 & n30341 ;
  assign n30343 = ( x648 & n30242 ) | ( x648 & ~n30342 ) | ( n30242 & ~n30342 ) ;
  assign n30344 = ~n30242 & n30343 ;
  assign n30345 = x789 & ~n30344 ;
  assign n30346 = n30339 & n30345 ;
  assign n30347 = ( n16519 & ~n30333 ) | ( n16519 & n30346 ) | ( ~n30333 & n30346 ) ;
  assign n30348 = n30333 | n30347 ;
  assign n30349 = n30348 ^ n30289 ^ 1'b0 ;
  assign n30350 = ( n30289 & n30348 ) | ( n30289 & n30349 ) | ( n30348 & n30349 ) ;
  assign n30351 = ( n18482 & ~n30289 ) | ( n18482 & n30350 ) | ( ~n30289 & n30350 ) ;
  assign n30352 = n19208 | n30266 ;
  assign n30353 = n16556 & ~n30247 ;
  assign n30354 = x629 & ~n30353 ;
  assign n30355 = n30352 & n30354 ;
  assign n30356 = n16557 & ~n30247 ;
  assign n30357 = n19212 & ~n30266 ;
  assign n30358 = n30356 | n30357 ;
  assign n30359 = ( x629 & ~n30355 ) | ( x629 & n30358 ) | ( ~n30355 & n30358 ) ;
  assign n30360 = ~n30355 & n30359 ;
  assign n30361 = ( x792 & ~n19206 ) | ( x792 & n30360 ) | ( ~n19206 & n30360 ) ;
  assign n30362 = ( n18484 & n19206 ) | ( n18484 & n30361 ) | ( n19206 & n30361 ) ;
  assign n30363 = ( n30276 & n30351 ) | ( n30276 & ~n30362 ) | ( n30351 & ~n30362 ) ;
  assign n30364 = n30363 ^ n30351 ^ 1'b0 ;
  assign n30365 = ( n30276 & n30363 ) | ( n30276 & ~n30364 ) | ( n30363 & ~n30364 ) ;
  assign n30366 = x790 | n30365 ;
  assign n30367 = x644 & ~n30365 ;
  assign n30368 = ( x787 & n30269 ) | ( x787 & ~n30272 ) | ( n30269 & ~n30272 ) ;
  assign n30369 = ~n30269 & n30368 ;
  assign n30370 = ( x787 & n30267 ) | ( x787 & ~n30369 ) | ( n30267 & ~n30369 ) ;
  assign n30371 = ~n30369 & n30370 ;
  assign n30372 = x644 | n30371 ;
  assign n30373 = ( x715 & n30367 ) | ( x715 & n30372 ) | ( n30367 & n30372 ) ;
  assign n30374 = ~n30367 & n30373 ;
  assign n30375 = x644 | n30222 ;
  assign n30376 = n30222 ^ n16376 ^ 1'b0 ;
  assign n30377 = ( n30222 & n30249 ) | ( n30222 & ~n30376 ) | ( n30249 & ~n30376 ) ;
  assign n30378 = x644 & ~n30377 ;
  assign n30379 = ( x715 & n30375 ) | ( x715 & ~n30378 ) | ( n30375 & ~n30378 ) ;
  assign n30380 = ~x715 & n30379 ;
  assign n30381 = ( x1160 & n30374 ) | ( x1160 & ~n30380 ) | ( n30374 & ~n30380 ) ;
  assign n30382 = ~n30374 & n30381 ;
  assign n30383 = x644 & ~n30222 ;
  assign n30384 = x715 & ~n30383 ;
  assign n30385 = ( n30377 & n30378 ) | ( n30377 & n30384 ) | ( n30378 & n30384 ) ;
  assign n30386 = x644 & ~n30371 ;
  assign n30387 = x715 | n30386 ;
  assign n30388 = ( n30365 & n30367 ) | ( n30365 & ~n30387 ) | ( n30367 & ~n30387 ) ;
  assign n30389 = ( x1160 & ~n30385 ) | ( x1160 & n30388 ) | ( ~n30385 & n30388 ) ;
  assign n30390 = n30385 | n30389 ;
  assign n30391 = x790 & ~n30390 ;
  assign n30392 = ( x790 & n30382 ) | ( x790 & n30391 ) | ( n30382 & n30391 ) ;
  assign n30393 = x832 & ~n30392 ;
  assign n30394 = n30366 & n30393 ;
  assign n30395 = ~x193 & n7318 ;
  assign n30396 = x832 | n30395 ;
  assign n30397 = ~n30394 & n30396 ;
  assign n30398 = ( n30221 & n30394 ) | ( n30221 & ~n30397 ) | ( n30394 & ~n30397 ) ;
  assign n30432 = x194 & n22651 ;
  assign n30433 = x748 | n30432 ;
  assign n30434 = ( x194 & n17893 ) | ( x194 & ~n30433 ) | ( n17893 & ~n30433 ) ;
  assign n30435 = ~n30433 & n30434 ;
  assign n30436 = x194 & n17910 ;
  assign n30437 = x194 | n17902 ;
  assign n30438 = ( x748 & n30436 ) | ( x748 & n30437 ) | ( n30436 & n30437 ) ;
  assign n30439 = ~n30436 & n30438 ;
  assign n30440 = ( x730 & n30435 ) | ( x730 & ~n30439 ) | ( n30435 & ~n30439 ) ;
  assign n30441 = ~n30435 & n30440 ;
  assign n30399 = n17843 ^ x194 ^ 1'b0 ;
  assign n30400 = ( n17843 & ~n22572 ) | ( n17843 & n30399 ) | ( ~n22572 & n30399 ) ;
  assign n30401 = x194 | n15655 ;
  assign n30402 = n30400 ^ x748 ^ 1'b0 ;
  assign n30403 = ( n30400 & n30401 ) | ( n30400 & ~n30402 ) | ( n30401 & ~n30402 ) ;
  assign n30442 = x730 | n30403 ;
  assign n30443 = ( n2069 & ~n30441 ) | ( n2069 & n30442 ) | ( ~n30441 & n30442 ) ;
  assign n30444 = ~n2069 & n30443 ;
  assign n30445 = n30444 ^ x194 ^ 1'b0 ;
  assign n30446 = ( ~x194 & n2069 ) | ( ~x194 & n30445 ) | ( n2069 & n30445 ) ;
  assign n30447 = ( x194 & n30444 ) | ( x194 & n30446 ) | ( n30444 & n30446 ) ;
  assign n30448 = x625 & ~n30447 ;
  assign n30404 = n30403 ^ n2069 ^ 1'b0 ;
  assign n30405 = ( x194 & n30403 ) | ( x194 & n30404 ) | ( n30403 & n30404 ) ;
  assign n30449 = x625 | n30405 ;
  assign n30450 = ( x1153 & n30448 ) | ( x1153 & n30449 ) | ( n30448 & n30449 ) ;
  assign n30451 = ~n30448 & n30450 ;
  assign n30406 = x194 | n15656 ;
  assign n30452 = x625 & ~n30406 ;
  assign n30453 = x1153 | n30452 ;
  assign n30454 = ~x194 & n22522 ;
  assign n30455 = x730 & ~n30454 ;
  assign n30456 = x730 | n30401 ;
  assign n30457 = ( n2069 & ~n30455 ) | ( n2069 & n30456 ) | ( ~n30455 & n30456 ) ;
  assign n30458 = ~n2069 & n30457 ;
  assign n30459 = n22530 & ~n30458 ;
  assign n30460 = ( x194 & n30458 ) | ( x194 & ~n30459 ) | ( n30458 & ~n30459 ) ;
  assign n30461 = ( x625 & ~n30453 ) | ( x625 & n30460 ) | ( ~n30453 & n30460 ) ;
  assign n30462 = ~n30453 & n30461 ;
  assign n30463 = ( x608 & n30451 ) | ( x608 & ~n30462 ) | ( n30451 & ~n30462 ) ;
  assign n30464 = ~n30451 & n30463 ;
  assign n30465 = x625 & ~n30460 ;
  assign n30466 = x625 | n30406 ;
  assign n30467 = ( x1153 & n30465 ) | ( x1153 & n30466 ) | ( n30465 & n30466 ) ;
  assign n30468 = ~n30465 & n30467 ;
  assign n30469 = x608 | n30468 ;
  assign n30470 = x625 & ~n30405 ;
  assign n30471 = x1153 | n30470 ;
  assign n30472 = ( n30447 & n30448 ) | ( n30447 & ~n30471 ) | ( n30448 & ~n30471 ) ;
  assign n30473 = ( ~n30464 & n30469 ) | ( ~n30464 & n30472 ) | ( n30469 & n30472 ) ;
  assign n30474 = ~n30464 & n30473 ;
  assign n30475 = n30447 ^ x778 ^ 1'b0 ;
  assign n30476 = ( n30447 & n30474 ) | ( n30447 & n30475 ) | ( n30474 & n30475 ) ;
  assign n30477 = x609 & ~n30476 ;
  assign n30478 = n30462 | n30468 ;
  assign n30479 = n30460 ^ x778 ^ 1'b0 ;
  assign n30480 = ( n30460 & n30478 ) | ( n30460 & n30479 ) | ( n30478 & n30479 ) ;
  assign n30481 = x609 | n30480 ;
  assign n30482 = ( x1155 & n30477 ) | ( x1155 & n30481 ) | ( n30477 & n30481 ) ;
  assign n30483 = ~n30477 & n30482 ;
  assign n30409 = ~n15659 & n30405 ;
  assign n30410 = x609 & n30409 ;
  assign n30411 = ~n15668 & n30406 ;
  assign n30412 = n30410 | n30411 ;
  assign n30407 = n30405 ^ n15659 ^ 1'b0 ;
  assign n30408 = ( n30405 & n30406 ) | ( n30405 & n30407 ) | ( n30406 & n30407 ) ;
  assign n30414 = n30412 ^ n30408 ^ n30406 ;
  assign n30484 = ~x1155 & n30414 ;
  assign n30485 = ( x660 & n30483 ) | ( x660 & ~n30484 ) | ( n30483 & ~n30484 ) ;
  assign n30486 = ~n30483 & n30485 ;
  assign n30487 = x1155 & n30412 ;
  assign n30488 = x660 | n30487 ;
  assign n30489 = x609 & ~n30480 ;
  assign n30490 = x1155 | n30489 ;
  assign n30491 = ( n30476 & n30477 ) | ( n30476 & ~n30490 ) | ( n30477 & ~n30490 ) ;
  assign n30492 = ( ~n30486 & n30488 ) | ( ~n30486 & n30491 ) | ( n30488 & n30491 ) ;
  assign n30493 = ~n30486 & n30492 ;
  assign n30494 = n30476 ^ x785 ^ 1'b0 ;
  assign n30495 = ( n30476 & n30493 ) | ( n30476 & n30494 ) | ( n30493 & n30494 ) ;
  assign n30496 = x618 & ~n30495 ;
  assign n30497 = n30406 ^ n16234 ^ 1'b0 ;
  assign n30498 = ( n30406 & n30480 ) | ( n30406 & ~n30497 ) | ( n30480 & ~n30497 ) ;
  assign n30499 = x618 | n30498 ;
  assign n30500 = ( x1154 & n30496 ) | ( x1154 & n30499 ) | ( n30496 & n30499 ) ;
  assign n30501 = ~n30496 & n30500 ;
  assign n30413 = n30412 ^ x1155 ^ 1'b0 ;
  assign n30415 = ( n30412 & ~n30413 ) | ( n30412 & n30414 ) | ( ~n30413 & n30414 ) ;
  assign n30416 = n30408 ^ x785 ^ 1'b0 ;
  assign n30417 = ( n30408 & n30415 ) | ( n30408 & n30416 ) | ( n30415 & n30416 ) ;
  assign n30418 = x618 & ~n30417 ;
  assign n30422 = x618 & ~n30406 ;
  assign n30423 = x1154 | n30422 ;
  assign n30424 = ( n30417 & n30418 ) | ( n30417 & ~n30423 ) | ( n30418 & ~n30423 ) ;
  assign n30502 = ( x627 & ~n30424 ) | ( x627 & n30501 ) | ( ~n30424 & n30501 ) ;
  assign n30503 = ~n30501 & n30502 ;
  assign n30419 = x618 | n30406 ;
  assign n30420 = ( x1154 & n30418 ) | ( x1154 & n30419 ) | ( n30418 & n30419 ) ;
  assign n30421 = ~n30418 & n30420 ;
  assign n30504 = x627 | n30421 ;
  assign n30505 = x618 & ~n30498 ;
  assign n30506 = x1154 | n30505 ;
  assign n30507 = ( n30495 & n30496 ) | ( n30495 & ~n30506 ) | ( n30496 & ~n30506 ) ;
  assign n30508 = ( ~n30503 & n30504 ) | ( ~n30503 & n30507 ) | ( n30504 & n30507 ) ;
  assign n30509 = ~n30503 & n30508 ;
  assign n30510 = n30495 ^ x781 ^ 1'b0 ;
  assign n30511 = ( n30495 & n30509 ) | ( n30495 & n30510 ) | ( n30509 & n30510 ) ;
  assign n30512 = x619 & ~n30511 ;
  assign n30513 = n30406 ^ n16254 ^ 1'b0 ;
  assign n30514 = ( n30406 & n30498 ) | ( n30406 & ~n30513 ) | ( n30498 & ~n30513 ) ;
  assign n30520 = x619 | n30514 ;
  assign n30521 = ( x1159 & n30512 ) | ( x1159 & n30520 ) | ( n30512 & n30520 ) ;
  assign n30522 = ~n30512 & n30521 ;
  assign n30425 = n30421 | n30424 ;
  assign n30426 = n30417 ^ x781 ^ 1'b0 ;
  assign n30427 = ( n30417 & n30425 ) | ( n30417 & n30426 ) | ( n30425 & n30426 ) ;
  assign n30428 = x619 & ~n30427 ;
  assign n30523 = x619 & ~n30406 ;
  assign n30524 = x1159 | n30523 ;
  assign n30525 = ( n30427 & n30428 ) | ( n30427 & ~n30524 ) | ( n30428 & ~n30524 ) ;
  assign n30526 = ( x648 & n30522 ) | ( x648 & ~n30525 ) | ( n30522 & ~n30525 ) ;
  assign n30527 = ~n30522 & n30526 ;
  assign n30429 = x619 | n30406 ;
  assign n30430 = ( x1159 & n30428 ) | ( x1159 & n30429 ) | ( n30428 & n30429 ) ;
  assign n30431 = ~n30428 & n30430 ;
  assign n30515 = x619 & ~n30514 ;
  assign n30516 = x1159 | n30515 ;
  assign n30517 = ( n30511 & n30512 ) | ( n30511 & ~n30516 ) | ( n30512 & ~n30516 ) ;
  assign n30518 = ( x648 & ~n30431 ) | ( x648 & n30517 ) | ( ~n30431 & n30517 ) ;
  assign n30519 = n30431 | n30518 ;
  assign n30528 = n30527 ^ n30519 ^ 1'b0 ;
  assign n30529 = ( x789 & ~n30519 ) | ( x789 & n30527 ) | ( ~n30519 & n30527 ) ;
  assign n30530 = ( x789 & ~n30528 ) | ( x789 & n30529 ) | ( ~n30528 & n30529 ) ;
  assign n30531 = ( x789 & n30511 ) | ( x789 & ~n30530 ) | ( n30511 & ~n30530 ) ;
  assign n30532 = ~n30530 & n30531 ;
  assign n30533 = ~x626 & n30532 ;
  assign n30534 = n30406 ^ n16279 ^ 1'b0 ;
  assign n30535 = ( n30406 & n30514 ) | ( n30406 & ~n30534 ) | ( n30514 & ~n30534 ) ;
  assign n30536 = x626 & n30535 ;
  assign n30537 = ( x641 & ~n30533 ) | ( x641 & n30536 ) | ( ~n30533 & n30536 ) ;
  assign n30538 = n30533 | n30537 ;
  assign n30539 = ~x626 & n30406 ;
  assign n30540 = n30431 | n30525 ;
  assign n30541 = n30427 ^ x789 ^ 1'b0 ;
  assign n30542 = ( n30427 & n30540 ) | ( n30427 & n30541 ) | ( n30540 & n30541 ) ;
  assign n30543 = x626 & n30542 ;
  assign n30544 = ( x641 & ~n30539 ) | ( x641 & n30543 ) | ( ~n30539 & n30543 ) ;
  assign n30545 = n30539 | n30544 ;
  assign n30546 = ~x626 & n30535 ;
  assign n30547 = x626 & n30532 ;
  assign n30548 = ( x641 & n30546 ) | ( x641 & ~n30547 ) | ( n30546 & ~n30547 ) ;
  assign n30549 = ~n30546 & n30548 ;
  assign n30550 = x1158 & ~n30549 ;
  assign n30551 = n30545 & n30550 ;
  assign n30552 = ~x626 & n30542 ;
  assign n30553 = x626 & n30406 ;
  assign n30554 = x641 & ~n30553 ;
  assign n30555 = n30554 ^ n30552 ^ 1'b0 ;
  assign n30556 = ( n30552 & n30554 ) | ( n30552 & n30555 ) | ( n30554 & n30555 ) ;
  assign n30557 = ( x1158 & ~n30552 ) | ( x1158 & n30556 ) | ( ~n30552 & n30556 ) ;
  assign n30558 = ~n30551 & n30557 ;
  assign n30559 = ( n30538 & n30551 ) | ( n30538 & ~n30558 ) | ( n30551 & ~n30558 ) ;
  assign n30560 = n30532 ^ x788 ^ 1'b0 ;
  assign n30561 = ( n30532 & n30559 ) | ( n30532 & n30560 ) | ( n30559 & n30560 ) ;
  assign n30562 = x628 & ~n30561 ;
  assign n30563 = n30406 ^ n16518 ^ 1'b0 ;
  assign n30564 = ( n30406 & n30542 ) | ( n30406 & ~n30563 ) | ( n30542 & ~n30563 ) ;
  assign n30565 = x628 | n30564 ;
  assign n30566 = ( x1156 & n30562 ) | ( x1156 & n30565 ) | ( n30562 & n30565 ) ;
  assign n30567 = ~n30562 & n30566 ;
  assign n30568 = x628 & ~n30406 ;
  assign n30569 = x1156 | n30568 ;
  assign n30570 = n30406 ^ n16318 ^ 1'b0 ;
  assign n30571 = ( n30406 & n30535 ) | ( n30406 & ~n30570 ) | ( n30535 & ~n30570 ) ;
  assign n30572 = x628 & ~n30571 ;
  assign n30573 = ( ~n30569 & n30571 ) | ( ~n30569 & n30572 ) | ( n30571 & n30572 ) ;
  assign n30574 = ( x629 & n30567 ) | ( x629 & ~n30573 ) | ( n30567 & ~n30573 ) ;
  assign n30575 = ~n30567 & n30574 ;
  assign n30576 = x628 | n30406 ;
  assign n30577 = ( x1156 & n30572 ) | ( x1156 & n30576 ) | ( n30572 & n30576 ) ;
  assign n30578 = ~n30572 & n30577 ;
  assign n30579 = x629 | n30578 ;
  assign n30580 = x628 & ~n30564 ;
  assign n30581 = x1156 | n30580 ;
  assign n30582 = ( n30561 & n30562 ) | ( n30561 & ~n30581 ) | ( n30562 & ~n30581 ) ;
  assign n30583 = ( ~n30575 & n30579 ) | ( ~n30575 & n30582 ) | ( n30579 & n30582 ) ;
  assign n30584 = ~n30575 & n30583 ;
  assign n30585 = n30561 ^ x792 ^ 1'b0 ;
  assign n30586 = ( n30561 & n30584 ) | ( n30561 & n30585 ) | ( n30584 & n30585 ) ;
  assign n30587 = x647 & ~n30586 ;
  assign n30588 = n30406 ^ n16339 ^ 1'b0 ;
  assign n30589 = ( n30406 & n30564 ) | ( n30406 & ~n30588 ) | ( n30564 & ~n30588 ) ;
  assign n30590 = x647 | n30589 ;
  assign n30591 = ( x1157 & n30587 ) | ( x1157 & n30590 ) | ( n30587 & n30590 ) ;
  assign n30592 = ~n30587 & n30591 ;
  assign n30593 = x647 & ~n30406 ;
  assign n30594 = x1157 | n30593 ;
  assign n30595 = n30573 | n30578 ;
  assign n30596 = n30571 ^ x792 ^ 1'b0 ;
  assign n30597 = ( n30571 & n30595 ) | ( n30571 & n30596 ) | ( n30595 & n30596 ) ;
  assign n30598 = x647 & ~n30597 ;
  assign n30599 = ( ~n30594 & n30597 ) | ( ~n30594 & n30598 ) | ( n30597 & n30598 ) ;
  assign n30600 = ( x630 & n30592 ) | ( x630 & ~n30599 ) | ( n30592 & ~n30599 ) ;
  assign n30601 = ~n30592 & n30600 ;
  assign n30602 = x647 | n30406 ;
  assign n30603 = ( x1157 & n30598 ) | ( x1157 & n30602 ) | ( n30598 & n30602 ) ;
  assign n30604 = ~n30598 & n30603 ;
  assign n30605 = x630 | n30604 ;
  assign n30606 = x647 & ~n30589 ;
  assign n30607 = x1157 | n30606 ;
  assign n30608 = ( n30586 & n30587 ) | ( n30586 & ~n30607 ) | ( n30587 & ~n30607 ) ;
  assign n30609 = ( ~n30601 & n30605 ) | ( ~n30601 & n30608 ) | ( n30605 & n30608 ) ;
  assign n30610 = ~n30601 & n30609 ;
  assign n30611 = n30586 ^ x787 ^ 1'b0 ;
  assign n30612 = ( n30586 & n30610 ) | ( n30586 & n30611 ) | ( n30610 & n30611 ) ;
  assign n30613 = x644 & ~n30612 ;
  assign n30614 = n30599 | n30604 ;
  assign n30615 = n30597 ^ x787 ^ 1'b0 ;
  assign n30616 = ( n30597 & n30614 ) | ( n30597 & n30615 ) | ( n30614 & n30615 ) ;
  assign n30617 = x644 | n30616 ;
  assign n30618 = ( x715 & n30613 ) | ( x715 & n30617 ) | ( n30613 & n30617 ) ;
  assign n30619 = ~n30613 & n30618 ;
  assign n30620 = x644 | n30406 ;
  assign n30621 = n30406 ^ n16376 ^ 1'b0 ;
  assign n30622 = ( n30406 & n30589 ) | ( n30406 & ~n30621 ) | ( n30589 & ~n30621 ) ;
  assign n30623 = x644 & ~n30622 ;
  assign n30624 = ( x715 & n30620 ) | ( x715 & ~n30623 ) | ( n30620 & ~n30623 ) ;
  assign n30625 = ~x715 & n30624 ;
  assign n30626 = ( x1160 & n30619 ) | ( x1160 & ~n30625 ) | ( n30619 & ~n30625 ) ;
  assign n30627 = ~n30619 & n30626 ;
  assign n30628 = x644 & ~n30406 ;
  assign n30629 = x715 & ~n30628 ;
  assign n30630 = ( n30622 & n30623 ) | ( n30622 & n30629 ) | ( n30623 & n30629 ) ;
  assign n30631 = x644 & ~n30616 ;
  assign n30632 = x715 | n30631 ;
  assign n30633 = ( n30612 & n30613 ) | ( n30612 & ~n30632 ) | ( n30613 & ~n30632 ) ;
  assign n30634 = ( x1160 & ~n30630 ) | ( x1160 & n30633 ) | ( ~n30630 & n30633 ) ;
  assign n30635 = n30630 | n30634 ;
  assign n30636 = ( x790 & n30627 ) | ( x790 & n30635 ) | ( n30627 & n30635 ) ;
  assign n30637 = ~n30627 & n30636 ;
  assign n30638 = ~x790 & n30612 ;
  assign n30639 = ( n7318 & ~n30637 ) | ( n7318 & n30638 ) | ( ~n30637 & n30638 ) ;
  assign n30640 = n30637 | n30639 ;
  assign n30641 = x194 | n1611 ;
  assign n30642 = x748 & n15591 ;
  assign n30643 = n30641 & ~n30642 ;
  assign n30644 = n16397 | n30643 ;
  assign n30645 = n16402 | n30643 ;
  assign n30646 = x1155 & n30645 ;
  assign n30647 = n16405 | n30644 ;
  assign n30648 = ~x1155 & n30647 ;
  assign n30649 = n30646 | n30648 ;
  assign n30650 = n30644 ^ x785 ^ 1'b0 ;
  assign n30651 = ( n30644 & n30649 ) | ( n30644 & n30650 ) | ( n30649 & n30650 ) ;
  assign n30652 = n16411 | n30651 ;
  assign n30653 = x1154 & n30652 ;
  assign n30654 = n16414 | n30651 ;
  assign n30655 = ~x1154 & n30654 ;
  assign n30656 = n30653 | n30655 ;
  assign n30657 = n30651 ^ x781 ^ 1'b0 ;
  assign n30658 = ( n30651 & n30656 ) | ( n30651 & n30657 ) | ( n30656 & n30657 ) ;
  assign n30659 = x619 & ~n30658 ;
  assign n30660 = x619 | n30641 ;
  assign n30661 = ( x1159 & n30659 ) | ( x1159 & n30660 ) | ( n30659 & n30660 ) ;
  assign n30662 = ~n30659 & n30661 ;
  assign n30663 = x619 & ~n30641 ;
  assign n30664 = x1159 | n30663 ;
  assign n30665 = ( n30658 & n30659 ) | ( n30658 & ~n30664 ) | ( n30659 & ~n30664 ) ;
  assign n30666 = n30662 | n30665 ;
  assign n30667 = n30658 ^ x789 ^ 1'b0 ;
  assign n30668 = ( n30658 & n30666 ) | ( n30658 & n30667 ) | ( n30666 & n30667 ) ;
  assign n30669 = n30641 ^ n16518 ^ 1'b0 ;
  assign n30670 = ( n30641 & n30668 ) | ( n30641 & ~n30669 ) | ( n30668 & ~n30669 ) ;
  assign n30671 = n30641 ^ n16339 ^ 1'b0 ;
  assign n30672 = ( n30641 & n30670 ) | ( n30641 & ~n30671 ) | ( n30670 & ~n30671 ) ;
  assign n30673 = n19055 & n30672 ;
  assign n30674 = x647 & ~n30641 ;
  assign n30675 = x1157 | n30674 ;
  assign n30676 = x730 & n15778 ;
  assign n30677 = n30641 & ~n30676 ;
  assign n30678 = ~x1153 & n30641 ;
  assign n30679 = ~x625 & n30676 ;
  assign n30680 = n30678 & ~n30679 ;
  assign n30681 = ( x1153 & n30677 ) | ( x1153 & n30679 ) | ( n30677 & n30679 ) ;
  assign n30682 = n30680 | n30681 ;
  assign n30683 = n30677 ^ x778 ^ 1'b0 ;
  assign n30684 = ( n30677 & n30682 ) | ( n30677 & n30683 ) | ( n30682 & n30683 ) ;
  assign n30685 = n16447 | n30684 ;
  assign n30686 = n16449 | n30685 ;
  assign n30687 = n16451 | n30686 ;
  assign n30688 = n16530 | n30687 ;
  assign n30689 = n16560 | n30688 ;
  assign n30690 = ( x647 & ~n30675 ) | ( x647 & n30689 ) | ( ~n30675 & n30689 ) ;
  assign n30691 = ~n30675 & n30690 ;
  assign n30692 = n30641 ^ x647 ^ 1'b0 ;
  assign n30693 = ( n30641 & n30689 ) | ( n30641 & n30692 ) | ( n30689 & n30692 ) ;
  assign n30694 = x1157 & n30693 ;
  assign n30695 = ( n16375 & n30691 ) | ( n16375 & n30694 ) | ( n30691 & n30694 ) ;
  assign n30696 = ( x787 & n30673 ) | ( x787 & n30695 ) | ( n30673 & n30695 ) ;
  assign n30697 = n30695 ^ n30673 ^ 1'b0 ;
  assign n30698 = ( x787 & n30696 ) | ( x787 & n30697 ) | ( n30696 & n30697 ) ;
  assign n30699 = ~x626 & n30641 ;
  assign n30700 = x626 & n30668 ;
  assign n30701 = ( n22317 & n30699 ) | ( n22317 & ~n30700 ) | ( n30699 & ~n30700 ) ;
  assign n30702 = ~n30699 & n30701 ;
  assign n30703 = ~x626 & n30668 ;
  assign n30704 = x626 & n30641 ;
  assign n30705 = ( n22322 & n30703 ) | ( n22322 & ~n30704 ) | ( n30703 & ~n30704 ) ;
  assign n30706 = ~n30703 & n30705 ;
  assign n30707 = n30687 & ~n30706 ;
  assign n30708 = ( n16459 & n30706 ) | ( n16459 & ~n30707 ) | ( n30706 & ~n30707 ) ;
  assign n30709 = ( x788 & n30702 ) | ( x788 & n30708 ) | ( n30702 & n30708 ) ;
  assign n30710 = n30708 ^ n30702 ^ 1'b0 ;
  assign n30711 = ( x788 & n30709 ) | ( x788 & n30710 ) | ( n30709 & n30710 ) ;
  assign n30712 = n15524 | n30677 ;
  assign n30713 = n30643 & n30712 ;
  assign n30714 = x625 & ~n30712 ;
  assign n30715 = ( n30678 & n30713 ) | ( n30678 & n30714 ) | ( n30713 & n30714 ) ;
  assign n30716 = ( x608 & n30681 ) | ( x608 & ~n30715 ) | ( n30681 & ~n30715 ) ;
  assign n30717 = n30715 | n30716 ;
  assign n30718 = x1153 & n30643 ;
  assign n30719 = ~n30714 & n30718 ;
  assign n30720 = x608 & ~n30680 ;
  assign n30721 = n30717 & ~n30720 ;
  assign n30722 = ( n30717 & n30719 ) | ( n30717 & n30721 ) | ( n30719 & n30721 ) ;
  assign n30723 = n30713 ^ x778 ^ 1'b0 ;
  assign n30724 = ( n30713 & n30722 ) | ( n30713 & n30723 ) | ( n30722 & n30723 ) ;
  assign n30725 = x609 & ~n30724 ;
  assign n30726 = x609 | n30684 ;
  assign n30727 = ( x1155 & n30725 ) | ( x1155 & n30726 ) | ( n30725 & n30726 ) ;
  assign n30728 = ~n30725 & n30727 ;
  assign n30729 = ( x660 & n30648 ) | ( x660 & ~n30728 ) | ( n30648 & ~n30728 ) ;
  assign n30730 = ~n30648 & n30729 ;
  assign n30731 = x660 | n30646 ;
  assign n30732 = x609 & ~n30684 ;
  assign n30733 = x1155 | n30732 ;
  assign n30734 = ( n30724 & n30725 ) | ( n30724 & ~n30733 ) | ( n30725 & ~n30733 ) ;
  assign n30735 = ( ~n30730 & n30731 ) | ( ~n30730 & n30734 ) | ( n30731 & n30734 ) ;
  assign n30736 = ~n30730 & n30735 ;
  assign n30737 = n30724 ^ x785 ^ 1'b0 ;
  assign n30738 = ( n30724 & n30736 ) | ( n30724 & n30737 ) | ( n30736 & n30737 ) ;
  assign n30739 = x618 & ~n30738 ;
  assign n30740 = x618 | n30685 ;
  assign n30741 = ( x1154 & n30739 ) | ( x1154 & n30740 ) | ( n30739 & n30740 ) ;
  assign n30742 = ~n30739 & n30741 ;
  assign n30743 = ( x627 & n30655 ) | ( x627 & ~n30742 ) | ( n30655 & ~n30742 ) ;
  assign n30744 = ~n30655 & n30743 ;
  assign n30745 = x627 | n30653 ;
  assign n30746 = x618 & ~n30685 ;
  assign n30747 = x1154 | n30746 ;
  assign n30748 = ( n30738 & n30739 ) | ( n30738 & ~n30747 ) | ( n30739 & ~n30747 ) ;
  assign n30749 = ( ~n30744 & n30745 ) | ( ~n30744 & n30748 ) | ( n30745 & n30748 ) ;
  assign n30750 = ~n30744 & n30749 ;
  assign n30751 = n30738 ^ x781 ^ 1'b0 ;
  assign n30752 = ( n30738 & n30750 ) | ( n30738 & n30751 ) | ( n30750 & n30751 ) ;
  assign n30753 = ~x789 & n30752 ;
  assign n30754 = x619 & ~n30686 ;
  assign n30755 = x1159 | n30754 ;
  assign n30756 = x619 & ~n30752 ;
  assign n30757 = ( n30752 & ~n30755 ) | ( n30752 & n30756 ) | ( ~n30755 & n30756 ) ;
  assign n30758 = ( x648 & n30662 ) | ( x648 & ~n30757 ) | ( n30662 & ~n30757 ) ;
  assign n30759 = n30757 | n30758 ;
  assign n30760 = x619 | n30686 ;
  assign n30761 = x1159 & ~n30756 ;
  assign n30762 = n30760 & n30761 ;
  assign n30763 = ( x648 & n30665 ) | ( x648 & ~n30762 ) | ( n30665 & ~n30762 ) ;
  assign n30764 = ~n30665 & n30763 ;
  assign n30765 = x789 & ~n30764 ;
  assign n30766 = n30759 & n30765 ;
  assign n30767 = ( n16519 & ~n30753 ) | ( n16519 & n30766 ) | ( ~n30753 & n30766 ) ;
  assign n30768 = n30753 | n30767 ;
  assign n30769 = n30768 ^ n30711 ^ 1'b0 ;
  assign n30770 = ( n30711 & n30768 ) | ( n30711 & n30769 ) | ( n30768 & n30769 ) ;
  assign n30771 = ( n18482 & ~n30711 ) | ( n18482 & n30770 ) | ( ~n30711 & n30770 ) ;
  assign n30772 = n19208 | n30688 ;
  assign n30773 = n16556 & ~n30670 ;
  assign n30774 = x629 & ~n30773 ;
  assign n30775 = n30772 & n30774 ;
  assign n30776 = n16557 & ~n30670 ;
  assign n30777 = n19212 & ~n30688 ;
  assign n30778 = n30776 | n30777 ;
  assign n30779 = ( x629 & ~n30775 ) | ( x629 & n30778 ) | ( ~n30775 & n30778 ) ;
  assign n30780 = ~n30775 & n30779 ;
  assign n30781 = ( x792 & ~n19206 ) | ( x792 & n30780 ) | ( ~n19206 & n30780 ) ;
  assign n30782 = ( n18484 & n19206 ) | ( n18484 & n30781 ) | ( n19206 & n30781 ) ;
  assign n30783 = ( n30698 & n30771 ) | ( n30698 & ~n30782 ) | ( n30771 & ~n30782 ) ;
  assign n30784 = n30783 ^ n30771 ^ 1'b0 ;
  assign n30785 = ( n30698 & n30783 ) | ( n30698 & ~n30784 ) | ( n30783 & ~n30784 ) ;
  assign n30786 = x790 | n30785 ;
  assign n30787 = x644 & ~n30785 ;
  assign n30788 = ( x787 & n30691 ) | ( x787 & ~n30694 ) | ( n30691 & ~n30694 ) ;
  assign n30789 = ~n30691 & n30788 ;
  assign n30790 = ( x787 & n30689 ) | ( x787 & ~n30789 ) | ( n30689 & ~n30789 ) ;
  assign n30791 = ~n30789 & n30790 ;
  assign n30792 = x644 | n30791 ;
  assign n30793 = ( x715 & n30787 ) | ( x715 & n30792 ) | ( n30787 & n30792 ) ;
  assign n30794 = ~n30787 & n30793 ;
  assign n30795 = x644 | n30641 ;
  assign n30796 = n30641 ^ n16376 ^ 1'b0 ;
  assign n30797 = ( n30641 & n30672 ) | ( n30641 & ~n30796 ) | ( n30672 & ~n30796 ) ;
  assign n30798 = x644 & ~n30797 ;
  assign n30799 = ( x715 & n30795 ) | ( x715 & ~n30798 ) | ( n30795 & ~n30798 ) ;
  assign n30800 = ~x715 & n30799 ;
  assign n30801 = ( x1160 & n30794 ) | ( x1160 & ~n30800 ) | ( n30794 & ~n30800 ) ;
  assign n30802 = ~n30794 & n30801 ;
  assign n30803 = x644 & ~n30641 ;
  assign n30804 = x715 & ~n30803 ;
  assign n30805 = ( n30797 & n30798 ) | ( n30797 & n30804 ) | ( n30798 & n30804 ) ;
  assign n30806 = x644 & ~n30791 ;
  assign n30807 = x715 | n30806 ;
  assign n30808 = ( n30785 & n30787 ) | ( n30785 & ~n30807 ) | ( n30787 & ~n30807 ) ;
  assign n30809 = ( x1160 & ~n30805 ) | ( x1160 & n30808 ) | ( ~n30805 & n30808 ) ;
  assign n30810 = n30805 | n30809 ;
  assign n30811 = x790 & ~n30810 ;
  assign n30812 = ( x790 & n30802 ) | ( x790 & n30811 ) | ( n30802 & n30811 ) ;
  assign n30813 = x832 & ~n30812 ;
  assign n30814 = n30786 & n30813 ;
  assign n30815 = ~x194 & n7318 ;
  assign n30816 = x832 | n30815 ;
  assign n30817 = ~n30814 & n30816 ;
  assign n30818 = ( n30640 & n30814 ) | ( n30640 & ~n30817 ) | ( n30814 & ~n30817 ) ;
  assign n30819 = x138 | n15187 ;
  assign n30820 = x196 | n30819 ;
  assign n30821 = x195 & n30820 ;
  assign n30822 = n8050 & ~n14750 ;
  assign n30823 = x171 & n7980 ;
  assign n30824 = ( x299 & n30822 ) | ( x299 & n30823 ) | ( n30822 & n30823 ) ;
  assign n30825 = n30823 ^ n30822 ^ 1'b0 ;
  assign n30826 = ( x299 & n30824 ) | ( x299 & n30825 ) | ( n30824 & n30825 ) ;
  assign n30827 = x192 & n15152 ;
  assign n30828 = ~x192 & n15139 ;
  assign n30829 = x232 & ~n30828 ;
  assign n30830 = ( n30826 & ~n30827 ) | ( n30826 & n30829 ) | ( ~n30827 & n30829 ) ;
  assign n30831 = ~n30826 & n30830 ;
  assign n30832 = ( x39 & n15142 ) | ( x39 & ~n30831 ) | ( n15142 & ~n30831 ) ;
  assign n30833 = ~x39 & n30832 ;
  assign n30834 = ~x192 & n15116 ;
  assign n30835 = x171 | n7699 ;
  assign n30836 = n7669 & ~n30835 ;
  assign n30837 = ( n7669 & ~n15124 ) | ( n7669 & n30836 ) | ( ~n15124 & n30836 ) ;
  assign n30838 = ~n30834 & n30837 ;
  assign n30839 = ( n7671 & n30834 ) | ( n7671 & ~n30838 ) | ( n30834 & ~n30838 ) ;
  assign n30840 = x192 & n15129 ;
  assign n30841 = ( x232 & n30839 ) | ( x232 & n30840 ) | ( n30839 & n30840 ) ;
  assign n30842 = n30840 ^ n30839 ^ 1'b0 ;
  assign n30843 = ( x232 & n30841 ) | ( x232 & n30842 ) | ( n30841 & n30842 ) ;
  assign n30844 = ( x39 & n15123 ) | ( x39 & n30843 ) | ( n15123 & n30843 ) ;
  assign n30845 = n30843 ^ n15123 ^ 1'b0 ;
  assign n30846 = ( x39 & n30844 ) | ( x39 & n30845 ) | ( n30844 & n30845 ) ;
  assign n30847 = ( x38 & x100 ) | ( x38 & ~n30846 ) | ( x100 & ~n30846 ) ;
  assign n30848 = n30846 | n30847 ;
  assign n30849 = ( ~x87 & n30833 ) | ( ~x87 & n30848 ) | ( n30833 & n30848 ) ;
  assign n30850 = ~x87 & n30849 ;
  assign n30851 = ( ~x92 & n15113 ) | ( ~x92 & n30850 ) | ( n15113 & n30850 ) ;
  assign n30852 = ~x92 & n30851 ;
  assign n30853 = ( ~x55 & n15112 ) | ( ~x55 & n30852 ) | ( n15112 & n30852 ) ;
  assign n30854 = ~x55 & n30853 ;
  assign n30855 = ( ~n2109 & n15196 ) | ( ~n2109 & n30854 ) | ( n15196 & n30854 ) ;
  assign n30856 = ~n2109 & n30855 ;
  assign n30857 = ( n8298 & n30821 ) | ( n8298 & ~n30856 ) | ( n30821 & ~n30856 ) ;
  assign n30858 = ~n8298 & n30857 ;
  assign n30862 = ~n5099 & n14780 ;
  assign n30863 = n10115 | n30862 ;
  assign n30859 = n14754 & ~n15173 ;
  assign n30860 = n10112 | n14757 ;
  assign n30861 = ~n30859 & n30860 ;
  assign n30864 = n30863 ^ n30861 ^ 1'b0 ;
  assign n30865 = ( x232 & ~n30861 ) | ( x232 & n30863 ) | ( ~n30861 & n30863 ) ;
  assign n30866 = ( x232 & ~n30864 ) | ( x232 & n30865 ) | ( ~n30864 & n30865 ) ;
  assign n30867 = x232 | n10116 ;
  assign n30868 = x39 & ~n30867 ;
  assign n30869 = ( x39 & n30866 ) | ( x39 & n30868 ) | ( n30866 & n30868 ) ;
  assign n30870 = n12242 & ~n14782 ;
  assign n30871 = x39 | n30870 ;
  assign n30872 = ( n9901 & ~n30821 ) | ( n9901 & n30871 ) | ( ~n30821 & n30871 ) ;
  assign n30873 = ~n9901 & n30872 ;
  assign n30874 = ( n30858 & ~n30869 ) | ( n30858 & n30873 ) | ( ~n30869 & n30873 ) ;
  assign n30875 = n30869 ^ n30858 ^ 1'b0 ;
  assign n30876 = ( n30858 & n30874 ) | ( n30858 & ~n30875 ) | ( n30874 & ~n30875 ) ;
  assign n30877 = x38 | x194 ;
  assign n30878 = n15122 ^ x232 ^ 1'b0 ;
  assign n30879 = x170 | n7699 ;
  assign n30880 = n7669 & ~n30879 ;
  assign n30881 = ( n7669 & ~n15124 ) | ( n7669 & n30880 ) | ( ~n15124 & n30880 ) ;
  assign n30882 = ( n7671 & n15116 ) | ( n7671 & ~n30881 ) | ( n15116 & ~n30881 ) ;
  assign n30883 = n30881 ^ n15116 ^ 1'b0 ;
  assign n30884 = ( n15116 & n30882 ) | ( n15116 & ~n30883 ) | ( n30882 & ~n30883 ) ;
  assign n30885 = ( n15122 & n30878 ) | ( n15122 & n30884 ) | ( n30878 & n30884 ) ;
  assign n30886 = x39 & n30885 ;
  assign n30887 = n30877 | n30886 ;
  assign n30888 = n15139 | n30887 ;
  assign n30889 = x232 & n15129 ;
  assign n30890 = n30885 | n30889 ;
  assign n30891 = x39 & n30890 ;
  assign n30892 = ( x38 & x194 ) | ( x38 & ~n30891 ) | ( x194 & ~n30891 ) ;
  assign n30893 = ~x38 & n30892 ;
  assign n30894 = ~n15152 & n30893 ;
  assign n30895 = n30888 & ~n30894 ;
  assign n30896 = n8050 & ~n14876 ;
  assign n30897 = x170 & n7980 ;
  assign n30898 = ( x299 & n30896 ) | ( x299 & n30897 ) | ( n30896 & n30897 ) ;
  assign n30899 = n30897 ^ n30896 ^ 1'b0 ;
  assign n30900 = ( x299 & n30898 ) | ( x299 & n30899 ) | ( n30898 & n30899 ) ;
  assign n30901 = ( x232 & n30895 ) | ( x232 & ~n30900 ) | ( n30895 & ~n30900 ) ;
  assign n30902 = ~n30895 & n30901 ;
  assign n30903 = ( ~x39 & n15139 ) | ( ~x39 & n15141 ) | ( n15139 & n15141 ) ;
  assign n30904 = ~x39 & n30903 ;
  assign n30905 = n30887 & ~n30893 ;
  assign n30906 = n30904 | n30905 ;
  assign n30907 = n30906 ^ n30902 ^ 1'b0 ;
  assign n30908 = ( n30902 & n30906 ) | ( n30902 & n30907 ) | ( n30906 & n30907 ) ;
  assign n30909 = ( x100 & ~n30902 ) | ( x100 & n30908 ) | ( ~n30902 & n30908 ) ;
  assign n30910 = x87 | n30909 ;
  assign n30911 = ( ~x87 & n15113 ) | ( ~x87 & n30910 ) | ( n15113 & n30910 ) ;
  assign n30912 = x92 | n30911 ;
  assign n30913 = ( ~x92 & n15112 ) | ( ~x92 & n30912 ) | ( n15112 & n30912 ) ;
  assign n30914 = x55 | n30913 ;
  assign n30915 = ( ~x55 & n15196 ) | ( ~x55 & n30914 ) | ( n15196 & n30914 ) ;
  assign n30916 = n2109 | n30915 ;
  assign n30917 = ( ~n2109 & n8298 ) | ( ~n2109 & n30916 ) | ( n8298 & n30916 ) ;
  assign n30918 = x195 & ~x196 ;
  assign n30919 = n30917 & n30918 ;
  assign n30923 = ~x170 & n8182 ;
  assign n30924 = n15172 | n30923 ;
  assign n30925 = n11620 & n30924 ;
  assign n30926 = n11618 & n15172 ;
  assign n30927 = x232 & ~n30926 ;
  assign n30928 = n30867 & ~n30927 ;
  assign n30929 = ( n30867 & n30925 ) | ( n30867 & n30928 ) | ( n30925 & n30928 ) ;
  assign n30930 = x39 & ~n30929 ;
  assign n30920 = n12242 & ~n14928 ;
  assign n30921 = ( ~x38 & x39 ) | ( ~x38 & n30920 ) | ( x39 & n30920 ) ;
  assign n30922 = ~x38 & n30921 ;
  assign n30931 = n30930 ^ n30922 ^ 1'b0 ;
  assign n30932 = ( x194 & ~n30922 ) | ( x194 & n30930 ) | ( ~n30922 & n30930 ) ;
  assign n30933 = ( x194 & ~n30931 ) | ( x194 & n30932 ) | ( ~n30931 & n30932 ) ;
  assign n30934 = n12242 & ~n14877 ;
  assign n30935 = ( ~x38 & x39 ) | ( ~x38 & n30934 ) | ( x39 & n30934 ) ;
  assign n30936 = ~x38 & n30935 ;
  assign n30937 = x299 & n30929 ;
  assign n30938 = ( x39 & n10113 ) | ( x39 & ~n30937 ) | ( n10113 & ~n30937 ) ;
  assign n30939 = ~n10113 & n30938 ;
  assign n30940 = ( x194 & n30936 ) | ( x194 & ~n30939 ) | ( n30936 & ~n30939 ) ;
  assign n30941 = n30940 ^ n30936 ^ 1'b0 ;
  assign n30942 = ( x194 & n30940 ) | ( x194 & ~n30941 ) | ( n30940 & ~n30941 ) ;
  assign n30943 = ( n8793 & ~n30933 ) | ( n8793 & n30942 ) | ( ~n30933 & n30942 ) ;
  assign n30944 = ~n8793 & n30943 ;
  assign n30945 = n30918 | n30944 ;
  assign n30946 = ( n30819 & ~n30919 ) | ( n30819 & n30945 ) | ( ~n30919 & n30945 ) ;
  assign n30947 = ~n30819 & n30946 ;
  assign n30948 = x196 & n30917 ;
  assign n30949 = x196 | n30944 ;
  assign n30950 = n30819 & n30949 ;
  assign n30951 = ( n30947 & ~n30948 ) | ( n30947 & n30950 ) | ( ~n30948 & n30950 ) ;
  assign n30952 = n30948 ^ n30947 ^ 1'b0 ;
  assign n30953 = ( n30947 & n30951 ) | ( n30947 & ~n30952 ) | ( n30951 & ~n30952 ) ;
  assign n30954 = x197 | n1611 ;
  assign n30955 = x832 & n30954 ;
  assign n30957 = ~x767 & x947 ;
  assign n30975 = n15644 & ~n30957 ;
  assign n30976 = x197 & ~n15653 ;
  assign n30977 = ( x38 & n30975 ) | ( x38 & ~n30976 ) | ( n30975 & ~n30976 ) ;
  assign n30978 = ~n30975 & n30977 ;
  assign n30956 = x197 | n15332 ;
  assign n30958 = n15332 & n30957 ;
  assign n30959 = ( x39 & n30956 ) | ( x39 & ~n30958 ) | ( n30956 & ~n30958 ) ;
  assign n30960 = ~x39 & n30959 ;
  assign n30961 = ~x197 & x767 ;
  assign n30962 = ~n15486 & n30961 ;
  assign n30963 = x39 & ~n30962 ;
  assign n30964 = x197 | n15484 ;
  assign n30965 = ~n19428 & n30964 ;
  assign n30966 = x197 & n19516 ;
  assign n30967 = x299 & ~n30966 ;
  assign n30968 = x197 | n19451 ;
  assign n30969 = n30967 & n30968 ;
  assign n30970 = ( x767 & ~n30965 ) | ( x767 & n30969 ) | ( ~n30965 & n30969 ) ;
  assign n30971 = n30965 | n30970 ;
  assign n30972 = n30963 & n30971 ;
  assign n30973 = ( x38 & ~n30960 ) | ( x38 & n30972 ) | ( ~n30960 & n30972 ) ;
  assign n30974 = n30960 | n30973 ;
  assign n30979 = n30978 ^ n30974 ^ 1'b0 ;
  assign n30980 = ( x698 & ~n30974 ) | ( x698 & n30978 ) | ( ~n30974 & n30978 ) ;
  assign n30981 = ( x698 & ~n30979 ) | ( x698 & n30980 ) | ( ~n30979 & n30980 ) ;
  assign n30982 = x767 & x947 ;
  assign n30983 = ( x39 & n19568 ) | ( x39 & ~n30982 ) | ( n19568 & ~n30982 ) ;
  assign n30984 = ~x39 & n30983 ;
  assign n30985 = x197 | n15644 ;
  assign n30986 = x38 & n30985 ;
  assign n30987 = n30986 ^ n30984 ^ 1'b0 ;
  assign n30988 = ( n30984 & n30986 ) | ( n30984 & n30987 ) | ( n30986 & n30987 ) ;
  assign n30989 = ( x698 & ~n30984 ) | ( x698 & n30988 ) | ( ~n30984 & n30988 ) ;
  assign n30990 = x197 & n19405 ;
  assign n30991 = x299 & ~n30990 ;
  assign n30992 = x197 | n19389 ;
  assign n30993 = n30991 & n30992 ;
  assign n30994 = ~n19409 & n30964 ;
  assign n30995 = ( x767 & n30993 ) | ( x767 & ~n30994 ) | ( n30993 & ~n30994 ) ;
  assign n30996 = ~n30993 & n30995 ;
  assign n30997 = ~x197 & n19378 ;
  assign n30998 = x197 & ~n19354 ;
  assign n30999 = ( x767 & ~n30997 ) | ( x767 & n30998 ) | ( ~n30997 & n30998 ) ;
  assign n31000 = n30997 | n30999 ;
  assign n31001 = ( x39 & n30996 ) | ( x39 & n31000 ) | ( n30996 & n31000 ) ;
  assign n31002 = ~n30996 & n31001 ;
  assign n31003 = ~n19397 & n30960 ;
  assign n31004 = ( ~x38 & n31002 ) | ( ~x38 & n31003 ) | ( n31002 & n31003 ) ;
  assign n31005 = ~x38 & n31004 ;
  assign n31006 = ( ~n30981 & n30989 ) | ( ~n30981 & n31005 ) | ( n30989 & n31005 ) ;
  assign n31007 = ~n30981 & n31006 ;
  assign n31008 = ( n2069 & n7318 ) | ( n2069 & ~n31007 ) | ( n7318 & ~n31007 ) ;
  assign n31009 = n31007 | n31008 ;
  assign n31010 = ~x197 & n8793 ;
  assign n31011 = ( x832 & n31009 ) | ( x832 & ~n31010 ) | ( n31009 & ~n31010 ) ;
  assign n31012 = ~x832 & n31011 ;
  assign n31013 = ~x698 & n19256 ;
  assign n31014 = n30957 | n31013 ;
  assign n31015 = n1611 & n31014 ;
  assign n31016 = ~n31012 & n31015 ;
  assign n31017 = ( n30955 & n31012 ) | ( n30955 & ~n31016 ) | ( n31012 & ~n31016 ) ;
  assign n31018 = x198 & ~n15337 ;
  assign n31019 = n5082 | n31018 ;
  assign n31020 = x198 & ~n15357 ;
  assign n31021 = n31019 & n31020 ;
  assign n31022 = n5081 & n15351 ;
  assign n31023 = x198 & ~n31022 ;
  assign n31024 = ~n5081 & n15353 ;
  assign n31025 = n31023 & ~n31024 ;
  assign n31026 = n5061 & n31025 ;
  assign n31027 = n31021 | n31026 ;
  assign n31028 = x215 & n31027 ;
  assign n31029 = x198 & ~n15445 ;
  assign n31030 = n31018 ^ n5082 ^ 1'b0 ;
  assign n31031 = ( n31018 & n31029 ) | ( n31018 & n31030 ) | ( n31029 & n31030 ) ;
  assign n31032 = ~n5061 & n31031 ;
  assign n31033 = x198 & ~n15433 ;
  assign n31034 = n5061 & n31033 ;
  assign n31035 = ( n2263 & n31032 ) | ( n2263 & ~n31034 ) | ( n31032 & ~n31034 ) ;
  assign n31036 = ~n31032 & n31035 ;
  assign n31037 = n2263 | n31018 ;
  assign n31038 = ( x215 & ~n31036 ) | ( x215 & n31037 ) | ( ~n31036 & n31037 ) ;
  assign n31039 = ~x215 & n31038 ;
  assign n31040 = ( x299 & n31028 ) | ( x299 & ~n31039 ) | ( n31028 & ~n31039 ) ;
  assign n31041 = ~n31028 & n31040 ;
  assign n31042 = ~n2069 & n9604 ;
  assign n31043 = n5114 & n31025 ;
  assign n31044 = n31021 | n31043 ;
  assign n31045 = x223 & n31044 ;
  assign n31046 = n1359 | n31018 ;
  assign n31047 = n5114 & n31033 ;
  assign n31048 = ~n5114 & n31031 ;
  assign n31049 = ( n1359 & n31047 ) | ( n1359 & ~n31048 ) | ( n31047 & ~n31048 ) ;
  assign n31050 = ~n31047 & n31049 ;
  assign n31051 = ( x223 & n31046 ) | ( x223 & ~n31050 ) | ( n31046 & ~n31050 ) ;
  assign n31052 = ~x223 & n31051 ;
  assign n31053 = ( x299 & ~n31045 ) | ( x299 & n31052 ) | ( ~n31045 & n31052 ) ;
  assign n31054 = n31045 | n31053 ;
  assign n31055 = ( n31041 & n31042 ) | ( n31041 & n31054 ) | ( n31042 & n31054 ) ;
  assign n31056 = ~n31041 & n31055 ;
  assign n31057 = n1994 | n15332 ;
  assign n31058 = ~n17328 & n31057 ;
  assign n31059 = ~n31056 & n31058 ;
  assign n31060 = ( x198 & n31056 ) | ( x198 & ~n31059 ) | ( n31056 & ~n31059 ) ;
  assign n31061 = x39 & x198 ;
  assign n31062 = x38 & ~n31061 ;
  assign n31063 = x633 & n15524 ;
  assign n31064 = n15340 ^ x198 ^ 1'b0 ;
  assign n31065 = ( x198 & n31063 ) | ( x198 & n31064 ) | ( n31063 & n31064 ) ;
  assign n31066 = ~x39 & n31065 ;
  assign n31067 = n31062 & ~n31066 ;
  assign n31068 = x198 & ~n15330 ;
  assign n31069 = n15635 ^ x198 ^ 1'b0 ;
  assign n31070 = ( ~n15493 & n15635 ) | ( ~n15493 & n31069 ) | ( n15635 & n31069 ) ;
  assign n31071 = x603 & x633 ;
  assign n31072 = n31071 ^ n31068 ^ 1'b0 ;
  assign n31073 = ( n31068 & n31070 ) | ( n31068 & n31072 ) | ( n31070 & n31072 ) ;
  assign n31074 = x299 & n31073 ;
  assign n31075 = n15501 & ~n15505 ;
  assign n31076 = x633 & n31075 ;
  assign n31077 = n15318 | n31076 ;
  assign n31078 = ~n15503 & n31077 ;
  assign n31079 = ~x299 & n31078 ;
  assign n31080 = ( x39 & ~n31074 ) | ( x39 & n31079 ) | ( ~n31074 & n31079 ) ;
  assign n31081 = n31074 | n31080 ;
  assign n31082 = n5078 & ~n15552 ;
  assign n31083 = x633 & n15337 ;
  assign n31084 = ~n15510 & n31083 ;
  assign n31085 = n15351 & n31084 ;
  assign n31086 = x198 & ~n15351 ;
  assign n31087 = n31085 | n31086 ;
  assign n31088 = n31082 & n31087 ;
  assign n31089 = x633 & n15610 ;
  assign n31090 = n31025 | n31089 ;
  assign n31091 = ( ~n5078 & n31088 ) | ( ~n5078 & n31090 ) | ( n31088 & n31090 ) ;
  assign n31092 = n31088 ^ n5078 ^ 1'b0 ;
  assign n31093 = ( n31088 & n31091 ) | ( n31088 & ~n31092 ) | ( n31091 & ~n31092 ) ;
  assign n31094 = n5061 & ~n31093 ;
  assign n31095 = x215 & ~n31094 ;
  assign n31096 = n31018 | n31084 ;
  assign n31097 = x603 & n31096 ;
  assign n31098 = ( n31018 & n31096 ) | ( n31018 & n31097 ) | ( n31096 & n31097 ) ;
  assign n31099 = n15527 & ~n31098 ;
  assign n31100 = ~n5075 & n31096 ;
  assign n31101 = n31020 | n31085 ;
  assign n31102 = ( x603 & n31100 ) | ( x603 & n31101 ) | ( n31100 & n31101 ) ;
  assign n31103 = n31101 ^ n31100 ^ 1'b0 ;
  assign n31104 = ( x603 & n31102 ) | ( x603 & n31103 ) | ( n31102 & n31103 ) ;
  assign n31105 = ~x603 & n31018 ;
  assign n31106 = n15527 | n31105 ;
  assign n31107 = ( ~n31099 & n31104 ) | ( ~n31099 & n31106 ) | ( n31104 & n31106 ) ;
  assign n31108 = ~n31099 & n31107 ;
  assign n31109 = n31020 | n31104 ;
  assign n31110 = n31108 ^ n5078 ^ 1'b0 ;
  assign n31111 = ( n31108 & n31109 ) | ( n31108 & n31110 ) | ( n31109 & n31110 ) ;
  assign n31112 = n5061 | n31111 ;
  assign n31113 = n31095 & n31112 ;
  assign n31114 = x198 & ~n15425 ;
  assign n31115 = ~x633 & n15425 ;
  assign n31116 = ( n15518 & n31114 ) | ( n15518 & ~n31115 ) | ( n31114 & ~n31115 ) ;
  assign n31117 = x603 & n31116 ;
  assign n31118 = n5078 & ~n31114 ;
  assign n31119 = ~n31117 & n31118 ;
  assign n31120 = x603 | n15427 ;
  assign n31121 = x198 & ~n31120 ;
  assign n31122 = x603 & n15527 ;
  assign n31123 = n5075 & ~n31096 ;
  assign n31124 = n31122 & ~n31123 ;
  assign n31125 = n5075 | n31116 ;
  assign n31126 = n31124 & n31125 ;
  assign n31127 = ~n15527 & n31117 ;
  assign n31128 = ( ~n31121 & n31126 ) | ( ~n31121 & n31127 ) | ( n31126 & n31127 ) ;
  assign n31129 = n31121 | n31128 ;
  assign n31130 = ( n5078 & ~n31119 ) | ( n5078 & n31129 ) | ( ~n31119 & n31129 ) ;
  assign n31131 = ~n31119 & n31130 ;
  assign n31132 = n5061 & n31131 ;
  assign n31133 = n31096 ^ n5075 ^ 1'b0 ;
  assign n31134 = ( n31096 & n31116 ) | ( n31096 & n31133 ) | ( n31116 & n31133 ) ;
  assign n31135 = x603 & n31134 ;
  assign n31136 = ~x603 & n31029 ;
  assign n31137 = ( n5078 & n31135 ) | ( n5078 & ~n31136 ) | ( n31135 & ~n31136 ) ;
  assign n31138 = ~n31135 & n31137 ;
  assign n31139 = n5080 & n31097 ;
  assign n31140 = x642 | n31135 ;
  assign n31141 = x642 & ~n31097 ;
  assign n31142 = ( n5080 & n31140 ) | ( n5080 & ~n31141 ) | ( n31140 & ~n31141 ) ;
  assign n31143 = ~n5080 & n31142 ;
  assign n31144 = ( n31105 & ~n31139 ) | ( n31105 & n31143 ) | ( ~n31139 & n31143 ) ;
  assign n31145 = n31139 | n31144 ;
  assign n31146 = ( n5078 & ~n31138 ) | ( n5078 & n31145 ) | ( ~n31138 & n31145 ) ;
  assign n31147 = ~n31138 & n31146 ;
  assign n31148 = ~n5061 & n31147 ;
  assign n31149 = ( n2263 & n31132 ) | ( n2263 & ~n31148 ) | ( n31132 & ~n31148 ) ;
  assign n31150 = ~n31132 & n31149 ;
  assign n31151 = n2263 | n31098 ;
  assign n31152 = ( x215 & ~n31150 ) | ( x215 & n31151 ) | ( ~n31150 & n31151 ) ;
  assign n31153 = ~x215 & n31152 ;
  assign n31154 = ( x299 & n31113 ) | ( x299 & n31153 ) | ( n31113 & n31153 ) ;
  assign n31155 = n31153 ^ n31113 ^ 1'b0 ;
  assign n31156 = ( x299 & n31154 ) | ( x299 & n31155 ) | ( n31154 & n31155 ) ;
  assign n31157 = n5114 & ~n31093 ;
  assign n31158 = x223 & ~n31157 ;
  assign n31159 = n5114 | n31111 ;
  assign n31160 = n31158 & n31159 ;
  assign n31161 = n5114 & n31131 ;
  assign n31162 = ~n5114 & n31147 ;
  assign n31163 = ( n1359 & n31161 ) | ( n1359 & ~n31162 ) | ( n31161 & ~n31162 ) ;
  assign n31164 = ~n31161 & n31163 ;
  assign n31165 = n1359 | n31098 ;
  assign n31166 = ( x223 & ~n31164 ) | ( x223 & n31165 ) | ( ~n31164 & n31165 ) ;
  assign n31167 = ~x223 & n31166 ;
  assign n31168 = ( ~x299 & n31160 ) | ( ~x299 & n31167 ) | ( n31160 & n31167 ) ;
  assign n31169 = ~x299 & n31168 ;
  assign n31170 = ( x39 & n31156 ) | ( x39 & ~n31169 ) | ( n31156 & ~n31169 ) ;
  assign n31171 = ~n31156 & n31170 ;
  assign n31172 = ( x38 & n31081 ) | ( x38 & ~n31171 ) | ( n31081 & ~n31171 ) ;
  assign n31173 = n31172 ^ n31081 ^ 1'b0 ;
  assign n31174 = ( x38 & n31172 ) | ( x38 & ~n31173 ) | ( n31172 & ~n31173 ) ;
  assign n31175 = ( n2069 & ~n31067 ) | ( n2069 & n31174 ) | ( ~n31067 & n31174 ) ;
  assign n31176 = ~n2069 & n31175 ;
  assign n31177 = n31176 ^ x198 ^ 1'b0 ;
  assign n31178 = ( ~x198 & n2069 ) | ( ~x198 & n31177 ) | ( n2069 & n31177 ) ;
  assign n31179 = ( x198 & n31176 ) | ( x198 & n31178 ) | ( n31176 & n31178 ) ;
  assign n31180 = n31060 ^ n15659 ^ 1'b0 ;
  assign n31181 = ( n31060 & n31179 ) | ( n31060 & ~n31180 ) | ( n31179 & ~n31180 ) ;
  assign n31182 = ~n15659 & n31179 ;
  assign n31183 = x609 & n31182 ;
  assign n31184 = ~n15668 & n31060 ;
  assign n31185 = n31183 | n31184 ;
  assign n31186 = ~x609 & n31182 ;
  assign n31187 = n15662 & n31060 ;
  assign n31188 = n31186 | n31187 ;
  assign n31189 = n31185 ^ x1155 ^ 1'b0 ;
  assign n31190 = ( n31185 & n31188 ) | ( n31185 & ~n31189 ) | ( n31188 & ~n31189 ) ;
  assign n31191 = n31181 ^ x785 ^ 1'b0 ;
  assign n31192 = ( n31181 & n31190 ) | ( n31181 & n31191 ) | ( n31190 & n31191 ) ;
  assign n31193 = x618 & ~n31192 ;
  assign n31194 = x618 | n31060 ;
  assign n31195 = ( x1154 & n31193 ) | ( x1154 & n31194 ) | ( n31193 & n31194 ) ;
  assign n31196 = ~n31193 & n31195 ;
  assign n31197 = x618 & ~n31060 ;
  assign n31198 = x1154 | n31197 ;
  assign n31199 = ( n31192 & n31193 ) | ( n31192 & ~n31198 ) | ( n31193 & ~n31198 ) ;
  assign n31200 = n31196 | n31199 ;
  assign n31201 = n31192 ^ x781 ^ 1'b0 ;
  assign n31202 = ( n31192 & n31200 ) | ( n31192 & n31201 ) | ( n31200 & n31201 ) ;
  assign n31203 = x619 & ~n31202 ;
  assign n31204 = x619 | n31060 ;
  assign n31205 = ( x1159 & n31203 ) | ( x1159 & n31204 ) | ( n31203 & n31204 ) ;
  assign n31206 = ~n31203 & n31205 ;
  assign n31207 = x619 & ~n31060 ;
  assign n31208 = x1159 | n31207 ;
  assign n31209 = ( n31202 & n31203 ) | ( n31202 & ~n31208 ) | ( n31203 & ~n31208 ) ;
  assign n31210 = n31206 | n31209 ;
  assign n31211 = n31202 ^ x789 ^ 1'b0 ;
  assign n31212 = ( n31202 & n31210 ) | ( n31202 & n31211 ) | ( n31210 & n31211 ) ;
  assign n31213 = n31060 ^ n16518 ^ 1'b0 ;
  assign n31214 = ( n31060 & n31212 ) | ( n31060 & ~n31213 ) | ( n31212 & ~n31213 ) ;
  assign n31215 = n31060 ^ n16339 ^ 1'b0 ;
  assign n31216 = ( n31060 & n31214 ) | ( n31060 & ~n31215 ) | ( n31214 & ~n31215 ) ;
  assign n31217 = n19055 & n31216 ;
  assign n31218 = x647 & ~n31060 ;
  assign n31219 = x1157 | n31218 ;
  assign n31220 = ( x634 & n15697 ) | ( x634 & n31018 ) | ( n15697 & n31018 ) ;
  assign n31221 = n31018 | n31220 ;
  assign n31222 = n5081 | n31221 ;
  assign n31223 = n15693 & n31222 ;
  assign n31228 = x198 & ~n15844 ;
  assign n31229 = ( ~n15394 & n31029 ) | ( ~n15394 & n31228 ) | ( n31029 & n31228 ) ;
  assign n31224 = n31221 ^ n5075 ^ 1'b0 ;
  assign n31225 = ~x634 & n15425 ;
  assign n31226 = ( n15724 & n31114 ) | ( n15724 & ~n31225 ) | ( n31114 & ~n31225 ) ;
  assign n31227 = ( n31221 & n31224 ) | ( n31221 & n31226 ) | ( n31224 & n31226 ) ;
  assign n31230 = n31229 ^ n5078 ^ 1'b0 ;
  assign n31231 = ( ~n5078 & n31227 ) | ( ~n5078 & n31230 ) | ( n31227 & n31230 ) ;
  assign n31232 = ( n5078 & n31229 ) | ( n5078 & n31231 ) | ( n31229 & n31231 ) ;
  assign n31233 = n5081 & ~n31227 ;
  assign n31234 = ~n31232 & n31233 ;
  assign n31235 = ( n31223 & n31232 ) | ( n31223 & ~n31234 ) | ( n31232 & ~n31234 ) ;
  assign n31236 = ~n5061 & n31235 ;
  assign n31237 = n5081 & ~n31226 ;
  assign n31238 = n15693 & ~n31237 ;
  assign n31239 = ( n31221 & ~n31224 ) | ( n31221 & n31226 ) | ( ~n31224 & n31226 ) ;
  assign n31240 = n5081 | n31239 ;
  assign n31241 = n31238 & n31240 ;
  assign n31242 = n5078 & n31226 ;
  assign n31243 = ( ~n31228 & n31241 ) | ( ~n31228 & n31242 ) | ( n31241 & n31242 ) ;
  assign n31244 = n31228 | n31243 ;
  assign n31245 = n5061 & n31244 ;
  assign n31246 = ( n2263 & n31236 ) | ( n2263 & ~n31245 ) | ( n31236 & ~n31245 ) ;
  assign n31247 = ~n31236 & n31246 ;
  assign n31248 = ( x680 & n31018 ) | ( x680 & n31221 ) | ( n31018 & n31221 ) ;
  assign n31249 = n2263 | n31248 ;
  assign n31250 = ( x215 & ~n31247 ) | ( x215 & n31249 ) | ( ~n31247 & n31249 ) ;
  assign n31251 = ~x215 & n31250 ;
  assign n31252 = x634 & n15351 ;
  assign n31253 = n15697 & n31252 ;
  assign n31254 = n31086 | n31253 ;
  assign n31255 = n5081 & ~n31254 ;
  assign n31256 = ( n31221 & ~n31224 ) | ( n31221 & n31254 ) | ( ~n31224 & n31254 ) ;
  assign n31257 = n5081 | n31256 ;
  assign n31258 = ( n15693 & n31255 ) | ( n15693 & n31257 ) | ( n31255 & n31257 ) ;
  assign n31259 = ~n31255 & n31258 ;
  assign n31260 = ~x680 & n31025 ;
  assign n31261 = n5078 & n31254 ;
  assign n31262 = ( ~n31259 & n31260 ) | ( ~n31259 & n31261 ) | ( n31260 & n31261 ) ;
  assign n31263 = n31259 | n31262 ;
  assign n31264 = n5061 & ~n31263 ;
  assign n31265 = ( n31221 & n31224 ) | ( n31221 & n31254 ) | ( n31224 & n31254 ) ;
  assign n31266 = n5078 & n31265 ;
  assign n31267 = n5081 & ~n31265 ;
  assign n31268 = n31223 & ~n31267 ;
  assign n31269 = n31020 & n31260 ;
  assign n31270 = ( ~n31266 & n31268 ) | ( ~n31266 & n31269 ) | ( n31268 & n31269 ) ;
  assign n31271 = n31266 | n31270 ;
  assign n31272 = n5061 | n31271 ;
  assign n31273 = ( x215 & n31264 ) | ( x215 & n31272 ) | ( n31264 & n31272 ) ;
  assign n31274 = ~n31264 & n31273 ;
  assign n31275 = ( x299 & n31251 ) | ( x299 & ~n31274 ) | ( n31251 & ~n31274 ) ;
  assign n31276 = ~n31251 & n31275 ;
  assign n31277 = n5114 & ~n31263 ;
  assign n31278 = n5114 | n31271 ;
  assign n31279 = ( x223 & n31277 ) | ( x223 & n31278 ) | ( n31277 & n31278 ) ;
  assign n31280 = ~n31277 & n31279 ;
  assign n31281 = ~n5114 & n31235 ;
  assign n31282 = n5114 & n31244 ;
  assign n31283 = ( n1359 & n31281 ) | ( n1359 & ~n31282 ) | ( n31281 & ~n31282 ) ;
  assign n31284 = ~n31281 & n31283 ;
  assign n31285 = n1359 | n31248 ;
  assign n31286 = ( x223 & ~n31284 ) | ( x223 & n31285 ) | ( ~n31284 & n31285 ) ;
  assign n31287 = ~x223 & n31286 ;
  assign n31288 = ( x299 & ~n31280 ) | ( x299 & n31287 ) | ( ~n31280 & n31287 ) ;
  assign n31289 = n31280 | n31288 ;
  assign n31290 = x39 & ~n31289 ;
  assign n31291 = ( x39 & n31276 ) | ( x39 & n31290 ) | ( n31276 & n31290 ) ;
  assign n31292 = n16024 ^ x198 ^ 1'b0 ;
  assign n31293 = ( n16024 & ~n16033 ) | ( n16024 & n31292 ) | ( ~n16033 & n31292 ) ;
  assign n31294 = x634 & x680 ;
  assign n31295 = n31294 ^ n31068 ^ 1'b0 ;
  assign n31296 = ( n31068 & n31293 ) | ( n31068 & n31295 ) | ( n31293 & n31295 ) ;
  assign n31297 = x299 & n31296 ;
  assign n31298 = x198 | n16014 ;
  assign n31299 = x198 & n16031 ;
  assign n31300 = n31294 & ~n31299 ;
  assign n31301 = n31298 & n31300 ;
  assign n31302 = n15317 & ~n31301 ;
  assign n31303 = ( x198 & n31301 ) | ( x198 & ~n31302 ) | ( n31301 & ~n31302 ) ;
  assign n31304 = ~x299 & n31303 ;
  assign n31305 = ( x39 & ~n31297 ) | ( x39 & n31304 ) | ( ~n31297 & n31304 ) ;
  assign n31306 = n31297 | n31305 ;
  assign n31307 = n31306 ^ n31291 ^ 1'b0 ;
  assign n31308 = ( n31291 & n31306 ) | ( n31291 & n31307 ) | ( n31306 & n31307 ) ;
  assign n31309 = ( x38 & ~n31291 ) | ( x38 & n31308 ) | ( ~n31291 & n31308 ) ;
  assign n31310 = n31062 ^ x39 ^ 1'b0 ;
  assign n31311 = x634 & n15777 ;
  assign n31312 = ( x198 & n31064 ) | ( x198 & n31311 ) | ( n31064 & n31311 ) ;
  assign n31313 = ( x39 & n31062 ) | ( x39 & ~n31312 ) | ( n31062 & ~n31312 ) ;
  assign n31314 = ( n31062 & ~n31310 ) | ( n31062 & n31313 ) | ( ~n31310 & n31313 ) ;
  assign n31315 = ( n2069 & n31309 ) | ( n2069 & ~n31314 ) | ( n31309 & ~n31314 ) ;
  assign n31316 = ~n2069 & n31315 ;
  assign n31317 = n31316 ^ x198 ^ 1'b0 ;
  assign n31318 = ( ~x198 & n2069 ) | ( ~x198 & n31317 ) | ( n2069 & n31317 ) ;
  assign n31319 = ( x198 & n31316 ) | ( x198 & n31318 ) | ( n31316 & n31318 ) ;
  assign n31320 = x625 & ~n31319 ;
  assign n31321 = x625 | n31060 ;
  assign n31322 = ( x1153 & n31320 ) | ( x1153 & n31321 ) | ( n31320 & n31321 ) ;
  assign n31323 = ~n31320 & n31322 ;
  assign n31324 = x625 & ~n31060 ;
  assign n31325 = x1153 | n31324 ;
  assign n31326 = ( n31319 & n31320 ) | ( n31319 & ~n31325 ) | ( n31320 & ~n31325 ) ;
  assign n31327 = n31323 | n31326 ;
  assign n31328 = n31319 ^ x778 ^ 1'b0 ;
  assign n31329 = ( n31319 & n31327 ) | ( n31319 & n31328 ) | ( n31327 & n31328 ) ;
  assign n31330 = n31060 ^ n16234 ^ 1'b0 ;
  assign n31331 = ( n31060 & n31329 ) | ( n31060 & ~n31330 ) | ( n31329 & ~n31330 ) ;
  assign n31332 = n31060 ^ n16254 ^ 1'b0 ;
  assign n31333 = ( n31060 & n31331 ) | ( n31060 & ~n31332 ) | ( n31331 & ~n31332 ) ;
  assign n31334 = n16279 | n31333 ;
  assign n31335 = n16318 | n31334 ;
  assign n31336 = n17086 & ~n31060 ;
  assign n31337 = n31335 & ~n31336 ;
  assign n31338 = n31060 ^ x628 ^ 1'b0 ;
  assign n31339 = ( n31060 & n31337 ) | ( n31060 & n31338 ) | ( n31337 & n31338 ) ;
  assign n31340 = x1156 & n31339 ;
  assign n31341 = x628 & ~n31060 ;
  assign n31342 = x1156 | n31341 ;
  assign n31343 = ( x628 & n31337 ) | ( x628 & ~n31342 ) | ( n31337 & ~n31342 ) ;
  assign n31344 = ~n31342 & n31343 ;
  assign n31345 = ( x792 & n31340 ) | ( x792 & ~n31344 ) | ( n31340 & ~n31344 ) ;
  assign n31346 = ~n31340 & n31345 ;
  assign n31347 = ( x792 & n31337 ) | ( x792 & ~n31346 ) | ( n31337 & ~n31346 ) ;
  assign n31348 = ~n31346 & n31347 ;
  assign n31349 = ( x647 & ~n31219 ) | ( x647 & n31348 ) | ( ~n31219 & n31348 ) ;
  assign n31350 = ~n31219 & n31349 ;
  assign n31351 = n31060 ^ x647 ^ 1'b0 ;
  assign n31352 = ( n31060 & n31348 ) | ( n31060 & n31351 ) | ( n31348 & n31351 ) ;
  assign n31353 = x1157 & n31352 ;
  assign n31354 = n31350 | n31353 ;
  assign n31355 = ( n16373 & n16374 ) | ( n16373 & n31354 ) | ( n16374 & n31354 ) ;
  assign n31356 = ( x787 & n31217 ) | ( x787 & n31355 ) | ( n31217 & n31355 ) ;
  assign n31357 = n31355 ^ n31217 ^ 1'b0 ;
  assign n31358 = ( x787 & n31356 ) | ( x787 & n31357 ) | ( n31356 & n31357 ) ;
  assign n31359 = ~x626 & n31060 ;
  assign n31360 = x626 & n31212 ;
  assign n31361 = ( n22317 & n31359 ) | ( n22317 & ~n31360 ) | ( n31359 & ~n31360 ) ;
  assign n31362 = ~n31359 & n31361 ;
  assign n31363 = ~x626 & n31212 ;
  assign n31364 = x626 & n31060 ;
  assign n31365 = ( n22322 & n31363 ) | ( n22322 & ~n31364 ) | ( n31363 & ~n31364 ) ;
  assign n31366 = ~n31363 & n31365 ;
  assign n31367 = n16279 & ~n31060 ;
  assign n31368 = n31334 & ~n31367 ;
  assign n31369 = ~n31366 & n31368 ;
  assign n31370 = ( n16459 & n31366 ) | ( n16459 & ~n31369 ) | ( n31366 & ~n31369 ) ;
  assign n31371 = ( x788 & n31362 ) | ( x788 & n31370 ) | ( n31362 & n31370 ) ;
  assign n31372 = n31370 ^ n31362 ^ 1'b0 ;
  assign n31373 = ( x788 & n31371 ) | ( x788 & n31372 ) | ( n31371 & n31372 ) ;
  assign n31374 = x198 | x665 ;
  assign n31375 = n15493 & ~n31374 ;
  assign n31376 = x198 & ~n16033 ;
  assign n31377 = ~n15635 & n31376 ;
  assign n31378 = ( x633 & ~n31375 ) | ( x633 & n31377 ) | ( ~n31375 & n31377 ) ;
  assign n31379 = n31375 | n31378 ;
  assign n31380 = x198 & ~x665 ;
  assign n31381 = x633 & ~n31380 ;
  assign n31382 = ~x198 & n16024 ;
  assign n31383 = ( n31070 & n31381 ) | ( n31070 & ~n31382 ) | ( n31381 & ~n31382 ) ;
  assign n31384 = ~n31070 & n31383 ;
  assign n31385 = x603 & ~n31384 ;
  assign n31386 = n31379 & n31385 ;
  assign n31387 = ( ~x603 & n31293 ) | ( ~x603 & n31386 ) | ( n31293 & n31386 ) ;
  assign n31388 = n31386 ^ x603 ^ 1'b0 ;
  assign n31389 = ( n31386 & n31387 ) | ( n31386 & ~n31388 ) | ( n31387 & ~n31388 ) ;
  assign n31390 = ( ~x634 & x680 ) | ( ~x634 & n31389 ) | ( x680 & n31389 ) ;
  assign n31391 = x634 & n31390 ;
  assign n31392 = n31073 & ~n31294 ;
  assign n31393 = ( x299 & n31391 ) | ( x299 & ~n31392 ) | ( n31391 & ~n31392 ) ;
  assign n31394 = ~n31391 & n31393 ;
  assign n31395 = ~x680 & n31078 ;
  assign n31396 = x603 | n31303 ;
  assign n31397 = x198 & ~x633 ;
  assign n31398 = x634 & ~x665 ;
  assign n31399 = ~n31397 & n31398 ;
  assign n31400 = x603 & ~n31399 ;
  assign n31401 = ( x603 & ~n15504 ) | ( x603 & n31400 ) | ( ~n15504 & n31400 ) ;
  assign n31402 = x634 & n16036 ;
  assign n31403 = ~n15497 & n31402 ;
  assign n31404 = ~x634 & n15318 ;
  assign n31405 = ( ~x633 & n31403 ) | ( ~x633 & n31404 ) | ( n31403 & n31404 ) ;
  assign n31406 = ~x633 & n31405 ;
  assign n31407 = ( n31076 & n31401 ) | ( n31076 & ~n31406 ) | ( n31401 & ~n31406 ) ;
  assign n31408 = ~n31076 & n31407 ;
  assign n31409 = x680 & ~n31408 ;
  assign n31410 = n31396 & n31409 ;
  assign n31411 = ( x299 & ~n31395 ) | ( x299 & n31410 ) | ( ~n31395 & n31410 ) ;
  assign n31412 = n31395 | n31411 ;
  assign n31413 = n31412 ^ n31394 ^ 1'b0 ;
  assign n31414 = ( n31394 & n31412 ) | ( n31394 & n31413 ) | ( n31412 & n31413 ) ;
  assign n31415 = ( x39 & ~n31394 ) | ( x39 & n31414 ) | ( ~n31394 & n31414 ) ;
  assign n31416 = ~x680 & n31090 ;
  assign n31417 = ~x634 & n31086 ;
  assign n31418 = n15557 & ~n31374 ;
  assign n31419 = n15510 & n31380 ;
  assign n31420 = n31086 | n31419 ;
  assign n31421 = ( x634 & n31418 ) | ( x634 & n31420 ) | ( n31418 & n31420 ) ;
  assign n31422 = n31420 ^ n31418 ^ 1'b0 ;
  assign n31423 = ( x634 & n31421 ) | ( x634 & n31422 ) | ( n31421 & n31422 ) ;
  assign n31424 = ( n31085 & ~n31417 ) | ( n31085 & n31423 ) | ( ~n31417 & n31423 ) ;
  assign n31425 = n31417 | n31424 ;
  assign n31426 = n15531 & n31398 ;
  assign n31427 = n31096 | n31426 ;
  assign n31428 = x603 & n31427 ;
  assign n31429 = ( n31122 & n31124 ) | ( n31122 & n31428 ) | ( n31124 & n31428 ) ;
  assign n31430 = n31425 & n31429 ;
  assign n31431 = n5075 & n31429 ;
  assign n31432 = ~x603 & n31256 ;
  assign n31433 = n31431 | n31432 ;
  assign n31434 = x603 & n31425 ;
  assign n31435 = ~n15527 & n31434 ;
  assign n31436 = ( ~n31430 & n31433 ) | ( ~n31430 & n31435 ) | ( n31433 & n31435 ) ;
  assign n31437 = n31430 | n31436 ;
  assign n31438 = ( ~x680 & n15383 ) | ( ~x680 & n31437 ) | ( n15383 & n31437 ) ;
  assign n31439 = x680 & n31438 ;
  assign n31440 = n31254 ^ x603 ^ 1'b0 ;
  assign n31441 = ( n31254 & n31425 ) | ( n31254 & n31440 ) | ( n31425 & n31440 ) ;
  assign n31442 = ( x681 & n5077 ) | ( x681 & n31441 ) | ( n5077 & n31441 ) ;
  assign n31443 = ~x681 & n31442 ;
  assign n31444 = ( ~n31416 & n31439 ) | ( ~n31416 & n31443 ) | ( n31439 & n31443 ) ;
  assign n31445 = n31416 | n31444 ;
  assign n31446 = n5061 & ~n31445 ;
  assign n31447 = ~x680 & n31108 ;
  assign n31448 = n31221 ^ x603 ^ 1'b0 ;
  assign n31449 = ( n31221 & n31427 ) | ( n31221 & n31448 ) | ( n31427 & n31448 ) ;
  assign n31450 = n15527 & ~n31449 ;
  assign n31451 = n5075 | n31427 ;
  assign n31452 = n5075 & ~n31425 ;
  assign n31453 = n31451 & ~n31452 ;
  assign n31454 = x603 & n31453 ;
  assign n31455 = ~x603 & n31221 ;
  assign n31456 = n15527 | n31455 ;
  assign n31457 = n31454 | n31456 ;
  assign n31458 = ( n15693 & n31450 ) | ( n15693 & n31457 ) | ( n31450 & n31457 ) ;
  assign n31459 = ~n31450 & n31458 ;
  assign n31460 = n31265 ^ x603 ^ 1'b0 ;
  assign n31461 = ( n31265 & n31453 ) | ( n31265 & n31460 ) | ( n31453 & n31460 ) ;
  assign n31462 = ( x681 & n5077 ) | ( x681 & n31461 ) | ( n5077 & n31461 ) ;
  assign n31463 = ~x681 & n31462 ;
  assign n31464 = ( ~n31447 & n31459 ) | ( ~n31447 & n31463 ) | ( n31459 & n31463 ) ;
  assign n31465 = n31447 | n31464 ;
  assign n31466 = n5061 | n31465 ;
  assign n31467 = ( x215 & n31446 ) | ( x215 & n31466 ) | ( n31446 & n31466 ) ;
  assign n31468 = ~n31446 & n31467 ;
  assign n31469 = ~x680 & n31129 ;
  assign n31470 = n5081 | n31429 ;
  assign n31471 = x634 & n15726 ;
  assign n31472 = n31116 | n31471 ;
  assign n31473 = n31431 | n31472 ;
  assign n31474 = n31470 & n31473 ;
  assign n31475 = ( ~x603 & n31239 ) | ( ~x603 & n31474 ) | ( n31239 & n31474 ) ;
  assign n31476 = n31474 ^ x603 ^ 1'b0 ;
  assign n31477 = ( n31474 & n31475 ) | ( n31474 & ~n31476 ) | ( n31475 & ~n31476 ) ;
  assign n31478 = ( ~x680 & n15383 ) | ( ~x680 & n31477 ) | ( n15383 & n31477 ) ;
  assign n31479 = x680 & n31478 ;
  assign n31480 = ~n15524 & n31226 ;
  assign n31481 = n31117 | n31480 ;
  assign n31482 = n5078 & n31481 ;
  assign n31483 = ( ~n31469 & n31479 ) | ( ~n31469 & n31482 ) | ( n31479 & n31482 ) ;
  assign n31484 = n31469 | n31483 ;
  assign n31485 = n5061 & n31484 ;
  assign n31486 = n5075 & ~n31472 ;
  assign n31487 = ( x603 & n31451 ) | ( x603 & n31486 ) | ( n31451 & n31486 ) ;
  assign n31488 = ~n31486 & n31487 ;
  assign n31489 = ~x642 & n31488 ;
  assign n31490 = ( x642 & n31449 ) | ( x642 & n31455 ) | ( n31449 & n31455 ) ;
  assign n31491 = ( ~n5080 & n31489 ) | ( ~n5080 & n31490 ) | ( n31489 & n31490 ) ;
  assign n31492 = ~n5080 & n31491 ;
  assign n31493 = n5080 & n31449 ;
  assign n31494 = ( n15383 & n31492 ) | ( n15383 & ~n31493 ) | ( n31492 & ~n31493 ) ;
  assign n31495 = ~n31492 & n31494 ;
  assign n31496 = ~x603 & n31227 ;
  assign n31497 = n15383 | n31496 ;
  assign n31498 = n31488 | n31497 ;
  assign n31499 = ~n31495 & n31498 ;
  assign n31500 = n31145 ^ x680 ^ 1'b0 ;
  assign n31501 = ( n31145 & n31499 ) | ( n31145 & n31500 ) | ( n31499 & n31500 ) ;
  assign n31502 = ~n5061 & n31501 ;
  assign n31503 = ( n2263 & n31485 ) | ( n2263 & ~n31502 ) | ( n31485 & ~n31502 ) ;
  assign n31504 = ~n31485 & n31503 ;
  assign n31505 = n15691 & n31220 ;
  assign n31506 = n31098 | n31505 ;
  assign n31507 = n2263 | n31506 ;
  assign n31508 = ( x215 & ~n31504 ) | ( x215 & n31507 ) | ( ~n31504 & n31507 ) ;
  assign n31509 = ~x215 & n31508 ;
  assign n31510 = ( x299 & n31468 ) | ( x299 & n31509 ) | ( n31468 & n31509 ) ;
  assign n31511 = n31509 ^ n31468 ^ 1'b0 ;
  assign n31512 = ( x299 & n31510 ) | ( x299 & n31511 ) | ( n31510 & n31511 ) ;
  assign n31513 = n5114 & ~n31445 ;
  assign n31514 = n5114 | n31465 ;
  assign n31515 = ( x223 & n31513 ) | ( x223 & n31514 ) | ( n31513 & n31514 ) ;
  assign n31516 = ~n31513 & n31515 ;
  assign n31517 = n5114 & n31484 ;
  assign n31518 = ~n5114 & n31501 ;
  assign n31519 = ( n1359 & n31517 ) | ( n1359 & ~n31518 ) | ( n31517 & ~n31518 ) ;
  assign n31520 = ~n31517 & n31519 ;
  assign n31521 = n1359 | n31506 ;
  assign n31522 = ( x223 & ~n31520 ) | ( x223 & n31521 ) | ( ~n31520 & n31521 ) ;
  assign n31523 = ~x223 & n31522 ;
  assign n31524 = ( ~x299 & n31516 ) | ( ~x299 & n31523 ) | ( n31516 & n31523 ) ;
  assign n31525 = ~x299 & n31524 ;
  assign n31526 = ( x39 & n31512 ) | ( x39 & ~n31525 ) | ( n31512 & ~n31525 ) ;
  assign n31527 = ~n31512 & n31526 ;
  assign n31528 = ( x38 & n31415 ) | ( x38 & ~n31527 ) | ( n31415 & ~n31527 ) ;
  assign n31529 = n31528 ^ n31415 ^ 1'b0 ;
  assign n31530 = ( x38 & n31528 ) | ( x38 & ~n31529 ) | ( n31528 & ~n31529 ) ;
  assign n31531 = x634 & n16068 ;
  assign n31532 = n31065 | n31531 ;
  assign n31533 = ( x39 & n31062 ) | ( x39 & ~n31532 ) | ( n31062 & ~n31532 ) ;
  assign n31534 = ( n31062 & ~n31310 ) | ( n31062 & n31533 ) | ( ~n31310 & n31533 ) ;
  assign n31535 = ( n2069 & n31530 ) | ( n2069 & ~n31534 ) | ( n31530 & ~n31534 ) ;
  assign n31536 = ~n2069 & n31535 ;
  assign n31537 = n31536 ^ x198 ^ 1'b0 ;
  assign n31538 = ( ~x198 & n2069 ) | ( ~x198 & n31537 ) | ( n2069 & n31537 ) ;
  assign n31539 = ( x198 & n31536 ) | ( x198 & n31538 ) | ( n31536 & n31538 ) ;
  assign n31540 = x625 & ~n31539 ;
  assign n31541 = x625 | n31179 ;
  assign n31542 = ( x1153 & n31540 ) | ( x1153 & n31541 ) | ( n31540 & n31541 ) ;
  assign n31543 = ~n31540 & n31542 ;
  assign n31544 = ( x608 & n31326 ) | ( x608 & ~n31543 ) | ( n31326 & ~n31543 ) ;
  assign n31545 = ~n31326 & n31544 ;
  assign n31546 = x625 & ~n31179 ;
  assign n31547 = x1153 | n31546 ;
  assign n31548 = ( x625 & n31539 ) | ( x625 & ~n31547 ) | ( n31539 & ~n31547 ) ;
  assign n31549 = ~n31547 & n31548 ;
  assign n31550 = x608 | n31323 ;
  assign n31551 = ( ~n31545 & n31549 ) | ( ~n31545 & n31550 ) | ( n31549 & n31550 ) ;
  assign n31552 = ~n31545 & n31551 ;
  assign n31553 = n31539 ^ x778 ^ 1'b0 ;
  assign n31554 = ( n31539 & n31552 ) | ( n31539 & n31553 ) | ( n31552 & n31553 ) ;
  assign n31555 = x609 & ~n31554 ;
  assign n31556 = x609 | n31329 ;
  assign n31557 = ( x1155 & n31555 ) | ( x1155 & n31556 ) | ( n31555 & n31556 ) ;
  assign n31558 = ~n31555 & n31557 ;
  assign n31559 = ~x1155 & n31188 ;
  assign n31560 = ( x660 & n31558 ) | ( x660 & ~n31559 ) | ( n31558 & ~n31559 ) ;
  assign n31561 = ~n31558 & n31560 ;
  assign n31562 = x1155 & n31185 ;
  assign n31563 = x660 | n31562 ;
  assign n31564 = x609 & ~n31329 ;
  assign n31565 = x1155 | n31564 ;
  assign n31566 = ( n31554 & n31555 ) | ( n31554 & ~n31565 ) | ( n31555 & ~n31565 ) ;
  assign n31567 = ( ~n31561 & n31563 ) | ( ~n31561 & n31566 ) | ( n31563 & n31566 ) ;
  assign n31568 = ~n31561 & n31567 ;
  assign n31569 = n31554 ^ x785 ^ 1'b0 ;
  assign n31570 = ( n31554 & n31568 ) | ( n31554 & n31569 ) | ( n31568 & n31569 ) ;
  assign n31571 = x618 & ~n31570 ;
  assign n31572 = x618 | n31331 ;
  assign n31573 = ( x1154 & n31571 ) | ( x1154 & n31572 ) | ( n31571 & n31572 ) ;
  assign n31574 = ~n31571 & n31573 ;
  assign n31575 = ( x627 & n31199 ) | ( x627 & ~n31574 ) | ( n31199 & ~n31574 ) ;
  assign n31576 = ~n31199 & n31575 ;
  assign n31577 = x627 | n31196 ;
  assign n31578 = x618 & ~n31331 ;
  assign n31579 = x1154 | n31578 ;
  assign n31580 = ( n31570 & n31571 ) | ( n31570 & ~n31579 ) | ( n31571 & ~n31579 ) ;
  assign n31581 = ( ~n31576 & n31577 ) | ( ~n31576 & n31580 ) | ( n31577 & n31580 ) ;
  assign n31582 = ~n31576 & n31581 ;
  assign n31583 = n31570 ^ x781 ^ 1'b0 ;
  assign n31584 = ( n31570 & n31582 ) | ( n31570 & n31583 ) | ( n31582 & n31583 ) ;
  assign n31585 = ~x789 & n31584 ;
  assign n31586 = n16519 | n31585 ;
  assign n31587 = x619 & ~n31333 ;
  assign n31588 = x1159 | n31587 ;
  assign n31589 = x619 & ~n31584 ;
  assign n31590 = ( n31584 & ~n31588 ) | ( n31584 & n31589 ) | ( ~n31588 & n31589 ) ;
  assign n31591 = ( x648 & n31206 ) | ( x648 & ~n31590 ) | ( n31206 & ~n31590 ) ;
  assign n31592 = n31590 | n31591 ;
  assign n31593 = x619 | n31333 ;
  assign n31594 = ( x1159 & n31589 ) | ( x1159 & n31593 ) | ( n31589 & n31593 ) ;
  assign n31595 = ~n31589 & n31594 ;
  assign n31596 = ( x648 & n31209 ) | ( x648 & ~n31595 ) | ( n31209 & ~n31595 ) ;
  assign n31597 = ~n31209 & n31596 ;
  assign n31598 = x789 & ~n31597 ;
  assign n31599 = n31592 & n31598 ;
  assign n31600 = ( ~n31373 & n31586 ) | ( ~n31373 & n31599 ) | ( n31586 & n31599 ) ;
  assign n31601 = ~n31373 & n31600 ;
  assign n31602 = n19046 & n31214 ;
  assign n31603 = x629 & n31344 ;
  assign n31604 = n16337 & n31339 ;
  assign n31605 = ( ~n31602 & n31603 ) | ( ~n31602 & n31604 ) | ( n31603 & n31604 ) ;
  assign n31606 = n31602 | n31605 ;
  assign n31607 = n31601 ^ x792 ^ 1'b0 ;
  assign n31608 = ( ~x792 & n31606 ) | ( ~x792 & n31607 ) | ( n31606 & n31607 ) ;
  assign n31609 = ( x792 & n31601 ) | ( x792 & n31608 ) | ( n31601 & n31608 ) ;
  assign n31610 = n18482 & ~n31606 ;
  assign n31611 = n18484 | n31610 ;
  assign n31612 = ( n31358 & n31609 ) | ( n31358 & ~n31611 ) | ( n31609 & ~n31611 ) ;
  assign n31613 = n31612 ^ n31609 ^ 1'b0 ;
  assign n31614 = ( n31358 & n31612 ) | ( n31358 & ~n31613 ) | ( n31612 & ~n31613 ) ;
  assign n31615 = x644 & ~n31614 ;
  assign n31616 = n31348 ^ x787 ^ 1'b0 ;
  assign n31617 = ( n31348 & n31354 ) | ( n31348 & n31616 ) | ( n31354 & n31616 ) ;
  assign n31618 = x644 | n31617 ;
  assign n31619 = ( x715 & n31615 ) | ( x715 & n31618 ) | ( n31615 & n31618 ) ;
  assign n31620 = ~n31615 & n31619 ;
  assign n31621 = x644 | n31060 ;
  assign n31622 = n31060 ^ n16376 ^ 1'b0 ;
  assign n31623 = ( n31060 & n31216 ) | ( n31060 & ~n31622 ) | ( n31216 & ~n31622 ) ;
  assign n31624 = x644 & ~n31623 ;
  assign n31625 = ( x715 & n31621 ) | ( x715 & ~n31624 ) | ( n31621 & ~n31624 ) ;
  assign n31626 = ~x715 & n31625 ;
  assign n31627 = ( x1160 & n31620 ) | ( x1160 & ~n31626 ) | ( n31620 & ~n31626 ) ;
  assign n31628 = ~n31620 & n31627 ;
  assign n31629 = x644 | n31614 ;
  assign n31630 = x644 & ~n31060 ;
  assign n31631 = x715 & ~n31630 ;
  assign n31632 = n31631 ^ x1160 ^ 1'b0 ;
  assign n31633 = x644 | n31623 ;
  assign n31634 = ( n31631 & ~n31632 ) | ( n31631 & n31633 ) | ( ~n31632 & n31633 ) ;
  assign n31635 = ( x1160 & n31632 ) | ( x1160 & n31634 ) | ( n31632 & n31634 ) ;
  assign n31636 = x644 & ~n31617 ;
  assign n31637 = x715 | n31636 ;
  assign n31638 = ~n31635 & n31637 ;
  assign n31639 = ( n31629 & n31635 ) | ( n31629 & ~n31638 ) | ( n31635 & ~n31638 ) ;
  assign n31640 = ( x790 & n31628 ) | ( x790 & n31639 ) | ( n31628 & n31639 ) ;
  assign n31641 = ~n31628 & n31640 ;
  assign n31642 = ( ~x790 & n31614 ) | ( ~x790 & n31641 ) | ( n31614 & n31641 ) ;
  assign n31643 = n31641 ^ x790 ^ 1'b0 ;
  assign n31644 = ( n31641 & n31642 ) | ( n31641 & ~n31643 ) | ( n31642 & ~n31643 ) ;
  assign n31645 = n31644 ^ n7318 ^ 1'b0 ;
  assign n31646 = ( x198 & n31644 ) | ( x198 & n31645 ) | ( n31644 & n31645 ) ;
  assign n31700 = x199 | n17838 ;
  assign n31701 = n17841 & n31700 ;
  assign n31702 = x199 | n15640 ;
  assign n31703 = x199 & n15587 ;
  assign n31704 = ( x38 & n31702 ) | ( x38 & ~n31703 ) | ( n31702 & ~n31703 ) ;
  assign n31705 = ~x38 & n31704 ;
  assign n31706 = ( ~n2069 & n31701 ) | ( ~n2069 & n31705 ) | ( n31701 & n31705 ) ;
  assign n31707 = ~n2069 & n31706 ;
  assign n31648 = x199 & n2069 ;
  assign n31708 = ( x617 & ~n31648 ) | ( x617 & n31707 ) | ( ~n31648 & n31707 ) ;
  assign n31709 = ~n31707 & n31708 ;
  assign n31647 = x199 & ~n15656 ;
  assign n31710 = ( x617 & n31647 ) | ( x617 & ~n31709 ) | ( n31647 & ~n31709 ) ;
  assign n31711 = ~n31709 & n31710 ;
  assign n31739 = x199 & n17902 ;
  assign n31740 = ~n2069 & n17910 ;
  assign n31741 = x199 | n31740 ;
  assign n31742 = ( x617 & n31739 ) | ( x617 & n31741 ) | ( n31739 & n31741 ) ;
  assign n31743 = ~n31739 & n31742 ;
  assign n31744 = x38 & n17889 ;
  assign n31745 = x617 | n31744 ;
  assign n31746 = ~n2069 & n22651 ;
  assign n31747 = ( x199 & ~n31745 ) | ( x199 & n31746 ) | ( ~n31745 & n31746 ) ;
  assign n31748 = ~n31745 & n31747 ;
  assign n31749 = ~x38 & n17891 ;
  assign n31750 = ( x199 & ~n31748 ) | ( x199 & n31749 ) | ( ~n31748 & n31749 ) ;
  assign n31751 = n31750 ^ n31748 ^ 1'b0 ;
  assign n31752 = ( n31748 & ~n31750 ) | ( n31748 & n31751 ) | ( ~n31750 & n31751 ) ;
  assign n31753 = ( n31648 & ~n31743 ) | ( n31648 & n31752 ) | ( ~n31743 & n31752 ) ;
  assign n31754 = n31743 | n31753 ;
  assign n31755 = n31711 ^ x637 ^ 1'b0 ;
  assign n31756 = ( n31711 & n31754 ) | ( n31711 & n31755 ) | ( n31754 & n31755 ) ;
  assign n31757 = x625 & ~n31756 ;
  assign n31758 = x625 | n31711 ;
  assign n31759 = ( x1153 & n31757 ) | ( x1153 & n31758 ) | ( n31757 & n31758 ) ;
  assign n31760 = ~n31757 & n31759 ;
  assign n31667 = x625 & ~n31647 ;
  assign n31668 = x1153 | n31667 ;
  assign n31649 = x199 | n15644 ;
  assign n31650 = n18524 & n31649 ;
  assign n31651 = x199 & ~n16141 ;
  assign n31652 = ~x199 & n16178 ;
  assign n31653 = ( x39 & n31651 ) | ( x39 & ~n31652 ) | ( n31651 & ~n31652 ) ;
  assign n31654 = ~n31651 & n31653 ;
  assign n31655 = x199 & ~n16041 ;
  assign n31656 = ~x199 & n16053 ;
  assign n31657 = ( x39 & ~n31655 ) | ( x39 & n31656 ) | ( ~n31655 & n31656 ) ;
  assign n31658 = n31655 | n31657 ;
  assign n31659 = ( x38 & ~n31654 ) | ( x38 & n31658 ) | ( ~n31654 & n31658 ) ;
  assign n31660 = ~x38 & n31659 ;
  assign n31661 = ( ~n2069 & n31650 ) | ( ~n2069 & n31660 ) | ( n31650 & n31660 ) ;
  assign n31662 = ~n2069 & n31661 ;
  assign n31663 = ( x637 & n31648 ) | ( x637 & ~n31662 ) | ( n31648 & ~n31662 ) ;
  assign n31664 = ~n31648 & n31663 ;
  assign n31665 = ( x637 & n31647 ) | ( x637 & ~n31664 ) | ( n31647 & ~n31664 ) ;
  assign n31666 = ~n31664 & n31665 ;
  assign n31669 = ( x625 & n31666 ) | ( x625 & ~n31668 ) | ( n31666 & ~n31668 ) ;
  assign n31670 = ~n31668 & n31669 ;
  assign n31761 = ( x608 & ~n31670 ) | ( x608 & n31760 ) | ( ~n31670 & n31760 ) ;
  assign n31762 = ~n31760 & n31761 ;
  assign n31671 = x625 & ~n31666 ;
  assign n31672 = x625 | n31647 ;
  assign n31673 = ( x1153 & n31671 ) | ( x1153 & n31672 ) | ( n31671 & n31672 ) ;
  assign n31674 = ~n31671 & n31673 ;
  assign n31763 = x608 | n31674 ;
  assign n31764 = x625 & ~n31711 ;
  assign n31765 = x1153 | n31764 ;
  assign n31766 = ( n31756 & n31757 ) | ( n31756 & ~n31765 ) | ( n31757 & ~n31765 ) ;
  assign n31767 = ( ~n31762 & n31763 ) | ( ~n31762 & n31766 ) | ( n31763 & n31766 ) ;
  assign n31768 = ~n31762 & n31767 ;
  assign n31769 = n31756 ^ x778 ^ 1'b0 ;
  assign n31770 = ( n31756 & n31768 ) | ( n31756 & n31769 ) | ( n31768 & n31769 ) ;
  assign n31771 = x609 & ~n31770 ;
  assign n31675 = n31670 | n31674 ;
  assign n31676 = n31666 ^ x778 ^ 1'b0 ;
  assign n31677 = ( n31666 & n31675 ) | ( n31666 & n31676 ) | ( n31675 & n31676 ) ;
  assign n31772 = x609 | n31677 ;
  assign n31773 = ( x1155 & n31771 ) | ( x1155 & n31772 ) | ( n31771 & n31772 ) ;
  assign n31774 = ~n31771 & n31773 ;
  assign n31714 = x609 & ~n31647 ;
  assign n31715 = x1155 | n31714 ;
  assign n31712 = n31647 ^ n15659 ^ 1'b0 ;
  assign n31713 = ( n31647 & n31711 ) | ( n31647 & ~n31712 ) | ( n31711 & ~n31712 ) ;
  assign n31716 = ( x609 & n31713 ) | ( x609 & ~n31715 ) | ( n31713 & ~n31715 ) ;
  assign n31717 = ~n31715 & n31716 ;
  assign n31775 = ( x660 & ~n31717 ) | ( x660 & n31774 ) | ( ~n31717 & n31774 ) ;
  assign n31776 = ~n31774 & n31775 ;
  assign n31718 = x609 & ~n31713 ;
  assign n31719 = x609 | n31647 ;
  assign n31720 = ( x1155 & n31718 ) | ( x1155 & n31719 ) | ( n31718 & n31719 ) ;
  assign n31721 = ~n31718 & n31720 ;
  assign n31777 = x660 | n31721 ;
  assign n31778 = x609 & ~n31677 ;
  assign n31779 = x1155 | n31778 ;
  assign n31780 = ( n31770 & n31771 ) | ( n31770 & ~n31779 ) | ( n31771 & ~n31779 ) ;
  assign n31781 = ( ~n31776 & n31777 ) | ( ~n31776 & n31780 ) | ( n31777 & n31780 ) ;
  assign n31782 = ~n31776 & n31781 ;
  assign n31783 = n31770 ^ x785 ^ 1'b0 ;
  assign n31784 = ( n31770 & n31782 ) | ( n31770 & n31783 ) | ( n31782 & n31783 ) ;
  assign n31785 = x618 & ~n31784 ;
  assign n31678 = n31647 ^ n16234 ^ 1'b0 ;
  assign n31679 = ( n31647 & n31677 ) | ( n31647 & ~n31678 ) | ( n31677 & ~n31678 ) ;
  assign n31786 = x618 | n31679 ;
  assign n31787 = ( x1154 & n31785 ) | ( x1154 & n31786 ) | ( n31785 & n31786 ) ;
  assign n31788 = ~n31785 & n31787 ;
  assign n31722 = n31717 | n31721 ;
  assign n31723 = n31713 ^ x785 ^ 1'b0 ;
  assign n31724 = ( n31713 & n31722 ) | ( n31713 & n31723 ) | ( n31722 & n31723 ) ;
  assign n31725 = x618 & ~n31724 ;
  assign n31729 = x618 & ~n31647 ;
  assign n31730 = x1154 | n31729 ;
  assign n31731 = ( n31724 & n31725 ) | ( n31724 & ~n31730 ) | ( n31725 & ~n31730 ) ;
  assign n31789 = ( x627 & ~n31731 ) | ( x627 & n31788 ) | ( ~n31731 & n31788 ) ;
  assign n31790 = ~n31788 & n31789 ;
  assign n31726 = x618 | n31647 ;
  assign n31727 = ( x1154 & n31725 ) | ( x1154 & n31726 ) | ( n31725 & n31726 ) ;
  assign n31728 = ~n31725 & n31727 ;
  assign n31791 = x627 | n31728 ;
  assign n31792 = x618 & ~n31679 ;
  assign n31793 = x1154 | n31792 ;
  assign n31794 = ( n31784 & n31785 ) | ( n31784 & ~n31793 ) | ( n31785 & ~n31793 ) ;
  assign n31795 = ( ~n31790 & n31791 ) | ( ~n31790 & n31794 ) | ( n31791 & n31794 ) ;
  assign n31796 = ~n31790 & n31795 ;
  assign n31797 = n31784 ^ x781 ^ 1'b0 ;
  assign n31798 = ( n31784 & n31796 ) | ( n31784 & n31797 ) | ( n31796 & n31797 ) ;
  assign n31799 = x619 & ~n31798 ;
  assign n31680 = n31647 ^ n16254 ^ 1'b0 ;
  assign n31681 = ( n31647 & n31679 ) | ( n31647 & ~n31680 ) | ( n31679 & ~n31680 ) ;
  assign n31805 = x619 | n31681 ;
  assign n31806 = ( x1159 & n31799 ) | ( x1159 & n31805 ) | ( n31799 & n31805 ) ;
  assign n31807 = ~n31799 & n31806 ;
  assign n31732 = n31728 | n31731 ;
  assign n31733 = n31724 ^ x781 ^ 1'b0 ;
  assign n31734 = ( n31724 & n31732 ) | ( n31724 & n31733 ) | ( n31732 & n31733 ) ;
  assign n31735 = x619 & ~n31734 ;
  assign n31808 = x619 & ~n31647 ;
  assign n31809 = x1159 | n31808 ;
  assign n31810 = ( n31734 & n31735 ) | ( n31734 & ~n31809 ) | ( n31735 & ~n31809 ) ;
  assign n31811 = ( x648 & n31807 ) | ( x648 & ~n31810 ) | ( n31807 & ~n31810 ) ;
  assign n31812 = ~n31807 & n31811 ;
  assign n31736 = x619 | n31647 ;
  assign n31737 = ( x1159 & n31735 ) | ( x1159 & n31736 ) | ( n31735 & n31736 ) ;
  assign n31738 = ~n31735 & n31737 ;
  assign n31800 = x619 & ~n31681 ;
  assign n31801 = x1159 | n31800 ;
  assign n31802 = ( n31798 & n31799 ) | ( n31798 & ~n31801 ) | ( n31799 & ~n31801 ) ;
  assign n31803 = ( x648 & ~n31738 ) | ( x648 & n31802 ) | ( ~n31738 & n31802 ) ;
  assign n31804 = n31738 | n31803 ;
  assign n31813 = n31812 ^ n31804 ^ 1'b0 ;
  assign n31814 = ( x789 & ~n31804 ) | ( x789 & n31812 ) | ( ~n31804 & n31812 ) ;
  assign n31815 = ( x789 & ~n31813 ) | ( x789 & n31814 ) | ( ~n31813 & n31814 ) ;
  assign n31816 = ( x789 & n31798 ) | ( x789 & ~n31815 ) | ( n31798 & ~n31815 ) ;
  assign n31817 = ~n31815 & n31816 ;
  assign n31818 = ~x626 & n31817 ;
  assign n31682 = n31647 ^ n16279 ^ 1'b0 ;
  assign n31683 = ( n31647 & n31681 ) | ( n31647 & ~n31682 ) | ( n31681 & ~n31682 ) ;
  assign n31819 = x626 & n31683 ;
  assign n31820 = ( x641 & ~n31818 ) | ( x641 & n31819 ) | ( ~n31818 & n31819 ) ;
  assign n31821 = n31818 | n31820 ;
  assign n31822 = ~x626 & n31647 ;
  assign n31823 = n31738 | n31810 ;
  assign n31824 = n31734 ^ x789 ^ 1'b0 ;
  assign n31825 = ( n31734 & n31823 ) | ( n31734 & n31824 ) | ( n31823 & n31824 ) ;
  assign n31826 = x626 & n31825 ;
  assign n31827 = ( x641 & ~n31822 ) | ( x641 & n31826 ) | ( ~n31822 & n31826 ) ;
  assign n31828 = n31822 | n31827 ;
  assign n31829 = ~x626 & n31683 ;
  assign n31830 = x626 & n31817 ;
  assign n31831 = ( x641 & n31829 ) | ( x641 & ~n31830 ) | ( n31829 & ~n31830 ) ;
  assign n31832 = ~n31829 & n31831 ;
  assign n31833 = x1158 & ~n31832 ;
  assign n31834 = n31828 & n31833 ;
  assign n31835 = ~x626 & n31825 ;
  assign n31836 = x626 & n31647 ;
  assign n31837 = x641 & ~n31836 ;
  assign n31838 = n31837 ^ n31835 ^ 1'b0 ;
  assign n31839 = ( n31835 & n31837 ) | ( n31835 & n31838 ) | ( n31837 & n31838 ) ;
  assign n31840 = ( x1158 & ~n31835 ) | ( x1158 & n31839 ) | ( ~n31835 & n31839 ) ;
  assign n31841 = ~n31834 & n31840 ;
  assign n31842 = ( n31821 & n31834 ) | ( n31821 & ~n31841 ) | ( n31834 & ~n31841 ) ;
  assign n31843 = n31817 ^ x788 ^ 1'b0 ;
  assign n31844 = ( n31817 & n31842 ) | ( n31817 & n31843 ) | ( n31842 & n31843 ) ;
  assign n31845 = x628 & ~n31844 ;
  assign n31846 = n31647 ^ n16518 ^ 1'b0 ;
  assign n31847 = ( n31647 & n31825 ) | ( n31647 & ~n31846 ) | ( n31825 & ~n31846 ) ;
  assign n31848 = x628 | n31847 ;
  assign n31849 = ( x1156 & n31845 ) | ( x1156 & n31848 ) | ( n31845 & n31848 ) ;
  assign n31850 = ~n31845 & n31849 ;
  assign n31684 = n31647 ^ n16318 ^ 1'b0 ;
  assign n31685 = ( n31647 & n31683 ) | ( n31647 & ~n31684 ) | ( n31683 & ~n31684 ) ;
  assign n31686 = x628 & ~n31685 ;
  assign n31690 = x628 & ~n31647 ;
  assign n31691 = x1156 | n31690 ;
  assign n31692 = ( n31685 & n31686 ) | ( n31685 & ~n31691 ) | ( n31686 & ~n31691 ) ;
  assign n31851 = ( x629 & ~n31692 ) | ( x629 & n31850 ) | ( ~n31692 & n31850 ) ;
  assign n31852 = ~n31850 & n31851 ;
  assign n31687 = x628 | n31647 ;
  assign n31688 = ( x1156 & n31686 ) | ( x1156 & n31687 ) | ( n31686 & n31687 ) ;
  assign n31689 = ~n31686 & n31688 ;
  assign n31853 = x629 | n31689 ;
  assign n31854 = x628 & ~n31847 ;
  assign n31855 = x1156 | n31854 ;
  assign n31856 = ( n31844 & n31845 ) | ( n31844 & ~n31855 ) | ( n31845 & ~n31855 ) ;
  assign n31857 = ( ~n31852 & n31853 ) | ( ~n31852 & n31856 ) | ( n31853 & n31856 ) ;
  assign n31858 = ~n31852 & n31857 ;
  assign n31859 = n31844 ^ x792 ^ 1'b0 ;
  assign n31860 = ( n31844 & n31858 ) | ( n31844 & n31859 ) | ( n31858 & n31859 ) ;
  assign n31861 = x647 & ~n31860 ;
  assign n31862 = n31647 ^ n16339 ^ 1'b0 ;
  assign n31863 = ( n31647 & n31847 ) | ( n31647 & ~n31862 ) | ( n31847 & ~n31862 ) ;
  assign n31869 = x647 | n31863 ;
  assign n31870 = ( x1157 & n31861 ) | ( x1157 & n31869 ) | ( n31861 & n31869 ) ;
  assign n31871 = ~n31861 & n31870 ;
  assign n31693 = n31689 | n31692 ;
  assign n31694 = n31685 ^ x792 ^ 1'b0 ;
  assign n31695 = ( n31685 & n31693 ) | ( n31685 & n31694 ) | ( n31693 & n31694 ) ;
  assign n31696 = x647 & ~n31695 ;
  assign n31872 = x647 & ~n31647 ;
  assign n31873 = x1157 | n31872 ;
  assign n31874 = ( n31695 & n31696 ) | ( n31695 & ~n31873 ) | ( n31696 & ~n31873 ) ;
  assign n31875 = ( x630 & n31871 ) | ( x630 & ~n31874 ) | ( n31871 & ~n31874 ) ;
  assign n31876 = ~n31871 & n31875 ;
  assign n31697 = x647 | n31647 ;
  assign n31698 = ( x1157 & n31696 ) | ( x1157 & n31697 ) | ( n31696 & n31697 ) ;
  assign n31699 = ~n31696 & n31698 ;
  assign n31864 = x647 & ~n31863 ;
  assign n31865 = x1157 | n31864 ;
  assign n31866 = ( n31860 & n31861 ) | ( n31860 & ~n31865 ) | ( n31861 & ~n31865 ) ;
  assign n31867 = ( x630 & ~n31699 ) | ( x630 & n31866 ) | ( ~n31699 & n31866 ) ;
  assign n31868 = n31699 | n31867 ;
  assign n31877 = n31876 ^ n31868 ^ 1'b0 ;
  assign n31878 = ( x787 & ~n31868 ) | ( x787 & n31876 ) | ( ~n31868 & n31876 ) ;
  assign n31879 = ( x787 & ~n31877 ) | ( x787 & n31878 ) | ( ~n31877 & n31878 ) ;
  assign n31880 = ( x787 & n31860 ) | ( x787 & ~n31879 ) | ( n31860 & ~n31879 ) ;
  assign n31881 = ~n31879 & n31880 ;
  assign n31882 = x644 & ~n31881 ;
  assign n31883 = n31699 | n31874 ;
  assign n31884 = n31695 ^ x787 ^ 1'b0 ;
  assign n31885 = ( n31695 & n31883 ) | ( n31695 & n31884 ) | ( n31883 & n31884 ) ;
  assign n31886 = x644 | n31885 ;
  assign n31887 = ( x715 & n31882 ) | ( x715 & n31886 ) | ( n31882 & n31886 ) ;
  assign n31888 = ~n31882 & n31887 ;
  assign n31889 = x644 | n31647 ;
  assign n31890 = n31647 ^ n16376 ^ 1'b0 ;
  assign n31891 = ( n31647 & n31863 ) | ( n31647 & ~n31890 ) | ( n31863 & ~n31890 ) ;
  assign n31892 = x644 & ~n31891 ;
  assign n31893 = ( x715 & n31889 ) | ( x715 & ~n31892 ) | ( n31889 & ~n31892 ) ;
  assign n31894 = ~x715 & n31893 ;
  assign n31895 = ( x1160 & n31888 ) | ( x1160 & ~n31894 ) | ( n31888 & ~n31894 ) ;
  assign n31896 = ~n31888 & n31895 ;
  assign n31897 = x644 | n31881 ;
  assign n31898 = x644 & ~n31647 ;
  assign n31899 = x715 & ~n31898 ;
  assign n31900 = n31899 ^ x1160 ^ 1'b0 ;
  assign n31901 = x644 | n31891 ;
  assign n31902 = ( n31899 & ~n31900 ) | ( n31899 & n31901 ) | ( ~n31900 & n31901 ) ;
  assign n31903 = ( x1160 & n31900 ) | ( x1160 & n31902 ) | ( n31900 & n31902 ) ;
  assign n31904 = x644 & ~n31885 ;
  assign n31905 = x715 | n31904 ;
  assign n31906 = ~n31903 & n31905 ;
  assign n31907 = ( n31897 & n31903 ) | ( n31897 & ~n31906 ) | ( n31903 & ~n31906 ) ;
  assign n31908 = ( x790 & n31896 ) | ( x790 & n31907 ) | ( n31896 & n31907 ) ;
  assign n31909 = ~n31896 & n31908 ;
  assign n31910 = ( ~x790 & n31881 ) | ( ~x790 & n31909 ) | ( n31881 & n31909 ) ;
  assign n31911 = n31909 ^ x790 ^ 1'b0 ;
  assign n31912 = ( n31909 & n31910 ) | ( n31909 & ~n31911 ) | ( n31910 & ~n31911 ) ;
  assign n31913 = n31912 ^ n7318 ^ 1'b0 ;
  assign n31914 = ( x199 & n31912 ) | ( x199 & n31913 ) | ( n31912 & n31913 ) ;
  assign n31915 = x200 & ~n15656 ;
  assign n31916 = x647 & ~n31915 ;
  assign n31917 = x1157 | n31916 ;
  assign n31918 = x200 & n2069 ;
  assign n31919 = x200 | n15644 ;
  assign n31920 = n18524 & n31919 ;
  assign n31921 = x200 | n16163 ;
  assign n31922 = x200 & n16127 ;
  assign n31923 = ( x299 & n31921 ) | ( x299 & ~n31922 ) | ( n31921 & ~n31922 ) ;
  assign n31924 = ~x299 & n31923 ;
  assign n31925 = x200 & n16139 ;
  assign n31926 = x200 | n16176 ;
  assign n31927 = ( x299 & n31925 ) | ( x299 & n31926 ) | ( n31925 & n31926 ) ;
  assign n31928 = ~n31925 & n31927 ;
  assign n31929 = ( x39 & n31924 ) | ( x39 & n31928 ) | ( n31924 & n31928 ) ;
  assign n31930 = n31928 ^ n31924 ^ 1'b0 ;
  assign n31931 = ( x39 & n31929 ) | ( x39 & n31930 ) | ( n31929 & n31930 ) ;
  assign n31932 = x200 | n16053 ;
  assign n31933 = x200 & n16041 ;
  assign n31934 = ( x39 & n31932 ) | ( x39 & ~n31933 ) | ( n31932 & ~n31933 ) ;
  assign n31935 = ~x39 & n31934 ;
  assign n31936 = ( ~x38 & n31931 ) | ( ~x38 & n31935 ) | ( n31931 & n31935 ) ;
  assign n31937 = ~x38 & n31936 ;
  assign n31938 = ( ~n2069 & n31920 ) | ( ~n2069 & n31937 ) | ( n31920 & n31937 ) ;
  assign n31939 = ~n2069 & n31938 ;
  assign n31940 = ( x643 & n31918 ) | ( x643 & ~n31939 ) | ( n31918 & ~n31939 ) ;
  assign n31941 = ~n31918 & n31940 ;
  assign n31942 = ( x643 & n31915 ) | ( x643 & ~n31941 ) | ( n31915 & ~n31941 ) ;
  assign n31943 = ~n31941 & n31942 ;
  assign n31944 = x625 & ~n31943 ;
  assign n31945 = x625 | n31915 ;
  assign n31946 = ( x1153 & n31944 ) | ( x1153 & n31945 ) | ( n31944 & n31945 ) ;
  assign n31947 = ~n31944 & n31946 ;
  assign n31948 = x625 & ~n31915 ;
  assign n31949 = x1153 | n31948 ;
  assign n31950 = ( x625 & n31943 ) | ( x625 & ~n31949 ) | ( n31943 & ~n31949 ) ;
  assign n31951 = ~n31949 & n31950 ;
  assign n31952 = n31947 | n31951 ;
  assign n31953 = n31943 ^ x778 ^ 1'b0 ;
  assign n31954 = ( n31943 & n31952 ) | ( n31943 & n31953 ) | ( n31952 & n31953 ) ;
  assign n31955 = n31915 ^ n16234 ^ 1'b0 ;
  assign n31956 = ( n31915 & n31954 ) | ( n31915 & ~n31955 ) | ( n31954 & ~n31955 ) ;
  assign n31957 = n31915 ^ n16254 ^ 1'b0 ;
  assign n31958 = ( n31915 & n31956 ) | ( n31915 & ~n31957 ) | ( n31956 & ~n31957 ) ;
  assign n31959 = n31915 ^ n16279 ^ 1'b0 ;
  assign n31960 = ( n31915 & n31958 ) | ( n31915 & ~n31959 ) | ( n31958 & ~n31959 ) ;
  assign n31961 = n31915 ^ n16318 ^ 1'b0 ;
  assign n31962 = ( n31915 & n31960 ) | ( n31915 & ~n31961 ) | ( n31960 & ~n31961 ) ;
  assign n31963 = x628 & ~n31962 ;
  assign n31964 = x628 | n31915 ;
  assign n31965 = ( x1156 & n31963 ) | ( x1156 & n31964 ) | ( n31963 & n31964 ) ;
  assign n31966 = ~n31963 & n31965 ;
  assign n31967 = x628 & ~n31915 ;
  assign n31968 = x1156 | n31967 ;
  assign n31969 = ( n31962 & n31963 ) | ( n31962 & ~n31968 ) | ( n31963 & ~n31968 ) ;
  assign n31970 = n31966 | n31969 ;
  assign n31971 = n31962 ^ x792 ^ 1'b0 ;
  assign n31972 = ( n31962 & n31970 ) | ( n31962 & n31971 ) | ( n31970 & n31971 ) ;
  assign n31973 = ( x647 & ~n31917 ) | ( x647 & n31972 ) | ( ~n31917 & n31972 ) ;
  assign n31974 = ~n31917 & n31973 ;
  assign n31975 = x630 & n31974 ;
  assign n31976 = x200 | n17838 ;
  assign n31977 = n17841 & n31976 ;
  assign n31978 = x200 | n15640 ;
  assign n31979 = x200 & n15587 ;
  assign n31980 = ( x38 & n31978 ) | ( x38 & ~n31979 ) | ( n31978 & ~n31979 ) ;
  assign n31981 = ~x38 & n31980 ;
  assign n31982 = ( ~n2069 & n31977 ) | ( ~n2069 & n31981 ) | ( n31977 & n31981 ) ;
  assign n31983 = ~n2069 & n31982 ;
  assign n31984 = ( x606 & ~n31918 ) | ( x606 & n31983 ) | ( ~n31918 & n31983 ) ;
  assign n31985 = ~n31983 & n31984 ;
  assign n31986 = ( x606 & n31915 ) | ( x606 & ~n31985 ) | ( n31915 & ~n31985 ) ;
  assign n31987 = ~n31985 & n31986 ;
  assign n31988 = n31915 ^ n15659 ^ 1'b0 ;
  assign n31989 = ( n31915 & n31987 ) | ( n31915 & ~n31988 ) | ( n31987 & ~n31988 ) ;
  assign n31990 = x609 & ~n31989 ;
  assign n31991 = x609 | n31915 ;
  assign n31992 = ( x1155 & n31990 ) | ( x1155 & n31991 ) | ( n31990 & n31991 ) ;
  assign n31993 = ~n31990 & n31992 ;
  assign n31994 = x609 & ~n31915 ;
  assign n31995 = x1155 | n31994 ;
  assign n31996 = ( x609 & n31989 ) | ( x609 & ~n31995 ) | ( n31989 & ~n31995 ) ;
  assign n31997 = ~n31995 & n31996 ;
  assign n31998 = n31993 | n31997 ;
  assign n31999 = n31989 ^ x785 ^ 1'b0 ;
  assign n32000 = ( n31989 & n31998 ) | ( n31989 & n31999 ) | ( n31998 & n31999 ) ;
  assign n32001 = x618 & ~n32000 ;
  assign n32002 = x618 | n31915 ;
  assign n32003 = ( x1154 & n32001 ) | ( x1154 & n32002 ) | ( n32001 & n32002 ) ;
  assign n32004 = ~n32001 & n32003 ;
  assign n32005 = x618 & ~n31915 ;
  assign n32006 = x1154 | n32005 ;
  assign n32007 = ( n32000 & n32001 ) | ( n32000 & ~n32006 ) | ( n32001 & ~n32006 ) ;
  assign n32008 = n32004 | n32007 ;
  assign n32009 = n32000 ^ x781 ^ 1'b0 ;
  assign n32010 = ( n32000 & n32008 ) | ( n32000 & n32009 ) | ( n32008 & n32009 ) ;
  assign n32011 = x619 | n31915 ;
  assign n32012 = x619 & ~n32010 ;
  assign n32013 = x1159 & ~n32012 ;
  assign n32014 = n32011 & n32013 ;
  assign n32015 = x619 & ~n31915 ;
  assign n32016 = x1159 | n32015 ;
  assign n32017 = ( n32010 & n32012 ) | ( n32010 & ~n32016 ) | ( n32012 & ~n32016 ) ;
  assign n32018 = n32014 | n32017 ;
  assign n32019 = n32010 ^ x789 ^ 1'b0 ;
  assign n32020 = ( n32010 & n32018 ) | ( n32010 & n32019 ) | ( n32018 & n32019 ) ;
  assign n32021 = n31915 ^ n16518 ^ 1'b0 ;
  assign n32022 = ( n31915 & n32020 ) | ( n31915 & ~n32021 ) | ( n32020 & ~n32021 ) ;
  assign n32023 = n31915 ^ n16339 ^ 1'b0 ;
  assign n32024 = ( n31915 & n32022 ) | ( n31915 & ~n32023 ) | ( n32022 & ~n32023 ) ;
  assign n32025 = n19055 & n32024 ;
  assign n32026 = n31975 | n32025 ;
  assign n32027 = n31915 ^ x647 ^ 1'b0 ;
  assign n32028 = ( n31915 & n31972 ) | ( n31915 & n32027 ) | ( n31972 & n32027 ) ;
  assign n32029 = n16373 & n32028 ;
  assign n32030 = ( x787 & n32026 ) | ( x787 & n32029 ) | ( n32026 & n32029 ) ;
  assign n32031 = n32029 ^ n32026 ^ 1'b0 ;
  assign n32032 = ( x787 & n32030 ) | ( x787 & n32031 ) | ( n32030 & n32031 ) ;
  assign n32033 = x200 & n17891 ;
  assign n32034 = x200 | n17885 ;
  assign n32035 = ( x38 & ~n32033 ) | ( x38 & n32034 ) | ( ~n32033 & n32034 ) ;
  assign n32036 = ~x38 & n32035 ;
  assign n32037 = n15691 | n16185 ;
  assign n32038 = n32036 ^ n31920 ^ 1'b0 ;
  assign n32039 = ( ~n31920 & n32037 ) | ( ~n31920 & n32038 ) | ( n32037 & n32038 ) ;
  assign n32040 = ( n31920 & n32036 ) | ( n31920 & n32039 ) | ( n32036 & n32039 ) ;
  assign n32041 = ( x606 & ~n2069 ) | ( x606 & n32040 ) | ( ~n2069 & n32040 ) ;
  assign n32042 = ~x606 & n32041 ;
  assign n32043 = ~x200 & n17907 ;
  assign n32044 = x38 | n32043 ;
  assign n32045 = n22969 & ~n32044 ;
  assign n32046 = ( x200 & n32044 ) | ( x200 & ~n32045 ) | ( n32044 & ~n32045 ) ;
  assign n32047 = n32046 ^ n31918 ^ 1'b0 ;
  assign n32048 = x38 & x200 ;
  assign n32049 = n17897 & n32048 ;
  assign n32050 = ( x606 & n2069 ) | ( x606 & ~n32049 ) | ( n2069 & ~n32049 ) ;
  assign n32051 = ~n2069 & n32050 ;
  assign n32052 = n32051 ^ x200 ^ 1'b0 ;
  assign n32053 = n17905 | n17906 ;
  assign n32054 = ( x200 & n32052 ) | ( x200 & ~n32053 ) | ( n32052 & ~n32053 ) ;
  assign n32055 = ( n32051 & ~n32052 ) | ( n32051 & n32054 ) | ( ~n32052 & n32054 ) ;
  assign n32056 = ( n32046 & ~n32047 ) | ( n32046 & n32055 ) | ( ~n32047 & n32055 ) ;
  assign n32057 = ( n31918 & n32047 ) | ( n31918 & n32056 ) | ( n32047 & n32056 ) ;
  assign n32058 = ( x643 & n32042 ) | ( x643 & ~n32057 ) | ( n32042 & ~n32057 ) ;
  assign n32059 = ~n32042 & n32058 ;
  assign n32060 = ( x643 & n31987 ) | ( x643 & ~n32059 ) | ( n31987 & ~n32059 ) ;
  assign n32061 = ~n32059 & n32060 ;
  assign n32062 = x625 & ~n32061 ;
  assign n32063 = x625 | n31987 ;
  assign n32064 = ( x1153 & n32062 ) | ( x1153 & n32063 ) | ( n32062 & n32063 ) ;
  assign n32065 = ~n32062 & n32064 ;
  assign n32066 = ( x608 & n31951 ) | ( x608 & ~n32065 ) | ( n31951 & ~n32065 ) ;
  assign n32067 = ~n31951 & n32066 ;
  assign n32068 = x608 | n31947 ;
  assign n32069 = x625 & ~n31987 ;
  assign n32070 = x1153 | n32069 ;
  assign n32071 = ( n32061 & n32062 ) | ( n32061 & ~n32070 ) | ( n32062 & ~n32070 ) ;
  assign n32072 = ( ~n32067 & n32068 ) | ( ~n32067 & n32071 ) | ( n32068 & n32071 ) ;
  assign n32073 = ~n32067 & n32072 ;
  assign n32074 = n32061 ^ x778 ^ 1'b0 ;
  assign n32075 = ( n32061 & n32073 ) | ( n32061 & n32074 ) | ( n32073 & n32074 ) ;
  assign n32076 = x609 | n32075 ;
  assign n32077 = x609 & ~n31954 ;
  assign n32078 = ( x1155 & n32076 ) | ( x1155 & ~n32077 ) | ( n32076 & ~n32077 ) ;
  assign n32079 = ~x1155 & n32078 ;
  assign n32080 = ( x660 & n31993 ) | ( x660 & ~n32079 ) | ( n31993 & ~n32079 ) ;
  assign n32081 = n32079 | n32080 ;
  assign n32082 = x609 | n31954 ;
  assign n32083 = x609 & ~n32075 ;
  assign n32084 = x1155 & ~n32083 ;
  assign n32085 = n32082 & n32084 ;
  assign n32086 = x660 & ~n31997 ;
  assign n32087 = n32081 & ~n32086 ;
  assign n32088 = ( n32081 & n32085 ) | ( n32081 & n32087 ) | ( n32085 & n32087 ) ;
  assign n32089 = n32075 ^ x785 ^ 1'b0 ;
  assign n32090 = ( n32075 & n32088 ) | ( n32075 & n32089 ) | ( n32088 & n32089 ) ;
  assign n32091 = x618 & ~n32090 ;
  assign n32092 = x618 | n31956 ;
  assign n32093 = ( x1154 & n32091 ) | ( x1154 & n32092 ) | ( n32091 & n32092 ) ;
  assign n32094 = ~n32091 & n32093 ;
  assign n32095 = ( x627 & n32007 ) | ( x627 & ~n32094 ) | ( n32007 & ~n32094 ) ;
  assign n32096 = ~n32007 & n32095 ;
  assign n32097 = x627 | n32004 ;
  assign n32098 = x618 & ~n31956 ;
  assign n32099 = x1154 | n32098 ;
  assign n32100 = ( n32090 & n32091 ) | ( n32090 & ~n32099 ) | ( n32091 & ~n32099 ) ;
  assign n32101 = ( ~n32096 & n32097 ) | ( ~n32096 & n32100 ) | ( n32097 & n32100 ) ;
  assign n32102 = ~n32096 & n32101 ;
  assign n32103 = n32090 ^ x781 ^ 1'b0 ;
  assign n32104 = ( n32090 & n32102 ) | ( n32090 & n32103 ) | ( n32102 & n32103 ) ;
  assign n32105 = x619 | n32104 ;
  assign n32106 = x619 & ~n31958 ;
  assign n32107 = ( x1159 & n32105 ) | ( x1159 & ~n32106 ) | ( n32105 & ~n32106 ) ;
  assign n32108 = ~x1159 & n32107 ;
  assign n32109 = ( x648 & n32014 ) | ( x648 & ~n32108 ) | ( n32014 & ~n32108 ) ;
  assign n32110 = n32108 | n32109 ;
  assign n32111 = x619 & ~n32104 ;
  assign n32112 = x619 | n31958 ;
  assign n32113 = ( x1159 & n32111 ) | ( x1159 & n32112 ) | ( n32111 & n32112 ) ;
  assign n32114 = ~n32111 & n32113 ;
  assign n32115 = ( x648 & n32017 ) | ( x648 & ~n32114 ) | ( n32017 & ~n32114 ) ;
  assign n32116 = ~n32017 & n32115 ;
  assign n32117 = x789 & ~n32116 ;
  assign n32118 = n32110 & n32117 ;
  assign n32119 = ~x789 & n32104 ;
  assign n32120 = ( n16519 & ~n32118 ) | ( n16519 & n32119 ) | ( ~n32118 & n32119 ) ;
  assign n32121 = n32118 | n32120 ;
  assign n32122 = n31966 ^ x629 ^ 1'b0 ;
  assign n32123 = ( n31966 & n31969 ) | ( n31966 & n32122 ) | ( n31969 & n32122 ) ;
  assign n32124 = n19046 & n32022 ;
  assign n32125 = ( x792 & n32123 ) | ( x792 & n32124 ) | ( n32123 & n32124 ) ;
  assign n32126 = n32124 ^ n32123 ^ 1'b0 ;
  assign n32127 = ( x792 & n32125 ) | ( x792 & n32126 ) | ( n32125 & n32126 ) ;
  assign n32128 = ~x626 & n32020 ;
  assign n32129 = x626 & n31915 ;
  assign n32130 = ( n22322 & n32128 ) | ( n22322 & ~n32129 ) | ( n32128 & ~n32129 ) ;
  assign n32131 = ~n32128 & n32130 ;
  assign n32132 = ~x626 & n31915 ;
  assign n32133 = x626 & n32020 ;
  assign n32134 = ( n22317 & n32132 ) | ( n22317 & ~n32133 ) | ( n32132 & ~n32133 ) ;
  assign n32135 = ~n32132 & n32134 ;
  assign n32136 = n16459 & ~n31960 ;
  assign n32137 = ( ~n32131 & n32135 ) | ( ~n32131 & n32136 ) | ( n32135 & n32136 ) ;
  assign n32138 = n32131 | n32137 ;
  assign n32139 = ( x788 & ~n22314 ) | ( x788 & n32138 ) | ( ~n22314 & n32138 ) ;
  assign n32140 = ( n18482 & n22314 ) | ( n18482 & n32139 ) | ( n22314 & n32139 ) ;
  assign n32141 = ~n32127 & n32140 ;
  assign n32142 = ( n32121 & n32127 ) | ( n32121 & ~n32141 ) | ( n32127 & ~n32141 ) ;
  assign n32143 = ( ~n18484 & n32032 ) | ( ~n18484 & n32142 ) | ( n32032 & n32142 ) ;
  assign n32144 = n32032 ^ n18484 ^ 1'b0 ;
  assign n32145 = ( n32032 & n32143 ) | ( n32032 & ~n32144 ) | ( n32143 & ~n32144 ) ;
  assign n32146 = x644 & ~n32145 ;
  assign n32147 = x1157 & n32028 ;
  assign n32148 = ( x787 & n31974 ) | ( x787 & ~n32147 ) | ( n31974 & ~n32147 ) ;
  assign n32149 = ~n31974 & n32148 ;
  assign n32150 = ( x787 & n31972 ) | ( x787 & ~n32149 ) | ( n31972 & ~n32149 ) ;
  assign n32151 = ~n32149 & n32150 ;
  assign n32152 = x644 | n32151 ;
  assign n32153 = ( x715 & n32146 ) | ( x715 & n32152 ) | ( n32146 & n32152 ) ;
  assign n32154 = ~n32146 & n32153 ;
  assign n32155 = x644 | n31915 ;
  assign n32156 = n31915 ^ n16376 ^ 1'b0 ;
  assign n32157 = ( n31915 & n32024 ) | ( n31915 & ~n32156 ) | ( n32024 & ~n32156 ) ;
  assign n32158 = x644 & ~n32157 ;
  assign n32159 = ( x715 & n32155 ) | ( x715 & ~n32158 ) | ( n32155 & ~n32158 ) ;
  assign n32160 = ~x715 & n32159 ;
  assign n32161 = ( x1160 & n32154 ) | ( x1160 & ~n32160 ) | ( n32154 & ~n32160 ) ;
  assign n32162 = ~n32154 & n32161 ;
  assign n32163 = x644 & ~n31915 ;
  assign n32164 = x715 & ~n32163 ;
  assign n32165 = n32164 ^ x1160 ^ 1'b0 ;
  assign n32166 = x644 | n32157 ;
  assign n32167 = ( n32164 & ~n32165 ) | ( n32164 & n32166 ) | ( ~n32165 & n32166 ) ;
  assign n32168 = ( x1160 & n32165 ) | ( x1160 & n32167 ) | ( n32165 & n32167 ) ;
  assign n32169 = x644 & ~n32151 ;
  assign n32170 = x715 | n32169 ;
  assign n32171 = ( n32145 & n32146 ) | ( n32145 & ~n32170 ) | ( n32146 & ~n32170 ) ;
  assign n32172 = ( ~n32162 & n32168 ) | ( ~n32162 & n32171 ) | ( n32168 & n32171 ) ;
  assign n32173 = ~n32162 & n32172 ;
  assign n32174 = n32145 ^ x790 ^ 1'b0 ;
  assign n32175 = ( n32145 & n32173 ) | ( n32145 & n32174 ) | ( n32173 & n32174 ) ;
  assign n32176 = n32175 ^ n7318 ^ 1'b0 ;
  assign n32177 = ( x200 & n32175 ) | ( x200 & n32176 ) | ( n32175 & n32176 ) ;
  assign n32178 = ~n1292 & n5539 ;
  assign n32179 = ( x332 & n14201 ) | ( x332 & n32178 ) | ( n14201 & n32178 ) ;
  assign n32180 = n14201 & n32179 ;
  assign n32181 = x332 & n2056 ;
  assign n32182 = n32180 | n32181 ;
  assign n32183 = n1397 & ~n9713 ;
  assign n32184 = n5538 & n32183 ;
  assign n32185 = x332 | n32184 ;
  assign n32186 = ~n6336 & n32185 ;
  assign n32187 = ( ~x74 & n32182 ) | ( ~x74 & n32186 ) | ( n32182 & n32186 ) ;
  assign n32188 = ~x74 & n32187 ;
  assign n32189 = x74 & x332 ;
  assign n32190 = ( x55 & ~n32188 ) | ( x55 & n32189 ) | ( ~n32188 & n32189 ) ;
  assign n32191 = n32188 | n32190 ;
  assign n32192 = ~n2070 & n5497 ;
  assign n32193 = ~n1292 & n32192 ;
  assign n32194 = x332 | n32193 ;
  assign n32195 = x55 & ~n32194 ;
  assign n32196 = ( n2109 & n32191 ) | ( n2109 & ~n32195 ) | ( n32191 & ~n32195 ) ;
  assign n32197 = ~n2109 & n32196 ;
  assign n32198 = x332 & n2109 ;
  assign n32199 = ( x59 & ~n32197 ) | ( x59 & n32198 ) | ( ~n32197 & n32198 ) ;
  assign n32200 = n32197 | n32199 ;
  assign n32201 = x332 & n5192 ;
  assign n32202 = x59 & ~n32201 ;
  assign n32203 = ~n5192 & n32194 ;
  assign n32204 = n32202 & ~n32203 ;
  assign n32205 = ( x57 & n32200 ) | ( x57 & ~n32204 ) | ( n32200 & ~n32204 ) ;
  assign n32206 = ~x57 & n32205 ;
  assign n32207 = n32206 ^ x57 ^ 1'b0 ;
  assign n32208 = ( ~x57 & x332 ) | ( ~x57 & n32207 ) | ( x332 & n32207 ) ;
  assign n32209 = ( x57 & n32206 ) | ( x57 & n32208 ) | ( n32206 & n32208 ) ;
  assign n32210 = x332 | n5081 ;
  assign n32211 = ~x947 & n32210 ;
  assign n32212 = x96 & x210 ;
  assign n32213 = x332 & n32212 ;
  assign n32214 = x32 | x96 ;
  assign n32215 = x70 & ~n32214 ;
  assign n32216 = x332 | n32215 ;
  assign n32217 = x70 | x841 ;
  assign n32218 = x32 & n32217 ;
  assign n32219 = x32 | x70 ;
  assign n32220 = ~n32218 & n32219 ;
  assign n32221 = ~x210 & n32220 ;
  assign n32222 = n32216 | n32221 ;
  assign n32223 = ~n32213 & n32222 ;
  assign n32224 = n5081 & ~n32223 ;
  assign n32225 = x947 & ~n32224 ;
  assign n32226 = n5075 & n32223 ;
  assign n32227 = n32226 ^ n32223 ^ x332 ;
  assign n32228 = n5081 | n32227 ;
  assign n32229 = n32225 & n32228 ;
  assign n32230 = n5081 & ~n32226 ;
  assign n32231 = ~n32229 & n32230 ;
  assign n32232 = ( n32211 & n32229 ) | ( n32211 & ~n32231 ) | ( n32229 & ~n32231 ) ;
  assign n32233 = n5192 & ~n32232 ;
  assign n32234 = x59 & ~n32233 ;
  assign n32235 = n2109 & ~n32232 ;
  assign n32236 = x95 | n1652 ;
  assign n32237 = n32218 | n32236 ;
  assign n32238 = n1376 | n32237 ;
  assign n32239 = n1399 | n32238 ;
  assign n32240 = ~n32220 & n32239 ;
  assign n32241 = x210 | n32240 ;
  assign n32242 = x95 | n1430 ;
  assign n32243 = x70 | n32242 ;
  assign n32244 = ( ~x70 & n32214 ) | ( ~x70 & n32243 ) | ( n32214 & n32243 ) ;
  assign n32245 = x210 & ~n32244 ;
  assign n32246 = ( x332 & n32241 ) | ( x332 & ~n32245 ) | ( n32241 & ~n32245 ) ;
  assign n32247 = ~x332 & n32246 ;
  assign n32248 = ( ~x332 & x468 ) | ( ~x332 & n32247 ) | ( x468 & n32247 ) ;
  assign n32249 = ~n5081 & n32248 ;
  assign n32250 = n32213 | n32247 ;
  assign n32251 = n5081 & n32250 ;
  assign n32252 = ( x947 & n32249 ) | ( x947 & ~n32251 ) | ( n32249 & ~n32251 ) ;
  assign n32253 = ~n32249 & n32252 ;
  assign n32254 = n5075 & ~n32250 ;
  assign n32255 = n5081 & ~n32254 ;
  assign n32256 = ~n32253 & n32255 ;
  assign n32257 = ( n32211 & n32253 ) | ( n32211 & ~n32256 ) | ( n32253 & ~n32256 ) ;
  assign n32258 = n32232 ^ n2070 ^ 1'b0 ;
  assign n32259 = ( n32232 & n32257 ) | ( n32232 & ~n32258 ) | ( n32257 & ~n32258 ) ;
  assign n32260 = x55 & n32259 ;
  assign n32261 = x96 & x198 ;
  assign n32262 = x332 & n32261 ;
  assign n32263 = ~x198 & n32220 ;
  assign n32264 = n32216 | n32263 ;
  assign n32265 = ~n32262 & n32264 ;
  assign n32266 = n5081 & ~n32265 ;
  assign n32267 = n5493 & n32264 ;
  assign n32268 = n32210 | n32267 ;
  assign n32269 = ~x299 & n5569 ;
  assign n32270 = ( n32266 & n32268 ) | ( n32266 & n32269 ) | ( n32268 & n32269 ) ;
  assign n32271 = ~n32266 & n32270 ;
  assign n32272 = ( x74 & n2056 ) | ( x74 & ~n32271 ) | ( n2056 & ~n32271 ) ;
  assign n32273 = ~n32271 & n32272 ;
  assign n32274 = x299 & n32232 ;
  assign n32275 = ( x55 & n32273 ) | ( x55 & ~n32274 ) | ( n32273 & ~n32274 ) ;
  assign n32276 = n32275 ^ n32273 ^ 1'b0 ;
  assign n32277 = ( x55 & n32275 ) | ( x55 & ~n32276 ) | ( n32275 & ~n32276 ) ;
  assign n32278 = x198 | n32240 ;
  assign n32279 = x198 & ~n32244 ;
  assign n32280 = ( x332 & n32278 ) | ( x332 & ~n32279 ) | ( n32278 & ~n32279 ) ;
  assign n32281 = ~x332 & n32280 ;
  assign n32282 = x468 | n32281 ;
  assign n32283 = ( n5081 & n5537 ) | ( n5081 & n32210 ) | ( n5537 & n32210 ) ;
  assign n32284 = n32282 & ~n32283 ;
  assign n32285 = n32262 | n32281 ;
  assign n32286 = n5081 & n32285 ;
  assign n32287 = ( x587 & n32284 ) | ( x587 & ~n32286 ) | ( n32284 & ~n32286 ) ;
  assign n32288 = ~n32284 & n32287 ;
  assign n32289 = ~x587 & n32210 ;
  assign n32290 = n5075 & ~n32285 ;
  assign n32291 = n5081 & ~n32290 ;
  assign n32292 = n32289 & ~n32291 ;
  assign n32293 = ( ~x299 & n32288 ) | ( ~x299 & n32292 ) | ( n32288 & n32292 ) ;
  assign n32294 = ~x299 & n32293 ;
  assign n32295 = x299 & n32257 ;
  assign n32296 = ( n14201 & n32294 ) | ( n14201 & ~n32295 ) | ( n32294 & ~n32295 ) ;
  assign n32297 = ~n32294 & n32296 ;
  assign n32298 = n1397 & ~n1411 ;
  assign n32299 = x95 | n1288 ;
  assign n32300 = n32298 & ~n32299 ;
  assign n32301 = x70 | n32300 ;
  assign n32302 = ~n32214 & n32301 ;
  assign n32303 = x210 & n32302 ;
  assign n32304 = ~n32237 & n32298 ;
  assign n32305 = n32220 | n32304 ;
  assign n32306 = ~x210 & n32305 ;
  assign n32307 = ( x332 & ~n32303 ) | ( x332 & n32306 ) | ( ~n32303 & n32306 ) ;
  assign n32308 = n32303 | n32307 ;
  assign n32309 = ~n32213 & n32308 ;
  assign n32310 = n5081 & ~n32309 ;
  assign n32311 = x947 & ~n32310 ;
  assign n32312 = n32308 ^ x468 ^ 1'b0 ;
  assign n32313 = ( x332 & n32308 ) | ( x332 & n32312 ) | ( n32308 & n32312 ) ;
  assign n32314 = n5081 | n32313 ;
  assign n32315 = n32311 & n32314 ;
  assign n32316 = n5075 & n32309 ;
  assign n32317 = n5081 & ~n32316 ;
  assign n32318 = n32211 & ~n32317 ;
  assign n32319 = ( x299 & n32315 ) | ( x299 & ~n32318 ) | ( n32315 & ~n32318 ) ;
  assign n32320 = ~n32315 & n32319 ;
  assign n32321 = x198 & n32302 ;
  assign n32322 = ~x198 & n32305 ;
  assign n32323 = ( x332 & ~n32321 ) | ( x332 & n32322 ) | ( ~n32321 & n32322 ) ;
  assign n32324 = n32321 | n32323 ;
  assign n32325 = ~n32262 & n32324 ;
  assign n32326 = n5081 & ~n32325 ;
  assign n32327 = ~x468 & n32324 ;
  assign n32328 = n32283 | n32327 ;
  assign n32329 = ( x587 & n32326 ) | ( x587 & n32328 ) | ( n32326 & n32328 ) ;
  assign n32330 = ~n32326 & n32329 ;
  assign n32331 = ( ~n5075 & n5081 ) | ( ~n5075 & n32326 ) | ( n5081 & n32326 ) ;
  assign n32332 = ( x299 & n32289 ) | ( x299 & ~n32331 ) | ( n32289 & ~n32331 ) ;
  assign n32333 = n32332 ^ n32289 ^ 1'b0 ;
  assign n32334 = ( x299 & n32332 ) | ( x299 & ~n32333 ) | ( n32332 & ~n32333 ) ;
  assign n32335 = ( ~n32320 & n32330 ) | ( ~n32320 & n32334 ) | ( n32330 & n32334 ) ;
  assign n32336 = ~n32320 & n32335 ;
  assign n32337 = ( n6336 & ~n32297 ) | ( n6336 & n32336 ) | ( ~n32297 & n32336 ) ;
  assign n32338 = ~n32297 & n32337 ;
  assign n32339 = ( x74 & ~n32277 ) | ( x74 & n32338 ) | ( ~n32277 & n32338 ) ;
  assign n32340 = ~n32277 & n32339 ;
  assign n32341 = ( n2109 & ~n32260 ) | ( n2109 & n32340 ) | ( ~n32260 & n32340 ) ;
  assign n32342 = n32260 | n32341 ;
  assign n32343 = ( x59 & ~n32235 ) | ( x59 & n32342 ) | ( ~n32235 & n32342 ) ;
  assign n32344 = ~x59 & n32343 ;
  assign n32345 = n5192 | n32259 ;
  assign n32346 = n32344 ^ n32234 ^ 1'b0 ;
  assign n32347 = ( ~n32234 & n32345 ) | ( ~n32234 & n32346 ) | ( n32345 & n32346 ) ;
  assign n32348 = ( n32234 & n32344 ) | ( n32234 & n32347 ) | ( n32344 & n32347 ) ;
  assign n32349 = n32232 ^ x57 ^ 1'b0 ;
  assign n32350 = ( n32232 & n32348 ) | ( n32232 & ~n32349 ) | ( n32348 & ~n32349 ) ;
  assign n32351 = x233 & x237 ;
  assign n32352 = n32351 ^ n32209 ^ 1'b0 ;
  assign n32353 = ( n32209 & n32350 ) | ( n32209 & n32352 ) | ( n32350 & n32352 ) ;
  assign n32354 = n5493 & n32261 ;
  assign n32355 = n32354 ^ n15098 ^ 1'b0 ;
  assign n32356 = ( n5497 & n32354 ) | ( n5497 & n32355 ) | ( n32354 & n32355 ) ;
  assign n32357 = n32356 ^ n32212 ^ 1'b0 ;
  assign n32358 = ( ~n15098 & n32212 ) | ( ~n15098 & n32357 ) | ( n32212 & n32357 ) ;
  assign n32359 = ( n32356 & ~n32357 ) | ( n32356 & n32358 ) | ( ~n32357 & n32358 ) ;
  assign n32360 = n32351 & n32359 ;
  assign n32361 = n32353 ^ x201 ^ 1'b0 ;
  assign n32362 = ( n32353 & ~n32360 ) | ( n32353 & n32361 ) | ( ~n32360 & n32361 ) ;
  assign n32363 = ~x233 & x237 ;
  assign n32364 = n32363 ^ n32350 ^ 1'b0 ;
  assign n32365 = ( n32209 & n32350 ) | ( n32209 & ~n32364 ) | ( n32350 & ~n32364 ) ;
  assign n32366 = n32359 & n32363 ;
  assign n32367 = n32365 ^ x202 ^ 1'b0 ;
  assign n32368 = ( n32365 & ~n32366 ) | ( n32365 & n32367 ) | ( ~n32366 & n32367 ) ;
  assign n32369 = x233 | x237 ;
  assign n32370 = n32369 ^ n32209 ^ 1'b0 ;
  assign n32371 = ( n32209 & n32350 ) | ( n32209 & ~n32370 ) | ( n32350 & ~n32370 ) ;
  assign n32372 = n32359 & ~n32369 ;
  assign n32373 = n32371 ^ x203 ^ 1'b0 ;
  assign n32374 = ( n32371 & ~n32372 ) | ( n32371 & n32373 ) | ( ~n32372 & n32373 ) ;
  assign n32375 = x299 & ~x907 ;
  assign n32376 = ( x299 & ~x468 ) | ( x299 & n5199 ) | ( ~x468 & n5199 ) ;
  assign n32377 = ( n5198 & ~n32375 ) | ( n5198 & n32376 ) | ( ~n32375 & n32376 ) ;
  assign n32378 = n32377 ^ n32376 ^ 1'b0 ;
  assign n32379 = ( n5198 & n32377 ) | ( n5198 & ~n32378 ) | ( n32377 & ~n32378 ) ;
  assign n32380 = n32183 & n32379 ;
  assign n32381 = x332 | n32380 ;
  assign n32382 = ~n6336 & n32381 ;
  assign n32383 = ( n5200 & n5292 ) | ( n5200 & ~n5400 ) | ( n5292 & ~n5400 ) ;
  assign n32384 = n32383 ^ n1292 ^ 1'b0 ;
  assign n32385 = ( n1292 & n32383 ) | ( n1292 & n32384 ) | ( n32383 & n32384 ) ;
  assign n32386 = ( x332 & ~n1292 ) | ( x332 & n32385 ) | ( ~n1292 & n32385 ) ;
  assign n32387 = n14201 & n32386 ;
  assign n32388 = ( ~x74 & n32382 ) | ( ~x74 & n32387 ) | ( n32382 & n32387 ) ;
  assign n32389 = ~x74 & n32388 ;
  assign n32390 = x55 | n32189 ;
  assign n32391 = ( n32181 & ~n32389 ) | ( n32181 & n32390 ) | ( ~n32389 & n32390 ) ;
  assign n32392 = n32389 | n32391 ;
  assign n32393 = ~n2070 & n5292 ;
  assign n32394 = ~n1292 & n32393 ;
  assign n32395 = x332 | n32394 ;
  assign n32396 = x55 & ~n32395 ;
  assign n32397 = ( n2109 & n32392 ) | ( n2109 & ~n32396 ) | ( n32392 & ~n32396 ) ;
  assign n32398 = ~n2109 & n32397 ;
  assign n32399 = ( x59 & n32198 ) | ( x59 & ~n32398 ) | ( n32198 & ~n32398 ) ;
  assign n32400 = n32398 | n32399 ;
  assign n32401 = ~n5192 & n32395 ;
  assign n32402 = n32202 & ~n32401 ;
  assign n32403 = ( x57 & n32400 ) | ( x57 & ~n32402 ) | ( n32400 & ~n32402 ) ;
  assign n32404 = ~x57 & n32403 ;
  assign n32405 = n32404 ^ x57 ^ 1'b0 ;
  assign n32406 = ( ~x57 & x332 ) | ( ~x57 & n32405 ) | ( x332 & n32405 ) ;
  assign n32407 = ( x57 & n32404 ) | ( x57 & n32406 ) | ( n32404 & n32406 ) ;
  assign n32408 = x332 | n5078 ;
  assign n32409 = ~x907 & n32408 ;
  assign n32410 = n5078 & ~n32223 ;
  assign n32411 = x907 & ~n32410 ;
  assign n32412 = n5078 | n32227 ;
  assign n32413 = n32411 & n32412 ;
  assign n32414 = n5078 & ~n32226 ;
  assign n32415 = ~n32413 & n32414 ;
  assign n32416 = ( n32409 & n32413 ) | ( n32409 & ~n32415 ) | ( n32413 & ~n32415 ) ;
  assign n32417 = n5192 & ~n32416 ;
  assign n32418 = x59 & ~n32417 ;
  assign n32419 = n2109 & ~n32416 ;
  assign n32420 = ~n5078 & n32248 ;
  assign n32421 = n5078 & n32250 ;
  assign n32422 = ( x907 & n32420 ) | ( x907 & ~n32421 ) | ( n32420 & ~n32421 ) ;
  assign n32423 = ~n32420 & n32422 ;
  assign n32424 = x332 & n15383 ;
  assign n32425 = ( x680 & n32254 ) | ( x680 & ~n32424 ) | ( n32254 & ~n32424 ) ;
  assign n32426 = ~n32254 & n32425 ;
  assign n32427 = ~n32423 & n32426 ;
  assign n32428 = ( n32409 & n32423 ) | ( n32409 & ~n32427 ) | ( n32423 & ~n32427 ) ;
  assign n32429 = n32416 ^ n2070 ^ 1'b0 ;
  assign n32430 = ( n32416 & n32428 ) | ( n32416 & ~n32429 ) | ( n32428 & ~n32429 ) ;
  assign n32431 = x55 & n32430 ;
  assign n32432 = n5078 & n32261 ;
  assign n32433 = x332 & ~n32432 ;
  assign n32434 = n5200 & n32265 ;
  assign n32435 = ( ~x299 & n32433 ) | ( ~x299 & n32434 ) | ( n32433 & n32434 ) ;
  assign n32436 = ~x299 & n32435 ;
  assign n32437 = ( x74 & n2056 ) | ( x74 & ~n32436 ) | ( n2056 & ~n32436 ) ;
  assign n32438 = ~n32436 & n32437 ;
  assign n32439 = x299 & n32416 ;
  assign n32440 = ( x55 & n32438 ) | ( x55 & ~n32439 ) | ( n32438 & ~n32439 ) ;
  assign n32441 = n32440 ^ n32438 ^ 1'b0 ;
  assign n32442 = ( x55 & n32440 ) | ( x55 & ~n32441 ) | ( n32440 & ~n32441 ) ;
  assign n32443 = x299 & ~n32428 ;
  assign n32444 = x299 | n32433 ;
  assign n32445 = n5201 & ~n32285 ;
  assign n32446 = n32444 | n32445 ;
  assign n32447 = n14201 & ~n32446 ;
  assign n32448 = ( n14201 & n32443 ) | ( n14201 & n32447 ) | ( n32443 & n32447 ) ;
  assign n32449 = n5078 & ~n32309 ;
  assign n32450 = x907 & ~n32449 ;
  assign n32451 = n5078 | n32313 ;
  assign n32452 = n32450 & n32451 ;
  assign n32453 = n5078 & ~n32316 ;
  assign n32454 = n32409 & ~n32453 ;
  assign n32455 = ( x299 & n32452 ) | ( x299 & ~n32454 ) | ( n32452 & ~n32454 ) ;
  assign n32456 = ~n32452 & n32455 ;
  assign n32457 = n5201 & n32325 ;
  assign n32458 = ( n32444 & ~n32456 ) | ( n32444 & n32457 ) | ( ~n32456 & n32457 ) ;
  assign n32459 = ~n32456 & n32458 ;
  assign n32460 = ( n6336 & ~n32448 ) | ( n6336 & n32459 ) | ( ~n32448 & n32459 ) ;
  assign n32461 = ~n32448 & n32460 ;
  assign n32462 = ( x74 & ~n32442 ) | ( x74 & n32461 ) | ( ~n32442 & n32461 ) ;
  assign n32463 = ~n32442 & n32462 ;
  assign n32464 = ( n2109 & ~n32431 ) | ( n2109 & n32463 ) | ( ~n32431 & n32463 ) ;
  assign n32465 = n32431 | n32464 ;
  assign n32466 = ( x59 & ~n32419 ) | ( x59 & n32465 ) | ( ~n32419 & n32465 ) ;
  assign n32467 = ~x59 & n32466 ;
  assign n32468 = n5192 | n32430 ;
  assign n32469 = n32467 ^ n32418 ^ 1'b0 ;
  assign n32470 = ( ~n32418 & n32468 ) | ( ~n32418 & n32469 ) | ( n32468 & n32469 ) ;
  assign n32471 = ( n32418 & n32467 ) | ( n32418 & n32470 ) | ( n32467 & n32470 ) ;
  assign n32472 = n32416 ^ x57 ^ 1'b0 ;
  assign n32473 = ( n32416 & n32471 ) | ( n32416 & ~n32472 ) | ( n32471 & ~n32472 ) ;
  assign n32474 = n32407 ^ n32351 ^ 1'b0 ;
  assign n32475 = ( n32407 & n32473 ) | ( n32407 & n32474 ) | ( n32473 & n32474 ) ;
  assign n32476 = n5201 & n32261 ;
  assign n32477 = n5292 & n32212 ;
  assign n32478 = n32476 ^ n15098 ^ 1'b0 ;
  assign n32479 = ( n32476 & n32477 ) | ( n32476 & n32478 ) | ( n32477 & n32478 ) ;
  assign n32480 = n32351 & n32479 ;
  assign n32481 = n32475 ^ x204 ^ 1'b0 ;
  assign n32482 = ( n32475 & ~n32480 ) | ( n32475 & n32481 ) | ( ~n32480 & n32481 ) ;
  assign n32483 = n32407 ^ n32363 ^ 1'b0 ;
  assign n32484 = ( n32407 & n32473 ) | ( n32407 & n32483 ) | ( n32473 & n32483 ) ;
  assign n32485 = n32363 & n32479 ;
  assign n32486 = n32484 ^ x205 ^ 1'b0 ;
  assign n32487 = ( n32484 & ~n32485 ) | ( n32484 & n32486 ) | ( ~n32485 & n32486 ) ;
  assign n32488 = x233 & ~x237 ;
  assign n32489 = n32488 ^ n32473 ^ 1'b0 ;
  assign n32490 = ( n32407 & n32473 ) | ( n32407 & ~n32489 ) | ( n32473 & ~n32489 ) ;
  assign n32491 = n32479 & n32488 ;
  assign n32492 = n32490 ^ x206 ^ 1'b0 ;
  assign n32493 = ( n32490 & ~n32491 ) | ( n32490 & n32492 ) | ( ~n32491 & n32492 ) ;
  assign n32494 = ~n2069 & n22572 ;
  assign n32495 = ~n15659 & n32494 ;
  assign n32496 = ~n18309 & n32495 ;
  assign n32497 = ~n18315 & n32496 ;
  assign n32500 = x1159 & ~n32497 ;
  assign n32501 = ~n17083 & n22530 ;
  assign n32502 = ~n17087 & n32501 ;
  assign n32503 = x1159 | n32502 ;
  assign n32504 = x619 & ~x648 ;
  assign n32505 = ( n32500 & n32503 ) | ( n32500 & n32504 ) | ( n32503 & n32504 ) ;
  assign n32506 = ~n32500 & n32505 ;
  assign n32507 = x1159 & ~n32502 ;
  assign n32508 = ~x619 & x648 ;
  assign n32509 = x1159 | n32497 ;
  assign n32510 = ( n32507 & n32508 ) | ( n32507 & n32509 ) | ( n32508 & n32509 ) ;
  assign n32511 = ~n32507 & n32510 ;
  assign n32512 = ( x789 & n32506 ) | ( x789 & ~n32511 ) | ( n32506 & ~n32511 ) ;
  assign n32513 = ~n32506 & n32512 ;
  assign n32514 = n21704 & n32513 ;
  assign n32516 = ~x625 & n22530 ;
  assign n32517 = ( x608 & x1153 ) | ( x608 & n32516 ) | ( x1153 & n32516 ) ;
  assign n32518 = ( x608 & ~n15658 ) | ( x608 & n32517 ) | ( ~n15658 & n32517 ) ;
  assign n32519 = x625 & n31740 ;
  assign n32520 = ~x625 & n32494 ;
  assign n32521 = x1153 & ~n32520 ;
  assign n32522 = n32518 & ~n32521 ;
  assign n32523 = ( n32518 & n32519 ) | ( n32518 & n32522 ) | ( n32519 & n32522 ) ;
  assign n32524 = x625 & n22530 ;
  assign n32525 = x1153 & ~n32524 ;
  assign n32526 = x608 | n32525 ;
  assign n32527 = x625 & n32494 ;
  assign n32528 = x1153 | n32527 ;
  assign n32529 = ~x625 & n31740 ;
  assign n32530 = ( ~n32526 & n32528 ) | ( ~n32526 & n32529 ) | ( n32528 & n32529 ) ;
  assign n32531 = ~n32526 & n32530 ;
  assign n32532 = ( x778 & n32523 ) | ( x778 & ~n32531 ) | ( n32523 & ~n32531 ) ;
  assign n32533 = ~n32523 & n32532 ;
  assign n32534 = ( x778 & n31740 ) | ( x778 & ~n32533 ) | ( n31740 & ~n32533 ) ;
  assign n32535 = ~n32533 & n32534 ;
  assign n32536 = x609 & ~n32535 ;
  assign n32542 = x609 | n32501 ;
  assign n32543 = x1155 & n32542 ;
  assign n32544 = ~n32536 & n32543 ;
  assign n32545 = ~n18307 & n32495 ;
  assign n32546 = ( x660 & n32544 ) | ( x660 & ~n32545 ) | ( n32544 & ~n32545 ) ;
  assign n32547 = ~n32544 & n32546 ;
  assign n32515 = n18306 & n32495 ;
  assign n32537 = x609 & ~n32501 ;
  assign n32538 = x1155 | n32537 ;
  assign n32539 = ( n32535 & n32536 ) | ( n32535 & ~n32538 ) | ( n32536 & ~n32538 ) ;
  assign n32540 = ( x660 & ~n32515 ) | ( x660 & n32539 ) | ( ~n32515 & n32539 ) ;
  assign n32541 = n32515 | n32540 ;
  assign n32548 = n32547 ^ n32541 ^ 1'b0 ;
  assign n32549 = ( x785 & ~n32541 ) | ( x785 & n32547 ) | ( ~n32541 & n32547 ) ;
  assign n32550 = ( x785 & ~n32548 ) | ( x785 & n32549 ) | ( ~n32548 & n32549 ) ;
  assign n32551 = ( x785 & n32535 ) | ( x785 & ~n32550 ) | ( n32535 & ~n32550 ) ;
  assign n32552 = ~n32550 & n32551 ;
  assign n32553 = x618 | x627 ;
  assign n32554 = x781 & n32553 ;
  assign n32555 = n32552 | n32554 ;
  assign n32556 = n18312 & n32496 ;
  assign n32557 = x627 | n32556 ;
  assign n32558 = ~n16234 & n32501 ;
  assign n32559 = x618 & ~n32558 ;
  assign n32560 = ( x1154 & ~n32557 ) | ( x1154 & n32559 ) | ( ~n32557 & n32559 ) ;
  assign n32561 = ~n32557 & n32560 ;
  assign n32562 = x618 | n32558 ;
  assign n32563 = x1154 & n32562 ;
  assign n32564 = x618 & ~n32552 ;
  assign n32565 = n32563 & ~n32564 ;
  assign n32566 = ~n18313 & n32496 ;
  assign n32567 = ( x627 & n32565 ) | ( x627 & ~n32566 ) | ( n32565 & ~n32566 ) ;
  assign n32568 = ~n32565 & n32567 ;
  assign n32569 = ( x781 & n32561 ) | ( x781 & n32568 ) | ( n32561 & n32568 ) ;
  assign n32570 = n32568 ^ n32561 ^ 1'b0 ;
  assign n32571 = ( x781 & n32569 ) | ( x781 & n32570 ) | ( n32569 & n32570 ) ;
  assign n32572 = ( n32514 & n32555 ) | ( n32514 & ~n32571 ) | ( n32555 & ~n32571 ) ;
  assign n32573 = ~n32514 & n32572 ;
  assign n32574 = n32513 & ~n32573 ;
  assign n32575 = ( x789 & n32573 ) | ( x789 & ~n32574 ) | ( n32573 & ~n32574 ) ;
  assign n32576 = x626 & ~n32575 ;
  assign n32577 = ~n16279 & n32502 ;
  assign n32578 = x626 & ~n32577 ;
  assign n32583 = ( x641 & n32577 ) | ( x641 & n32578 ) | ( n32577 & n32578 ) ;
  assign n32584 = ~n32576 & n32583 ;
  assign n32498 = ~n18319 & n32497 ;
  assign n32585 = n16457 & n32498 ;
  assign n32586 = ( x1158 & n32584 ) | ( x1158 & ~n32585 ) | ( n32584 & ~n32585 ) ;
  assign n32587 = ~n32584 & n32586 ;
  assign n32499 = n16456 & n32498 ;
  assign n32579 = x641 | n32578 ;
  assign n32580 = ( n32575 & n32576 ) | ( n32575 & ~n32579 ) | ( n32576 & ~n32579 ) ;
  assign n32581 = ( x1158 & ~n32499 ) | ( x1158 & n32580 ) | ( ~n32499 & n32580 ) ;
  assign n32582 = n32499 | n32581 ;
  assign n32588 = n32587 ^ n32582 ^ 1'b0 ;
  assign n32589 = ( x788 & ~n32582 ) | ( x788 & n32587 ) | ( ~n32582 & n32587 ) ;
  assign n32590 = ( x788 & ~n32588 ) | ( x788 & n32589 ) | ( ~n32588 & n32589 ) ;
  assign n32591 = x788 | n32575 ;
  assign n32592 = ( n18482 & ~n32590 ) | ( n18482 & n32591 ) | ( ~n32590 & n32591 ) ;
  assign n32593 = ~n18482 & n32592 ;
  assign n32594 = ~n16518 & n32498 ;
  assign n32595 = x1156 & ~n32594 ;
  assign n32596 = ~x628 & x629 ;
  assign n32597 = ~n17088 & n32501 ;
  assign n32598 = x1156 | n32597 ;
  assign n32599 = ( n32595 & n32596 ) | ( n32595 & n32598 ) | ( n32596 & n32598 ) ;
  assign n32600 = ~n32595 & n32599 ;
  assign n32601 = x628 & ~x629 ;
  assign n32602 = x1156 & ~n32597 ;
  assign n32603 = n32601 & ~n32602 ;
  assign n32604 = n32603 ^ n32600 ^ 1'b0 ;
  assign n32605 = x1156 | n32594 ;
  assign n32606 = ( n32603 & ~n32604 ) | ( n32603 & n32605 ) | ( ~n32604 & n32605 ) ;
  assign n32607 = ( n32600 & n32604 ) | ( n32600 & n32606 ) | ( n32604 & n32606 ) ;
  assign n32608 = n32593 ^ x792 ^ 1'b0 ;
  assign n32609 = ( ~x792 & n32607 ) | ( ~x792 & n32608 ) | ( n32607 & n32608 ) ;
  assign n32610 = ( x792 & n32593 ) | ( x792 & n32609 ) | ( n32593 & n32609 ) ;
  assign n32611 = x207 & n32610 ;
  assign n32612 = x623 & ~n32611 ;
  assign n32613 = ~n2069 & n22522 ;
  assign n32614 = n15656 ^ x625 ^ 1'b0 ;
  assign n32615 = ( n15656 & n32613 ) | ( n15656 & n32614 ) | ( n32613 & n32614 ) ;
  assign n32616 = x1153 & ~n32615 ;
  assign n32617 = ( n15656 & n32613 ) | ( n15656 & ~n32614 ) | ( n32613 & ~n32614 ) ;
  assign n32618 = x1153 | n32617 ;
  assign n32619 = ~n32616 & n32618 ;
  assign n32620 = n32613 ^ x778 ^ 1'b0 ;
  assign n32621 = ( n32613 & n32619 ) | ( n32613 & n32620 ) | ( n32619 & n32620 ) ;
  assign n32622 = n32621 ^ n16234 ^ 1'b0 ;
  assign n32623 = ( n15656 & n32621 ) | ( n15656 & n32622 ) | ( n32621 & n32622 ) ;
  assign n32624 = n32623 ^ n16254 ^ 1'b0 ;
  assign n32625 = ( n15656 & n32623 ) | ( n15656 & n32624 ) | ( n32623 & n32624 ) ;
  assign n32626 = n32625 ^ n16279 ^ 1'b0 ;
  assign n32627 = ( n15656 & n32625 ) | ( n15656 & n32626 ) | ( n32625 & n32626 ) ;
  assign n32628 = n32627 ^ n16318 ^ 1'b0 ;
  assign n32629 = ( n15656 & n32627 ) | ( n15656 & n32628 ) | ( n32627 & n32628 ) ;
  assign n32630 = n15656 ^ x628 ^ 1'b0 ;
  assign n32631 = ( n15656 & n32629 ) | ( n15656 & n32630 ) | ( n32629 & n32630 ) ;
  assign n32632 = x629 | n32631 ;
  assign n32633 = x1156 & ~n32632 ;
  assign n32634 = ( n15656 & n32629 ) | ( n15656 & ~n32630 ) | ( n32629 & ~n32630 ) ;
  assign n32635 = ( x629 & x1156 ) | ( x629 & ~n32634 ) | ( x1156 & ~n32634 ) ;
  assign n32636 = ~x1156 & n32635 ;
  assign n32637 = ~n2069 & n17843 ;
  assign n32638 = n32637 ^ n15659 ^ 1'b0 ;
  assign n32639 = ( n15656 & n32637 ) | ( n15656 & n32638 ) | ( n32637 & n32638 ) ;
  assign n32640 = ~n15656 & n15662 ;
  assign n32641 = n15659 | n32637 ;
  assign n32642 = x609 | n32641 ;
  assign n32643 = n32642 ^ n32640 ^ 1'b0 ;
  assign n32644 = ( n32640 & n32642 ) | ( n32640 & n32643 ) | ( n32642 & n32643 ) ;
  assign n32645 = ( x1155 & ~n32640 ) | ( x1155 & n32644 ) | ( ~n32640 & n32644 ) ;
  assign n32646 = x609 & ~n32641 ;
  assign n32647 = n15656 | n15668 ;
  assign n32648 = x1155 & ~n32647 ;
  assign n32649 = ( x1155 & n32646 ) | ( x1155 & n32648 ) | ( n32646 & n32648 ) ;
  assign n32650 = n32645 & ~n32649 ;
  assign n32651 = n32639 ^ x785 ^ 1'b0 ;
  assign n32652 = ( n32639 & n32650 ) | ( n32639 & n32651 ) | ( n32650 & n32651 ) ;
  assign n32653 = ~x618 & n32652 ;
  assign n32654 = x618 & n15656 ;
  assign n32655 = ( x1154 & ~n32653 ) | ( x1154 & n32654 ) | ( ~n32653 & n32654 ) ;
  assign n32656 = n32653 | n32655 ;
  assign n32657 = ~x618 & n15656 ;
  assign n32658 = x618 & n32652 ;
  assign n32659 = ( x1154 & n32657 ) | ( x1154 & ~n32658 ) | ( n32657 & ~n32658 ) ;
  assign n32660 = ~n32657 & n32659 ;
  assign n32661 = n32656 & ~n32660 ;
  assign n32662 = n32652 ^ x781 ^ 1'b0 ;
  assign n32663 = ( n32652 & n32661 ) | ( n32652 & n32662 ) | ( n32661 & n32662 ) ;
  assign n32664 = ~x619 & n32663 ;
  assign n32665 = x619 & n15656 ;
  assign n32666 = ( x1159 & ~n32664 ) | ( x1159 & n32665 ) | ( ~n32664 & n32665 ) ;
  assign n32667 = n32664 | n32666 ;
  assign n32668 = ~x619 & n15656 ;
  assign n32669 = x619 & n32663 ;
  assign n32670 = ( x1159 & n32668 ) | ( x1159 & ~n32669 ) | ( n32668 & ~n32669 ) ;
  assign n32671 = ~n32668 & n32670 ;
  assign n32672 = n32667 & ~n32671 ;
  assign n32673 = n32663 ^ x789 ^ 1'b0 ;
  assign n32674 = ( n32663 & n32672 ) | ( n32663 & n32673 ) | ( n32672 & n32673 ) ;
  assign n32675 = n32674 ^ n16518 ^ 1'b0 ;
  assign n32676 = ( n15656 & n32674 ) | ( n15656 & n32675 ) | ( n32674 & n32675 ) ;
  assign n32677 = n19046 & ~n32676 ;
  assign n32678 = n32636 | n32677 ;
  assign n32679 = ( x792 & n32633 ) | ( x792 & n32678 ) | ( n32633 & n32678 ) ;
  assign n32680 = n32678 ^ n32633 ^ 1'b0 ;
  assign n32681 = ( x792 & n32679 ) | ( x792 & n32680 ) | ( n32679 & n32680 ) ;
  assign n32682 = n32625 ^ x619 ^ 1'b0 ;
  assign n32683 = x660 | n32649 ;
  assign n32702 = x609 & ~n32621 ;
  assign n32684 = x608 | n32616 ;
  assign n32685 = ~n2069 & n17902 ;
  assign n32686 = ~x625 & n32685 ;
  assign n32687 = x1153 | n32686 ;
  assign n32688 = x625 & n32637 ;
  assign n32689 = ( ~n32684 & n32687 ) | ( ~n32684 & n32688 ) | ( n32687 & n32688 ) ;
  assign n32690 = ~n32684 & n32689 ;
  assign n32691 = x625 & n32685 ;
  assign n32692 = ~x625 & n32637 ;
  assign n32693 = ( x1153 & n32691 ) | ( x1153 & ~n32692 ) | ( n32691 & ~n32692 ) ;
  assign n32694 = ~n32691 & n32693 ;
  assign n32695 = ( x608 & n32618 ) | ( x608 & n32694 ) | ( n32618 & n32694 ) ;
  assign n32696 = ~n32694 & n32695 ;
  assign n32697 = ( x778 & n32690 ) | ( x778 & ~n32696 ) | ( n32690 & ~n32696 ) ;
  assign n32698 = ~n32690 & n32697 ;
  assign n32699 = ( x778 & n32685 ) | ( x778 & ~n32698 ) | ( n32685 & ~n32698 ) ;
  assign n32700 = ~n32698 & n32699 ;
  assign n32701 = x609 & ~n32700 ;
  assign n32703 = n32702 ^ n32701 ^ n32700 ;
  assign n32704 = ( x1155 & ~n32683 ) | ( x1155 & n32703 ) | ( ~n32683 & n32703 ) ;
  assign n32705 = ~n32683 & n32704 ;
  assign n32706 = x609 | n32621 ;
  assign n32707 = x1155 & ~n32706 ;
  assign n32708 = ( x1155 & n32701 ) | ( x1155 & n32707 ) | ( n32701 & n32707 ) ;
  assign n32709 = ( x660 & n32645 ) | ( x660 & n32708 ) | ( n32645 & n32708 ) ;
  assign n32710 = ~n32708 & n32709 ;
  assign n32711 = ( x785 & n32705 ) | ( x785 & ~n32710 ) | ( n32705 & ~n32710 ) ;
  assign n32712 = ~n32705 & n32711 ;
  assign n32713 = ( x785 & n32700 ) | ( x785 & ~n32712 ) | ( n32700 & ~n32712 ) ;
  assign n32714 = ~n32712 & n32713 ;
  assign n32715 = x627 | n32660 ;
  assign n32717 = x618 & ~n32623 ;
  assign n32716 = x618 & ~n32714 ;
  assign n32718 = n32717 ^ n32716 ^ n32714 ;
  assign n32719 = ( x1154 & ~n32715 ) | ( x1154 & n32718 ) | ( ~n32715 & n32718 ) ;
  assign n32720 = ~n32715 & n32719 ;
  assign n32721 = x627 & n32656 ;
  assign n32722 = x618 | n32623 ;
  assign n32723 = x1154 & ~n32722 ;
  assign n32724 = ( x1154 & n32716 ) | ( x1154 & n32723 ) | ( n32716 & n32723 ) ;
  assign n32725 = ( n32720 & n32721 ) | ( n32720 & ~n32724 ) | ( n32721 & ~n32724 ) ;
  assign n32726 = n32725 ^ n32721 ^ 1'b0 ;
  assign n32727 = ( n32720 & n32725 ) | ( n32720 & ~n32726 ) | ( n32725 & ~n32726 ) ;
  assign n32728 = n32714 ^ x781 ^ 1'b0 ;
  assign n32729 = ( n32714 & n32727 ) | ( n32714 & n32728 ) | ( n32727 & n32728 ) ;
  assign n32730 = ( n32625 & n32682 ) | ( n32625 & n32729 ) | ( n32682 & n32729 ) ;
  assign n32731 = x1159 & ~n32730 ;
  assign n32732 = ( x648 & n32667 ) | ( x648 & n32731 ) | ( n32667 & n32731 ) ;
  assign n32733 = ~n32731 & n32732 ;
  assign n32734 = x648 | n32671 ;
  assign n32735 = ( n32625 & ~n32682 ) | ( n32625 & n32729 ) | ( ~n32682 & n32729 ) ;
  assign n32736 = ( x1159 & ~n32734 ) | ( x1159 & n32735 ) | ( ~n32734 & n32735 ) ;
  assign n32737 = ~n32734 & n32736 ;
  assign n32738 = ( x789 & n32733 ) | ( x789 & ~n32737 ) | ( n32733 & ~n32737 ) ;
  assign n32739 = ~n32733 & n32738 ;
  assign n32740 = x789 | n32729 ;
  assign n32741 = ( n16519 & ~n32739 ) | ( n16519 & n32740 ) | ( ~n32739 & n32740 ) ;
  assign n32742 = ~n16519 & n32741 ;
  assign n32743 = x641 | n15656 ;
  assign n32744 = n16453 & n32743 ;
  assign n32745 = x641 & ~n32627 ;
  assign n32746 = x641 & ~n15656 ;
  assign n32747 = n16454 & ~n32746 ;
  assign n32748 = ( n32627 & n32745 ) | ( n32627 & n32747 ) | ( n32745 & n32747 ) ;
  assign n32749 = n32745 & ~n32748 ;
  assign n32750 = ( n32744 & n32748 ) | ( n32744 & ~n32749 ) | ( n32748 & ~n32749 ) ;
  assign n32751 = n16317 & n16458 ;
  assign n32752 = n32750 ^ n32674 ^ 1'b0 ;
  assign n32753 = ( ~n32674 & n32751 ) | ( ~n32674 & n32752 ) | ( n32751 & n32752 ) ;
  assign n32754 = ( n32674 & n32750 ) | ( n32674 & n32753 ) | ( n32750 & n32753 ) ;
  assign n32755 = ( x788 & ~n22314 ) | ( x788 & n32754 ) | ( ~n22314 & n32754 ) ;
  assign n32756 = ( n18482 & n22314 ) | ( n18482 & n32755 ) | ( n22314 & n32755 ) ;
  assign n32757 = ( ~n32681 & n32742 ) | ( ~n32681 & n32756 ) | ( n32742 & n32756 ) ;
  assign n32758 = ~n32681 & n32757 ;
  assign n32759 = x207 | n32758 ;
  assign n32760 = n32612 & n32759 ;
  assign n32761 = x628 | n15656 ;
  assign n32762 = ( x1156 & n32633 ) | ( x1156 & ~n32761 ) | ( n32633 & ~n32761 ) ;
  assign n32763 = x628 & ~n15656 ;
  assign n32764 = ( ~x1156 & n32636 ) | ( ~x1156 & n32763 ) | ( n32636 & n32763 ) ;
  assign n32765 = ( x792 & n32762 ) | ( x792 & n32764 ) | ( n32762 & n32764 ) ;
  assign n32766 = n32764 ^ n32762 ^ 1'b0 ;
  assign n32767 = ( x792 & n32765 ) | ( x792 & n32766 ) | ( n32765 & n32766 ) ;
  assign n32768 = x626 & n32627 ;
  assign n32769 = x1159 & ~n15656 ;
  assign n32770 = x648 | n32769 ;
  assign n32771 = x1154 & ~n15656 ;
  assign n32772 = x627 | n32771 ;
  assign n32773 = x1155 & ~n15656 ;
  assign n32774 = x660 | n32773 ;
  assign n32775 = ~n2069 & n17893 ;
  assign n32776 = ( n15656 & n32614 ) | ( n15656 & n32775 ) | ( n32614 & n32775 ) ;
  assign n32777 = x1153 & ~n32776 ;
  assign n32778 = ( x608 & n32618 ) | ( x608 & n32777 ) | ( n32618 & n32777 ) ;
  assign n32779 = ~n32777 & n32778 ;
  assign n32780 = ( n15656 & ~n32614 ) | ( n15656 & n32775 ) | ( ~n32614 & n32775 ) ;
  assign n32781 = x1153 | n32780 ;
  assign n32782 = ( x608 & ~n32616 ) | ( x608 & n32781 ) | ( ~n32616 & n32781 ) ;
  assign n32783 = ~x608 & n32782 ;
  assign n32784 = ( x778 & n32779 ) | ( x778 & ~n32783 ) | ( n32779 & ~n32783 ) ;
  assign n32785 = ~n32779 & n32784 ;
  assign n32786 = ( x778 & n32775 ) | ( x778 & ~n32785 ) | ( n32775 & ~n32785 ) ;
  assign n32787 = ~n32785 & n32786 ;
  assign n32788 = x609 & ~n32787 ;
  assign n32789 = n32706 & ~n32788 ;
  assign n32790 = n32789 ^ n32787 ^ n32621 ;
  assign n32791 = ( x1155 & ~n32774 ) | ( x1155 & n32790 ) | ( ~n32774 & n32790 ) ;
  assign n32792 = ~n32774 & n32791 ;
  assign n32793 = x1155 & ~n32789 ;
  assign n32794 = x1155 | n15656 ;
  assign n32795 = ( x660 & n32793 ) | ( x660 & n32794 ) | ( n32793 & n32794 ) ;
  assign n32796 = ~n32793 & n32795 ;
  assign n32797 = ( x785 & n32792 ) | ( x785 & ~n32796 ) | ( n32792 & ~n32796 ) ;
  assign n32798 = ~n32792 & n32797 ;
  assign n32799 = ( x785 & n32787 ) | ( x785 & ~n32798 ) | ( n32787 & ~n32798 ) ;
  assign n32800 = ~n32798 & n32799 ;
  assign n32801 = x618 & ~n32800 ;
  assign n32802 = n32722 & ~n32801 ;
  assign n32803 = n32802 ^ n32800 ^ n32623 ;
  assign n32804 = ( x1154 & ~n32772 ) | ( x1154 & n32803 ) | ( ~n32772 & n32803 ) ;
  assign n32805 = ~n32772 & n32804 ;
  assign n32806 = x1154 & ~n32802 ;
  assign n32807 = x1154 | n15656 ;
  assign n32808 = ( x627 & n32806 ) | ( x627 & n32807 ) | ( n32806 & n32807 ) ;
  assign n32809 = ~n32806 & n32808 ;
  assign n32810 = ( x781 & n32805 ) | ( x781 & ~n32809 ) | ( n32805 & ~n32809 ) ;
  assign n32811 = ~n32805 & n32810 ;
  assign n32812 = ( x781 & n32800 ) | ( x781 & ~n32811 ) | ( n32800 & ~n32811 ) ;
  assign n32813 = ~n32811 & n32812 ;
  assign n32814 = ( n32625 & ~n32682 ) | ( n32625 & n32813 ) | ( ~n32682 & n32813 ) ;
  assign n32815 = ( x1159 & ~n32770 ) | ( x1159 & n32814 ) | ( ~n32770 & n32814 ) ;
  assign n32816 = ~n32770 & n32815 ;
  assign n32817 = ( n32625 & n32682 ) | ( n32625 & n32813 ) | ( n32682 & n32813 ) ;
  assign n32818 = x1159 & ~n32817 ;
  assign n32819 = x1159 | n15656 ;
  assign n32820 = ( x648 & n32818 ) | ( x648 & n32819 ) | ( n32818 & n32819 ) ;
  assign n32821 = ~n32818 & n32820 ;
  assign n32822 = ( x789 & n32816 ) | ( x789 & ~n32821 ) | ( n32816 & ~n32821 ) ;
  assign n32823 = ~n32816 & n32822 ;
  assign n32824 = ( x789 & n32813 ) | ( x789 & ~n32823 ) | ( n32813 & ~n32823 ) ;
  assign n32825 = ~n32823 & n32824 ;
  assign n32826 = ~x626 & n32825 ;
  assign n32827 = ( x641 & ~n32768 ) | ( x641 & n32826 ) | ( ~n32768 & n32826 ) ;
  assign n32828 = n32768 | n32827 ;
  assign n32829 = ( x1158 & ~n32746 ) | ( x1158 & n32828 ) | ( ~n32746 & n32828 ) ;
  assign n32830 = ~x1158 & n32829 ;
  assign n32831 = x626 & n32825 ;
  assign n32832 = ~x626 & n32627 ;
  assign n32833 = ( x641 & n32831 ) | ( x641 & ~n32832 ) | ( n32831 & ~n32832 ) ;
  assign n32834 = ~n32831 & n32833 ;
  assign n32835 = ( x1158 & n32743 ) | ( x1158 & n32834 ) | ( n32743 & n32834 ) ;
  assign n32836 = ~n32834 & n32835 ;
  assign n32837 = ( x788 & n32830 ) | ( x788 & n32836 ) | ( n32830 & n32836 ) ;
  assign n32838 = n32836 ^ n32830 ^ 1'b0 ;
  assign n32839 = ( x788 & n32837 ) | ( x788 & n32838 ) | ( n32837 & n32838 ) ;
  assign n32840 = ~x788 & n32825 ;
  assign n32841 = n18482 | n32840 ;
  assign n32842 = ( ~n32767 & n32839 ) | ( ~n32767 & n32841 ) | ( n32839 & n32841 ) ;
  assign n32843 = ~n32767 & n32842 ;
  assign n32844 = x207 | n32843 ;
  assign n32845 = x1158 & n32583 ;
  assign n32847 = x625 & n31746 ;
  assign n32848 = x1153 & ~n32847 ;
  assign n32849 = n32518 & ~n32848 ;
  assign n32850 = ~x625 & n31746 ;
  assign n32851 = x1153 | n32850 ;
  assign n32852 = ~n32526 & n32851 ;
  assign n32853 = ( x778 & n32849 ) | ( x778 & ~n32852 ) | ( n32849 & ~n32852 ) ;
  assign n32854 = ~n32849 & n32853 ;
  assign n32855 = ( x778 & n31746 ) | ( x778 & ~n32854 ) | ( n31746 & ~n32854 ) ;
  assign n32856 = ~n32854 & n32855 ;
  assign n32857 = x609 & ~n32856 ;
  assign n32859 = n16231 | n32537 ;
  assign n32860 = ( n32856 & n32857 ) | ( n32856 & ~n32859 ) | ( n32857 & ~n32859 ) ;
  assign n32846 = n16232 & n32542 ;
  assign n32858 = n32846 & ~n32857 ;
  assign n32861 = ( x785 & ~n32858 ) | ( x785 & n32860 ) | ( ~n32858 & n32860 ) ;
  assign n32862 = ~n32860 & n32861 ;
  assign n32863 = ( x785 & n32856 ) | ( x785 & ~n32862 ) | ( n32856 & ~n32862 ) ;
  assign n32864 = ~n32862 & n32863 ;
  assign n32865 = x781 | n32864 ;
  assign n32866 = n16252 & n32562 ;
  assign n32867 = x618 & ~n32864 ;
  assign n32868 = n32866 & ~n32867 ;
  assign n32869 = n16251 | n32559 ;
  assign n32870 = ( n32864 & n32867 ) | ( n32864 & ~n32869 ) | ( n32867 & ~n32869 ) ;
  assign n32871 = ( x781 & n32868 ) | ( x781 & ~n32870 ) | ( n32868 & ~n32870 ) ;
  assign n32872 = ~n32868 & n32871 ;
  assign n32873 = ( n21705 & n32865 ) | ( n21705 & ~n32872 ) | ( n32865 & ~n32872 ) ;
  assign n32874 = ~n21705 & n32873 ;
  assign n32875 = n32874 ^ n32502 ^ 1'b0 ;
  assign n32876 = ~n16278 & n18319 ;
  assign n32877 = ( n32502 & ~n32875 ) | ( n32502 & n32876 ) | ( ~n32875 & n32876 ) ;
  assign n32878 = ( n32874 & n32875 ) | ( n32874 & n32877 ) | ( n32875 & n32877 ) ;
  assign n32879 = x626 & ~n32878 ;
  assign n32880 = n32845 & ~n32879 ;
  assign n32881 = x1158 | n32579 ;
  assign n32882 = ( n32878 & n32879 ) | ( n32878 & ~n32881 ) | ( n32879 & ~n32881 ) ;
  assign n32883 = ( x788 & n32880 ) | ( x788 & ~n32882 ) | ( n32880 & ~n32882 ) ;
  assign n32884 = ~n32880 & n32883 ;
  assign n32885 = x788 | n32878 ;
  assign n32886 = ( n18482 & ~n32884 ) | ( n18482 & n32885 ) | ( ~n32884 & n32885 ) ;
  assign n32887 = ~n18482 & n32886 ;
  assign n32888 = n16339 & ~n16558 ;
  assign n32889 = n32887 ^ n32597 ^ 1'b0 ;
  assign n32890 = ( ~n32597 & n32888 ) | ( ~n32597 & n32889 ) | ( n32888 & n32889 ) ;
  assign n32891 = ( n32597 & n32887 ) | ( n32597 & n32890 ) | ( n32887 & n32890 ) ;
  assign n32892 = x207 & n32891 ;
  assign n32893 = ( x623 & n32844 ) | ( x623 & ~n32892 ) | ( n32844 & ~n32892 ) ;
  assign n32894 = ~x623 & n32893 ;
  assign n32895 = ( x710 & n32760 ) | ( x710 & ~n32894 ) | ( n32760 & ~n32894 ) ;
  assign n32896 = ~n32760 & n32895 ;
  assign n32897 = ~n16339 & n32594 ;
  assign n32898 = x207 & ~n32897 ;
  assign n32899 = n32676 ^ n16339 ^ 1'b0 ;
  assign n32900 = ( n15656 & n32676 ) | ( n15656 & n32899 ) | ( n32676 & n32899 ) ;
  assign n32901 = ~x207 & n32900 ;
  assign n32902 = ( x623 & n32898 ) | ( x623 & ~n32901 ) | ( n32898 & ~n32901 ) ;
  assign n32903 = ~n32898 & n32902 ;
  assign n32904 = x207 | n15656 ;
  assign n32905 = ( x623 & ~n32903 ) | ( x623 & n32904 ) | ( ~n32903 & n32904 ) ;
  assign n32906 = ~n32903 & n32905 ;
  assign n32907 = x710 | n32906 ;
  assign n32908 = ( n18484 & ~n32896 ) | ( n18484 & n32907 ) | ( ~n32896 & n32907 ) ;
  assign n32909 = ~n18484 & n32908 ;
  assign n32910 = x647 & ~n32904 ;
  assign n32911 = x1157 | n32910 ;
  assign n32912 = ~n17093 & n32597 ;
  assign n32913 = ~n17093 & n32629 ;
  assign n32914 = n15656 & n16559 ;
  assign n32915 = n32913 | n32914 ;
  assign n32916 = n32915 ^ x207 ^ 1'b0 ;
  assign n32917 = ( ~n32912 & n32915 ) | ( ~n32912 & n32916 ) | ( n32915 & n32916 ) ;
  assign n32918 = n32917 ^ x710 ^ 1'b0 ;
  assign n32919 = ( n32904 & n32917 ) | ( n32904 & ~n32918 ) | ( n32917 & ~n32918 ) ;
  assign n32920 = x647 & ~n32919 ;
  assign n32921 = ( ~n32911 & n32919 ) | ( ~n32911 & n32920 ) | ( n32919 & n32920 ) ;
  assign n32922 = x630 & n32921 ;
  assign n32923 = n19055 & n32906 ;
  assign n32924 = x647 | n32904 ;
  assign n32925 = ( x1157 & n32920 ) | ( x1157 & n32924 ) | ( n32920 & n32924 ) ;
  assign n32926 = ~n32920 & n32925 ;
  assign n32927 = ~x630 & n32926 ;
  assign n32928 = ( ~n32922 & n32923 ) | ( ~n32922 & n32927 ) | ( n32923 & n32927 ) ;
  assign n32929 = n32922 | n32928 ;
  assign n32930 = n32909 ^ x787 ^ 1'b0 ;
  assign n32931 = ( ~x787 & n32929 ) | ( ~x787 & n32930 ) | ( n32929 & n32930 ) ;
  assign n32932 = ( x787 & n32909 ) | ( x787 & n32931 ) | ( n32909 & n32931 ) ;
  assign n32933 = x644 & ~n32932 ;
  assign n32934 = n32921 | n32926 ;
  assign n32935 = n32919 ^ x787 ^ 1'b0 ;
  assign n32936 = ( n32919 & n32934 ) | ( n32919 & n32935 ) | ( n32934 & n32935 ) ;
  assign n32937 = x644 | n32936 ;
  assign n32938 = ( x715 & n32933 ) | ( x715 & n32937 ) | ( n32933 & n32937 ) ;
  assign n32939 = ~n32933 & n32938 ;
  assign n32940 = x644 | n32904 ;
  assign n32941 = n32904 ^ n16376 ^ 1'b0 ;
  assign n32942 = ( n32904 & n32906 ) | ( n32904 & ~n32941 ) | ( n32906 & ~n32941 ) ;
  assign n32943 = x644 & ~n32942 ;
  assign n32944 = ( x715 & n32940 ) | ( x715 & ~n32943 ) | ( n32940 & ~n32943 ) ;
  assign n32945 = ~x715 & n32944 ;
  assign n32946 = ( x1160 & n32939 ) | ( x1160 & ~n32945 ) | ( n32939 & ~n32945 ) ;
  assign n32947 = ~n32939 & n32946 ;
  assign n32948 = x644 & ~n32904 ;
  assign n32949 = x715 & ~n32948 ;
  assign n32950 = ( n32942 & n32943 ) | ( n32942 & n32949 ) | ( n32943 & n32949 ) ;
  assign n32951 = x644 & ~n32936 ;
  assign n32952 = x715 | n32951 ;
  assign n32953 = ( n32932 & n32933 ) | ( n32932 & ~n32952 ) | ( n32933 & ~n32952 ) ;
  assign n32954 = ( x1160 & ~n32950 ) | ( x1160 & n32953 ) | ( ~n32950 & n32953 ) ;
  assign n32955 = n32950 | n32954 ;
  assign n32956 = x790 & ~n32955 ;
  assign n32957 = ( x790 & n32947 ) | ( x790 & n32956 ) | ( n32947 & n32956 ) ;
  assign n32958 = ( x790 & n32932 ) | ( x790 & ~n32957 ) | ( n32932 & ~n32957 ) ;
  assign n32959 = ~n32957 & n32958 ;
  assign n32960 = n32959 ^ n7318 ^ 1'b0 ;
  assign n32961 = ( x207 & n32959 ) | ( x207 & n32960 ) | ( n32959 & n32960 ) ;
  assign n32962 = x208 & n32610 ;
  assign n32963 = x607 & ~n32962 ;
  assign n32964 = x208 | n32758 ;
  assign n32965 = n32963 & n32964 ;
  assign n32966 = x208 | n32843 ;
  assign n32967 = x208 & n32891 ;
  assign n32968 = ( x607 & n32966 ) | ( x607 & ~n32967 ) | ( n32966 & ~n32967 ) ;
  assign n32969 = ~x607 & n32968 ;
  assign n32970 = ( x638 & n32965 ) | ( x638 & ~n32969 ) | ( n32965 & ~n32969 ) ;
  assign n32971 = ~n32965 & n32970 ;
  assign n32972 = x208 & ~n32897 ;
  assign n32973 = ~x208 & n32900 ;
  assign n32974 = ( x607 & n32972 ) | ( x607 & ~n32973 ) | ( n32972 & ~n32973 ) ;
  assign n32975 = ~n32972 & n32974 ;
  assign n32976 = x208 | n15656 ;
  assign n32977 = ( x607 & ~n32975 ) | ( x607 & n32976 ) | ( ~n32975 & n32976 ) ;
  assign n32978 = ~n32975 & n32977 ;
  assign n32979 = x638 | n32978 ;
  assign n32980 = ( n18484 & ~n32971 ) | ( n18484 & n32979 ) | ( ~n32971 & n32979 ) ;
  assign n32981 = ~n18484 & n32980 ;
  assign n32982 = x647 & ~n32976 ;
  assign n32983 = x1157 | n32982 ;
  assign n32984 = n32915 ^ x208 ^ 1'b0 ;
  assign n32985 = ( ~n32912 & n32915 ) | ( ~n32912 & n32984 ) | ( n32915 & n32984 ) ;
  assign n32986 = n32985 ^ x638 ^ 1'b0 ;
  assign n32987 = ( n32976 & n32985 ) | ( n32976 & ~n32986 ) | ( n32985 & ~n32986 ) ;
  assign n32988 = x647 & ~n32987 ;
  assign n32989 = ( ~n32983 & n32987 ) | ( ~n32983 & n32988 ) | ( n32987 & n32988 ) ;
  assign n32990 = x630 & n32989 ;
  assign n32991 = n19055 & n32978 ;
  assign n32992 = x647 | n32976 ;
  assign n32993 = ( x1157 & n32988 ) | ( x1157 & n32992 ) | ( n32988 & n32992 ) ;
  assign n32994 = ~n32988 & n32993 ;
  assign n32995 = ~x630 & n32994 ;
  assign n32996 = ( ~n32990 & n32991 ) | ( ~n32990 & n32995 ) | ( n32991 & n32995 ) ;
  assign n32997 = n32990 | n32996 ;
  assign n32998 = n32981 ^ x787 ^ 1'b0 ;
  assign n32999 = ( ~x787 & n32997 ) | ( ~x787 & n32998 ) | ( n32997 & n32998 ) ;
  assign n33000 = ( x787 & n32981 ) | ( x787 & n32999 ) | ( n32981 & n32999 ) ;
  assign n33001 = x644 & ~n33000 ;
  assign n33002 = n32989 | n32994 ;
  assign n33003 = n32987 ^ x787 ^ 1'b0 ;
  assign n33004 = ( n32987 & n33002 ) | ( n32987 & n33003 ) | ( n33002 & n33003 ) ;
  assign n33005 = x644 | n33004 ;
  assign n33006 = ( x715 & n33001 ) | ( x715 & n33005 ) | ( n33001 & n33005 ) ;
  assign n33007 = ~n33001 & n33006 ;
  assign n33008 = x644 | n32976 ;
  assign n33009 = n32976 ^ n16376 ^ 1'b0 ;
  assign n33010 = ( n32976 & n32978 ) | ( n32976 & ~n33009 ) | ( n32978 & ~n33009 ) ;
  assign n33011 = x644 & ~n33010 ;
  assign n33012 = ( x715 & n33008 ) | ( x715 & ~n33011 ) | ( n33008 & ~n33011 ) ;
  assign n33013 = ~x715 & n33012 ;
  assign n33014 = ( x1160 & n33007 ) | ( x1160 & ~n33013 ) | ( n33007 & ~n33013 ) ;
  assign n33015 = ~n33007 & n33014 ;
  assign n33016 = x644 & ~n32976 ;
  assign n33017 = x715 & ~n33016 ;
  assign n33018 = ( n33010 & n33011 ) | ( n33010 & n33017 ) | ( n33011 & n33017 ) ;
  assign n33019 = x644 & ~n33004 ;
  assign n33020 = x715 | n33019 ;
  assign n33021 = ( n33000 & n33001 ) | ( n33000 & ~n33020 ) | ( n33001 & ~n33020 ) ;
  assign n33022 = ( x1160 & ~n33018 ) | ( x1160 & n33021 ) | ( ~n33018 & n33021 ) ;
  assign n33023 = n33018 | n33022 ;
  assign n33024 = x790 & ~n33023 ;
  assign n33025 = ( x790 & n33015 ) | ( x790 & n33024 ) | ( n33015 & n33024 ) ;
  assign n33026 = ( x790 & n33000 ) | ( x790 & ~n33025 ) | ( n33000 & ~n33025 ) ;
  assign n33027 = ~n33025 & n33026 ;
  assign n33028 = n33027 ^ n7318 ^ 1'b0 ;
  assign n33029 = ( x208 & n33027 ) | ( x208 & n33028 ) | ( n33027 & n33028 ) ;
  assign n33030 = ~x647 & n32912 ;
  assign n33031 = x1157 | n33030 ;
  assign n33032 = ~x647 & n32897 ;
  assign n33033 = x647 & n32610 ;
  assign n33034 = ( x1157 & n33032 ) | ( x1157 & ~n33033 ) | ( n33032 & ~n33033 ) ;
  assign n33035 = ~n33032 & n33034 ;
  assign n33036 = x630 & ~n33035 ;
  assign n33037 = n33031 & n33036 ;
  assign n33038 = ~x647 & n32610 ;
  assign n33039 = x647 & n32897 ;
  assign n33040 = ( x1157 & ~n33038 ) | ( x1157 & n33039 ) | ( ~n33038 & n33039 ) ;
  assign n33041 = n33038 | n33040 ;
  assign n33042 = x647 & n32912 ;
  assign n33043 = x1157 & ~n33042 ;
  assign n33044 = ( x630 & n33041 ) | ( x630 & ~n33043 ) | ( n33041 & ~n33043 ) ;
  assign n33045 = ~x630 & n33044 ;
  assign n33046 = ( x787 & n33037 ) | ( x787 & ~n33045 ) | ( n33037 & ~n33045 ) ;
  assign n33047 = ~n33037 & n33046 ;
  assign n33048 = ( x787 & n32610 ) | ( x787 & ~n33047 ) | ( n32610 & ~n33047 ) ;
  assign n33049 = ~n33047 & n33048 ;
  assign n33050 = x790 | n33049 ;
  assign n33054 = x644 & ~n33049 ;
  assign n33055 = ~n17273 & n32912 ;
  assign n33056 = x644 & ~n33055 ;
  assign n33061 = ( x715 & n33055 ) | ( x715 & n33056 ) | ( n33055 & n33056 ) ;
  assign n33062 = ~n33054 & n33061 ;
  assign n33051 = ~n21755 & n32594 ;
  assign n33063 = x644 & ~x715 ;
  assign n33064 = n33051 & n33063 ;
  assign n33065 = ( x1160 & n33062 ) | ( x1160 & ~n33064 ) | ( n33062 & ~n33064 ) ;
  assign n33066 = ~n33062 & n33065 ;
  assign n33052 = ~x644 & x715 ;
  assign n33053 = n33051 & n33052 ;
  assign n33057 = x715 | n33056 ;
  assign n33058 = ( n33049 & n33054 ) | ( n33049 & ~n33057 ) | ( n33054 & ~n33057 ) ;
  assign n33059 = ( x1160 & ~n33053 ) | ( x1160 & n33058 ) | ( ~n33053 & n33058 ) ;
  assign n33060 = n33053 | n33059 ;
  assign n33067 = n33066 ^ n33060 ^ 1'b0 ;
  assign n33068 = ( x790 & ~n33060 ) | ( x790 & n33066 ) | ( ~n33060 & n33066 ) ;
  assign n33069 = ( x790 & ~n33067 ) | ( x790 & n33068 ) | ( ~n33067 & n33068 ) ;
  assign n33070 = ( n7318 & n33050 ) | ( n7318 & ~n33069 ) | ( n33050 & ~n33069 ) ;
  assign n33071 = ~n7318 & n33070 ;
  assign n33072 = x622 & x639 ;
  assign n33073 = ~n33071 & n33072 ;
  assign n33074 = x1160 ^ x644 ^ 1'b0 ;
  assign n33075 = x790 & n33074 ;
  assign n33076 = n7318 | n33075 ;
  assign n33077 = n33051 & ~n33076 ;
  assign n33078 = x622 & n33077 ;
  assign n33079 = x639 | n33078 ;
  assign n33080 = x209 & n33079 ;
  assign n33081 = n16376 & ~n17272 ;
  assign n33082 = n32912 & n33081 ;
  assign n33083 = ~n18484 & n32891 ;
  assign n33084 = n33082 | n33083 ;
  assign n33085 = x790 | n33084 ;
  assign n33086 = x644 & ~n33084 ;
  assign n33089 = x1160 | n33057 ;
  assign n33090 = ( n33084 & n33086 ) | ( n33084 & ~n33089 ) | ( n33086 & ~n33089 ) ;
  assign n33087 = x1160 & n33061 ;
  assign n33088 = ~n33086 & n33087 ;
  assign n33091 = ( x790 & ~n33088 ) | ( x790 & n33090 ) | ( ~n33088 & n33090 ) ;
  assign n33092 = ~n33090 & n33091 ;
  assign n33093 = ( n7318 & n33085 ) | ( n7318 & ~n33092 ) | ( n33085 & ~n33092 ) ;
  assign n33094 = ~n7318 & n33093 ;
  assign n33095 = x622 | n33094 ;
  assign n33096 = ( n33073 & n33080 ) | ( n33073 & n33095 ) | ( n33080 & n33095 ) ;
  assign n33097 = ~n33073 & n33096 ;
  assign n33098 = x647 & ~n15656 ;
  assign n33099 = x647 | n32915 ;
  assign n33100 = ~n33098 & n33099 ;
  assign n33101 = n33100 ^ n32915 ^ n15656 ;
  assign n33102 = x630 | n33101 ;
  assign n33103 = ( x647 & n33101 ) | ( x647 & n33102 ) | ( n33101 & n33102 ) ;
  assign n33104 = x1157 & ~n33103 ;
  assign n33105 = n16374 & ~n33100 ;
  assign n33106 = ~x1157 & n33098 ;
  assign n33107 = n33105 | n33106 ;
  assign n33108 = ( x787 & n33104 ) | ( x787 & n33107 ) | ( n33104 & n33107 ) ;
  assign n33109 = n33107 ^ n33104 ^ 1'b0 ;
  assign n33110 = ( x787 & n33108 ) | ( x787 & n33109 ) | ( n33108 & n33109 ) ;
  assign n33111 = ( n18484 & n32843 ) | ( n18484 & ~n33110 ) | ( n32843 & ~n33110 ) ;
  assign n33112 = ~n33110 & n33111 ;
  assign n33113 = x790 | n33112 ;
  assign n33115 = x644 & ~n33112 ;
  assign n33116 = n32915 ^ n17273 ^ 1'b0 ;
  assign n33117 = ( n15656 & n32915 ) | ( n15656 & n33116 ) | ( n32915 & n33116 ) ;
  assign n33118 = x644 & ~n33117 ;
  assign n33123 = ( x715 & n33117 ) | ( x715 & n33118 ) | ( n33117 & n33118 ) ;
  assign n33124 = ~n33115 & n33123 ;
  assign n33125 = ~x715 & n15656 ;
  assign n33126 = ( x1160 & n33124 ) | ( x1160 & ~n33125 ) | ( n33124 & ~n33125 ) ;
  assign n33127 = ~n33124 & n33126 ;
  assign n33114 = x715 & n15656 ;
  assign n33119 = x715 | n33118 ;
  assign n33120 = ( n33112 & n33115 ) | ( n33112 & ~n33119 ) | ( n33115 & ~n33119 ) ;
  assign n33121 = ( x1160 & ~n33114 ) | ( x1160 & n33120 ) | ( ~n33114 & n33120 ) ;
  assign n33122 = n33114 | n33121 ;
  assign n33128 = n33127 ^ n33122 ^ 1'b0 ;
  assign n33129 = ( x790 & ~n33122 ) | ( x790 & n33127 ) | ( ~n33122 & n33127 ) ;
  assign n33130 = ( x790 & ~n33128 ) | ( x790 & n33129 ) | ( ~n33128 & n33129 ) ;
  assign n33131 = ( n7318 & n33113 ) | ( n7318 & ~n33130 ) | ( n33113 & ~n33130 ) ;
  assign n33132 = ~n7318 & n33131 ;
  assign n33133 = x639 & n33132 ;
  assign n33134 = ~n8793 & n15655 ;
  assign n33135 = ~x639 & n33134 ;
  assign n33136 = ( x622 & ~n33133 ) | ( x622 & n33135 ) | ( ~n33133 & n33135 ) ;
  assign n33137 = n33133 | n33136 ;
  assign n33138 = x1157 & ~n33102 ;
  assign n33139 = n19055 & ~n32900 ;
  assign n33140 = n33105 | n33139 ;
  assign n33141 = ( x787 & n33138 ) | ( x787 & n33140 ) | ( n33138 & n33140 ) ;
  assign n33142 = n33140 ^ n33138 ^ 1'b0 ;
  assign n33143 = ( x787 & n33141 ) | ( x787 & n33142 ) | ( n33141 & n33142 ) ;
  assign n33144 = ( n18484 & n32758 ) | ( n18484 & ~n33143 ) | ( n32758 & ~n33143 ) ;
  assign n33145 = ~n33143 & n33144 ;
  assign n33146 = x790 | n33145 ;
  assign n33152 = x644 & ~n33145 ;
  assign n33156 = n33123 & ~n33152 ;
  assign n33147 = n32900 ^ n16376 ^ 1'b0 ;
  assign n33148 = ( n15656 & n32900 ) | ( n15656 & n33147 ) | ( n32900 & n33147 ) ;
  assign n33149 = n15656 ^ x644 ^ 1'b0 ;
  assign n33157 = ( n15656 & n33148 ) | ( n15656 & n33149 ) | ( n33148 & n33149 ) ;
  assign n33158 = ~x715 & n33157 ;
  assign n33159 = ( x1160 & n33156 ) | ( x1160 & ~n33158 ) | ( n33156 & ~n33158 ) ;
  assign n33160 = ~n33156 & n33159 ;
  assign n33150 = ( n15656 & n33148 ) | ( n15656 & ~n33149 ) | ( n33148 & ~n33149 ) ;
  assign n33151 = x715 & n33150 ;
  assign n33153 = ( ~n33119 & n33145 ) | ( ~n33119 & n33152 ) | ( n33145 & n33152 ) ;
  assign n33154 = ( x1160 & ~n33151 ) | ( x1160 & n33153 ) | ( ~n33151 & n33153 ) ;
  assign n33155 = n33151 | n33154 ;
  assign n33161 = n33160 ^ n33155 ^ 1'b0 ;
  assign n33162 = ( x790 & ~n33155 ) | ( x790 & n33160 ) | ( ~n33155 & n33160 ) ;
  assign n33163 = ( x790 & ~n33161 ) | ( x790 & n33162 ) | ( ~n33161 & n33162 ) ;
  assign n33164 = ( n7318 & n33146 ) | ( n7318 & ~n33163 ) | ( n33146 & ~n33163 ) ;
  assign n33165 = ~n7318 & n33164 ;
  assign n33166 = x639 & n33165 ;
  assign n33167 = x790 | n33148 ;
  assign n33168 = ~x1160 & n33150 ;
  assign n33169 = x1160 & n33157 ;
  assign n33170 = ( x790 & n33168 ) | ( x790 & ~n33169 ) | ( n33168 & ~n33169 ) ;
  assign n33171 = ~n33168 & n33170 ;
  assign n33172 = ( n7318 & n33167 ) | ( n7318 & ~n33171 ) | ( n33167 & ~n33171 ) ;
  assign n33173 = ~n7318 & n33172 ;
  assign n33174 = ~x639 & n33173 ;
  assign n33175 = x622 & ~n33174 ;
  assign n33176 = n33137 & ~n33175 ;
  assign n33177 = ( n33137 & n33166 ) | ( n33137 & n33176 ) | ( n33166 & n33176 ) ;
  assign n33178 = ( x209 & ~n33097 ) | ( x209 & n33177 ) | ( ~n33097 & n33177 ) ;
  assign n33179 = ~n33097 & n33178 ;
  assign n33180 = x210 & ~n15644 ;
  assign n33181 = x634 & n19256 ;
  assign n33182 = x633 & x947 ;
  assign n33183 = n33181 | n33182 ;
  assign n33184 = n15644 & n33183 ;
  assign n33185 = ( x38 & n33180 ) | ( x38 & ~n33184 ) | ( n33180 & ~n33184 ) ;
  assign n33186 = ~n33180 & n33185 ;
  assign n33187 = x210 | n15337 ;
  assign n33188 = x210 & ~n15337 ;
  assign n33189 = ( x634 & n33187 ) | ( x634 & n33188 ) | ( n33187 & n33188 ) ;
  assign n33190 = n5083 & ~n33189 ;
  assign n33191 = x907 & ~n33190 ;
  assign n33192 = x210 | n15351 ;
  assign n33193 = n33192 ^ n31252 ^ n15351 ;
  assign n33194 = n5083 | n33193 ;
  assign n33195 = n33191 & n33194 ;
  assign n33196 = n5083 & ~n15336 ;
  assign n33197 = n1611 & n33196 ;
  assign n33198 = ( x210 & n15351 ) | ( x210 & ~n33197 ) | ( n15351 & ~n33197 ) ;
  assign n33199 = ~n15351 & n33198 ;
  assign n33200 = n33195 | n33199 ;
  assign n33201 = ~x947 & n33200 ;
  assign n33202 = ( x633 & n33187 ) | ( x633 & n33188 ) | ( n33187 & n33188 ) ;
  assign n33203 = n5083 & ~n33202 ;
  assign n33204 = x947 & ~n33203 ;
  assign n33205 = ~x633 & n15351 ;
  assign n33206 = n33192 & ~n33205 ;
  assign n33207 = n5083 | n33206 ;
  assign n33208 = n33204 & n33207 ;
  assign n33209 = ( n5114 & n33201 ) | ( n5114 & ~n33208 ) | ( n33201 & ~n33208 ) ;
  assign n33210 = ~n33201 & n33209 ;
  assign n33211 = n5082 | n33202 ;
  assign n33212 = x947 & n33211 ;
  assign n33213 = ~n5075 & n33202 ;
  assign n33214 = n5082 & ~n33213 ;
  assign n33215 = n33212 & ~n33214 ;
  assign n33216 = n5075 & n33206 ;
  assign n33217 = ( n33212 & n33215 ) | ( n33212 & n33216 ) | ( n33215 & n33216 ) ;
  assign n33218 = ~n5099 & n33189 ;
  assign n33219 = x907 & ~n33218 ;
  assign n33220 = n5099 & n33193 ;
  assign n33221 = n33219 & ~n33220 ;
  assign n33222 = x947 | n33221 ;
  assign n33223 = ~n5082 & n33188 ;
  assign n33224 = x210 & n5082 ;
  assign n33225 = ~n15357 & n33224 ;
  assign n33226 = n33223 | n33225 ;
  assign n33227 = ( x907 & ~n33222 ) | ( x907 & n33226 ) | ( ~n33222 & n33226 ) ;
  assign n33228 = ~n33222 & n33227 ;
  assign n33229 = ( n5114 & ~n33217 ) | ( n5114 & n33228 ) | ( ~n33217 & n33228 ) ;
  assign n33230 = n33217 | n33229 ;
  assign n33231 = ( x223 & n33210 ) | ( x223 & n33230 ) | ( n33210 & n33230 ) ;
  assign n33232 = ~n33210 & n33231 ;
  assign n33233 = ( n33183 & n33187 ) | ( n33183 & n33188 ) | ( n33187 & n33188 ) ;
  assign n33234 = n1359 | n33233 ;
  assign n33235 = x210 | n15425 ;
  assign n33236 = ~n31115 & n33235 ;
  assign n33237 = n5083 | n33236 ;
  assign n33238 = n33204 & n33237 ;
  assign n33239 = ~n31225 & n33235 ;
  assign n33240 = n5083 | n33239 ;
  assign n33241 = n33191 & n33240 ;
  assign n33242 = x210 & ~n15433 ;
  assign n33243 = ~x907 & n33242 ;
  assign n33244 = ( ~x947 & n33241 ) | ( ~x947 & n33243 ) | ( n33241 & n33243 ) ;
  assign n33245 = ~x947 & n33244 ;
  assign n33246 = ( n5114 & n33238 ) | ( n5114 & ~n33245 ) | ( n33238 & ~n33245 ) ;
  assign n33247 = ~n33238 & n33246 ;
  assign n33248 = n5099 & n33239 ;
  assign n33249 = n33219 & ~n33248 ;
  assign n33250 = x947 | n33249 ;
  assign n33251 = ~n15445 & n33224 ;
  assign n33252 = n33223 | n33251 ;
  assign n33253 = ( x907 & ~n33250 ) | ( x907 & n33252 ) | ( ~n33250 & n33252 ) ;
  assign n33254 = ~n33250 & n33253 ;
  assign n33255 = n5075 & n33236 ;
  assign n33256 = n33214 & ~n33255 ;
  assign n33257 = ( n5114 & n33212 ) | ( n5114 & ~n33256 ) | ( n33212 & ~n33256 ) ;
  assign n33258 = n33257 ^ n33212 ^ 1'b0 ;
  assign n33259 = ( n5114 & n33257 ) | ( n5114 & ~n33258 ) | ( n33257 & ~n33258 ) ;
  assign n33260 = ( ~n33247 & n33254 ) | ( ~n33247 & n33259 ) | ( n33254 & n33259 ) ;
  assign n33261 = ~n33247 & n33260 ;
  assign n33262 = ( x222 & x224 ) | ( x222 & ~n33261 ) | ( x224 & ~n33261 ) ;
  assign n33263 = ~n33261 & n33262 ;
  assign n33264 = ( x223 & n33234 ) | ( x223 & ~n33263 ) | ( n33234 & ~n33263 ) ;
  assign n33265 = ~x223 & n33264 ;
  assign n33266 = ( x299 & ~n33232 ) | ( x299 & n33265 ) | ( ~n33232 & n33265 ) ;
  assign n33267 = n33232 | n33266 ;
  assign n33268 = n2263 | n33233 ;
  assign n33269 = n5060 | n33252 ;
  assign n33270 = n5060 & ~n33242 ;
  assign n33271 = ( x907 & n33269 ) | ( x907 & ~n33270 ) | ( n33269 & ~n33270 ) ;
  assign n33272 = ~x907 & n33271 ;
  assign n33273 = ( ~x947 & n33241 ) | ( ~x947 & n33272 ) | ( n33241 & n33272 ) ;
  assign n33274 = ~x947 & n33273 ;
  assign n33275 = ( n2263 & n33238 ) | ( n2263 & ~n33274 ) | ( n33238 & ~n33274 ) ;
  assign n33276 = ~n33238 & n33275 ;
  assign n33277 = ( x215 & n33268 ) | ( x215 & ~n33276 ) | ( n33268 & ~n33276 ) ;
  assign n33278 = ~x215 & n33277 ;
  assign n33279 = n5060 | n33226 ;
  assign n33280 = n5060 & ~n33199 ;
  assign n33281 = ( x907 & n33279 ) | ( x907 & ~n33280 ) | ( n33279 & ~n33280 ) ;
  assign n33282 = ~x907 & n33281 ;
  assign n33283 = ( ~x947 & n33195 ) | ( ~x947 & n33282 ) | ( n33195 & n33282 ) ;
  assign n33284 = ~x947 & n33283 ;
  assign n33285 = ( x215 & n33208 ) | ( x215 & n33284 ) | ( n33208 & n33284 ) ;
  assign n33286 = n33284 ^ n33208 ^ 1'b0 ;
  assign n33287 = ( x215 & n33285 ) | ( x215 & n33286 ) | ( n33285 & n33286 ) ;
  assign n33288 = ( x299 & n33278 ) | ( x299 & ~n33287 ) | ( n33278 & ~n33287 ) ;
  assign n33289 = ~n33278 & n33288 ;
  assign n33290 = x39 & ~n33289 ;
  assign n33291 = n33267 & n33290 ;
  assign n33292 = n15327 & n33183 ;
  assign n33293 = x210 & ~n15327 ;
  assign n33294 = ( x299 & ~n33292 ) | ( x299 & n33293 ) | ( ~n33292 & n33293 ) ;
  assign n33295 = n33292 | n33294 ;
  assign n33296 = n15329 & n33183 ;
  assign n33297 = ( x299 & n15328 ) | ( x299 & ~n33296 ) | ( n15328 & ~n33296 ) ;
  assign n33298 = ~n15328 & n33297 ;
  assign n33299 = x39 | n33298 ;
  assign n33300 = ( x38 & n33295 ) | ( x38 & ~n33299 ) | ( n33295 & ~n33299 ) ;
  assign n33301 = n33300 ^ n33295 ^ 1'b0 ;
  assign n33302 = ( x38 & n33300 ) | ( x38 & ~n33301 ) | ( n33300 & ~n33301 ) ;
  assign n33303 = ( ~n33186 & n33291 ) | ( ~n33186 & n33302 ) | ( n33291 & n33302 ) ;
  assign n33304 = ~n33186 & n33303 ;
  assign n33305 = n33304 ^ n8793 ^ 1'b0 ;
  assign n33306 = ( x210 & n33304 ) | ( x210 & n33305 ) | ( n33304 & n33305 ) ;
  assign n33307 = ~n2069 & n20002 ;
  assign n33308 = x606 & ~n33307 ;
  assign n33309 = ~n2069 & n19999 ;
  assign n33310 = x606 | n33309 ;
  assign n33311 = ( x643 & n33308 ) | ( x643 & n33310 ) | ( n33308 & n33310 ) ;
  assign n33312 = ~n33308 & n33311 ;
  assign n33313 = ~n2069 & n19440 ;
  assign n33314 = n33313 ^ n33312 ^ 1'b0 ;
  assign n33315 = x606 & ~x643 ;
  assign n33316 = ( n33313 & ~n33314 ) | ( n33313 & n33315 ) | ( ~n33314 & n33315 ) ;
  assign n33317 = ( n33312 & n33314 ) | ( n33312 & n33316 ) | ( n33314 & n33316 ) ;
  assign n33318 = ( x211 & ~n7318 ) | ( x211 & n33317 ) | ( ~n7318 & n33317 ) ;
  assign n33319 = ~x211 & n33318 ;
  assign n33320 = ~n2069 & n20011 ;
  assign n33321 = ~x606 & n33320 ;
  assign n33322 = ~n2069 & n20014 ;
  assign n33323 = x606 & n33322 ;
  assign n33324 = ( x643 & n33321 ) | ( x643 & ~n33323 ) | ( n33321 & ~n33323 ) ;
  assign n33325 = ~n33321 & n33324 ;
  assign n33326 = ~n2069 & n19459 ;
  assign n33327 = x606 & n33326 ;
  assign n33328 = ~x606 & n15656 ;
  assign n33329 = ( x643 & ~n33327 ) | ( x643 & n33328 ) | ( ~n33327 & n33328 ) ;
  assign n33330 = n33327 | n33329 ;
  assign n33331 = ( n7318 & ~n33325 ) | ( n7318 & n33330 ) | ( ~n33325 & n33330 ) ;
  assign n33332 = ~n7318 & n33331 ;
  assign n33333 = ~n33319 & n33332 ;
  assign n33334 = ( x211 & n33319 ) | ( x211 & ~n33333 ) | ( n33319 & ~n33333 ) ;
  assign n33335 = ~x607 & n33320 ;
  assign n33336 = x607 & n33322 ;
  assign n33337 = ( x638 & n33335 ) | ( x638 & ~n33336 ) | ( n33335 & ~n33336 ) ;
  assign n33338 = ~n33335 & n33337 ;
  assign n33339 = ~x607 & n15656 ;
  assign n33340 = x638 | n33339 ;
  assign n33341 = x607 & n33326 ;
  assign n33342 = ( ~n7318 & n33340 ) | ( ~n7318 & n33341 ) | ( n33340 & n33341 ) ;
  assign n33343 = ~n7318 & n33342 ;
  assign n33344 = n33343 ^ n33338 ^ 1'b0 ;
  assign n33345 = ( n33338 & n33343 ) | ( n33338 & n33344 ) | ( n33343 & n33344 ) ;
  assign n33346 = ( x212 & ~n33338 ) | ( x212 & n33345 ) | ( ~n33338 & n33345 ) ;
  assign n33347 = x212 & ~n7318 ;
  assign n33348 = x607 & ~n33307 ;
  assign n33349 = x638 & ~n33348 ;
  assign n33350 = x607 | n33309 ;
  assign n33351 = n33349 & n33350 ;
  assign n33352 = n33351 ^ n33313 ^ 1'b0 ;
  assign n33353 = x607 & ~x638 ;
  assign n33354 = ( n33313 & ~n33352 ) | ( n33313 & n33353 ) | ( ~n33352 & n33353 ) ;
  assign n33355 = ( n33351 & n33352 ) | ( n33351 & n33354 ) | ( n33352 & n33354 ) ;
  assign n33356 = n33346 & ~n33355 ;
  assign n33357 = ( n33346 & ~n33347 ) | ( n33346 & n33356 ) | ( ~n33347 & n33356 ) ;
  assign n33358 = x213 & ~n7318 ;
  assign n33359 = x622 & ~n33307 ;
  assign n33360 = x639 & ~n33359 ;
  assign n33361 = x622 | n33309 ;
  assign n33362 = n33360 & n33361 ;
  assign n33363 = n33362 ^ n33313 ^ 1'b0 ;
  assign n33364 = x622 & ~x639 ;
  assign n33365 = ( n33313 & ~n33363 ) | ( n33313 & n33364 ) | ( ~n33363 & n33364 ) ;
  assign n33366 = ( n33362 & n33363 ) | ( n33362 & n33365 ) | ( n33363 & n33365 ) ;
  assign n33367 = n33358 & n33366 ;
  assign n33368 = x639 & n33320 ;
  assign n33369 = ~x639 & n15656 ;
  assign n33370 = ( x622 & ~n33368 ) | ( x622 & n33369 ) | ( ~n33368 & n33369 ) ;
  assign n33371 = n33368 | n33370 ;
  assign n33372 = x639 & n33322 ;
  assign n33373 = ~x639 & n33326 ;
  assign n33374 = ( x622 & n33372 ) | ( x622 & ~n33373 ) | ( n33372 & ~n33373 ) ;
  assign n33375 = ~n33372 & n33374 ;
  assign n33376 = ( n7318 & n33371 ) | ( n7318 & ~n33375 ) | ( n33371 & ~n33375 ) ;
  assign n33377 = ~n7318 & n33376 ;
  assign n33378 = x213 | n33377 ;
  assign n33379 = ~n33367 & n33378 ;
  assign n33380 = ~x623 & n33320 ;
  assign n33381 = x623 & n33322 ;
  assign n33382 = ( x710 & n33380 ) | ( x710 & ~n33381 ) | ( n33380 & ~n33381 ) ;
  assign n33383 = ~n33380 & n33382 ;
  assign n33384 = ~x623 & n15656 ;
  assign n33385 = x710 | n33384 ;
  assign n33386 = x623 & n33326 ;
  assign n33387 = ( ~n7318 & n33385 ) | ( ~n7318 & n33386 ) | ( n33385 & n33386 ) ;
  assign n33388 = ~n7318 & n33387 ;
  assign n33389 = n33388 ^ n33383 ^ 1'b0 ;
  assign n33390 = ( n33383 & n33388 ) | ( n33383 & n33389 ) | ( n33388 & n33389 ) ;
  assign n33391 = ( x214 & ~n33383 ) | ( x214 & n33390 ) | ( ~n33383 & n33390 ) ;
  assign n33392 = x214 & ~n7318 ;
  assign n33393 = x623 & ~n33307 ;
  assign n33394 = x710 & ~n33393 ;
  assign n33395 = x623 | n33309 ;
  assign n33396 = n33394 & n33395 ;
  assign n33397 = n33396 ^ n33313 ^ 1'b0 ;
  assign n33398 = x623 & ~x710 ;
  assign n33399 = ( n33313 & ~n33397 ) | ( n33313 & n33398 ) | ( ~n33397 & n33398 ) ;
  assign n33400 = ( n33396 & n33397 ) | ( n33396 & n33399 ) | ( n33397 & n33399 ) ;
  assign n33401 = n33391 & ~n33400 ;
  assign n33402 = ( n33391 & ~n33392 ) | ( n33391 & n33401 ) | ( ~n33392 & n33401 ) ;
  assign n33418 = x681 & x907 ;
  assign n33423 = x947 | n33418 ;
  assign n33430 = n15364 & ~n15382 ;
  assign n33431 = x642 | n33430 ;
  assign n33432 = n5078 | n15361 ;
  assign n33433 = ~n33431 & n33432 ;
  assign n33449 = x947 & n33433 ;
  assign n33450 = n33423 & ~n33449 ;
  assign n33451 = x947 | n19673 ;
  assign n33452 = x299 & ~n33451 ;
  assign n33453 = ( x299 & n33450 ) | ( x299 & n33452 ) | ( n33450 & n33452 ) ;
  assign n33403 = ~x642 & n15445 ;
  assign n33404 = n5078 & ~n33403 ;
  assign n33405 = n15446 & ~n15527 ;
  assign n33406 = n5080 & n15337 ;
  assign n33407 = ~x642 & n33406 ;
  assign n33408 = ( n5078 & ~n33405 ) | ( n5078 & n33407 ) | ( ~n33405 & n33407 ) ;
  assign n33409 = n33405 | n33408 ;
  assign n33410 = n33409 ^ n33404 ^ 1'b0 ;
  assign n33411 = ( n33404 & n33409 ) | ( n33404 & n33410 ) | ( n33409 & n33410 ) ;
  assign n33412 = ( n5114 & ~n33404 ) | ( n5114 & n33411 ) | ( ~n33404 & n33411 ) ;
  assign n33413 = ~x642 & n15433 ;
  assign n33414 = n5114 & ~n33413 ;
  assign n33415 = x947 & ~n33414 ;
  assign n33416 = n1359 & ~n33415 ;
  assign n33417 = ( n1359 & ~n33412 ) | ( n1359 & n33416 ) | ( ~n33412 & n33416 ) ;
  assign n33419 = n33418 ^ n33417 ^ 1'b0 ;
  assign n33420 = ( ~n19765 & n33418 ) | ( ~n19765 & n33419 ) | ( n33418 & n33419 ) ;
  assign n33421 = ( n33417 & ~n33419 ) | ( n33417 & n33420 ) | ( ~n33419 & n33420 ) ;
  assign n33422 = n1359 | n15337 ;
  assign n33424 = ~x947 & n33418 ;
  assign n33425 = ( x642 & n33423 ) | ( x642 & n33424 ) | ( n33423 & n33424 ) ;
  assign n33426 = ~n1359 & n33425 ;
  assign n33427 = x223 | n33426 ;
  assign n33428 = ( n33421 & n33422 ) | ( n33421 & ~n33427 ) | ( n33422 & ~n33427 ) ;
  assign n33429 = ~n33421 & n33428 ;
  assign n33434 = n5114 & ~n33433 ;
  assign n33435 = x947 & ~n33434 ;
  assign n33436 = n33435 ^ n19361 ^ 1'b0 ;
  assign n33437 = n5078 & ~n15357 ;
  assign n33438 = x642 | n33437 ;
  assign n33439 = n5078 | n15371 ;
  assign n33440 = n33439 ^ n33438 ^ 1'b0 ;
  assign n33441 = ( n33438 & n33439 ) | ( n33438 & n33440 ) | ( n33439 & n33440 ) ;
  assign n33442 = ( n5114 & ~n33438 ) | ( n5114 & n33441 ) | ( ~n33438 & n33441 ) ;
  assign n33443 = ( n33435 & ~n33436 ) | ( n33435 & n33442 ) | ( ~n33436 & n33442 ) ;
  assign n33444 = ( n19361 & n33436 ) | ( n19361 & n33443 ) | ( n33436 & n33443 ) ;
  assign n33445 = ( x223 & n33424 ) | ( x223 & n33444 ) | ( n33424 & n33444 ) ;
  assign n33446 = ~n33424 & n33445 ;
  assign n33447 = ( x299 & ~n33429 ) | ( x299 & n33446 ) | ( ~n33429 & n33446 ) ;
  assign n33448 = n33429 | n33447 ;
  assign n33454 = n33453 ^ n33448 ^ 1'b0 ;
  assign n33455 = ( x215 & ~n33448 ) | ( x215 & n33453 ) | ( ~n33448 & n33453 ) ;
  assign n33456 = ( x215 & ~n33454 ) | ( x215 & n33455 ) | ( ~n33454 & n33455 ) ;
  assign n33457 = x642 & ~n15383 ;
  assign n33458 = n15432 & n33457 ;
  assign n33459 = x642 & n15383 ;
  assign n33460 = n15427 & n33459 ;
  assign n33461 = x947 & ~n33460 ;
  assign n33462 = ~n33458 & n33461 ;
  assign n33463 = n15429 & n33418 ;
  assign n33464 = ( x947 & ~n33462 ) | ( x947 & n33463 ) | ( ~n33462 & n33463 ) ;
  assign n33465 = ~n33462 & n33464 ;
  assign n33466 = n5114 & ~n33465 ;
  assign n33467 = n5114 ^ x947 ^ 1'b0 ;
  assign n33468 = n15337 & n33459 ;
  assign n33469 = n15394 & n33457 ;
  assign n33470 = ~n15454 & n33469 ;
  assign n33471 = n33468 | n33470 ;
  assign n33472 = ( x947 & ~n33467 ) | ( x947 & n33471 ) | ( ~n33467 & n33471 ) ;
  assign n33473 = ( n5114 & n33467 ) | ( n5114 & n33472 ) | ( n33467 & n33472 ) ;
  assign n33474 = n33473 ^ n15466 ^ 1'b0 ;
  assign n33475 = ( ~n15466 & n33424 ) | ( ~n15466 & n33474 ) | ( n33424 & n33474 ) ;
  assign n33476 = ( n15466 & n33473 ) | ( n15466 & n33475 ) | ( n33473 & n33475 ) ;
  assign n33477 = ( n1359 & n33466 ) | ( n1359 & n33476 ) | ( n33466 & n33476 ) ;
  assign n33478 = ~n33466 & n33477 ;
  assign n33479 = n15337 & n33426 ;
  assign n33480 = ( x223 & ~n33478 ) | ( x223 & n33479 ) | ( ~n33478 & n33479 ) ;
  assign n33481 = n33478 | n33480 ;
  assign n33482 = ~n15381 & n33469 ;
  assign n33483 = x947 & ~n33468 ;
  assign n33484 = ~n33482 & n33483 ;
  assign n33485 = ( x947 & n15353 ) | ( x947 & n15361 ) | ( n15353 & n15361 ) ;
  assign n33486 = ~n33484 & n33485 ;
  assign n33487 = ( n5114 & n33484 ) | ( n5114 & ~n33486 ) | ( n33484 & ~n33486 ) ;
  assign n33488 = n5114 | n15371 ;
  assign n33489 = ( x947 & n33423 ) | ( x947 & n33488 ) | ( n33423 & n33488 ) ;
  assign n33490 = x223 & ~n33489 ;
  assign n33491 = ( x223 & n33487 ) | ( x223 & n33490 ) | ( n33487 & n33490 ) ;
  assign n33492 = ( x299 & n33481 ) | ( x299 & ~n33491 ) | ( n33481 & ~n33491 ) ;
  assign n33493 = n33492 ^ n33481 ^ 1'b0 ;
  assign n33494 = ( x299 & n33492 ) | ( x299 & ~n33493 ) | ( n33492 & ~n33493 ) ;
  assign n33495 = n15436 & n33425 ;
  assign n33496 = n2263 & n33465 ;
  assign n33497 = ( x299 & n33495 ) | ( x299 & ~n33496 ) | ( n33495 & ~n33496 ) ;
  assign n33498 = ~n33495 & n33497 ;
  assign n33499 = ( x215 & n33494 ) | ( x215 & ~n33498 ) | ( n33494 & ~n33498 ) ;
  assign n33500 = ~x215 & n33499 ;
  assign n33501 = ( x39 & n33456 ) | ( x39 & n33500 ) | ( n33456 & n33500 ) ;
  assign n33502 = n33500 ^ n33456 ^ 1'b0 ;
  assign n33503 = ( x39 & n33501 ) | ( x39 & n33502 ) | ( n33501 & n33502 ) ;
  assign n33504 = n15327 & n33425 ;
  assign n33505 = x299 | n33504 ;
  assign n33506 = n15327 & ~n33505 ;
  assign n33507 = ( x215 & n33505 ) | ( x215 & ~n33506 ) | ( n33505 & ~n33506 ) ;
  assign n33508 = n15330 & n33425 ;
  assign n33509 = x215 & ~n15330 ;
  assign n33510 = ( x299 & n33508 ) | ( x299 & ~n33509 ) | ( n33508 & ~n33509 ) ;
  assign n33511 = ~n33508 & n33510 ;
  assign n33512 = ( x39 & n33507 ) | ( x39 & ~n33511 ) | ( n33507 & ~n33511 ) ;
  assign n33513 = ~x39 & n33512 ;
  assign n33514 = ( x38 & ~n33503 ) | ( x38 & n33513 ) | ( ~n33503 & n33513 ) ;
  assign n33515 = n33503 | n33514 ;
  assign n33516 = x215 & ~n15644 ;
  assign n33517 = n15644 & n33425 ;
  assign n33518 = ( x38 & n33516 ) | ( x38 & ~n33517 ) | ( n33516 & ~n33517 ) ;
  assign n33519 = ~n33516 & n33518 ;
  assign n33520 = ( n8793 & n33515 ) | ( n8793 & ~n33519 ) | ( n33515 & ~n33519 ) ;
  assign n33521 = ~n8793 & n33520 ;
  assign n33522 = n33521 ^ x215 ^ 1'b0 ;
  assign n33523 = ( ~x215 & n8793 ) | ( ~x215 & n33522 ) | ( n8793 & n33522 ) ;
  assign n33524 = ( x215 & n33521 ) | ( x215 & n33523 ) | ( n33521 & n33523 ) ;
  assign n33525 = x662 & x907 ;
  assign n33526 = ~x947 & n33525 ;
  assign n33527 = x614 & x947 ;
  assign n33528 = n33526 | n33527 ;
  assign n33529 = n15644 & n33528 ;
  assign n33530 = x216 & ~n15644 ;
  assign n33531 = ( x38 & n33529 ) | ( x38 & ~n33530 ) | ( n33529 & ~n33530 ) ;
  assign n33532 = ~n33529 & n33531 ;
  assign n33533 = n15327 & n33528 ;
  assign n33534 = x299 | n33533 ;
  assign n33535 = n15327 & ~n33534 ;
  assign n33536 = ( x216 & n33534 ) | ( x216 & ~n33535 ) | ( n33534 & ~n33535 ) ;
  assign n33537 = n15330 & n33528 ;
  assign n33538 = x216 & ~n15330 ;
  assign n33539 = x299 & ~n33538 ;
  assign n33540 = n33539 ^ n33537 ^ 1'b0 ;
  assign n33541 = ( n33537 & n33539 ) | ( n33537 & n33540 ) | ( n33539 & n33540 ) ;
  assign n33542 = ( x39 & ~n33537 ) | ( x39 & n33541 ) | ( ~n33537 & n33541 ) ;
  assign n33543 = ( x38 & n33536 ) | ( x38 & ~n33542 ) | ( n33536 & ~n33542 ) ;
  assign n33544 = n33543 ^ n33536 ^ 1'b0 ;
  assign n33545 = ( x38 & n33543 ) | ( x38 & ~n33544 ) | ( n33543 & ~n33544 ) ;
  assign n33546 = n15432 & n33527 ;
  assign n33547 = n15429 & n33526 ;
  assign n33548 = n33546 | n33547 ;
  assign n33549 = n5114 & ~n33548 ;
  assign n33550 = n15466 & n33526 ;
  assign n33551 = x947 & n15460 ;
  assign n33552 = ( n5114 & ~n33550 ) | ( n5114 & n33551 ) | ( ~n33550 & n33551 ) ;
  assign n33553 = n33550 | n33552 ;
  assign n33554 = ( n1359 & n33549 ) | ( n1359 & n33553 ) | ( n33549 & n33553 ) ;
  assign n33555 = ~n33549 & n33554 ;
  assign n33556 = ~n1359 & n33528 ;
  assign n33557 = n15337 & n33556 ;
  assign n33558 = ( x223 & ~n33555 ) | ( x223 & n33557 ) | ( ~n33555 & n33557 ) ;
  assign n33559 = n33555 | n33558 ;
  assign n33560 = n5114 & ~n33485 ;
  assign n33561 = ~n15381 & n15456 ;
  assign n33562 = x947 & ~n15459 ;
  assign n33563 = ~n33561 & n33562 ;
  assign n33564 = n33560 | n33563 ;
  assign n33565 = n33488 & n33525 ;
  assign n33566 = x947 | n33565 ;
  assign n33567 = x223 & ~n33566 ;
  assign n33568 = ( x223 & n33564 ) | ( x223 & n33567 ) | ( n33564 & n33567 ) ;
  assign n33569 = ( x216 & n33559 ) | ( x216 & ~n33568 ) | ( n33559 & ~n33568 ) ;
  assign n33570 = ~x216 & n33569 ;
  assign n33571 = ~x616 & n15358 ;
  assign n33572 = n5078 | n15392 ;
  assign n33573 = n33571 | n33572 ;
  assign n33574 = x614 | n33437 ;
  assign n33575 = ( n5114 & n33573 ) | ( n5114 & ~n33574 ) | ( n33573 & ~n33574 ) ;
  assign n33576 = n33575 ^ n33573 ^ 1'b0 ;
  assign n33577 = ( n5114 & n33575 ) | ( n5114 & ~n33576 ) | ( n33575 & ~n33576 ) ;
  assign n33578 = n33577 ^ n19361 ^ 1'b0 ;
  assign n33579 = n5078 & n15368 ;
  assign n33580 = n15762 | n31022 ;
  assign n33581 = n31024 | n33580 ;
  assign n33582 = ~n15441 & n33581 ;
  assign n33583 = n33579 | n33582 ;
  assign n33584 = n5114 & ~n33583 ;
  assign n33585 = x947 & ~n33584 ;
  assign n33586 = ( n33577 & ~n33578 ) | ( n33577 & n33585 ) | ( ~n33578 & n33585 ) ;
  assign n33587 = ( n19361 & n33578 ) | ( n19361 & n33586 ) | ( n33578 & n33586 ) ;
  assign n33588 = x223 & ~n33526 ;
  assign n33589 = n33587 & n33588 ;
  assign n33590 = x947 | n15433 ;
  assign n33591 = ~x614 & n15433 ;
  assign n33592 = x947 & ~n33591 ;
  assign n33593 = n5114 & ~n33526 ;
  assign n33594 = ~n33592 & n33593 ;
  assign n33595 = n33590 & n33594 ;
  assign n33596 = ~x947 & n15468 ;
  assign n33597 = ~n33525 & n33596 ;
  assign n33598 = x947 & n15453 ;
  assign n33599 = ( ~n5114 & n33597 ) | ( ~n5114 & n33598 ) | ( n33597 & n33598 ) ;
  assign n33600 = ~n5114 & n33599 ;
  assign n33601 = ( n1359 & n33595 ) | ( n1359 & ~n33600 ) | ( n33595 & ~n33600 ) ;
  assign n33602 = ~n33595 & n33601 ;
  assign n33603 = x223 | n33556 ;
  assign n33604 = ( n33422 & n33602 ) | ( n33422 & ~n33603 ) | ( n33602 & ~n33603 ) ;
  assign n33605 = ~n33602 & n33604 ;
  assign n33606 = ( x216 & n33589 ) | ( x216 & ~n33605 ) | ( n33589 & ~n33605 ) ;
  assign n33607 = ~n33589 & n33606 ;
  assign n33608 = ( x299 & ~n33570 ) | ( x299 & n33607 ) | ( ~n33570 & n33607 ) ;
  assign n33609 = n33570 | n33608 ;
  assign n33610 = n15361 & n33525 ;
  assign n33611 = x947 | n33610 ;
  assign n33612 = x947 & ~n15353 ;
  assign n33613 = n33563 | n33612 ;
  assign n33614 = ( x216 & n33611 ) | ( x216 & ~n33613 ) | ( n33611 & ~n33613 ) ;
  assign n33615 = n33614 ^ n33611 ^ 1'b0 ;
  assign n33616 = ( x216 & n33614 ) | ( x216 & ~n33615 ) | ( n33614 & ~n33615 ) ;
  assign n33617 = x947 & ~n33583 ;
  assign n33618 = x216 & ~n33526 ;
  assign n33619 = ( n33451 & n33617 ) | ( n33451 & n33618 ) | ( n33617 & n33618 ) ;
  assign n33620 = ~n33617 & n33619 ;
  assign n33621 = x215 & ~n33620 ;
  assign n33622 = n33616 & n33621 ;
  assign n33623 = n4652 & n33548 ;
  assign n33624 = n15436 & n33528 ;
  assign n33625 = n33623 | n33624 ;
  assign n33626 = n33526 | n33592 ;
  assign n33627 = x947 | n19447 ;
  assign n33628 = x216 & ~n33627 ;
  assign n33629 = ( x216 & n33626 ) | ( x216 & n33628 ) | ( n33626 & n33628 ) ;
  assign n33630 = ( ~x215 & n33625 ) | ( ~x215 & n33629 ) | ( n33625 & n33629 ) ;
  assign n33631 = ~x215 & n33630 ;
  assign n33632 = ( x299 & n33622 ) | ( x299 & ~n33631 ) | ( n33622 & ~n33631 ) ;
  assign n33633 = ~n33622 & n33632 ;
  assign n33634 = x39 & ~n33633 ;
  assign n33635 = n33609 & n33634 ;
  assign n33636 = ( ~n33532 & n33545 ) | ( ~n33532 & n33635 ) | ( n33545 & n33635 ) ;
  assign n33637 = ~n33532 & n33636 ;
  assign n33638 = n33637 ^ n8793 ^ 1'b0 ;
  assign n33639 = ( x216 & n33637 ) | ( x216 & n33638 ) | ( n33637 & n33638 ) ;
  assign n33640 = x695 & ~n33173 ;
  assign n33641 = x217 | n33640 ;
  assign n33642 = ( x695 & n33165 ) | ( x695 & ~n33641 ) | ( n33165 & ~n33641 ) ;
  assign n33643 = ~n33641 & n33642 ;
  assign n33644 = x695 & n33077 ;
  assign n33645 = ~x695 & n33071 ;
  assign n33646 = ( x217 & n33644 ) | ( x217 & ~n33645 ) | ( n33644 & ~n33645 ) ;
  assign n33647 = ~n33644 & n33646 ;
  assign n33648 = ( x612 & n33643 ) | ( x612 & ~n33647 ) | ( n33643 & ~n33647 ) ;
  assign n33649 = ~n33643 & n33648 ;
  assign n33650 = x695 & ~n33134 ;
  assign n33651 = x217 | n33650 ;
  assign n33652 = ( x695 & n33132 ) | ( x695 & ~n33651 ) | ( n33132 & ~n33651 ) ;
  assign n33653 = ~n33651 & n33652 ;
  assign n33654 = ~x695 & n33094 ;
  assign n33655 = x217 & ~n33654 ;
  assign n33656 = x612 | n33655 ;
  assign n33657 = ( ~n33649 & n33653 ) | ( ~n33649 & n33656 ) | ( n33653 & n33656 ) ;
  assign n33658 = ~n33649 & n33657 ;
  assign n33659 = n32407 ^ n32369 ^ 1'b0 ;
  assign n33660 = ( n32407 & n32473 ) | ( n32407 & ~n33659 ) | ( n32473 & ~n33659 ) ;
  assign n33661 = ~n32369 & n32479 ;
  assign n33662 = n33660 ^ x218 ^ 1'b0 ;
  assign n33663 = ( n33660 & ~n33661 ) | ( n33660 & n33662 ) | ( ~n33661 & n33662 ) ;
  assign n33664 = x617 & ~n33307 ;
  assign n33665 = x637 & ~n33664 ;
  assign n33666 = x617 | n33309 ;
  assign n33667 = n33665 & n33666 ;
  assign n33668 = n33667 ^ n33313 ^ 1'b0 ;
  assign n33669 = x617 & ~x637 ;
  assign n33670 = ( n33313 & ~n33668 ) | ( n33313 & n33669 ) | ( ~n33668 & n33669 ) ;
  assign n33671 = ( n33667 & n33668 ) | ( n33667 & n33670 ) | ( n33668 & n33670 ) ;
  assign n33672 = ( x219 & ~n7318 ) | ( x219 & n33671 ) | ( ~n7318 & n33671 ) ;
  assign n33673 = ~x219 & n33672 ;
  assign n33674 = ~x617 & n33320 ;
  assign n33675 = x617 & n33322 ;
  assign n33676 = ( x637 & n33674 ) | ( x637 & ~n33675 ) | ( n33674 & ~n33675 ) ;
  assign n33677 = ~n33674 & n33676 ;
  assign n33678 = x617 & n33326 ;
  assign n33679 = ~x617 & n15656 ;
  assign n33680 = ( x637 & ~n33678 ) | ( x637 & n33679 ) | ( ~n33678 & n33679 ) ;
  assign n33681 = n33678 | n33680 ;
  assign n33682 = ( n7318 & ~n33677 ) | ( n7318 & n33681 ) | ( ~n33677 & n33681 ) ;
  assign n33683 = ~n7318 & n33682 ;
  assign n33684 = ( x219 & n33673 ) | ( x219 & ~n33683 ) | ( n33673 & ~n33683 ) ;
  assign n33685 = n33683 ^ n33673 ^ 1'b0 ;
  assign n33686 = ( n33673 & n33684 ) | ( n33673 & ~n33685 ) | ( n33684 & ~n33685 ) ;
  assign n33687 = n32488 ^ n32350 ^ 1'b0 ;
  assign n33688 = ( n32209 & n32350 ) | ( n32209 & ~n33687 ) | ( n32350 & ~n33687 ) ;
  assign n33689 = n32359 & n32488 ;
  assign n33690 = n33688 ^ x220 ^ 1'b0 ;
  assign n33691 = ( n33688 & ~n33689 ) | ( n33688 & n33690 ) | ( ~n33689 & n33690 ) ;
  assign n33692 = x661 & x907 ;
  assign n33693 = ~x947 & n33692 ;
  assign n33694 = x616 & x947 ;
  assign n33695 = n33693 | n33694 ;
  assign n33696 = n15644 & n33695 ;
  assign n33697 = x221 & ~n15644 ;
  assign n33698 = ( x38 & n33696 ) | ( x38 & ~n33697 ) | ( n33696 & ~n33697 ) ;
  assign n33699 = ~n33696 & n33698 ;
  assign n33700 = n15432 & n33694 ;
  assign n33701 = n15429 & n33693 ;
  assign n33702 = n33700 | n33701 ;
  assign n33703 = x216 & n33702 ;
  assign n33704 = n15337 & n33695 ;
  assign n33705 = ~x216 & n33704 ;
  assign n33706 = ( x221 & ~n33703 ) | ( x221 & n33705 ) | ( ~n33703 & n33705 ) ;
  assign n33707 = n33703 | n33706 ;
  assign n33708 = n15464 ^ n15427 ^ n15337 ;
  assign n33709 = n15388 & n33708 ;
  assign n33710 = ( ~n15384 & n33413 ) | ( ~n15384 & n33458 ) | ( n33413 & n33458 ) ;
  assign n33711 = ( x947 & n33709 ) | ( x947 & ~n33710 ) | ( n33709 & ~n33710 ) ;
  assign n33712 = ~n33709 & n33711 ;
  assign n33713 = n19447 & ~n33692 ;
  assign n33714 = x947 | n33713 ;
  assign n33715 = ( x221 & n33712 ) | ( x221 & n33714 ) | ( n33712 & n33714 ) ;
  assign n33716 = ~n33712 & n33715 ;
  assign n33717 = ( x215 & n33707 ) | ( x215 & ~n33716 ) | ( n33707 & ~n33716 ) ;
  assign n33718 = ~x215 & n33717 ;
  assign n33719 = x947 & n15398 ;
  assign n33720 = n33693 | n33719 ;
  assign n33721 = n33485 & n33720 ;
  assign n33722 = x221 | n33721 ;
  assign n33723 = x221 & ~n33693 ;
  assign n33724 = x616 | n33430 ;
  assign n33725 = n5078 | n15360 ;
  assign n33726 = x947 & ~n33725 ;
  assign n33727 = ( x947 & n33724 ) | ( x947 & n33726 ) | ( n33724 & n33726 ) ;
  assign n33728 = n33451 & ~n33727 ;
  assign n33729 = n33723 & n33728 ;
  assign n33730 = x215 & ~n33729 ;
  assign n33731 = n33722 & n33730 ;
  assign n33732 = ( x299 & n33718 ) | ( x299 & ~n33731 ) | ( n33718 & ~n33731 ) ;
  assign n33733 = ~n33718 & n33732 ;
  assign n33734 = ~n33560 & n33720 ;
  assign n33735 = n33488 | n33719 ;
  assign n33736 = n33734 & n33735 ;
  assign n33737 = ( x221 & x223 ) | ( x221 & ~n33736 ) | ( x223 & ~n33736 ) ;
  assign n33738 = n33737 ^ x223 ^ 1'b0 ;
  assign n33739 = ( x221 & n33737 ) | ( x221 & ~n33738 ) | ( n33737 & ~n33738 ) ;
  assign n33740 = n5114 & ~n33702 ;
  assign n33741 = n15396 & ~n15454 ;
  assign n33742 = n15393 | n33741 ;
  assign n33743 = ( x947 & ~n33467 ) | ( x947 & n33742 ) | ( ~n33467 & n33742 ) ;
  assign n33744 = ( n5114 & n33467 ) | ( n5114 & n33743 ) | ( n33467 & n33743 ) ;
  assign n33745 = n33744 ^ n15466 ^ 1'b0 ;
  assign n33746 = ( ~n15466 & n33693 ) | ( ~n15466 & n33745 ) | ( n33693 & n33745 ) ;
  assign n33747 = ( n15466 & n33744 ) | ( n15466 & n33746 ) | ( n33744 & n33746 ) ;
  assign n33748 = ( n1359 & n33740 ) | ( n1359 & n33747 ) | ( n33740 & n33747 ) ;
  assign n33749 = ~n33740 & n33748 ;
  assign n33750 = ( x223 & n15479 ) | ( x223 & n33695 ) | ( n15479 & n33695 ) ;
  assign n33751 = ( ~n33739 & n33749 ) | ( ~n33739 & n33750 ) | ( n33749 & n33750 ) ;
  assign n33752 = ~n33739 & n33751 ;
  assign n33753 = x947 | n15378 ;
  assign n33754 = ~n33727 & n33753 ;
  assign n33755 = n5114 & ~n33754 ;
  assign n33756 = x223 & ~n33693 ;
  assign n33757 = x947 & n15391 ;
  assign n33758 = ~x947 & n15402 ;
  assign n33759 = ( n5114 & ~n33757 ) | ( n5114 & n33758 ) | ( ~n33757 & n33758 ) ;
  assign n33760 = n33757 | n33759 ;
  assign n33761 = ( n33755 & n33756 ) | ( n33755 & n33760 ) | ( n33756 & n33760 ) ;
  assign n33762 = ~n33755 & n33761 ;
  assign n33763 = n33590 & ~n33712 ;
  assign n33764 = n5114 & ~n33763 ;
  assign n33765 = n33693 | n33764 ;
  assign n33766 = n15453 | n15457 ;
  assign n33767 = ~n15384 & n33766 ;
  assign n33768 = n15388 & n15464 ;
  assign n33769 = ( x947 & n33767 ) | ( x947 & n33768 ) | ( n33767 & n33768 ) ;
  assign n33770 = n33768 ^ n33767 ^ 1'b0 ;
  assign n33771 = ( x947 & n33769 ) | ( x947 & n33770 ) | ( n33769 & n33770 ) ;
  assign n33772 = ( n5114 & n33596 ) | ( n5114 & ~n33771 ) | ( n33596 & ~n33771 ) ;
  assign n33773 = n33771 | n33772 ;
  assign n33774 = n1359 & ~n33773 ;
  assign n33775 = ( n1359 & n33765 ) | ( n1359 & n33774 ) | ( n33765 & n33774 ) ;
  assign n33776 = ( n33422 & ~n33750 ) | ( n33422 & n33775 ) | ( ~n33750 & n33775 ) ;
  assign n33777 = ~n33775 & n33776 ;
  assign n33778 = ( x221 & n33762 ) | ( x221 & ~n33777 ) | ( n33762 & ~n33777 ) ;
  assign n33779 = ~n33762 & n33778 ;
  assign n33780 = ( x299 & ~n33752 ) | ( x299 & n33779 ) | ( ~n33752 & n33779 ) ;
  assign n33781 = n33752 | n33780 ;
  assign n33782 = ( x39 & n33733 ) | ( x39 & n33781 ) | ( n33733 & n33781 ) ;
  assign n33783 = ~n33733 & n33782 ;
  assign n33784 = n15327 & n33695 ;
  assign n33785 = x221 & ~n15327 ;
  assign n33786 = ( x299 & ~n33784 ) | ( x299 & n33785 ) | ( ~n33784 & n33785 ) ;
  assign n33787 = n33784 | n33786 ;
  assign n33788 = n15330 & n33695 ;
  assign n33789 = x221 & ~n15330 ;
  assign n33790 = x299 & ~n33789 ;
  assign n33791 = n33790 ^ n33788 ^ 1'b0 ;
  assign n33792 = ( n33788 & n33790 ) | ( n33788 & n33791 ) | ( n33790 & n33791 ) ;
  assign n33793 = ( x39 & ~n33788 ) | ( x39 & n33792 ) | ( ~n33788 & n33792 ) ;
  assign n33794 = ( x38 & n33787 ) | ( x38 & ~n33793 ) | ( n33787 & ~n33793 ) ;
  assign n33795 = n33794 ^ n33787 ^ 1'b0 ;
  assign n33796 = ( x38 & n33794 ) | ( x38 & ~n33795 ) | ( n33794 & ~n33795 ) ;
  assign n33797 = ( ~n33699 & n33783 ) | ( ~n33699 & n33796 ) | ( n33783 & n33796 ) ;
  assign n33798 = ~n33699 & n33797 ;
  assign n33799 = n33798 ^ n8793 ^ 1'b0 ;
  assign n33800 = ( x221 & n33798 ) | ( x221 & n33799 ) | ( n33798 & n33799 ) ;
  assign n33801 = x38 | n15487 ;
  assign n33802 = x223 | n15476 ;
  assign n33803 = ~n15483 & n33802 ;
  assign n33804 = x299 | n33803 ;
  assign n33805 = x39 & ~n15474 ;
  assign n33806 = n33804 & n33805 ;
  assign n33807 = ( ~n17328 & n33801 ) | ( ~n17328 & n33806 ) | ( n33801 & n33806 ) ;
  assign n33808 = ~n17328 & n33807 ;
  assign n33809 = x222 & ~n33808 ;
  assign n33810 = n15392 & n15524 ;
  assign n33811 = x222 & ~n15337 ;
  assign n33812 = n2263 | n33811 ;
  assign n33813 = n33810 | n33812 ;
  assign n33814 = x616 & n15525 ;
  assign n33815 = n33814 ^ n15466 ^ n15392 ;
  assign n33816 = ~n5076 & n33815 ;
  assign n33817 = x616 & n15524 ;
  assign n33818 = n5076 & ~n33817 ;
  assign n33819 = n15445 & n33818 ;
  assign n33820 = ( n15382 & ~n33816 ) | ( n15382 & n33819 ) | ( ~n33816 & n33819 ) ;
  assign n33821 = n33816 | n33820 ;
  assign n33822 = n15382 & ~n33815 ;
  assign n33823 = n33821 & ~n33822 ;
  assign n33824 = ~n5061 & n33823 ;
  assign n33825 = n15382 ^ n5076 ^ 1'b0 ;
  assign n33826 = n15518 & ~n33817 ;
  assign n33827 = n15512 | n33826 ;
  assign n33828 = ( n5076 & ~n33825 ) | ( n5076 & n33827 ) | ( ~n33825 & n33827 ) ;
  assign n33829 = ( n15382 & n33825 ) | ( n15382 & n33828 ) | ( n33825 & n33828 ) ;
  assign n33830 = n15516 ^ x616 ^ 1'b0 ;
  assign n33831 = ( n15516 & n33708 ) | ( n15516 & ~n33830 ) | ( n33708 & ~n33830 ) ;
  assign n33832 = ( ~n5076 & n33829 ) | ( ~n5076 & n33831 ) | ( n33829 & n33831 ) ;
  assign n33833 = n33829 ^ n5076 ^ 1'b0 ;
  assign n33834 = ( n33829 & n33832 ) | ( n33829 & ~n33833 ) | ( n33832 & ~n33833 ) ;
  assign n33835 = n15382 & ~n33831 ;
  assign n33836 = n33834 & ~n33835 ;
  assign n33837 = n5061 & n33836 ;
  assign n33838 = ( x222 & n33824 ) | ( x222 & ~n33837 ) | ( n33824 & ~n33837 ) ;
  assign n33839 = ~n33824 & n33838 ;
  assign n33840 = x616 & n5076 ;
  assign n33841 = n15845 & n33840 ;
  assign n33842 = n15427 & n33817 ;
  assign n33843 = ~n5076 & n33842 ;
  assign n33844 = ( n15382 & ~n33841 ) | ( n15382 & n33843 ) | ( ~n33841 & n33843 ) ;
  assign n33845 = n33841 | n33844 ;
  assign n33846 = n15382 & ~n33842 ;
  assign n33847 = n33845 & ~n33846 ;
  assign n33848 = n5061 & ~n33847 ;
  assign n33849 = ( n15594 & n15595 ) | ( n15594 & ~n15598 ) | ( n15595 & ~n15598 ) ;
  assign n33850 = x616 & n33849 ;
  assign n33851 = n5061 | n33850 ;
  assign n33852 = ( x222 & ~n33848 ) | ( x222 & n33851 ) | ( ~n33848 & n33851 ) ;
  assign n33853 = ~x222 & n33852 ;
  assign n33854 = ( n2263 & n33839 ) | ( n2263 & ~n33853 ) | ( n33839 & ~n33853 ) ;
  assign n33855 = ~n33839 & n33854 ;
  assign n33856 = ( x215 & n33813 ) | ( x215 & ~n33855 ) | ( n33813 & ~n33855 ) ;
  assign n33857 = ~x215 & n33856 ;
  assign n33858 = n33814 ^ n15392 ^ n15371 ;
  assign n33859 = ~n5076 & n33858 ;
  assign n33860 = n15357 & n33818 ;
  assign n33861 = ( n15382 & ~n33859 ) | ( n15382 & n33860 ) | ( ~n33859 & n33860 ) ;
  assign n33862 = n33859 | n33861 ;
  assign n33863 = n15382 & ~n33858 ;
  assign n33864 = n33862 & ~n33863 ;
  assign n33865 = ~n5061 & n33864 ;
  assign n33866 = x616 & ~n15547 ;
  assign n33867 = n15361 & ~n33866 ;
  assign n33868 = n15364 | n33866 ;
  assign n33869 = n5076 | n15361 ;
  assign n33870 = ~n33868 & n33869 ;
  assign n33871 = n33867 ^ n15382 ^ 1'b0 ;
  assign n33872 = ( n33867 & n33870 ) | ( n33867 & ~n33871 ) | ( n33870 & ~n33871 ) ;
  assign n33873 = n5061 & n33872 ;
  assign n33874 = ( x222 & n33865 ) | ( x222 & ~n33873 ) | ( n33865 & ~n33873 ) ;
  assign n33875 = ~n33865 & n33874 ;
  assign n33876 = ( n5197 & n15595 ) | ( n5197 & n15607 ) | ( n15595 & n15607 ) ;
  assign n33877 = x616 & n33876 ;
  assign n33878 = ~x222 & n33877 ;
  assign n33879 = ~n15613 & n33878 ;
  assign n33880 = ( x215 & n33875 ) | ( x215 & n33879 ) | ( n33875 & n33879 ) ;
  assign n33881 = n33879 ^ n33875 ^ 1'b0 ;
  assign n33882 = ( x215 & n33880 ) | ( x215 & n33881 ) | ( n33880 & n33881 ) ;
  assign n33883 = ( x299 & n33857 ) | ( x299 & ~n33882 ) | ( n33857 & ~n33882 ) ;
  assign n33884 = ~n33857 & n33883 ;
  assign n33885 = n5114 & n33872 ;
  assign n33886 = ~n5114 & n33864 ;
  assign n33887 = ( x222 & n33885 ) | ( x222 & ~n33886 ) | ( n33885 & ~n33886 ) ;
  assign n33888 = ~n33885 & n33887 ;
  assign n33889 = ~n15618 & n33878 ;
  assign n33890 = ( x223 & n33888 ) | ( x223 & ~n33889 ) | ( n33888 & ~n33889 ) ;
  assign n33891 = ~n33888 & n33890 ;
  assign n33892 = n5114 & n33847 ;
  assign n33893 = ~n5114 & n33850 ;
  assign n33894 = ( x224 & n33892 ) | ( x224 & ~n33893 ) | ( n33892 & ~n33893 ) ;
  assign n33895 = ~n33892 & n33894 ;
  assign n33896 = x224 | n33810 ;
  assign n33897 = ( x222 & ~n33895 ) | ( x222 & n33896 ) | ( ~n33895 & n33896 ) ;
  assign n33898 = ~x222 & n33897 ;
  assign n33899 = ~n5114 & n33823 ;
  assign n33900 = n5114 & n33836 ;
  assign n33901 = ( x222 & n33899 ) | ( x222 & ~n33900 ) | ( n33899 & ~n33900 ) ;
  assign n33902 = ~n33899 & n33901 ;
  assign n33903 = ( x223 & ~n33898 ) | ( x223 & n33902 ) | ( ~n33898 & n33902 ) ;
  assign n33904 = n33898 | n33903 ;
  assign n33905 = n33904 ^ n33891 ^ 1'b0 ;
  assign n33906 = ( n33891 & n33904 ) | ( n33891 & n33905 ) | ( n33904 & n33905 ) ;
  assign n33907 = ( x299 & ~n33891 ) | ( x299 & n33906 ) | ( ~n33891 & n33906 ) ;
  assign n33908 = ( x39 & n33884 ) | ( x39 & n33907 ) | ( n33884 & n33907 ) ;
  assign n33909 = ~n33884 & n33908 ;
  assign n33910 = x222 & n15509 ;
  assign n33911 = ~x616 & n15638 ;
  assign n33912 = x39 | n33911 ;
  assign n33913 = x222 | n15638 ;
  assign n33914 = ( n33910 & ~n33912 ) | ( n33910 & n33913 ) | ( ~n33912 & n33913 ) ;
  assign n33915 = ~n33910 & n33914 ;
  assign n33916 = ( x38 & ~n33909 ) | ( x38 & n33915 ) | ( ~n33909 & n33915 ) ;
  assign n33917 = n33909 | n33916 ;
  assign n33918 = x222 & ~n15644 ;
  assign n33919 = x38 & ~n33918 ;
  assign n33920 = x616 & n15646 ;
  assign n33921 = n33919 & ~n33920 ;
  assign n33922 = ( n2069 & n33917 ) | ( n2069 & ~n33921 ) | ( n33917 & ~n33921 ) ;
  assign n33923 = ~n2069 & n33922 ;
  assign n33924 = n33923 ^ x222 ^ 1'b0 ;
  assign n33925 = ( ~x222 & n2069 ) | ( ~x222 & n33924 ) | ( n2069 & n33924 ) ;
  assign n33926 = ( x222 & n33923 ) | ( x222 & n33925 ) | ( n33923 & n33925 ) ;
  assign n33927 = n33809 ^ n15659 ^ 1'b0 ;
  assign n33928 = ( n33809 & n33926 ) | ( n33809 & ~n33927 ) | ( n33926 & ~n33927 ) ;
  assign n33929 = x609 & ~n33928 ;
  assign n33930 = x609 | n33809 ;
  assign n33931 = ( x1155 & n33929 ) | ( x1155 & n33930 ) | ( n33929 & n33930 ) ;
  assign n33932 = ~n33929 & n33931 ;
  assign n33933 = x609 & ~n33809 ;
  assign n33934 = x1155 | n33933 ;
  assign n33935 = ( n33928 & n33929 ) | ( n33928 & ~n33934 ) | ( n33929 & ~n33934 ) ;
  assign n33936 = n33932 | n33935 ;
  assign n33937 = n33928 ^ x785 ^ 1'b0 ;
  assign n33938 = ( n33928 & n33936 ) | ( n33928 & n33937 ) | ( n33936 & n33937 ) ;
  assign n33939 = x618 & ~n33938 ;
  assign n33940 = x618 | n33809 ;
  assign n33941 = ( x1154 & n33939 ) | ( x1154 & n33940 ) | ( n33939 & n33940 ) ;
  assign n33942 = ~n33939 & n33941 ;
  assign n33943 = x618 & ~n33809 ;
  assign n33944 = x1154 | n33943 ;
  assign n33945 = ( n33938 & n33939 ) | ( n33938 & ~n33944 ) | ( n33939 & ~n33944 ) ;
  assign n33946 = n33942 | n33945 ;
  assign n33947 = n33938 ^ x781 ^ 1'b0 ;
  assign n33948 = ( n33938 & n33946 ) | ( n33938 & n33947 ) | ( n33946 & n33947 ) ;
  assign n33949 = x619 & ~n33948 ;
  assign n33950 = x619 | n33809 ;
  assign n33951 = ( x1159 & n33949 ) | ( x1159 & n33950 ) | ( n33949 & n33950 ) ;
  assign n33952 = ~n33949 & n33951 ;
  assign n33953 = x619 & ~n33809 ;
  assign n33954 = x1159 | n33953 ;
  assign n33955 = ( n33948 & n33949 ) | ( n33948 & ~n33954 ) | ( n33949 & ~n33954 ) ;
  assign n33956 = n33952 | n33955 ;
  assign n33957 = n33948 ^ x789 ^ 1'b0 ;
  assign n33958 = ( n33948 & n33956 ) | ( n33948 & n33957 ) | ( n33956 & n33957 ) ;
  assign n33959 = n33809 ^ n16518 ^ 1'b0 ;
  assign n33960 = ( n33809 & n33958 ) | ( n33809 & ~n33959 ) | ( n33958 & ~n33959 ) ;
  assign n33961 = n33809 ^ n16339 ^ 1'b0 ;
  assign n33962 = ( n33809 & n33960 ) | ( n33809 & ~n33961 ) | ( n33960 & ~n33961 ) ;
  assign n33963 = n19055 & n33962 ;
  assign n33964 = x661 & n16184 ;
  assign n33965 = n33919 & ~n33964 ;
  assign n33988 = x661 & n16164 ;
  assign n34016 = n33812 | n33988 ;
  assign n33992 = n15429 ^ x680 ^ 1'b0 ;
  assign n33993 = ( n15429 & n15949 ) | ( n15429 & n33992 ) | ( n15949 & n33992 ) ;
  assign n33994 = n15433 ^ x661 ^ 1'b0 ;
  assign n33995 = ( n15433 & n33993 ) | ( n15433 & n33994 ) | ( n33993 & n33994 ) ;
  assign n34017 = n5061 & n33995 ;
  assign n33997 = ~x662 & n15454 ;
  assign n33998 = n5076 | n15466 ;
  assign n33999 = n33998 ^ n33997 ^ 1'b0 ;
  assign n34000 = ( n33997 & n33998 ) | ( n33997 & n33999 ) | ( n33998 & n33999 ) ;
  assign n34001 = ( n15382 & ~n33997 ) | ( n15382 & n34000 ) | ( ~n33997 & n34000 ) ;
  assign n34002 = n34001 ^ x661 ^ 1'b0 ;
  assign n34003 = ( x661 & ~n15467 ) | ( x661 & n34002 ) | ( ~n15467 & n34002 ) ;
  assign n34004 = ( n34001 & ~n34002 ) | ( n34001 & n34003 ) | ( ~n34002 & n34003 ) ;
  assign n34005 = n34004 ^ n16119 ^ 1'b0 ;
  assign n34006 = ( ~x661 & n16119 ) | ( ~x661 & n34005 ) | ( n16119 & n34005 ) ;
  assign n34007 = ( n34004 & ~n34005 ) | ( n34004 & n34006 ) | ( ~n34005 & n34006 ) ;
  assign n34018 = ~n5061 & n34007 ;
  assign n34019 = ( x222 & n34017 ) | ( x222 & ~n34018 ) | ( n34017 & ~n34018 ) ;
  assign n34020 = ~n34017 & n34019 ;
  assign n33981 = x661 & x680 ;
  assign n33982 = n16146 & n33981 ;
  assign n34021 = n5061 | n33982 ;
  assign n33984 = x661 & n16152 ;
  assign n34022 = n5061 & ~n33984 ;
  assign n34023 = ( x222 & n34021 ) | ( x222 & ~n34022 ) | ( n34021 & ~n34022 ) ;
  assign n34024 = ~x222 & n34023 ;
  assign n34025 = ( n2263 & n34020 ) | ( n2263 & ~n34024 ) | ( n34020 & ~n34024 ) ;
  assign n34026 = ~n34020 & n34025 ;
  assign n34027 = ( x215 & n34016 ) | ( x215 & ~n34026 ) | ( n34016 & ~n34026 ) ;
  assign n34028 = ~x215 & n34027 ;
  assign n33966 = n15817 & ~n16097 ;
  assign n33967 = n15402 ^ x661 ^ 1'b0 ;
  assign n33968 = ( n15402 & n33966 ) | ( n15402 & n33967 ) | ( n33966 & n33967 ) ;
  assign n34029 = ~n5061 & n33968 ;
  assign n33970 = n15362 ^ x661 ^ 1'b0 ;
  assign n33971 = ( n15362 & ~n16100 ) | ( n15362 & n33970 ) | ( ~n16100 & n33970 ) ;
  assign n33972 = ( n15374 & n15382 ) | ( n15374 & ~n33971 ) | ( n15382 & ~n33971 ) ;
  assign n33973 = ~n33971 & n33972 ;
  assign n34030 = n5061 & n33973 ;
  assign n34031 = ( x222 & n34029 ) | ( x222 & ~n34030 ) | ( n34029 & ~n34030 ) ;
  assign n34032 = ~n34029 & n34031 ;
  assign n33977 = ~x222 & x661 ;
  assign n34033 = n16172 & n33977 ;
  assign n34034 = ( x215 & n34032 ) | ( x215 & n34033 ) | ( n34032 & n34033 ) ;
  assign n34035 = n34033 ^ n34032 ^ 1'b0 ;
  assign n34036 = ( x215 & n34034 ) | ( x215 & n34035 ) | ( n34034 & n34035 ) ;
  assign n34037 = ( x299 & n34028 ) | ( x299 & ~n34036 ) | ( n34028 & ~n34036 ) ;
  assign n34038 = ~n34028 & n34037 ;
  assign n33969 = ~n5114 & n33968 ;
  assign n33974 = n5114 & n33973 ;
  assign n33975 = ( x222 & n33969 ) | ( x222 & ~n33974 ) | ( n33969 & ~n33974 ) ;
  assign n33976 = ~n33969 & n33975 ;
  assign n33978 = n16144 & n33977 ;
  assign n33979 = ( x223 & n33976 ) | ( x223 & ~n33978 ) | ( n33976 & ~n33978 ) ;
  assign n33980 = ~n33976 & n33979 ;
  assign n33983 = ~n5114 & n33982 ;
  assign n33985 = n5114 & n33984 ;
  assign n33986 = ( x224 & n33983 ) | ( x224 & ~n33985 ) | ( n33983 & ~n33985 ) ;
  assign n33987 = ~n33983 & n33986 ;
  assign n33989 = x224 | n33988 ;
  assign n33990 = ( x222 & ~n33987 ) | ( x222 & n33989 ) | ( ~n33987 & n33989 ) ;
  assign n33991 = ~x222 & n33990 ;
  assign n33996 = n5114 & n33995 ;
  assign n34008 = ~n5114 & n34007 ;
  assign n34009 = ( x222 & n33996 ) | ( x222 & ~n34008 ) | ( n33996 & ~n34008 ) ;
  assign n34010 = ~n33996 & n34009 ;
  assign n34011 = ( x223 & ~n33991 ) | ( x223 & n34010 ) | ( ~n33991 & n34010 ) ;
  assign n34012 = n33991 | n34011 ;
  assign n34013 = n34012 ^ n33980 ^ 1'b0 ;
  assign n34014 = ( n33980 & n34012 ) | ( n33980 & n34013 ) | ( n34012 & n34013 ) ;
  assign n34015 = ( x299 & ~n33980 ) | ( x299 & n34014 ) | ( ~n33980 & n34014 ) ;
  assign n34039 = n34038 ^ n34015 ^ 1'b0 ;
  assign n34040 = ( x39 & ~n34015 ) | ( x39 & n34038 ) | ( ~n34015 & n34038 ) ;
  assign n34041 = ( x39 & ~n34039 ) | ( x39 & n34040 ) | ( ~n34039 & n34040 ) ;
  assign n34042 = x222 & n16038 ;
  assign n34043 = x299 | n34042 ;
  assign n34044 = n33981 & ~n34043 ;
  assign n34045 = ( n16018 & n34043 ) | ( n16018 & ~n34044 ) | ( n34043 & ~n34044 ) ;
  assign n34046 = ( x222 & n16018 ) | ( x222 & ~n34045 ) | ( n16018 & ~n34045 ) ;
  assign n34047 = ~n34045 & n34046 ;
  assign n34048 = x222 & n16033 ;
  assign n34049 = n16024 & ~n33981 ;
  assign n34050 = ( x299 & n34048 ) | ( x299 & ~n34049 ) | ( n34048 & ~n34049 ) ;
  assign n34051 = ~n34048 & n34050 ;
  assign n34052 = n16024 ^ x222 ^ 1'b0 ;
  assign n34053 = ( x222 & n16024 ) | ( x222 & ~n34052 ) | ( n16024 & ~n34052 ) ;
  assign n34054 = ( n34051 & n34052 ) | ( n34051 & n34053 ) | ( n34052 & n34053 ) ;
  assign n34055 = ( x39 & ~n34047 ) | ( x39 & n34054 ) | ( ~n34047 & n34054 ) ;
  assign n34056 = n34047 | n34055 ;
  assign n34057 = n34056 ^ n34041 ^ 1'b0 ;
  assign n34058 = ( n34041 & n34056 ) | ( n34041 & n34057 ) | ( n34056 & n34057 ) ;
  assign n34059 = ( x38 & ~n34041 ) | ( x38 & n34058 ) | ( ~n34041 & n34058 ) ;
  assign n34060 = ( n2069 & ~n33965 ) | ( n2069 & n34059 ) | ( ~n33965 & n34059 ) ;
  assign n34061 = ~n2069 & n34060 ;
  assign n34062 = n34061 ^ x222 ^ 1'b0 ;
  assign n34063 = ( ~x222 & n2069 ) | ( ~x222 & n34062 ) | ( n2069 & n34062 ) ;
  assign n34064 = ( x222 & n34061 ) | ( x222 & n34063 ) | ( n34061 & n34063 ) ;
  assign n34065 = x625 & ~n34064 ;
  assign n34066 = x625 | n33809 ;
  assign n34067 = ( x1153 & n34065 ) | ( x1153 & n34066 ) | ( n34065 & n34066 ) ;
  assign n34068 = ~n34065 & n34067 ;
  assign n34069 = x625 & ~n33809 ;
  assign n34070 = x1153 | n34069 ;
  assign n34071 = ( n34064 & n34065 ) | ( n34064 & ~n34070 ) | ( n34065 & ~n34070 ) ;
  assign n34072 = n34068 | n34071 ;
  assign n34073 = n34064 ^ x778 ^ 1'b0 ;
  assign n34074 = ( n34064 & n34072 ) | ( n34064 & n34073 ) | ( n34072 & n34073 ) ;
  assign n34075 = n33809 ^ n16234 ^ 1'b0 ;
  assign n34076 = ( n33809 & n34074 ) | ( n33809 & ~n34075 ) | ( n34074 & ~n34075 ) ;
  assign n34077 = n33809 ^ n16254 ^ 1'b0 ;
  assign n34078 = ( n33809 & n34076 ) | ( n33809 & ~n34077 ) | ( n34076 & ~n34077 ) ;
  assign n34079 = n16279 | n34078 ;
  assign n34080 = n16318 | n34079 ;
  assign n34081 = n17086 & ~n33809 ;
  assign n34082 = n34080 & ~n34081 ;
  assign n34083 = n17093 | n34082 ;
  assign n34084 = n16559 & ~n33809 ;
  assign n34085 = n34083 & ~n34084 ;
  assign n34086 = x647 & ~n34085 ;
  assign n34087 = x647 | n33809 ;
  assign n34088 = ( x1157 & n34086 ) | ( x1157 & n34087 ) | ( n34086 & n34087 ) ;
  assign n34089 = ~n34086 & n34088 ;
  assign n34090 = x647 & ~n33809 ;
  assign n34091 = x1157 | n34090 ;
  assign n34092 = ( n34085 & n34086 ) | ( n34085 & ~n34091 ) | ( n34086 & ~n34091 ) ;
  assign n34093 = ( n16375 & n34089 ) | ( n16375 & n34092 ) | ( n34089 & n34092 ) ;
  assign n34094 = ( x787 & n33963 ) | ( x787 & n34093 ) | ( n33963 & n34093 ) ;
  assign n34095 = n34093 ^ n33963 ^ 1'b0 ;
  assign n34096 = ( x787 & n34094 ) | ( x787 & n34095 ) | ( n34094 & n34095 ) ;
  assign n34097 = n16279 & ~n33809 ;
  assign n34098 = ( n16459 & n34079 ) | ( n16459 & n34097 ) | ( n34079 & n34097 ) ;
  assign n34099 = ~n34097 & n34098 ;
  assign n34100 = x626 | n33809 ;
  assign n34101 = x626 & ~n33958 ;
  assign n34102 = n22317 & ~n34101 ;
  assign n34103 = n34100 & n34102 ;
  assign n34104 = x626 & ~n33809 ;
  assign n34105 = n22322 & ~n34104 ;
  assign n34106 = ( n33958 & n34101 ) | ( n33958 & n34105 ) | ( n34101 & n34105 ) ;
  assign n34107 = ( ~n34099 & n34103 ) | ( ~n34099 & n34106 ) | ( n34103 & n34106 ) ;
  assign n34108 = n34099 | n34107 ;
  assign n34109 = n16519 & ~n34108 ;
  assign n34114 = n16026 & ~n33981 ;
  assign n34115 = x603 | n16033 ;
  assign n34116 = n15494 | n15698 ;
  assign n34117 = n34115 & ~n34116 ;
  assign n34118 = ~x616 & n15636 ;
  assign n34119 = n34117 | n34118 ;
  assign n34120 = ( x222 & n34114 ) | ( x222 & n34119 ) | ( n34114 & n34119 ) ;
  assign n34121 = n34119 ^ n34114 ^ 1'b0 ;
  assign n34122 = ( x222 & n34120 ) | ( x222 & n34121 ) | ( n34120 & n34121 ) ;
  assign n34110 = x661 & n16027 ;
  assign n34111 = x616 & n15636 ;
  assign n34112 = ( x222 & ~n34110 ) | ( x222 & n34111 ) | ( ~n34110 & n34111 ) ;
  assign n34113 = n34110 | n34112 ;
  assign n34123 = n34122 ^ n34113 ^ 1'b0 ;
  assign n34124 = ( x299 & ~n34113 ) | ( x299 & n34122 ) | ( ~n34113 & n34122 ) ;
  assign n34125 = ( x299 & ~n34123 ) | ( x299 & n34124 ) | ( ~n34123 & n34124 ) ;
  assign n34126 = x661 & n16021 ;
  assign n34127 = x616 & n15633 ;
  assign n34128 = ( x222 & ~n34126 ) | ( x222 & n34127 ) | ( ~n34126 & n34127 ) ;
  assign n34129 = n34126 | n34128 ;
  assign n34130 = n16020 & ~n33981 ;
  assign n34131 = n15698 | n16011 ;
  assign n34132 = x603 | n16038 ;
  assign n34133 = ~n34131 & n34132 ;
  assign n34134 = ~x616 & n15633 ;
  assign n34135 = n34133 | n34134 ;
  assign n34136 = ( x222 & n34130 ) | ( x222 & n34135 ) | ( n34130 & n34135 ) ;
  assign n34137 = n34135 ^ n34130 ^ 1'b0 ;
  assign n34138 = ( x222 & n34136 ) | ( x222 & n34137 ) | ( n34136 & n34137 ) ;
  assign n34139 = ( x299 & n34129 ) | ( x299 & ~n34138 ) | ( n34129 & ~n34138 ) ;
  assign n34140 = n34139 ^ n34129 ^ 1'b0 ;
  assign n34141 = ( x299 & n34139 ) | ( x299 & ~n34140 ) | ( n34139 & ~n34140 ) ;
  assign n34142 = ( x39 & ~n34125 ) | ( x39 & n34141 ) | ( ~n34125 & n34141 ) ;
  assign n34143 = ~x39 & n34142 ;
  assign n34144 = x616 & n15609 ;
  assign n34145 = ~x680 & n34144 ;
  assign n34146 = n15609 | n15880 ;
  assign n34147 = x616 & ~n34146 ;
  assign n34148 = ( x680 & n15764 ) | ( x680 & n34147 ) | ( n15764 & n34147 ) ;
  assign n34149 = ~n34147 & n34148 ;
  assign n34150 = ( x661 & n34145 ) | ( x661 & ~n34149 ) | ( n34145 & ~n34149 ) ;
  assign n34151 = ~n34145 & n34150 ;
  assign n34152 = n15351 & n33810 ;
  assign n34153 = n5078 & ~n34152 ;
  assign n34154 = x661 | n34144 ;
  assign n34155 = ( n34151 & ~n34153 ) | ( n34151 & n34154 ) | ( ~n34153 & n34154 ) ;
  assign n34156 = ~n34151 & n34155 ;
  assign n34157 = n5114 & n34156 ;
  assign n34158 = n15751 & n33981 ;
  assign n34159 = n33877 | n34158 ;
  assign n34160 = ~n5114 & n34159 ;
  assign n34161 = ( x222 & ~n34157 ) | ( x222 & n34160 ) | ( ~n34157 & n34160 ) ;
  assign n34162 = n34157 | n34161 ;
  assign n34163 = ~x661 & x681 ;
  assign n34164 = ~n33867 & n34163 ;
  assign n34165 = n15382 | n33870 ;
  assign n34166 = ~x680 & n33867 ;
  assign n34167 = n15802 & n15890 ;
  assign n34168 = x616 & ~n34167 ;
  assign n34169 = ( x680 & n15805 ) | ( x680 & n34168 ) | ( n15805 & n34168 ) ;
  assign n34170 = ~n34168 & n34169 ;
  assign n34171 = ( x661 & n34166 ) | ( x661 & ~n34170 ) | ( n34166 & ~n34170 ) ;
  assign n34172 = ~n34166 & n34171 ;
  assign n34173 = ( n34164 & n34165 ) | ( n34164 & ~n34172 ) | ( n34165 & ~n34172 ) ;
  assign n34174 = ~n34164 & n34173 ;
  assign n34175 = n5114 & ~n34174 ;
  assign n34176 = x616 & ~n15954 ;
  assign n34177 = x680 & ~n34176 ;
  assign n34178 = n15828 & n34177 ;
  assign n34179 = ~x680 & n33858 ;
  assign n34180 = ( x661 & n34178 ) | ( x661 & ~n34179 ) | ( n34178 & ~n34179 ) ;
  assign n34181 = ~n34178 & n34180 ;
  assign n34182 = ~n33858 & n34163 ;
  assign n34183 = ( n33862 & n34181 ) | ( n33862 & ~n34182 ) | ( n34181 & ~n34182 ) ;
  assign n34184 = ~n34181 & n34183 ;
  assign n34185 = n5114 | n34184 ;
  assign n34186 = ( x222 & n34175 ) | ( x222 & n34185 ) | ( n34175 & n34185 ) ;
  assign n34187 = ~n34175 & n34186 ;
  assign n34188 = x223 & ~n34187 ;
  assign n34189 = n34162 & n34188 ;
  assign n34190 = ~x680 & n33842 ;
  assign n34191 = x616 & ~n15905 ;
  assign n34192 = x680 & ~n34191 ;
  assign n34193 = n15741 & n34192 ;
  assign n34194 = ( x661 & n34190 ) | ( x661 & ~n34193 ) | ( n34190 & ~n34193 ) ;
  assign n34195 = ~n34190 & n34194 ;
  assign n34196 = ~n33842 & n34163 ;
  assign n34197 = ( n33845 & n34195 ) | ( n33845 & ~n34196 ) | ( n34195 & ~n34196 ) ;
  assign n34198 = ~n34195 & n34197 ;
  assign n34199 = n5114 & n34198 ;
  assign n34200 = ~n33810 & n34163 ;
  assign n34201 = n15594 & n33840 ;
  assign n34202 = ~n5076 & n33810 ;
  assign n34203 = ( n15382 & ~n34201 ) | ( n15382 & n34202 ) | ( ~n34201 & n34202 ) ;
  assign n34204 = n34201 | n34203 ;
  assign n34205 = x616 & ~n15891 ;
  assign n34206 = x680 & n15704 ;
  assign n34207 = ~n34205 & n34206 ;
  assign n34208 = ~x680 & n33810 ;
  assign n34209 = ( x661 & n34207 ) | ( x661 & ~n34208 ) | ( n34207 & ~n34208 ) ;
  assign n34210 = ~n34207 & n34209 ;
  assign n34211 = ( n34200 & n34204 ) | ( n34200 & ~n34210 ) | ( n34204 & ~n34210 ) ;
  assign n34212 = ~n34200 & n34211 ;
  assign n34213 = ~n5114 & n34212 ;
  assign n34214 = ( x224 & n34199 ) | ( x224 & ~n34213 ) | ( n34199 & ~n34213 ) ;
  assign n34215 = ~n34199 & n34214 ;
  assign n34216 = ( n15392 & n15694 ) | ( n15392 & n15891 ) | ( n15694 & n15891 ) ;
  assign n34217 = n33981 & ~n34216 ;
  assign n34218 = n33810 | n33981 ;
  assign n34219 = ( x222 & ~n34217 ) | ( x222 & n34218 ) | ( ~n34217 & n34218 ) ;
  assign n34220 = ~x222 & n34219 ;
  assign n34221 = ( n2161 & ~n34215 ) | ( n2161 & n34220 ) | ( ~n34215 & n34220 ) ;
  assign n34222 = ~n34215 & n34221 ;
  assign n34223 = n15712 | n15904 ;
  assign n34224 = x642 & n34223 ;
  assign n34225 = x603 & ~n15425 ;
  assign n34226 = n15706 | n34225 ;
  assign n34227 = ( x603 & n15712 ) | ( x603 & ~n34226 ) | ( n15712 & ~n34226 ) ;
  assign n34228 = ~n34226 & n34227 ;
  assign n34229 = ~x642 & n34228 ;
  assign n34230 = ( n5080 & ~n34224 ) | ( n5080 & n34229 ) | ( ~n34224 & n34229 ) ;
  assign n34231 = n34224 | n34230 ;
  assign n34232 = n15762 & ~n34223 ;
  assign n34233 = n15712 & n15890 ;
  assign n34234 = x616 & ~n34233 ;
  assign n34235 = ( x680 & n34232 ) | ( x680 & ~n34234 ) | ( n34232 & ~n34234 ) ;
  assign n34236 = ~n34232 & n34235 ;
  assign n34237 = x661 & ~n34236 ;
  assign n34238 = ( x661 & ~n34231 ) | ( x661 & n34237 ) | ( ~n34231 & n34237 ) ;
  assign n34239 = n34238 ^ x680 ^ 1'b0 ;
  assign n34240 = ( x680 & ~n33831 ) | ( x680 & n34239 ) | ( ~n33831 & n34239 ) ;
  assign n34241 = ( n34238 & ~n34239 ) | ( n34238 & n34240 ) | ( ~n34239 & n34240 ) ;
  assign n34242 = ~n33831 & n34163 ;
  assign n34243 = ( n33834 & n34241 ) | ( n33834 & ~n34242 ) | ( n34241 & ~n34242 ) ;
  assign n34244 = ~n34241 & n34243 ;
  assign n34245 = n5114 & n34244 ;
  assign n34246 = n15836 & n34177 ;
  assign n34247 = ~x680 & n33815 ;
  assign n34248 = ( x661 & n34246 ) | ( x661 & ~n34247 ) | ( n34246 & ~n34247 ) ;
  assign n34249 = ~n34246 & n34248 ;
  assign n34250 = ~n33815 & n34163 ;
  assign n34251 = ( n33821 & n34249 ) | ( n33821 & ~n34250 ) | ( n34249 & ~n34250 ) ;
  assign n34252 = ~n34249 & n34251 ;
  assign n34253 = ~n5114 & n34252 ;
  assign n34254 = ( x222 & n34245 ) | ( x222 & ~n34253 ) | ( n34245 & ~n34253 ) ;
  assign n34255 = ~n34245 & n34254 ;
  assign n34256 = ( ~x223 & n34222 ) | ( ~x223 & n34255 ) | ( n34222 & n34255 ) ;
  assign n34257 = ~x223 & n34256 ;
  assign n34258 = ( x299 & ~n34189 ) | ( x299 & n34257 ) | ( ~n34189 & n34257 ) ;
  assign n34259 = n34189 | n34258 ;
  assign n34260 = n5061 & ~n34244 ;
  assign n34261 = n5061 | n34252 ;
  assign n34262 = ( x222 & n34260 ) | ( x222 & n34261 ) | ( n34260 & n34261 ) ;
  assign n34263 = ~n34260 & n34262 ;
  assign n34264 = n5061 & n34198 ;
  assign n34265 = ~n5061 & n34212 ;
  assign n34266 = x222 | n34265 ;
  assign n34267 = ( ~n34263 & n34264 ) | ( ~n34263 & n34266 ) | ( n34264 & n34266 ) ;
  assign n34268 = ~n34263 & n34267 ;
  assign n34269 = ( x216 & x221 ) | ( x216 & ~n34268 ) | ( x221 & ~n34268 ) ;
  assign n34270 = ~n34268 & n34269 ;
  assign n34271 = n33817 | n33981 ;
  assign n34272 = n34216 & n34271 ;
  assign n34273 = n33812 | n34272 ;
  assign n34274 = ( x215 & ~n34270 ) | ( x215 & n34273 ) | ( ~n34270 & n34273 ) ;
  assign n34275 = ~x215 & n34274 ;
  assign n34276 = n5061 & n34156 ;
  assign n34277 = ~n5061 & n34159 ;
  assign n34278 = ( x222 & ~n34276 ) | ( x222 & n34277 ) | ( ~n34276 & n34277 ) ;
  assign n34279 = n34276 | n34278 ;
  assign n34280 = n5061 & ~n34174 ;
  assign n34281 = n5061 | n34184 ;
  assign n34282 = ( x222 & n34280 ) | ( x222 & n34281 ) | ( n34280 & n34281 ) ;
  assign n34283 = ~n34280 & n34282 ;
  assign n34284 = x215 & ~n34283 ;
  assign n34285 = n34279 & n34284 ;
  assign n34286 = ( x299 & n34275 ) | ( x299 & ~n34285 ) | ( n34275 & ~n34285 ) ;
  assign n34287 = ~n34275 & n34286 ;
  assign n34288 = x39 & ~n34287 ;
  assign n34289 = n34259 & n34288 ;
  assign n34290 = ( x38 & ~n34143 ) | ( x38 & n34289 ) | ( ~n34143 & n34289 ) ;
  assign n34291 = n34143 | n34290 ;
  assign n34292 = ~x39 & x616 ;
  assign n34293 = n33981 & n34292 ;
  assign n34294 = ( x222 & x616 ) | ( x222 & ~n34293 ) | ( x616 & ~n34293 ) ;
  assign n34295 = ~n34293 & n34294 ;
  assign n34296 = ( n15340 & n15890 ) | ( n15340 & n34295 ) | ( n15890 & n34295 ) ;
  assign n34297 = ~n34295 & n34296 ;
  assign n34298 = x616 | n15691 ;
  assign n34299 = ( ~n15644 & n34271 ) | ( ~n15644 & n34298 ) | ( n34271 & n34298 ) ;
  assign n34300 = n15644 & n34299 ;
  assign n34301 = n15644 & ~n34300 ;
  assign n34302 = ( x222 & n34300 ) | ( x222 & ~n34301 ) | ( n34300 & ~n34301 ) ;
  assign n34303 = x38 & ~n34302 ;
  assign n34304 = ( x38 & n34297 ) | ( x38 & n34303 ) | ( n34297 & n34303 ) ;
  assign n34305 = ( n2069 & n34291 ) | ( n2069 & ~n34304 ) | ( n34291 & ~n34304 ) ;
  assign n34306 = ~n2069 & n34305 ;
  assign n34307 = n34306 ^ x222 ^ 1'b0 ;
  assign n34308 = ( ~x222 & n2069 ) | ( ~x222 & n34307 ) | ( n2069 & n34307 ) ;
  assign n34309 = ( x222 & n34306 ) | ( x222 & n34308 ) | ( n34306 & n34308 ) ;
  assign n34310 = x625 & ~n34309 ;
  assign n34311 = x625 | n33926 ;
  assign n34312 = ( x1153 & n34310 ) | ( x1153 & n34311 ) | ( n34310 & n34311 ) ;
  assign n34313 = ~n34310 & n34312 ;
  assign n34314 = ( x608 & n34071 ) | ( x608 & ~n34313 ) | ( n34071 & ~n34313 ) ;
  assign n34315 = ~n34071 & n34314 ;
  assign n34316 = x625 & ~n33926 ;
  assign n34317 = x1153 | n34316 ;
  assign n34318 = ( x625 & n34309 ) | ( x625 & ~n34317 ) | ( n34309 & ~n34317 ) ;
  assign n34319 = ~n34317 & n34318 ;
  assign n34320 = x608 | n34068 ;
  assign n34321 = ( ~n34315 & n34319 ) | ( ~n34315 & n34320 ) | ( n34319 & n34320 ) ;
  assign n34322 = ~n34315 & n34321 ;
  assign n34323 = n34309 ^ x778 ^ 1'b0 ;
  assign n34324 = ( n34309 & n34322 ) | ( n34309 & n34323 ) | ( n34322 & n34323 ) ;
  assign n34325 = x609 & ~n34324 ;
  assign n34326 = x609 | n34074 ;
  assign n34327 = ( x1155 & n34325 ) | ( x1155 & n34326 ) | ( n34325 & n34326 ) ;
  assign n34328 = ~n34325 & n34327 ;
  assign n34329 = ( x660 & n33935 ) | ( x660 & ~n34328 ) | ( n33935 & ~n34328 ) ;
  assign n34330 = ~n33935 & n34329 ;
  assign n34331 = x609 & ~n34074 ;
  assign n34332 = x1155 | n34331 ;
  assign n34333 = ( x609 & n34324 ) | ( x609 & ~n34332 ) | ( n34324 & ~n34332 ) ;
  assign n34334 = ~n34332 & n34333 ;
  assign n34335 = x660 | n33932 ;
  assign n34336 = ( ~n34330 & n34334 ) | ( ~n34330 & n34335 ) | ( n34334 & n34335 ) ;
  assign n34337 = ~n34330 & n34336 ;
  assign n34338 = n34324 ^ x785 ^ 1'b0 ;
  assign n34339 = ( n34324 & n34337 ) | ( n34324 & n34338 ) | ( n34337 & n34338 ) ;
  assign n34340 = x618 & ~n34339 ;
  assign n34341 = x618 | n34076 ;
  assign n34342 = ( x1154 & n34340 ) | ( x1154 & n34341 ) | ( n34340 & n34341 ) ;
  assign n34343 = ~n34340 & n34342 ;
  assign n34344 = ( x627 & n33945 ) | ( x627 & ~n34343 ) | ( n33945 & ~n34343 ) ;
  assign n34345 = ~n33945 & n34344 ;
  assign n34346 = x627 | n33942 ;
  assign n34347 = x618 & ~n34076 ;
  assign n34348 = x1154 | n34347 ;
  assign n34349 = ( n34339 & n34340 ) | ( n34339 & ~n34348 ) | ( n34340 & ~n34348 ) ;
  assign n34350 = ( ~n34345 & n34346 ) | ( ~n34345 & n34349 ) | ( n34346 & n34349 ) ;
  assign n34351 = ~n34345 & n34350 ;
  assign n34352 = n34339 ^ x781 ^ 1'b0 ;
  assign n34353 = ( n34339 & n34351 ) | ( n34339 & n34352 ) | ( n34351 & n34352 ) ;
  assign n34354 = ~x789 & n34353 ;
  assign n34355 = x619 | n34078 ;
  assign n34356 = x619 & ~n34353 ;
  assign n34357 = x1159 & ~n34356 ;
  assign n34358 = n34355 & n34357 ;
  assign n34359 = ( x648 & n33955 ) | ( x648 & ~n34358 ) | ( n33955 & ~n34358 ) ;
  assign n34360 = ~n33955 & n34359 ;
  assign n34361 = x619 & ~n34078 ;
  assign n34362 = x1159 | n34361 ;
  assign n34363 = ( n34353 & n34356 ) | ( n34353 & ~n34362 ) | ( n34356 & ~n34362 ) ;
  assign n34364 = ( x648 & n33952 ) | ( x648 & ~n34363 ) | ( n33952 & ~n34363 ) ;
  assign n34365 = n34363 | n34364 ;
  assign n34366 = ( x789 & n34360 ) | ( x789 & n34365 ) | ( n34360 & n34365 ) ;
  assign n34367 = ~n34360 & n34366 ;
  assign n34368 = x788 & n34108 ;
  assign n34369 = ( ~n34354 & n34367 ) | ( ~n34354 & n34368 ) | ( n34367 & n34368 ) ;
  assign n34370 = n34354 | n34369 ;
  assign n34371 = ( n18482 & ~n34109 ) | ( n18482 & n34370 ) | ( ~n34109 & n34370 ) ;
  assign n34372 = ~n18482 & n34371 ;
  assign n34373 = x628 | n34082 ;
  assign n34374 = x628 | n33809 ;
  assign n34375 = x628 & ~n34082 ;
  assign n34376 = n16337 & ~n34375 ;
  assign n34377 = n34374 & n34376 ;
  assign n34378 = x628 & ~n33809 ;
  assign n34379 = n16338 & ~n34378 ;
  assign n34380 = n34377 ^ n34373 ^ 1'b0 ;
  assign n34381 = ( ~n34373 & n34379 ) | ( ~n34373 & n34380 ) | ( n34379 & n34380 ) ;
  assign n34382 = ( n34373 & n34377 ) | ( n34373 & n34381 ) | ( n34377 & n34381 ) ;
  assign n34383 = n34382 ^ n19046 ^ 1'b0 ;
  assign n34384 = ( ~n19046 & n33960 ) | ( ~n19046 & n34383 ) | ( n33960 & n34383 ) ;
  assign n34385 = ( n19046 & n34382 ) | ( n19046 & n34384 ) | ( n34382 & n34384 ) ;
  assign n34386 = n34372 ^ x792 ^ 1'b0 ;
  assign n34387 = ( ~x792 & n34385 ) | ( ~x792 & n34386 ) | ( n34385 & n34386 ) ;
  assign n34388 = ( x792 & n34372 ) | ( x792 & n34387 ) | ( n34372 & n34387 ) ;
  assign n34389 = ( ~n18484 & n34096 ) | ( ~n18484 & n34388 ) | ( n34096 & n34388 ) ;
  assign n34390 = n34096 ^ n18484 ^ 1'b0 ;
  assign n34391 = ( n34096 & n34389 ) | ( n34096 & ~n34390 ) | ( n34389 & ~n34390 ) ;
  assign n34392 = x644 & ~n34391 ;
  assign n34393 = n34089 | n34092 ;
  assign n34394 = n34085 ^ x787 ^ 1'b0 ;
  assign n34395 = ( n34085 & n34393 ) | ( n34085 & n34394 ) | ( n34393 & n34394 ) ;
  assign n34396 = x644 | n34395 ;
  assign n34397 = ( x715 & n34392 ) | ( x715 & n34396 ) | ( n34392 & n34396 ) ;
  assign n34398 = ~n34392 & n34397 ;
  assign n34399 = x644 | n33809 ;
  assign n34400 = n33809 ^ n16376 ^ 1'b0 ;
  assign n34401 = ( n33809 & n33962 ) | ( n33809 & ~n34400 ) | ( n33962 & ~n34400 ) ;
  assign n34402 = x644 & ~n34401 ;
  assign n34403 = ( x715 & n34399 ) | ( x715 & ~n34402 ) | ( n34399 & ~n34402 ) ;
  assign n34404 = ~x715 & n34403 ;
  assign n34405 = ( x1160 & n34398 ) | ( x1160 & ~n34404 ) | ( n34398 & ~n34404 ) ;
  assign n34406 = ~n34398 & n34405 ;
  assign n34407 = x644 & ~n33809 ;
  assign n34408 = x715 & ~n34407 ;
  assign n34409 = n34408 ^ x1160 ^ 1'b0 ;
  assign n34410 = x644 | n34401 ;
  assign n34411 = ( n34408 & ~n34409 ) | ( n34408 & n34410 ) | ( ~n34409 & n34410 ) ;
  assign n34412 = ( x1160 & n34409 ) | ( x1160 & n34411 ) | ( n34409 & n34411 ) ;
  assign n34413 = x644 & ~n34395 ;
  assign n34414 = x715 | n34413 ;
  assign n34415 = ( n34391 & n34392 ) | ( n34391 & ~n34414 ) | ( n34392 & ~n34414 ) ;
  assign n34416 = ( ~n34406 & n34412 ) | ( ~n34406 & n34415 ) | ( n34412 & n34415 ) ;
  assign n34417 = ~n34406 & n34416 ;
  assign n34418 = n34391 ^ x790 ^ 1'b0 ;
  assign n34419 = ( n34391 & n34417 ) | ( n34391 & n34418 ) | ( n34417 & n34418 ) ;
  assign n34420 = n34419 ^ n7318 ^ 1'b0 ;
  assign n34421 = ( x222 & n34419 ) | ( x222 & n34420 ) | ( n34419 & n34420 ) ;
  assign n34422 = x299 | n15482 ;
  assign n34423 = n33805 & n34422 ;
  assign n34424 = ( n15102 & n15487 ) | ( n15102 & ~n34423 ) | ( n15487 & ~n34423 ) ;
  assign n34425 = n34423 | n34424 ;
  assign n34426 = n34425 ^ n17328 ^ 1'b0 ;
  assign n34427 = ( x223 & n17328 ) | ( x223 & ~n34425 ) | ( n17328 & ~n34425 ) ;
  assign n34428 = ( x223 & ~n34426 ) | ( x223 & n34427 ) | ( ~n34426 & n34427 ) ;
  assign n34429 = x626 & n34428 ;
  assign n34430 = x642 & n15524 ;
  assign n34431 = n33406 & ~n34430 ;
  assign n34432 = x642 & ~n15525 ;
  assign n34433 = n33858 & ~n34432 ;
  assign n34434 = n34431 | n34433 ;
  assign n34435 = x681 & ~n34434 ;
  assign n34436 = ~n5077 & n34434 ;
  assign n34437 = n15340 & ~n34430 ;
  assign n34438 = n5077 & n34437 ;
  assign n34439 = n15357 & n34438 ;
  assign n34440 = ( x681 & ~n34436 ) | ( x681 & n34439 ) | ( ~n34436 & n34439 ) ;
  assign n34441 = n34436 | n34440 ;
  assign n34442 = ~n34435 & n34441 ;
  assign n34443 = ~n5114 & n34442 ;
  assign n34444 = x642 & ~n15547 ;
  assign n34445 = ( n5077 & n15351 ) | ( n5077 & n34444 ) | ( n15351 & n34444 ) ;
  assign n34446 = ~n34444 & n34445 ;
  assign n34447 = x681 | n34446 ;
  assign n34448 = n15361 ^ x642 ^ 1'b0 ;
  assign n34449 = ( n15361 & n15548 ) | ( n15361 & n34448 ) | ( n15548 & n34448 ) ;
  assign n34450 = ~n5077 & n34449 ;
  assign n34451 = n34447 | n34450 ;
  assign n34452 = x681 & ~n34449 ;
  assign n34453 = n34451 & ~n34452 ;
  assign n34454 = n5114 & n34453 ;
  assign n34455 = ( x223 & n34443 ) | ( x223 & ~n34454 ) | ( n34443 & ~n34454 ) ;
  assign n34456 = ~n34443 & n34455 ;
  assign n34457 = x642 & n15595 ;
  assign n34458 = n1359 | n34457 ;
  assign n34459 = n15427 & n34430 ;
  assign n34460 = x681 & ~n34459 ;
  assign n34461 = x642 & n5077 ;
  assign n34462 = n15845 & n34461 ;
  assign n34463 = ~n5077 & n34459 ;
  assign n34464 = ( x681 & ~n34462 ) | ( x681 & n34463 ) | ( ~n34462 & n34463 ) ;
  assign n34465 = n34462 | n34464 ;
  assign n34466 = ~n34460 & n34465 ;
  assign n34467 = n5114 & n34466 ;
  assign n34468 = ~n5077 & n34457 ;
  assign n34469 = x681 | n34468 ;
  assign n34470 = n15594 & n34461 ;
  assign n34471 = n34469 | n34470 ;
  assign n34472 = x681 & ~n34457 ;
  assign n34473 = n34471 & ~n34472 ;
  assign n34474 = ~n5114 & n34473 ;
  assign n34475 = ( n1359 & n34467 ) | ( n1359 & ~n34474 ) | ( n34467 & ~n34474 ) ;
  assign n34476 = ~n34467 & n34475 ;
  assign n34477 = ( x223 & n34458 ) | ( x223 & ~n34476 ) | ( n34458 & ~n34476 ) ;
  assign n34478 = ~x223 & n34477 ;
  assign n34479 = ( x299 & ~n34456 ) | ( x299 & n34478 ) | ( ~n34456 & n34478 ) ;
  assign n34480 = n34456 | n34479 ;
  assign n34481 = ~n5061 & n34442 ;
  assign n34482 = n5061 & n34453 ;
  assign n34483 = ( x223 & n34481 ) | ( x223 & ~n34482 ) | ( n34481 & ~n34482 ) ;
  assign n34484 = ~n34481 & n34483 ;
  assign n34485 = n15607 & n34461 ;
  assign n34486 = n34469 | n34485 ;
  assign n34487 = n15353 | n34447 ;
  assign n34488 = n34486 & n34487 ;
  assign n34489 = x642 & n15609 ;
  assign n34490 = x681 & ~n34489 ;
  assign n34491 = n34488 & ~n34490 ;
  assign n34492 = n19292 & n34491 ;
  assign n34493 = ~n5061 & n34486 ;
  assign n34494 = n34457 & n34493 ;
  assign n34495 = ( x947 & ~n34492 ) | ( x947 & n34494 ) | ( ~n34492 & n34494 ) ;
  assign n34496 = n34492 | n34495 ;
  assign n34497 = x947 & ~n34491 ;
  assign n34498 = ( x223 & n34496 ) | ( x223 & ~n34497 ) | ( n34496 & ~n34497 ) ;
  assign n34499 = ~x223 & n34498 ;
  assign n34500 = ( x215 & n34484 ) | ( x215 & n34499 ) | ( n34484 & n34499 ) ;
  assign n34501 = n34499 ^ n34484 ^ 1'b0 ;
  assign n34502 = ( x215 & n34500 ) | ( x215 & n34501 ) | ( n34500 & n34501 ) ;
  assign n34503 = n19292 & n34466 ;
  assign n34504 = ~n19292 & n34473 ;
  assign n34505 = ( x947 & ~n34503 ) | ( x947 & n34504 ) | ( ~n34503 & n34504 ) ;
  assign n34506 = n34503 | n34505 ;
  assign n34507 = x947 & ~n34466 ;
  assign n34508 = ( x223 & n34506 ) | ( x223 & ~n34507 ) | ( n34506 & ~n34507 ) ;
  assign n34509 = ~x223 & n34508 ;
  assign n34510 = x642 | n15446 ;
  assign n34511 = n5080 | n34432 ;
  assign n34512 = n34510 & ~n34511 ;
  assign n34513 = n34431 | n34512 ;
  assign n34514 = x681 & ~n34513 ;
  assign n34515 = ~n5077 & n34513 ;
  assign n34516 = n15538 | n33403 ;
  assign n34517 = n5077 & n34516 ;
  assign n34518 = x681 | n34517 ;
  assign n34519 = ( ~n5061 & n34515 ) | ( ~n5061 & n34518 ) | ( n34515 & n34518 ) ;
  assign n34520 = ~n5061 & n34519 ;
  assign n34521 = ~n34514 & n34520 ;
  assign n34522 = n15429 ^ x642 ^ 1'b0 ;
  assign n34523 = ( n15429 & n15516 ) | ( n15429 & n34522 ) | ( n15516 & n34522 ) ;
  assign n34524 = x681 & ~n34523 ;
  assign n34525 = n5077 & n15425 ;
  assign n34526 = ~n34430 & n34525 ;
  assign n34527 = x681 | n34526 ;
  assign n34528 = ~n5077 & n34523 ;
  assign n34529 = ( n5061 & n34527 ) | ( n5061 & n34528 ) | ( n34527 & n34528 ) ;
  assign n34530 = n34528 ^ n34527 ^ 1'b0 ;
  assign n34531 = ( n5061 & n34529 ) | ( n5061 & n34530 ) | ( n34529 & n34530 ) ;
  assign n34532 = ~n34524 & n34531 ;
  assign n34533 = ( x223 & n34521 ) | ( x223 & ~n34532 ) | ( n34521 & ~n34532 ) ;
  assign n34534 = ~n34521 & n34533 ;
  assign n34535 = ( n2263 & n34509 ) | ( n2263 & ~n34534 ) | ( n34509 & ~n34534 ) ;
  assign n34536 = ~n34509 & n34535 ;
  assign n34537 = x223 & ~n15337 ;
  assign n34538 = n2263 | n34537 ;
  assign n34539 = n34457 | n34538 ;
  assign n34540 = ( x215 & ~n34536 ) | ( x215 & n34539 ) | ( ~n34536 & n34539 ) ;
  assign n34541 = ~x215 & n34540 ;
  assign n34542 = ( x299 & n34502 ) | ( x299 & ~n34541 ) | ( n34502 & ~n34541 ) ;
  assign n34543 = ~n34502 & n34542 ;
  assign n34544 = x39 & ~n34543 ;
  assign n34545 = n34480 & n34544 ;
  assign n34546 = ~x223 & x642 ;
  assign n34547 = n15636 & n34546 ;
  assign n34548 = x299 & ~n34547 ;
  assign n34549 = n5079 & n15635 ;
  assign n34550 = x223 & ~n15495 ;
  assign n34551 = ~n34549 & n34550 ;
  assign n34552 = ( x39 & n34548 ) | ( x39 & ~n34551 ) | ( n34548 & ~n34551 ) ;
  assign n34553 = n34552 ^ n34548 ^ 1'b0 ;
  assign n34554 = ( x39 & n34552 ) | ( x39 & ~n34553 ) | ( n34552 & ~n34553 ) ;
  assign n34555 = n15633 & n34546 ;
  assign n34556 = x299 | n34555 ;
  assign n34557 = ~x642 & n15633 ;
  assign n34558 = x223 & ~n34557 ;
  assign n34559 = ~n15507 & n34558 ;
  assign n34560 = ( ~n34554 & n34556 ) | ( ~n34554 & n34559 ) | ( n34556 & n34559 ) ;
  assign n34561 = ~n34554 & n34560 ;
  assign n34562 = ( x38 & ~n34545 ) | ( x38 & n34561 ) | ( ~n34545 & n34561 ) ;
  assign n34563 = n34545 | n34562 ;
  assign n34564 = x39 & x223 ;
  assign n34565 = x38 & ~n34564 ;
  assign n34566 = ( ~x39 & x223 ) | ( ~x39 & n15644 ) | ( x223 & n15644 ) ;
  assign n34567 = ~n34437 & n34566 ;
  assign n34568 = n34565 & ~n34567 ;
  assign n34569 = ( n2069 & n34563 ) | ( n2069 & ~n34568 ) | ( n34563 & ~n34568 ) ;
  assign n34570 = ~n2069 & n34569 ;
  assign n34571 = n34570 ^ x223 ^ 1'b0 ;
  assign n34572 = ( ~x223 & n2069 ) | ( ~x223 & n34571 ) | ( n2069 & n34571 ) ;
  assign n34573 = ( x223 & n34570 ) | ( x223 & n34572 ) | ( n34570 & n34572 ) ;
  assign n34574 = n34428 ^ n15659 ^ 1'b0 ;
  assign n34575 = ( n34428 & n34573 ) | ( n34428 & ~n34574 ) | ( n34573 & ~n34574 ) ;
  assign n34576 = x609 & ~n34575 ;
  assign n34577 = x609 | n34428 ;
  assign n34578 = ( x1155 & n34576 ) | ( x1155 & n34577 ) | ( n34576 & n34577 ) ;
  assign n34579 = ~n34576 & n34578 ;
  assign n34580 = x609 & ~n34428 ;
  assign n34581 = x1155 | n34580 ;
  assign n34582 = ( n34575 & n34576 ) | ( n34575 & ~n34581 ) | ( n34576 & ~n34581 ) ;
  assign n34583 = n34579 | n34582 ;
  assign n34584 = n34575 ^ x785 ^ 1'b0 ;
  assign n34585 = ( n34575 & n34583 ) | ( n34575 & n34584 ) | ( n34583 & n34584 ) ;
  assign n34586 = x618 & ~n34585 ;
  assign n34587 = x618 | n34428 ;
  assign n34588 = ( x1154 & n34586 ) | ( x1154 & n34587 ) | ( n34586 & n34587 ) ;
  assign n34589 = ~n34586 & n34588 ;
  assign n34590 = x618 & ~n34428 ;
  assign n34591 = x1154 | n34590 ;
  assign n34592 = ( n34585 & n34586 ) | ( n34585 & ~n34591 ) | ( n34586 & ~n34591 ) ;
  assign n34593 = n34589 | n34592 ;
  assign n34594 = n34585 ^ x781 ^ 1'b0 ;
  assign n34595 = ( n34585 & n34593 ) | ( n34585 & n34594 ) | ( n34593 & n34594 ) ;
  assign n34596 = x619 & ~n34595 ;
  assign n34597 = x619 | n34428 ;
  assign n34598 = ( x1159 & n34596 ) | ( x1159 & n34597 ) | ( n34596 & n34597 ) ;
  assign n34599 = ~n34596 & n34598 ;
  assign n34600 = x619 & ~n34428 ;
  assign n34601 = x1159 | n34600 ;
  assign n34602 = ( n34595 & n34596 ) | ( n34595 & ~n34601 ) | ( n34596 & ~n34601 ) ;
  assign n34603 = n34599 | n34602 ;
  assign n34604 = n34595 ^ x789 ^ 1'b0 ;
  assign n34605 = ( n34595 & n34603 ) | ( n34595 & n34604 ) | ( n34603 & n34604 ) ;
  assign n34606 = ~x626 & n34605 ;
  assign n34607 = ( n22322 & n34429 ) | ( n22322 & ~n34606 ) | ( n34429 & ~n34606 ) ;
  assign n34608 = ~n34429 & n34607 ;
  assign n34609 = x626 & n34605 ;
  assign n34610 = ~x626 & n34428 ;
  assign n34611 = ( n22317 & n34609 ) | ( n22317 & ~n34610 ) | ( n34609 & ~n34610 ) ;
  assign n34612 = ~n34609 & n34611 ;
  assign n34613 = x223 & n16038 ;
  assign n34614 = x299 | n34613 ;
  assign n34615 = x680 & x681 ;
  assign n34616 = ~n34614 & n34615 ;
  assign n34617 = ( n16018 & n34614 ) | ( n16018 & ~n34616 ) | ( n34614 & ~n34616 ) ;
  assign n34618 = ( x223 & n16018 ) | ( x223 & ~n34617 ) | ( n16018 & ~n34617 ) ;
  assign n34619 = ~n34617 & n34618 ;
  assign n34620 = x223 & n16033 ;
  assign n34621 = n16024 & ~n34615 ;
  assign n34622 = ( x299 & n34620 ) | ( x299 & ~n34621 ) | ( n34620 & ~n34621 ) ;
  assign n34623 = ~n34620 & n34622 ;
  assign n34624 = n16024 ^ x223 ^ 1'b0 ;
  assign n34625 = ( x223 & n16024 ) | ( x223 & ~n34624 ) | ( n16024 & ~n34624 ) ;
  assign n34626 = ( n34623 & n34624 ) | ( n34623 & n34625 ) | ( n34624 & n34625 ) ;
  assign n34627 = ( x39 & ~n34619 ) | ( x39 & n34626 ) | ( ~n34619 & n34626 ) ;
  assign n34628 = n34619 | n34627 ;
  assign n34629 = ~x223 & x681 ;
  assign n34630 = n16172 & n34629 ;
  assign n34631 = x681 & ~n16100 ;
  assign n34632 = n15377 & ~n34631 ;
  assign n34633 = n5061 & n34632 ;
  assign n34634 = x681 & ~n33966 ;
  assign n34635 = n15400 & ~n34634 ;
  assign n34636 = ~n5061 & n34635 ;
  assign n34637 = ( x223 & n34633 ) | ( x223 & ~n34636 ) | ( n34633 & ~n34636 ) ;
  assign n34638 = ~n34633 & n34637 ;
  assign n34639 = ( x215 & n34630 ) | ( x215 & ~n34638 ) | ( n34630 & ~n34638 ) ;
  assign n34640 = ~n34630 & n34639 ;
  assign n34641 = x681 & n16164 ;
  assign n34642 = n34538 | n34641 ;
  assign n34643 = ~n5061 & n15462 ;
  assign n34644 = x681 & ~n16119 ;
  assign n34645 = n34643 & ~n34644 ;
  assign n34646 = x681 & ~n33993 ;
  assign n34647 = ~n5077 & n15429 ;
  assign n34648 = ( x681 & n34525 ) | ( x681 & ~n34647 ) | ( n34525 & ~n34647 ) ;
  assign n34649 = n34647 | n34648 ;
  assign n34650 = n5061 & n34649 ;
  assign n34651 = ~n34646 & n34650 ;
  assign n34652 = ( x223 & n34645 ) | ( x223 & ~n34651 ) | ( n34645 & ~n34651 ) ;
  assign n34653 = ~n34645 & n34652 ;
  assign n34654 = n16146 & n34615 ;
  assign n34655 = n5061 | n34654 ;
  assign n34656 = x681 & n16152 ;
  assign n34657 = n5061 & ~n34656 ;
  assign n34658 = ( x223 & n34655 ) | ( x223 & ~n34657 ) | ( n34655 & ~n34657 ) ;
  assign n34659 = ~x223 & n34658 ;
  assign n34660 = ( n2263 & n34653 ) | ( n2263 & ~n34659 ) | ( n34653 & ~n34659 ) ;
  assign n34661 = ~n34653 & n34660 ;
  assign n34662 = ( x215 & n34642 ) | ( x215 & ~n34661 ) | ( n34642 & ~n34661 ) ;
  assign n34663 = n34662 ^ n34642 ^ 1'b0 ;
  assign n34664 = ( x215 & n34662 ) | ( x215 & ~n34663 ) | ( n34662 & ~n34663 ) ;
  assign n34665 = ( x299 & n34640 ) | ( x299 & n34664 ) | ( n34640 & n34664 ) ;
  assign n34666 = ~n34640 & n34665 ;
  assign n34667 = n5114 & ~n34632 ;
  assign n34668 = n5114 | n34635 ;
  assign n34669 = x223 & n34668 ;
  assign n34670 = n34669 ^ n34667 ^ 1'b0 ;
  assign n34671 = ( n34667 & n34669 ) | ( n34667 & n34670 ) | ( n34669 & n34670 ) ;
  assign n34672 = ( x299 & ~n34667 ) | ( x299 & n34671 ) | ( ~n34667 & n34671 ) ;
  assign n34673 = n5114 & n34656 ;
  assign n34674 = ~n5114 & n34654 ;
  assign n34675 = ( n1359 & n34673 ) | ( n1359 & ~n34674 ) | ( n34673 & ~n34674 ) ;
  assign n34676 = ~n34673 & n34675 ;
  assign n34677 = ( n1359 & n34641 ) | ( n1359 & ~n34676 ) | ( n34641 & ~n34676 ) ;
  assign n34678 = ~n34676 & n34677 ;
  assign n34679 = ( x223 & ~n34672 ) | ( x223 & n34678 ) | ( ~n34672 & n34678 ) ;
  assign n34680 = ~n34672 & n34679 ;
  assign n34681 = ( x39 & n34666 ) | ( x39 & ~n34680 ) | ( n34666 & ~n34680 ) ;
  assign n34682 = ~n34666 & n34681 ;
  assign n34683 = ( x38 & n34628 ) | ( x38 & ~n34682 ) | ( n34628 & ~n34682 ) ;
  assign n34684 = n34683 ^ n34628 ^ 1'b0 ;
  assign n34685 = ( x38 & n34683 ) | ( x38 & ~n34684 ) | ( n34683 & ~n34684 ) ;
  assign n34686 = x223 & ~n15644 ;
  assign n34687 = ( x38 & ~x681 ) | ( x38 & n16185 ) | ( ~x681 & n16185 ) ;
  assign n34688 = ~n34686 & n34687 ;
  assign n34689 = ( n2069 & n34685 ) | ( n2069 & ~n34688 ) | ( n34685 & ~n34688 ) ;
  assign n34690 = ~n2069 & n34689 ;
  assign n34691 = n34690 ^ x223 ^ 1'b0 ;
  assign n34692 = ( ~x223 & n2069 ) | ( ~x223 & n34691 ) | ( n2069 & n34691 ) ;
  assign n34693 = ( x223 & n34690 ) | ( x223 & n34692 ) | ( n34690 & n34692 ) ;
  assign n34694 = x625 & ~n34693 ;
  assign n34695 = x625 | n34428 ;
  assign n34696 = ( x1153 & n34694 ) | ( x1153 & n34695 ) | ( n34694 & n34695 ) ;
  assign n34697 = ~n34694 & n34696 ;
  assign n34698 = x625 & ~n34428 ;
  assign n34699 = x1153 | n34698 ;
  assign n34700 = ( n34693 & n34694 ) | ( n34693 & ~n34699 ) | ( n34694 & ~n34699 ) ;
  assign n34701 = n34697 | n34700 ;
  assign n34702 = n34693 ^ x778 ^ 1'b0 ;
  assign n34703 = ( n34693 & n34701 ) | ( n34693 & n34702 ) | ( n34701 & n34702 ) ;
  assign n34704 = n34428 ^ n16234 ^ 1'b0 ;
  assign n34705 = ( n34428 & n34703 ) | ( n34428 & ~n34704 ) | ( n34703 & ~n34704 ) ;
  assign n34706 = n34428 ^ n16254 ^ 1'b0 ;
  assign n34707 = ( n34428 & n34705 ) | ( n34428 & ~n34706 ) | ( n34705 & ~n34706 ) ;
  assign n34708 = n16279 | n34707 ;
  assign n34709 = n16279 & ~n34428 ;
  assign n34710 = n34708 & ~n34709 ;
  assign n34711 = ~n34612 & n34710 ;
  assign n34712 = ( n16459 & n34612 ) | ( n16459 & ~n34711 ) | ( n34612 & ~n34711 ) ;
  assign n34713 = ( x788 & n34608 ) | ( x788 & n34712 ) | ( n34608 & n34712 ) ;
  assign n34714 = n34712 ^ n34608 ^ 1'b0 ;
  assign n34715 = ( x788 & n34713 ) | ( x788 & n34714 ) | ( n34713 & n34714 ) ;
  assign n34716 = n15340 & n15890 ;
  assign n34717 = ~x642 & n15690 ;
  assign n34718 = n34615 & ~n34717 ;
  assign n34719 = ~n34716 & n34718 ;
  assign n34720 = n34615 & ~n34719 ;
  assign n34721 = ( n34430 & n34719 ) | ( n34430 & ~n34720 ) | ( n34719 & ~n34720 ) ;
  assign n34722 = n15690 ^ x642 ^ 1'b0 ;
  assign n34723 = ( n15690 & n15890 ) | ( n15690 & n34722 ) | ( n15890 & n34722 ) ;
  assign n34724 = ( n1292 & n1611 ) | ( n1292 & n34723 ) | ( n1611 & n34723 ) ;
  assign n34725 = ~n1292 & n34724 ;
  assign n34726 = n34615 & n34725 ;
  assign n34727 = n34437 & ~n34615 ;
  assign n34728 = ( x223 & n34726 ) | ( x223 & ~n34727 ) | ( n34726 & ~n34727 ) ;
  assign n34729 = ~n34726 & n34728 ;
  assign n34730 = n34721 | n34729 ;
  assign n34731 = n34565 & ~n34730 ;
  assign n34732 = ( n34565 & ~n34566 ) | ( n34565 & n34731 ) | ( ~n34566 & n34731 ) ;
  assign n34733 = x223 & ~n34549 ;
  assign n34734 = n16026 & ~n34615 ;
  assign n34735 = ( n34117 & n34733 ) | ( n34117 & ~n34734 ) | ( n34733 & ~n34734 ) ;
  assign n34736 = ~n34117 & n34735 ;
  assign n34737 = n16027 & n34629 ;
  assign n34738 = ( n34548 & n34736 ) | ( n34548 & ~n34737 ) | ( n34736 & ~n34737 ) ;
  assign n34739 = ~n34736 & n34738 ;
  assign n34740 = n16021 & n34629 ;
  assign n34741 = ~n34133 & n34558 ;
  assign n34742 = n16020 & ~n34615 ;
  assign n34743 = n34741 & ~n34742 ;
  assign n34744 = ( n34556 & ~n34740 ) | ( n34556 & n34743 ) | ( ~n34740 & n34743 ) ;
  assign n34745 = n34740 | n34744 ;
  assign n34746 = ( x39 & ~n34739 ) | ( x39 & n34745 ) | ( ~n34739 & n34745 ) ;
  assign n34747 = ~x39 & n34746 ;
  assign n34748 = n15337 & n34721 ;
  assign n34749 = ~x223 & n34748 ;
  assign n34750 = n34538 | n34729 ;
  assign n34751 = n34749 | n34750 ;
  assign n34752 = x642 & ~n15954 ;
  assign n34753 = n15690 & ~n34752 ;
  assign n34754 = x680 & ~n33406 ;
  assign n34755 = ( x680 & n34753 ) | ( x680 & n34754 ) | ( n34753 & n34754 ) ;
  assign n34756 = x642 & ~n15891 ;
  assign n34757 = n5080 | n34756 ;
  assign n34758 = x642 | n15700 ;
  assign n34759 = ~n34757 & n34758 ;
  assign n34760 = n34755 & ~n34759 ;
  assign n34761 = x680 | n34457 ;
  assign n34762 = x681 & ~n34761 ;
  assign n34763 = ( x681 & n34760 ) | ( x681 & n34762 ) | ( n34760 & n34762 ) ;
  assign n34764 = ( n34469 & n34470 ) | ( n34469 & ~n34763 ) | ( n34470 & ~n34763 ) ;
  assign n34765 = ~n34763 & n34764 ;
  assign n34766 = n5061 | n34765 ;
  assign n34767 = x642 & ~n15905 ;
  assign n34768 = x680 & ~n34767 ;
  assign n34769 = ~x642 & n5080 ;
  assign n34770 = ( n15738 & n15739 ) | ( n15738 & ~n34769 ) | ( n15739 & ~n34769 ) ;
  assign n34771 = n34768 & n34770 ;
  assign n34772 = n34460 | n34615 ;
  assign n34773 = n34465 & ~n34772 ;
  assign n34774 = ( n34465 & n34771 ) | ( n34465 & n34773 ) | ( n34771 & n34773 ) ;
  assign n34775 = n5061 & ~n34774 ;
  assign n34776 = ( x223 & n34766 ) | ( x223 & ~n34775 ) | ( n34766 & ~n34775 ) ;
  assign n34777 = ~x223 & n34776 ;
  assign n34778 = ~n15335 & n34725 ;
  assign n34779 = x680 & ~n5080 ;
  assign n34780 = ( x680 & n34778 ) | ( x680 & n34779 ) | ( n34778 & n34779 ) ;
  assign n34781 = ( x642 & n34510 ) | ( x642 & n34722 ) | ( n34510 & n34722 ) ;
  assign n34782 = ~n34752 & n34781 ;
  assign n34783 = n5080 | n34782 ;
  assign n34784 = n34780 & n34783 ;
  assign n34785 = n34514 | n34615 ;
  assign n34786 = n34520 & ~n34785 ;
  assign n34787 = ( n34520 & n34784 ) | ( n34520 & n34786 ) | ( n34784 & n34786 ) ;
  assign n34789 = ~n34223 & n34769 ;
  assign n34790 = n15527 | n34228 ;
  assign n34791 = x642 & ~n34233 ;
  assign n34792 = x680 & ~n34791 ;
  assign n34793 = ( n34789 & n34790 ) | ( n34789 & n34792 ) | ( n34790 & n34792 ) ;
  assign n34794 = ~n34789 & n34793 ;
  assign n34788 = n34524 | n34615 ;
  assign n34795 = n34794 ^ n34788 ^ 1'b0 ;
  assign n34796 = ( n34531 & ~n34788 ) | ( n34531 & n34794 ) | ( ~n34788 & n34794 ) ;
  assign n34797 = ( n34531 & ~n34795 ) | ( n34531 & n34796 ) | ( ~n34795 & n34796 ) ;
  assign n34798 = ( x223 & n34787 ) | ( x223 & ~n34797 ) | ( n34787 & ~n34797 ) ;
  assign n34799 = ~n34787 & n34798 ;
  assign n34800 = ( n2263 & n34777 ) | ( n2263 & ~n34799 ) | ( n34777 & ~n34799 ) ;
  assign n34801 = ~n34777 & n34800 ;
  assign n34802 = ( x215 & n34751 ) | ( x215 & ~n34801 ) | ( n34751 & ~n34801 ) ;
  assign n34803 = ~x215 & n34802 ;
  assign n34804 = n15759 & ~n34757 ;
  assign n34805 = n34755 & ~n34804 ;
  assign n34806 = ( x681 & n34762 ) | ( x681 & n34805 ) | ( n34762 & n34805 ) ;
  assign n34807 = ( n5061 & n34486 ) | ( n5061 & ~n34806 ) | ( n34486 & ~n34806 ) ;
  assign n34808 = ~n5061 & n34807 ;
  assign n34809 = x642 & ~n34146 ;
  assign n34810 = n15758 & n15880 ;
  assign n34811 = n15527 | n34810 ;
  assign n34812 = ~n15756 & n34769 ;
  assign n34813 = x680 & ~n34812 ;
  assign n34814 = ( n34809 & n34811 ) | ( n34809 & n34813 ) | ( n34811 & n34813 ) ;
  assign n34815 = ~n34809 & n34814 ;
  assign n34816 = ( n34490 & n34615 ) | ( n34490 & ~n34815 ) | ( n34615 & ~n34815 ) ;
  assign n34817 = ~n34815 & n34816 ;
  assign n34818 = ( n5061 & n34488 ) | ( n5061 & n34817 ) | ( n34488 & n34817 ) ;
  assign n34819 = ~n34817 & n34818 ;
  assign n34820 = ( x223 & ~n34808 ) | ( x223 & n34819 ) | ( ~n34808 & n34819 ) ;
  assign n34821 = n34808 | n34820 ;
  assign n34822 = ~x680 & n34449 ;
  assign n34823 = n5080 & ~n15803 ;
  assign n34824 = n15527 | n15801 ;
  assign n34825 = x680 & n34824 ;
  assign n34826 = x642 & ~n34167 ;
  assign n34827 = ( n34823 & n34825 ) | ( n34823 & ~n34826 ) | ( n34825 & ~n34826 ) ;
  assign n34828 = ~n34823 & n34827 ;
  assign n34829 = ( x681 & n34822 ) | ( x681 & ~n34828 ) | ( n34822 & ~n34828 ) ;
  assign n34830 = ~n34822 & n34829 ;
  assign n34831 = ( n34447 & n34450 ) | ( n34447 & ~n34830 ) | ( n34450 & ~n34830 ) ;
  assign n34832 = ~n34830 & n34831 ;
  assign n34833 = n5061 & ~n34832 ;
  assign n34834 = x223 & ~n34833 ;
  assign n34835 = x614 | n15824 ;
  assign n34836 = ~n34752 & n34835 ;
  assign n34837 = ( x616 & n34780 ) | ( x616 & n34836 ) | ( n34780 & n34836 ) ;
  assign n34838 = n34780 & n34837 ;
  assign n34839 = n34435 | n34615 ;
  assign n34840 = n34441 & ~n34839 ;
  assign n34841 = ( n34441 & n34838 ) | ( n34441 & n34840 ) | ( n34838 & n34840 ) ;
  assign n34842 = n5061 | n34841 ;
  assign n34843 = n34834 & n34842 ;
  assign n34844 = x215 & ~n34843 ;
  assign n34845 = n34821 & n34844 ;
  assign n34846 = ( x299 & n34803 ) | ( x299 & ~n34845 ) | ( n34803 & ~n34845 ) ;
  assign n34847 = ~n34803 & n34846 ;
  assign n34848 = ~n5114 & n34841 ;
  assign n34849 = n5114 & n34832 ;
  assign n34850 = ( x223 & n34848 ) | ( x223 & ~n34849 ) | ( n34848 & ~n34849 ) ;
  assign n34851 = ~n34848 & n34850 ;
  assign n34852 = n1359 | n34748 ;
  assign n34853 = ~n5114 & n34765 ;
  assign n34854 = n5114 & n34774 ;
  assign n34855 = ( n1359 & n34853 ) | ( n1359 & ~n34854 ) | ( n34853 & ~n34854 ) ;
  assign n34856 = ~n34853 & n34855 ;
  assign n34857 = ( x223 & n34852 ) | ( x223 & ~n34856 ) | ( n34852 & ~n34856 ) ;
  assign n34858 = ~x223 & n34857 ;
  assign n34859 = ( x299 & ~n34851 ) | ( x299 & n34858 ) | ( ~n34851 & n34858 ) ;
  assign n34860 = n34851 | n34859 ;
  assign n34861 = ( x39 & n34847 ) | ( x39 & n34860 ) | ( n34847 & n34860 ) ;
  assign n34862 = ~n34847 & n34861 ;
  assign n34863 = ( x38 & ~n34747 ) | ( x38 & n34862 ) | ( ~n34747 & n34862 ) ;
  assign n34864 = n34747 | n34863 ;
  assign n34865 = ( n2069 & ~n34732 ) | ( n2069 & n34864 ) | ( ~n34732 & n34864 ) ;
  assign n34866 = ~n2069 & n34865 ;
  assign n34867 = n34866 ^ x223 ^ 1'b0 ;
  assign n34868 = ( ~x223 & n2069 ) | ( ~x223 & n34867 ) | ( n2069 & n34867 ) ;
  assign n34869 = ( x223 & n34866 ) | ( x223 & n34868 ) | ( n34866 & n34868 ) ;
  assign n34870 = x625 & ~n34869 ;
  assign n34871 = x625 | n34573 ;
  assign n34872 = ( x1153 & n34870 ) | ( x1153 & n34871 ) | ( n34870 & n34871 ) ;
  assign n34873 = ~n34870 & n34872 ;
  assign n34874 = ( x608 & n34700 ) | ( x608 & ~n34873 ) | ( n34700 & ~n34873 ) ;
  assign n34875 = ~n34700 & n34874 ;
  assign n34876 = x625 & ~n34573 ;
  assign n34877 = x1153 | n34876 ;
  assign n34878 = x625 | n34869 ;
  assign n34879 = n34878 ^ n34877 ^ 1'b0 ;
  assign n34880 = ( n34877 & n34878 ) | ( n34877 & n34879 ) | ( n34878 & n34879 ) ;
  assign n34881 = ( x608 & ~n34877 ) | ( x608 & n34880 ) | ( ~n34877 & n34880 ) ;
  assign n34882 = ( n34697 & ~n34875 ) | ( n34697 & n34881 ) | ( ~n34875 & n34881 ) ;
  assign n34883 = ~n34875 & n34882 ;
  assign n34884 = n34869 ^ x778 ^ 1'b0 ;
  assign n34885 = ( n34869 & n34883 ) | ( n34869 & n34884 ) | ( n34883 & n34884 ) ;
  assign n34886 = x609 & ~n34885 ;
  assign n34887 = x609 | n34703 ;
  assign n34888 = ( x1155 & n34886 ) | ( x1155 & n34887 ) | ( n34886 & n34887 ) ;
  assign n34889 = ~n34886 & n34888 ;
  assign n34890 = ( x660 & n34582 ) | ( x660 & ~n34889 ) | ( n34582 & ~n34889 ) ;
  assign n34891 = ~n34582 & n34890 ;
  assign n34892 = x609 & ~n34703 ;
  assign n34893 = x1155 | n34892 ;
  assign n34894 = ( x609 & n34885 ) | ( x609 & ~n34893 ) | ( n34885 & ~n34893 ) ;
  assign n34895 = ~n34893 & n34894 ;
  assign n34896 = x660 | n34579 ;
  assign n34897 = ( ~n34891 & n34895 ) | ( ~n34891 & n34896 ) | ( n34895 & n34896 ) ;
  assign n34898 = ~n34891 & n34897 ;
  assign n34899 = n34885 ^ x785 ^ 1'b0 ;
  assign n34900 = ( n34885 & n34898 ) | ( n34885 & n34899 ) | ( n34898 & n34899 ) ;
  assign n34901 = x618 & ~n34900 ;
  assign n34902 = x618 | n34705 ;
  assign n34903 = ( x1154 & n34901 ) | ( x1154 & n34902 ) | ( n34901 & n34902 ) ;
  assign n34904 = ~n34901 & n34903 ;
  assign n34905 = ( x627 & n34592 ) | ( x627 & ~n34904 ) | ( n34592 & ~n34904 ) ;
  assign n34906 = ~n34592 & n34905 ;
  assign n34907 = x627 | n34589 ;
  assign n34908 = x618 & ~n34705 ;
  assign n34909 = x1154 | n34908 ;
  assign n34910 = ( n34900 & n34901 ) | ( n34900 & ~n34909 ) | ( n34901 & ~n34909 ) ;
  assign n34911 = ( ~n34906 & n34907 ) | ( ~n34906 & n34910 ) | ( n34907 & n34910 ) ;
  assign n34912 = ~n34906 & n34911 ;
  assign n34913 = n34900 ^ x781 ^ 1'b0 ;
  assign n34914 = ( n34900 & n34912 ) | ( n34900 & n34913 ) | ( n34912 & n34913 ) ;
  assign n34915 = ~x789 & n34914 ;
  assign n34916 = n16519 | n34915 ;
  assign n34917 = x619 | n34914 ;
  assign n34918 = x619 & ~n34707 ;
  assign n34919 = ( x1159 & n34917 ) | ( x1159 & ~n34918 ) | ( n34917 & ~n34918 ) ;
  assign n34920 = ~x1159 & n34919 ;
  assign n34921 = ( x648 & n34599 ) | ( x648 & ~n34920 ) | ( n34599 & ~n34920 ) ;
  assign n34922 = n34920 | n34921 ;
  assign n34923 = x619 & ~n34914 ;
  assign n34924 = x619 | n34707 ;
  assign n34925 = ( x1159 & n34923 ) | ( x1159 & n34924 ) | ( n34923 & n34924 ) ;
  assign n34926 = ~n34923 & n34925 ;
  assign n34927 = ( x648 & n34602 ) | ( x648 & ~n34926 ) | ( n34602 & ~n34926 ) ;
  assign n34928 = ~n34602 & n34927 ;
  assign n34929 = x789 & ~n34928 ;
  assign n34930 = n34922 & n34929 ;
  assign n34931 = ( ~n34715 & n34916 ) | ( ~n34715 & n34930 ) | ( n34916 & n34930 ) ;
  assign n34932 = ~n34715 & n34931 ;
  assign n34933 = n16318 | n34708 ;
  assign n34934 = n17086 & ~n34428 ;
  assign n34935 = n34933 & ~n34934 ;
  assign n34936 = x628 | n34935 ;
  assign n34937 = x628 | n34428 ;
  assign n34938 = x628 & ~n34935 ;
  assign n34939 = n16337 & ~n34938 ;
  assign n34940 = n34937 & n34939 ;
  assign n34941 = x628 & ~n34428 ;
  assign n34942 = n16338 & ~n34941 ;
  assign n34943 = n34940 ^ n34936 ^ 1'b0 ;
  assign n34944 = ( ~n34936 & n34942 ) | ( ~n34936 & n34943 ) | ( n34942 & n34943 ) ;
  assign n34945 = ( n34936 & n34940 ) | ( n34936 & n34944 ) | ( n34940 & n34944 ) ;
  assign n34946 = n34428 ^ n16518 ^ 1'b0 ;
  assign n34947 = ( n34428 & n34605 ) | ( n34428 & ~n34946 ) | ( n34605 & ~n34946 ) ;
  assign n34948 = n34945 ^ n19046 ^ 1'b0 ;
  assign n34949 = ( ~n19046 & n34947 ) | ( ~n19046 & n34948 ) | ( n34947 & n34948 ) ;
  assign n34950 = ( n19046 & n34945 ) | ( n19046 & n34949 ) | ( n34945 & n34949 ) ;
  assign n34951 = n34932 ^ x792 ^ 1'b0 ;
  assign n34952 = ( ~x792 & n34950 ) | ( ~x792 & n34951 ) | ( n34950 & n34951 ) ;
  assign n34953 = ( x792 & n34932 ) | ( x792 & n34952 ) | ( n34932 & n34952 ) ;
  assign n34954 = n34428 ^ n16339 ^ 1'b0 ;
  assign n34955 = ( n34428 & n34947 ) | ( n34428 & ~n34954 ) | ( n34947 & ~n34954 ) ;
  assign n34956 = n19055 & n34955 ;
  assign n34957 = n17093 | n34935 ;
  assign n34958 = n16559 & ~n34428 ;
  assign n34959 = n34957 & ~n34958 ;
  assign n34960 = x647 & ~n34959 ;
  assign n34961 = x647 | n34428 ;
  assign n34962 = ( x1157 & n34960 ) | ( x1157 & n34961 ) | ( n34960 & n34961 ) ;
  assign n34963 = ~n34960 & n34962 ;
  assign n34964 = x647 & ~n34428 ;
  assign n34965 = x1157 | n34964 ;
  assign n34966 = ( n34959 & n34960 ) | ( n34959 & ~n34965 ) | ( n34960 & ~n34965 ) ;
  assign n34967 = ( n16375 & n34963 ) | ( n16375 & n34966 ) | ( n34963 & n34966 ) ;
  assign n34968 = ( x787 & n34956 ) | ( x787 & n34967 ) | ( n34956 & n34967 ) ;
  assign n34969 = n34967 ^ n34956 ^ 1'b0 ;
  assign n34970 = ( x787 & n34968 ) | ( x787 & n34969 ) | ( n34968 & n34969 ) ;
  assign n34971 = n18482 & ~n34950 ;
  assign n34972 = n18484 | n34971 ;
  assign n34973 = ~n34970 & n34972 ;
  assign n34974 = ( n34953 & n34970 ) | ( n34953 & ~n34973 ) | ( n34970 & ~n34973 ) ;
  assign n34975 = x644 & ~n34974 ;
  assign n34976 = n34963 | n34966 ;
  assign n34977 = n34959 ^ x787 ^ 1'b0 ;
  assign n34978 = ( n34959 & n34976 ) | ( n34959 & n34977 ) | ( n34976 & n34977 ) ;
  assign n34979 = x644 | n34978 ;
  assign n34980 = ( x715 & n34975 ) | ( x715 & n34979 ) | ( n34975 & n34979 ) ;
  assign n34981 = ~n34975 & n34980 ;
  assign n34982 = x644 | n34428 ;
  assign n34983 = n34428 ^ n16376 ^ 1'b0 ;
  assign n34984 = ( n34428 & n34955 ) | ( n34428 & ~n34983 ) | ( n34955 & ~n34983 ) ;
  assign n34985 = x644 & ~n34984 ;
  assign n34986 = ( x715 & n34982 ) | ( x715 & ~n34985 ) | ( n34982 & ~n34985 ) ;
  assign n34987 = ~x715 & n34986 ;
  assign n34988 = ( x1160 & n34981 ) | ( x1160 & ~n34987 ) | ( n34981 & ~n34987 ) ;
  assign n34989 = ~n34981 & n34988 ;
  assign n34990 = x644 & ~n34428 ;
  assign n34991 = x715 & ~n34990 ;
  assign n34992 = n34991 ^ x1160 ^ 1'b0 ;
  assign n34993 = x644 | n34984 ;
  assign n34994 = ( n34991 & ~n34992 ) | ( n34991 & n34993 ) | ( ~n34992 & n34993 ) ;
  assign n34995 = ( x1160 & n34992 ) | ( x1160 & n34994 ) | ( n34992 & n34994 ) ;
  assign n34996 = x644 & ~n34978 ;
  assign n34997 = x715 | n34996 ;
  assign n34998 = ( n34974 & n34975 ) | ( n34974 & ~n34997 ) | ( n34975 & ~n34997 ) ;
  assign n34999 = ( ~n34989 & n34995 ) | ( ~n34989 & n34998 ) | ( n34995 & n34998 ) ;
  assign n35000 = ~n34989 & n34999 ;
  assign n35001 = n34974 ^ x790 ^ 1'b0 ;
  assign n35002 = ( n34974 & n35000 ) | ( n34974 & n35001 ) | ( n35000 & n35001 ) ;
  assign n35003 = n35002 ^ n7318 ^ 1'b0 ;
  assign n35004 = ( x223 & n35002 ) | ( x223 & n35003 ) | ( n35002 & n35003 ) ;
  assign n35005 = x224 & ~n33808 ;
  assign n35006 = x224 & ~n15644 ;
  assign n35007 = x38 & ~n35006 ;
  assign n35008 = x614 & n15646 ;
  assign n35009 = n35007 & ~n35008 ;
  assign n35010 = x614 & n15636 ;
  assign n35011 = x224 & n15493 ;
  assign n35012 = n35010 & ~n35011 ;
  assign n35013 = n15330 & ~n35012 ;
  assign n35014 = ( x224 & n35012 ) | ( x224 & ~n35013 ) | ( n35012 & ~n35013 ) ;
  assign n35015 = x299 & ~n35014 ;
  assign n35016 = x614 & n15633 ;
  assign n35017 = ~x224 & n35016 ;
  assign n35018 = ~x614 & n15633 ;
  assign n35019 = x224 & ~n35018 ;
  assign n35020 = ~n15507 & n35019 ;
  assign n35021 = ( x299 & ~n35017 ) | ( x299 & n35020 ) | ( ~n35017 & n35020 ) ;
  assign n35022 = n35017 | n35021 ;
  assign n35023 = ( x39 & ~n35015 ) | ( x39 & n35022 ) | ( ~n35015 & n35022 ) ;
  assign n35024 = ~x39 & n35023 ;
  assign n35025 = x614 & n15845 ;
  assign n35026 = x680 & ~n35025 ;
  assign n35027 = x614 & n15524 ;
  assign n35028 = n15427 & n35027 ;
  assign n35029 = x680 | n35028 ;
  assign n35030 = ~n35026 & n35029 ;
  assign n35031 = n15383 | n35030 ;
  assign n35032 = n15383 & ~n35028 ;
  assign n35033 = n35031 & ~n35032 ;
  assign n35034 = n5061 & ~n35033 ;
  assign n35035 = x614 & n33849 ;
  assign n35036 = n5061 | n35035 ;
  assign n35037 = ( x224 & ~n35034 ) | ( x224 & n35036 ) | ( ~n35034 & n35036 ) ;
  assign n35038 = ~x224 & n35037 ;
  assign n35039 = n15337 & ~n35027 ;
  assign n35040 = n5081 | n35039 ;
  assign n35041 = n15465 & n35040 ;
  assign n35042 = x680 & n35027 ;
  assign n35043 = n15454 | n35042 ;
  assign n35044 = x680 | n35041 ;
  assign n35045 = ~n35043 & n35044 ;
  assign n35046 = n35041 ^ n15383 ^ 1'b0 ;
  assign n35047 = ( n35041 & n35045 ) | ( n35041 & ~n35046 ) | ( n35045 & ~n35046 ) ;
  assign n35048 = ~n5061 & n35047 ;
  assign n35049 = ~x614 & x616 ;
  assign n35050 = ~n15427 & n35049 ;
  assign n35051 = n5080 | n15426 ;
  assign n35052 = n5075 & n15447 ;
  assign n35053 = n35051 | n35052 ;
  assign n35054 = x614 & ~n15516 ;
  assign n35055 = ( n35050 & n35053 ) | ( n35050 & ~n35054 ) | ( n35053 & ~n35054 ) ;
  assign n35056 = ~n35050 & n35055 ;
  assign n35057 = x680 | n35056 ;
  assign n35058 = ~n15425 & n35026 ;
  assign n35059 = n35042 | n35058 ;
  assign n35060 = ( n15383 & n35057 ) | ( n15383 & ~n35059 ) | ( n35057 & ~n35059 ) ;
  assign n35061 = n35060 ^ n35057 ^ 1'b0 ;
  assign n35062 = ( n15383 & n35060 ) | ( n15383 & ~n35061 ) | ( n35060 & ~n35061 ) ;
  assign n35063 = n15383 & ~n35056 ;
  assign n35064 = n35062 & ~n35063 ;
  assign n35065 = n5061 & n35064 ;
  assign n35066 = ( x224 & n35048 ) | ( x224 & ~n35065 ) | ( n35048 & ~n35065 ) ;
  assign n35067 = ~n35048 & n35066 ;
  assign n35068 = ( n2263 & n35038 ) | ( n2263 & ~n35067 ) | ( n35038 & ~n35067 ) ;
  assign n35069 = ~n35038 & n35068 ;
  assign n35070 = x224 & ~n15337 ;
  assign n35071 = n2263 | n35070 ;
  assign n35072 = n15458 & n15524 ;
  assign n35073 = n35071 | n35072 ;
  assign n35074 = ( x215 & ~n35069 ) | ( x215 & n35073 ) | ( ~n35069 & n35073 ) ;
  assign n35075 = ~x215 & n35074 ;
  assign n35076 = n15370 & n35040 ;
  assign n35077 = n35076 ^ n15383 ^ 1'b0 ;
  assign n35078 = n15381 | n35042 ;
  assign n35079 = ~x680 & n35076 ;
  assign n35080 = ( x680 & ~n35078 ) | ( x680 & n35079 ) | ( ~n35078 & n35079 ) ;
  assign n35081 = ( n35076 & ~n35077 ) | ( n35076 & n35080 ) | ( ~n35077 & n35080 ) ;
  assign n35082 = ~n5061 & n35081 ;
  assign n35083 = x614 & ~n15548 ;
  assign n35084 = n33581 & ~n35083 ;
  assign n35085 = x680 | n35084 ;
  assign n35086 = x680 & ~n15552 ;
  assign n35087 = ~n15368 & n35086 ;
  assign n35088 = ( n15383 & n35085 ) | ( n15383 & ~n35087 ) | ( n35085 & ~n35087 ) ;
  assign n35089 = n35088 ^ n35085 ^ 1'b0 ;
  assign n35090 = ( n15383 & n35088 ) | ( n15383 & ~n35089 ) | ( n35088 & ~n35089 ) ;
  assign n35091 = n15383 & ~n35084 ;
  assign n35092 = n35090 & ~n35091 ;
  assign n35093 = n5061 & n35092 ;
  assign n35094 = ( x224 & n35082 ) | ( x224 & ~n35093 ) | ( n35082 & ~n35093 ) ;
  assign n35095 = ~n35082 & n35094 ;
  assign n35096 = x614 & n33876 ;
  assign n35097 = ~x224 & n35096 ;
  assign n35098 = ~n15613 & n35097 ;
  assign n35099 = ( x215 & n35095 ) | ( x215 & n35098 ) | ( n35095 & n35098 ) ;
  assign n35100 = n35098 ^ n35095 ^ 1'b0 ;
  assign n35101 = ( x215 & n35099 ) | ( x215 & n35100 ) | ( n35099 & n35100 ) ;
  assign n35102 = ( x299 & n35075 ) | ( x299 & ~n35101 ) | ( n35075 & ~n35101 ) ;
  assign n35103 = ~n35075 & n35102 ;
  assign n35104 = ~n15618 & n35097 ;
  assign n35105 = ~n5114 & n35081 ;
  assign n35106 = n5114 & n35092 ;
  assign n35107 = ( x224 & n35105 ) | ( x224 & ~n35106 ) | ( n35105 & ~n35106 ) ;
  assign n35108 = ~n35105 & n35107 ;
  assign n35109 = ( x223 & n35104 ) | ( x223 & ~n35108 ) | ( n35104 & ~n35108 ) ;
  assign n35110 = ~n35104 & n35109 ;
  assign n35119 = ( x223 & x614 ) | ( x223 & n15776 ) | ( x614 & n15776 ) ;
  assign n35111 = ~n5114 & n35047 ;
  assign n35112 = n5114 & n35064 ;
  assign n35113 = ( x224 & n35111 ) | ( x224 & ~n35112 ) | ( n35111 & ~n35112 ) ;
  assign n35114 = ~n35111 & n35113 ;
  assign n35115 = n5114 | n35035 ;
  assign n35116 = n5114 & ~n35033 ;
  assign n35117 = n4692 & ~n35116 ;
  assign n35118 = n35115 & n35117 ;
  assign n35120 = ( n35114 & n35118 ) | ( n35114 & ~n35119 ) | ( n35118 & ~n35119 ) ;
  assign n35121 = n35119 | n35120 ;
  assign n35122 = n35121 ^ n35110 ^ 1'b0 ;
  assign n35123 = ( n35110 & n35121 ) | ( n35110 & n35122 ) | ( n35121 & n35122 ) ;
  assign n35124 = ( x299 & ~n35110 ) | ( x299 & n35123 ) | ( ~n35110 & n35123 ) ;
  assign n35125 = ( x39 & n35103 ) | ( x39 & n35124 ) | ( n35103 & n35124 ) ;
  assign n35126 = ~n35103 & n35125 ;
  assign n35127 = ( x38 & ~n35024 ) | ( x38 & n35126 ) | ( ~n35024 & n35126 ) ;
  assign n35128 = n35024 | n35127 ;
  assign n35129 = ( n2069 & ~n35009 ) | ( n2069 & n35128 ) | ( ~n35009 & n35128 ) ;
  assign n35130 = ~n2069 & n35129 ;
  assign n35131 = n35130 ^ x224 ^ 1'b0 ;
  assign n35132 = ( ~x224 & n2069 ) | ( ~x224 & n35131 ) | ( n2069 & n35131 ) ;
  assign n35133 = ( x224 & n35130 ) | ( x224 & n35132 ) | ( n35130 & n35132 ) ;
  assign n35134 = n35005 ^ n15659 ^ 1'b0 ;
  assign n35135 = ( n35005 & n35133 ) | ( n35005 & ~n35134 ) | ( n35133 & ~n35134 ) ;
  assign n35136 = x609 & ~n35135 ;
  assign n35137 = x609 | n35005 ;
  assign n35138 = ( x1155 & n35136 ) | ( x1155 & n35137 ) | ( n35136 & n35137 ) ;
  assign n35139 = ~n35136 & n35138 ;
  assign n35140 = x609 & ~n35005 ;
  assign n35141 = x1155 | n35140 ;
  assign n35142 = ( n35135 & n35136 ) | ( n35135 & ~n35141 ) | ( n35136 & ~n35141 ) ;
  assign n35143 = n35139 | n35142 ;
  assign n35144 = n35135 ^ x785 ^ 1'b0 ;
  assign n35145 = ( n35135 & n35143 ) | ( n35135 & n35144 ) | ( n35143 & n35144 ) ;
  assign n35146 = x618 & ~n35145 ;
  assign n35147 = x618 | n35005 ;
  assign n35148 = ( x1154 & n35146 ) | ( x1154 & n35147 ) | ( n35146 & n35147 ) ;
  assign n35149 = ~n35146 & n35148 ;
  assign n35150 = x618 & ~n35005 ;
  assign n35151 = x1154 | n35150 ;
  assign n35152 = ( n35145 & n35146 ) | ( n35145 & ~n35151 ) | ( n35146 & ~n35151 ) ;
  assign n35153 = n35149 | n35152 ;
  assign n35154 = n35145 ^ x781 ^ 1'b0 ;
  assign n35155 = ( n35145 & n35153 ) | ( n35145 & n35154 ) | ( n35153 & n35154 ) ;
  assign n35156 = x619 & ~n35155 ;
  assign n35157 = x619 | n35005 ;
  assign n35158 = ( x1159 & n35156 ) | ( x1159 & n35157 ) | ( n35156 & n35157 ) ;
  assign n35159 = ~n35156 & n35158 ;
  assign n35160 = x619 & ~n35005 ;
  assign n35161 = x1159 | n35160 ;
  assign n35162 = ( n35155 & n35156 ) | ( n35155 & ~n35161 ) | ( n35156 & ~n35161 ) ;
  assign n35163 = n35159 | n35162 ;
  assign n35164 = n35155 ^ x789 ^ 1'b0 ;
  assign n35165 = ( n35155 & n35163 ) | ( n35155 & n35164 ) | ( n35163 & n35164 ) ;
  assign n35166 = n35005 ^ n16518 ^ 1'b0 ;
  assign n35167 = ( n35005 & n35165 ) | ( n35005 & ~n35166 ) | ( n35165 & ~n35166 ) ;
  assign n35168 = n35005 ^ n16339 ^ 1'b0 ;
  assign n35169 = ( n35005 & n35167 ) | ( n35005 & ~n35168 ) | ( n35167 & ~n35168 ) ;
  assign n35170 = n19055 & n35169 ;
  assign n35171 = x662 & n16184 ;
  assign n35172 = n35007 & ~n35171 ;
  assign n35173 = x662 & x680 ;
  assign n35174 = n15697 & n35173 ;
  assign n35175 = n35071 | n35174 ;
  assign n35176 = n5076 | n33993 ;
  assign n35177 = n15433 & n35176 ;
  assign n35178 = n5061 & n35177 ;
  assign n35179 = n15468 ^ x662 ^ 1'b0 ;
  assign n35180 = ( n15468 & n16119 ) | ( n15468 & n35179 ) | ( n16119 & n35179 ) ;
  assign n35181 = ~n5061 & n35180 ;
  assign n35182 = ( x224 & n35178 ) | ( x224 & ~n35181 ) | ( n35178 & ~n35181 ) ;
  assign n35183 = ~n35178 & n35182 ;
  assign n35184 = n16146 & n35173 ;
  assign n35185 = n5061 | n35184 ;
  assign n35186 = x662 & n16152 ;
  assign n35187 = n5061 & ~n35186 ;
  assign n35188 = ( x224 & n35185 ) | ( x224 & ~n35187 ) | ( n35185 & ~n35187 ) ;
  assign n35189 = ~x224 & n35188 ;
  assign n35190 = ( n2263 & n35183 ) | ( n2263 & ~n35189 ) | ( n35183 & ~n35189 ) ;
  assign n35191 = ~n35183 & n35190 ;
  assign n35192 = ( x215 & n35175 ) | ( x215 & ~n35191 ) | ( n35175 & ~n35191 ) ;
  assign n35193 = n35192 ^ n35175 ^ 1'b0 ;
  assign n35194 = ( x215 & n35192 ) | ( x215 & ~n35193 ) | ( n35192 & ~n35193 ) ;
  assign n35195 = n15402 ^ x662 ^ 1'b0 ;
  assign n35196 = ( n15402 & n33966 ) | ( n15402 & n35195 ) | ( n33966 & n35195 ) ;
  assign n35197 = ~n5061 & n35196 ;
  assign n35198 = n15378 ^ x662 ^ 1'b0 ;
  assign n35199 = ( n15378 & n16100 ) | ( n15378 & n35198 ) | ( n16100 & n35198 ) ;
  assign n35200 = n5061 & n35199 ;
  assign n35201 = ( x224 & n35197 ) | ( x224 & ~n35200 ) | ( n35197 & ~n35200 ) ;
  assign n35202 = ~n35197 & n35201 ;
  assign n35203 = ~x224 & x662 ;
  assign n35204 = n16172 & n35203 ;
  assign n35205 = ( x215 & n35202 ) | ( x215 & ~n35204 ) | ( n35202 & ~n35204 ) ;
  assign n35206 = ~n35202 & n35205 ;
  assign n35207 = x299 & ~n35206 ;
  assign n35208 = n35194 & n35207 ;
  assign n35209 = ~n5114 & n35196 ;
  assign n35210 = n5114 & n35199 ;
  assign n35211 = ( x224 & n35209 ) | ( x224 & ~n35210 ) | ( n35209 & ~n35210 ) ;
  assign n35212 = ~n35209 & n35211 ;
  assign n35213 = n16144 & n35203 ;
  assign n35214 = x223 & ~n35213 ;
  assign n35215 = n35214 ^ n35212 ^ 1'b0 ;
  assign n35216 = ( n35212 & n35214 ) | ( n35212 & n35215 ) | ( n35214 & n35215 ) ;
  assign n35217 = ( x299 & ~n35212 ) | ( x299 & n35216 ) | ( ~n35212 & n35216 ) ;
  assign n35218 = ~n5114 & n35180 ;
  assign n35219 = n5114 & n35177 ;
  assign n35220 = ( x224 & n35218 ) | ( x224 & ~n35219 ) | ( n35218 & ~n35219 ) ;
  assign n35221 = ~n35218 & n35220 ;
  assign n35222 = n5114 & ~n35186 ;
  assign n35223 = n5114 | n35184 ;
  assign n35224 = ( n4692 & n35222 ) | ( n4692 & n35223 ) | ( n35222 & n35223 ) ;
  assign n35225 = ~n35222 & n35224 ;
  assign n35226 = x662 & n16145 ;
  assign n35227 = ( x223 & ~n35225 ) | ( x223 & n35226 ) | ( ~n35225 & n35226 ) ;
  assign n35228 = n35225 | n35227 ;
  assign n35229 = ( ~n35217 & n35221 ) | ( ~n35217 & n35228 ) | ( n35221 & n35228 ) ;
  assign n35230 = ~n35217 & n35229 ;
  assign n35231 = ( x39 & n35208 ) | ( x39 & ~n35230 ) | ( n35208 & ~n35230 ) ;
  assign n35232 = ~n35208 & n35231 ;
  assign n35233 = x224 & n16038 ;
  assign n35234 = x299 | n35233 ;
  assign n35235 = n35173 & ~n35234 ;
  assign n35236 = ( n16018 & n35234 ) | ( n16018 & ~n35235 ) | ( n35234 & ~n35235 ) ;
  assign n35237 = ( x224 & n16018 ) | ( x224 & ~n35236 ) | ( n16018 & ~n35236 ) ;
  assign n35238 = ~n35236 & n35237 ;
  assign n35239 = x224 & n16033 ;
  assign n35240 = n16024 & ~n35173 ;
  assign n35241 = ( x299 & n35239 ) | ( x299 & ~n35240 ) | ( n35239 & ~n35240 ) ;
  assign n35242 = ~n35239 & n35241 ;
  assign n35243 = n16024 ^ x224 ^ 1'b0 ;
  assign n35244 = ( x224 & n16024 ) | ( x224 & ~n35243 ) | ( n16024 & ~n35243 ) ;
  assign n35245 = ( n35242 & n35243 ) | ( n35242 & n35244 ) | ( n35243 & n35244 ) ;
  assign n35246 = ( x39 & ~n35238 ) | ( x39 & n35245 ) | ( ~n35238 & n35245 ) ;
  assign n35247 = n35238 | n35246 ;
  assign n35248 = n35247 ^ n35232 ^ 1'b0 ;
  assign n35249 = ( n35232 & n35247 ) | ( n35232 & n35248 ) | ( n35247 & n35248 ) ;
  assign n35250 = ( x38 & ~n35232 ) | ( x38 & n35249 ) | ( ~n35232 & n35249 ) ;
  assign n35251 = ( n2069 & ~n35172 ) | ( n2069 & n35250 ) | ( ~n35172 & n35250 ) ;
  assign n35252 = ~n2069 & n35251 ;
  assign n35253 = n35252 ^ x224 ^ 1'b0 ;
  assign n35254 = ( ~x224 & n2069 ) | ( ~x224 & n35253 ) | ( n2069 & n35253 ) ;
  assign n35255 = ( x224 & n35252 ) | ( x224 & n35254 ) | ( n35252 & n35254 ) ;
  assign n35256 = x625 & ~n35255 ;
  assign n35257 = x625 | n35005 ;
  assign n35258 = ( x1153 & n35256 ) | ( x1153 & n35257 ) | ( n35256 & n35257 ) ;
  assign n35259 = ~n35256 & n35258 ;
  assign n35260 = x625 & ~n35005 ;
  assign n35261 = x1153 | n35260 ;
  assign n35262 = ( n35255 & n35256 ) | ( n35255 & ~n35261 ) | ( n35256 & ~n35261 ) ;
  assign n35263 = n35259 | n35262 ;
  assign n35264 = n35255 ^ x778 ^ 1'b0 ;
  assign n35265 = ( n35255 & n35263 ) | ( n35255 & n35264 ) | ( n35263 & n35264 ) ;
  assign n35266 = n35005 ^ n16234 ^ 1'b0 ;
  assign n35267 = ( n35005 & n35265 ) | ( n35005 & ~n35266 ) | ( n35265 & ~n35266 ) ;
  assign n35268 = n35005 ^ n16254 ^ 1'b0 ;
  assign n35269 = ( n35005 & n35267 ) | ( n35005 & ~n35268 ) | ( n35267 & ~n35268 ) ;
  assign n35270 = n16279 | n35269 ;
  assign n35271 = n16318 | n35270 ;
  assign n35272 = n17086 & ~n35005 ;
  assign n35273 = n35271 & ~n35272 ;
  assign n35274 = n17093 | n35273 ;
  assign n35275 = n16559 & ~n35005 ;
  assign n35276 = n35274 & ~n35275 ;
  assign n35277 = x647 & ~n35276 ;
  assign n35278 = x647 | n35005 ;
  assign n35279 = ( x1157 & n35277 ) | ( x1157 & n35278 ) | ( n35277 & n35278 ) ;
  assign n35280 = ~n35277 & n35279 ;
  assign n35281 = x647 & ~n35005 ;
  assign n35282 = x1157 | n35281 ;
  assign n35283 = ( n35276 & n35277 ) | ( n35276 & ~n35282 ) | ( n35277 & ~n35282 ) ;
  assign n35284 = ( n16375 & n35280 ) | ( n16375 & n35283 ) | ( n35280 & n35283 ) ;
  assign n35285 = ( x787 & n35170 ) | ( x787 & n35284 ) | ( n35170 & n35284 ) ;
  assign n35286 = n35284 ^ n35170 ^ 1'b0 ;
  assign n35287 = ( x787 & n35285 ) | ( x787 & n35286 ) | ( n35285 & n35286 ) ;
  assign n35288 = n35014 | n35173 ;
  assign n35289 = ~x614 & n15636 ;
  assign n35290 = n34117 | n35289 ;
  assign n35291 = x224 & n35290 ;
  assign n35292 = x224 | n16026 ;
  assign n35293 = n35010 | n35292 ;
  assign n35294 = n35173 & ~n35293 ;
  assign n35295 = ( n35173 & n35291 ) | ( n35173 & n35294 ) | ( n35291 & n35294 ) ;
  assign n35296 = x299 & ~n35295 ;
  assign n35297 = n35288 & n35296 ;
  assign n35298 = n16020 & n35173 ;
  assign n35299 = ( ~x224 & n35016 ) | ( ~x224 & n35298 ) | ( n35016 & n35298 ) ;
  assign n35300 = ~x224 & n35299 ;
  assign n35301 = ~n34133 & n35019 ;
  assign n35302 = n16020 & ~n35173 ;
  assign n35303 = n35301 & ~n35302 ;
  assign n35304 = ( ~x299 & n35300 ) | ( ~x299 & n35303 ) | ( n35300 & n35303 ) ;
  assign n35305 = ~x299 & n35304 ;
  assign n35306 = ( ~x39 & n35297 ) | ( ~x39 & n35305 ) | ( n35297 & n35305 ) ;
  assign n35307 = ~x39 & n35306 ;
  assign n35308 = ( n15695 & n34205 ) | ( n15695 & n35049 ) | ( n34205 & n35049 ) ;
  assign n35309 = x680 & n35308 ;
  assign n35310 = x680 & n15752 ;
  assign n35311 = n35072 | n35310 ;
  assign n35312 = ~n35309 & n35311 ;
  assign n35313 = n35096 ^ x662 ^ 1'b0 ;
  assign n35314 = ( n35096 & n35312 ) | ( n35096 & n35313 ) | ( n35312 & n35313 ) ;
  assign n35315 = x224 | n35314 ;
  assign n35316 = n22207 ^ x614 ^ 1'b0 ;
  assign n35317 = ( n22207 & n34716 ) | ( n22207 & n35316 ) | ( n34716 & n35316 ) ;
  assign n35318 = ~n15335 & n35317 ;
  assign n35319 = n35318 ^ x616 ^ 1'b0 ;
  assign n35320 = x614 & ~n15954 ;
  assign n35321 = n15826 & ~n35320 ;
  assign n35322 = ( n35318 & ~n35319 ) | ( n35318 & n35321 ) | ( ~n35319 & n35321 ) ;
  assign n35323 = x680 & n35322 ;
  assign n35324 = ( x662 & ~n35079 ) | ( x662 & n35323 ) | ( ~n35079 & n35323 ) ;
  assign n35325 = ~n35323 & n35324 ;
  assign n35326 = n15730 & ~n35076 ;
  assign n35327 = n15383 | n35080 ;
  assign n35328 = ( n35325 & ~n35326 ) | ( n35325 & n35327 ) | ( ~n35326 & n35327 ) ;
  assign n35329 = ~n35325 & n35328 ;
  assign n35330 = x224 & n35329 ;
  assign n35331 = ( n5114 & n35315 ) | ( n5114 & ~n35330 ) | ( n35315 & ~n35330 ) ;
  assign n35332 = ~n5114 & n35331 ;
  assign n35333 = x614 & ~n34167 ;
  assign n35334 = x680 & ~n15805 ;
  assign n35335 = ( x680 & n35333 ) | ( x680 & n35334 ) | ( n35333 & n35334 ) ;
  assign n35336 = x662 & ~n35085 ;
  assign n35337 = ( x662 & n35335 ) | ( x662 & n35336 ) | ( n35335 & n35336 ) ;
  assign n35338 = n15730 & ~n35084 ;
  assign n35339 = ( n35090 & n35337 ) | ( n35090 & ~n35338 ) | ( n35337 & ~n35338 ) ;
  assign n35340 = ~n35337 & n35339 ;
  assign n35341 = x224 & n35340 ;
  assign n35342 = x614 & ~x680 ;
  assign n35343 = n15609 & n35342 ;
  assign n35344 = ~x614 & n15757 ;
  assign n35345 = x614 & ~n34146 ;
  assign n35346 = x680 & ~n35345 ;
  assign n35347 = ( n15761 & n35344 ) | ( n15761 & n35346 ) | ( n35344 & n35346 ) ;
  assign n35348 = ~n35344 & n35347 ;
  assign n35349 = ( x662 & n35343 ) | ( x662 & ~n35348 ) | ( n35343 & ~n35348 ) ;
  assign n35350 = ~n35343 & n35349 ;
  assign n35351 = n15353 & n35096 ;
  assign n35352 = ( x662 & ~n35350 ) | ( x662 & n35351 ) | ( ~n35350 & n35351 ) ;
  assign n35353 = ~n35350 & n35352 ;
  assign n35354 = x224 | n35353 ;
  assign n35355 = ( n5114 & n35341 ) | ( n5114 & n35354 ) | ( n35341 & n35354 ) ;
  assign n35356 = ~n35341 & n35355 ;
  assign n35357 = ( x223 & n35332 ) | ( x223 & ~n35356 ) | ( n35332 & ~n35356 ) ;
  assign n35358 = ~n35332 & n35357 ;
  assign n35359 = n34206 | n35072 ;
  assign n35360 = ~n35309 & n35359 ;
  assign n35361 = n35035 ^ x662 ^ 1'b0 ;
  assign n35362 = ( n35035 & n35360 ) | ( n35035 & n35361 ) | ( n35360 & n35361 ) ;
  assign n35363 = n5114 | n35362 ;
  assign n35364 = x614 & n15905 ;
  assign n35365 = ~x614 & n15742 ;
  assign n35366 = ( x680 & n35364 ) | ( x680 & ~n35365 ) | ( n35364 & ~n35365 ) ;
  assign n35367 = ~n35364 & n35366 ;
  assign n35368 = x662 & ~n35029 ;
  assign n35369 = ( x662 & n35367 ) | ( x662 & n35368 ) | ( n35367 & n35368 ) ;
  assign n35370 = n15730 & ~n35028 ;
  assign n35371 = ( n35031 & n35369 ) | ( n35031 & ~n35370 ) | ( n35369 & ~n35370 ) ;
  assign n35372 = ~n35369 & n35371 ;
  assign n35373 = n5114 & ~n35372 ;
  assign n35374 = n4692 & ~n35373 ;
  assign n35375 = n35363 & n35374 ;
  assign n35376 = ~n34223 & n35049 ;
  assign n35377 = x614 & ~n34233 ;
  assign n35378 = n35376 | n35377 ;
  assign n35379 = x680 & ~n34231 ;
  assign n35380 = ( x680 & n35378 ) | ( x680 & n35379 ) | ( n35378 & n35379 ) ;
  assign n35381 = x662 & ~n35057 ;
  assign n35382 = ( x662 & n35380 ) | ( x662 & n35381 ) | ( n35380 & n35381 ) ;
  assign n35383 = ( x662 & n35062 ) | ( x662 & n35064 ) | ( n35062 & n35064 ) ;
  assign n35384 = ~n35382 & n35383 ;
  assign n35385 = n5114 & n35384 ;
  assign n35386 = n15730 & ~n35041 ;
  assign n35387 = n15383 | n35045 ;
  assign n35388 = ~n15821 & n34781 ;
  assign n35389 = x614 | n35388 ;
  assign n35390 = ~n35320 & n35389 ;
  assign n35391 = ( n35318 & ~n35319 ) | ( n35318 & n35390 ) | ( ~n35319 & n35390 ) ;
  assign n35392 = x680 & ~n35391 ;
  assign n35393 = x662 & ~n35044 ;
  assign n35394 = ( x662 & n35392 ) | ( x662 & n35393 ) | ( n35392 & n35393 ) ;
  assign n35395 = ( n35386 & n35387 ) | ( n35386 & ~n35394 ) | ( n35387 & ~n35394 ) ;
  assign n35396 = ~n35386 & n35395 ;
  assign n35397 = ~n5114 & n35396 ;
  assign n35398 = ( x224 & n35385 ) | ( x224 & ~n35397 ) | ( n35385 & ~n35397 ) ;
  assign n35399 = ~n35385 & n35398 ;
  assign n35400 = n15694 & n35173 ;
  assign n35401 = ( ~x224 & n35072 ) | ( ~x224 & n35400 ) | ( n35072 & n35400 ) ;
  assign n35402 = ~x224 & n35401 ;
  assign n35403 = ~x222 & n35402 ;
  assign n35404 = x223 | n35403 ;
  assign n35405 = ( ~n35375 & n35399 ) | ( ~n35375 & n35404 ) | ( n35399 & n35404 ) ;
  assign n35406 = n35375 | n35405 ;
  assign n35407 = n35406 ^ n35358 ^ 1'b0 ;
  assign n35408 = ( n35358 & n35406 ) | ( n35358 & n35407 ) | ( n35406 & n35407 ) ;
  assign n35409 = ( x299 & ~n35358 ) | ( x299 & n35408 ) | ( ~n35358 & n35408 ) ;
  assign n35410 = n35027 | n35173 ;
  assign n35411 = x224 & ~n15340 ;
  assign n35412 = ( x224 & n35410 ) | ( x224 & n35411 ) | ( n35410 & n35411 ) ;
  assign n35413 = ( n35173 & n35317 ) | ( n35173 & ~n35412 ) | ( n35317 & ~n35412 ) ;
  assign n35414 = n35413 ^ n35412 ^ 1'b0 ;
  assign n35415 = ( n35412 & ~n35413 ) | ( n35412 & n35414 ) | ( ~n35413 & n35414 ) ;
  assign n35416 = ( n35071 & n35402 ) | ( n35071 & ~n35415 ) | ( n35402 & ~n35415 ) ;
  assign n35417 = n35415 | n35416 ;
  assign n35418 = x224 | n35372 ;
  assign n35419 = x224 & n35384 ;
  assign n35420 = n5061 & ~n35419 ;
  assign n35421 = n35418 & n35420 ;
  assign n35422 = x224 | n35362 ;
  assign n35423 = x224 & n35396 ;
  assign n35424 = ( n5061 & n35422 ) | ( n5061 & ~n35423 ) | ( n35422 & ~n35423 ) ;
  assign n35425 = ~n5061 & n35424 ;
  assign n35426 = ( n2263 & n35421 ) | ( n2263 & ~n35425 ) | ( n35421 & ~n35425 ) ;
  assign n35427 = ~n35421 & n35426 ;
  assign n35428 = ( x215 & n35417 ) | ( x215 & ~n35427 ) | ( n35417 & ~n35427 ) ;
  assign n35429 = ~x215 & n35428 ;
  assign n35430 = n5061 & n35353 ;
  assign n35431 = ~n5061 & n35314 ;
  assign n35432 = ( x224 & ~n35430 ) | ( x224 & n35431 ) | ( ~n35430 & n35431 ) ;
  assign n35433 = n35430 | n35432 ;
  assign n35434 = n5061 & ~n35340 ;
  assign n35435 = n5061 | n35329 ;
  assign n35436 = ( x224 & n35434 ) | ( x224 & n35435 ) | ( n35434 & n35435 ) ;
  assign n35437 = ~n35434 & n35436 ;
  assign n35438 = x215 & ~n35437 ;
  assign n35439 = n35433 & n35438 ;
  assign n35440 = ( x299 & n35429 ) | ( x299 & ~n35439 ) | ( n35429 & ~n35439 ) ;
  assign n35441 = ~n35429 & n35440 ;
  assign n35442 = x39 & ~n35441 ;
  assign n35443 = n35409 & n35442 ;
  assign n35444 = ( x38 & ~n35307 ) | ( x38 & n35443 ) | ( ~n35307 & n35443 ) ;
  assign n35445 = n35307 | n35444 ;
  assign n35446 = x662 & n15691 ;
  assign n35447 = n15644 & n35446 ;
  assign n35448 = n35009 & ~n35447 ;
  assign n35449 = ( n2069 & n35445 ) | ( n2069 & ~n35448 ) | ( n35445 & ~n35448 ) ;
  assign n35450 = ~n2069 & n35449 ;
  assign n35451 = n35450 ^ x224 ^ 1'b0 ;
  assign n35452 = ( ~x224 & n2069 ) | ( ~x224 & n35451 ) | ( n2069 & n35451 ) ;
  assign n35453 = ( x224 & n35450 ) | ( x224 & n35452 ) | ( n35450 & n35452 ) ;
  assign n35454 = x625 & ~n35453 ;
  assign n35455 = x625 | n35133 ;
  assign n35456 = ( x1153 & n35454 ) | ( x1153 & n35455 ) | ( n35454 & n35455 ) ;
  assign n35457 = ~n35454 & n35456 ;
  assign n35458 = ( x608 & n35262 ) | ( x608 & ~n35457 ) | ( n35262 & ~n35457 ) ;
  assign n35459 = ~n35262 & n35458 ;
  assign n35460 = x625 & ~n35133 ;
  assign n35461 = x1153 | n35460 ;
  assign n35462 = ( x625 & n35453 ) | ( x625 & ~n35461 ) | ( n35453 & ~n35461 ) ;
  assign n35463 = ~n35461 & n35462 ;
  assign n35464 = x608 | n35259 ;
  assign n35465 = ( ~n35459 & n35463 ) | ( ~n35459 & n35464 ) | ( n35463 & n35464 ) ;
  assign n35466 = ~n35459 & n35465 ;
  assign n35467 = n35453 ^ x778 ^ 1'b0 ;
  assign n35468 = ( n35453 & n35466 ) | ( n35453 & n35467 ) | ( n35466 & n35467 ) ;
  assign n35469 = x609 & ~n35468 ;
  assign n35470 = x609 | n35265 ;
  assign n35471 = ( x1155 & n35469 ) | ( x1155 & n35470 ) | ( n35469 & n35470 ) ;
  assign n35472 = ~n35469 & n35471 ;
  assign n35473 = ( x660 & n35142 ) | ( x660 & ~n35472 ) | ( n35142 & ~n35472 ) ;
  assign n35474 = ~n35142 & n35473 ;
  assign n35475 = x609 & ~n35265 ;
  assign n35476 = x1155 | n35475 ;
  assign n35477 = ( x609 & n35468 ) | ( x609 & ~n35476 ) | ( n35468 & ~n35476 ) ;
  assign n35478 = ~n35476 & n35477 ;
  assign n35479 = x660 | n35139 ;
  assign n35480 = ( ~n35474 & n35478 ) | ( ~n35474 & n35479 ) | ( n35478 & n35479 ) ;
  assign n35481 = ~n35474 & n35480 ;
  assign n35482 = n35468 ^ x785 ^ 1'b0 ;
  assign n35483 = ( n35468 & n35481 ) | ( n35468 & n35482 ) | ( n35481 & n35482 ) ;
  assign n35484 = x618 & ~n35483 ;
  assign n35485 = x618 | n35267 ;
  assign n35486 = ( x1154 & n35484 ) | ( x1154 & n35485 ) | ( n35484 & n35485 ) ;
  assign n35487 = ~n35484 & n35486 ;
  assign n35488 = ( x627 & n35152 ) | ( x627 & ~n35487 ) | ( n35152 & ~n35487 ) ;
  assign n35489 = ~n35152 & n35488 ;
  assign n35490 = x627 | n35149 ;
  assign n35491 = x618 & ~n35267 ;
  assign n35492 = x1154 | n35491 ;
  assign n35493 = ( n35483 & n35484 ) | ( n35483 & ~n35492 ) | ( n35484 & ~n35492 ) ;
  assign n35494 = ( ~n35489 & n35490 ) | ( ~n35489 & n35493 ) | ( n35490 & n35493 ) ;
  assign n35495 = ~n35489 & n35494 ;
  assign n35496 = n35483 ^ x781 ^ 1'b0 ;
  assign n35497 = ( n35483 & n35495 ) | ( n35483 & n35496 ) | ( n35495 & n35496 ) ;
  assign n35498 = x619 | n35497 ;
  assign n35499 = x619 & ~n35269 ;
  assign n35500 = ( x1159 & n35498 ) | ( x1159 & ~n35499 ) | ( n35498 & ~n35499 ) ;
  assign n35501 = ~x1159 & n35500 ;
  assign n35502 = ( x648 & n35159 ) | ( x648 & ~n35501 ) | ( n35159 & ~n35501 ) ;
  assign n35503 = n35501 | n35502 ;
  assign n35504 = x619 & ~n35497 ;
  assign n35505 = x619 | n35269 ;
  assign n35506 = ( x1159 & n35504 ) | ( x1159 & n35505 ) | ( n35504 & n35505 ) ;
  assign n35507 = ~n35504 & n35506 ;
  assign n35508 = ( x648 & n35162 ) | ( x648 & ~n35507 ) | ( n35162 & ~n35507 ) ;
  assign n35509 = ~n35162 & n35508 ;
  assign n35510 = x789 & ~n35509 ;
  assign n35511 = n35503 & n35510 ;
  assign n35512 = ~x789 & n35497 ;
  assign n35513 = ( n16519 & ~n35511 ) | ( n16519 & n35512 ) | ( ~n35511 & n35512 ) ;
  assign n35514 = n35511 | n35513 ;
  assign n35515 = x628 | n35273 ;
  assign n35516 = x628 | n35005 ;
  assign n35517 = x628 & ~n35273 ;
  assign n35518 = n16337 & ~n35517 ;
  assign n35519 = n35516 & n35518 ;
  assign n35520 = x628 & ~n35005 ;
  assign n35521 = n16338 & ~n35520 ;
  assign n35522 = n35519 ^ n35515 ^ 1'b0 ;
  assign n35523 = ( ~n35515 & n35521 ) | ( ~n35515 & n35522 ) | ( n35521 & n35522 ) ;
  assign n35524 = ( n35515 & n35519 ) | ( n35515 & n35523 ) | ( n35519 & n35523 ) ;
  assign n35525 = n19046 & n35167 ;
  assign n35526 = ( x792 & n35524 ) | ( x792 & n35525 ) | ( n35524 & n35525 ) ;
  assign n35527 = n35525 ^ n35524 ^ 1'b0 ;
  assign n35528 = ( x792 & n35526 ) | ( x792 & n35527 ) | ( n35526 & n35527 ) ;
  assign n35529 = n16279 & ~n35005 ;
  assign n35530 = n16459 & ~n35270 ;
  assign n35531 = ( n16459 & n35529 ) | ( n16459 & n35530 ) | ( n35529 & n35530 ) ;
  assign n35532 = x626 & n35005 ;
  assign n35533 = ~x626 & n35165 ;
  assign n35534 = ( n22322 & n35532 ) | ( n22322 & ~n35533 ) | ( n35532 & ~n35533 ) ;
  assign n35535 = ~n35532 & n35534 ;
  assign n35536 = x626 & n35165 ;
  assign n35537 = ~x626 & n35005 ;
  assign n35538 = ( n22317 & n35536 ) | ( n22317 & ~n35537 ) | ( n35536 & ~n35537 ) ;
  assign n35539 = ~n35536 & n35538 ;
  assign n35540 = ( ~n35531 & n35535 ) | ( ~n35531 & n35539 ) | ( n35535 & n35539 ) ;
  assign n35541 = n35531 | n35540 ;
  assign n35542 = ( x788 & ~n22314 ) | ( x788 & n35541 ) | ( ~n22314 & n35541 ) ;
  assign n35543 = ( n18482 & n22314 ) | ( n18482 & n35542 ) | ( n22314 & n35542 ) ;
  assign n35544 = ~n35528 & n35543 ;
  assign n35545 = ( n35514 & n35528 ) | ( n35514 & ~n35544 ) | ( n35528 & ~n35544 ) ;
  assign n35546 = ( ~n18484 & n35287 ) | ( ~n18484 & n35545 ) | ( n35287 & n35545 ) ;
  assign n35547 = n35287 ^ n18484 ^ 1'b0 ;
  assign n35548 = ( n35287 & n35546 ) | ( n35287 & ~n35547 ) | ( n35546 & ~n35547 ) ;
  assign n35549 = x644 & ~n35548 ;
  assign n35550 = n35280 | n35283 ;
  assign n35551 = n35276 ^ x787 ^ 1'b0 ;
  assign n35552 = ( n35276 & n35550 ) | ( n35276 & n35551 ) | ( n35550 & n35551 ) ;
  assign n35553 = x644 | n35552 ;
  assign n35554 = ( x715 & n35549 ) | ( x715 & n35553 ) | ( n35549 & n35553 ) ;
  assign n35555 = ~n35549 & n35554 ;
  assign n35556 = x644 | n35005 ;
  assign n35557 = n35005 ^ n16376 ^ 1'b0 ;
  assign n35558 = ( n35005 & n35169 ) | ( n35005 & ~n35557 ) | ( n35169 & ~n35557 ) ;
  assign n35559 = x644 & ~n35558 ;
  assign n35560 = ( x715 & n35556 ) | ( x715 & ~n35559 ) | ( n35556 & ~n35559 ) ;
  assign n35561 = ~x715 & n35560 ;
  assign n35562 = ( x1160 & n35555 ) | ( x1160 & ~n35561 ) | ( n35555 & ~n35561 ) ;
  assign n35563 = ~n35555 & n35562 ;
  assign n35564 = x644 & ~n35005 ;
  assign n35565 = x715 & ~n35564 ;
  assign n35566 = n35565 ^ x1160 ^ 1'b0 ;
  assign n35567 = x644 | n35558 ;
  assign n35568 = ( n35565 & ~n35566 ) | ( n35565 & n35567 ) | ( ~n35566 & n35567 ) ;
  assign n35569 = ( x1160 & n35566 ) | ( x1160 & n35568 ) | ( n35566 & n35568 ) ;
  assign n35570 = x644 & ~n35552 ;
  assign n35571 = x715 | n35570 ;
  assign n35572 = ( n35548 & n35549 ) | ( n35548 & ~n35571 ) | ( n35549 & ~n35571 ) ;
  assign n35573 = ( ~n35563 & n35569 ) | ( ~n35563 & n35572 ) | ( n35569 & n35572 ) ;
  assign n35574 = ~n35563 & n35573 ;
  assign n35575 = n35548 ^ x790 ^ 1'b0 ;
  assign n35576 = ( n35548 & n35574 ) | ( n35548 & n35575 ) | ( n35574 & n35575 ) ;
  assign n35577 = n35576 ^ n7318 ^ 1'b0 ;
  assign n35578 = ( x224 & n35576 ) | ( x224 & n35577 ) | ( n35576 & n35577 ) ;
  assign n35579 = n1979 & ~n2036 ;
  assign n35580 = ~n2150 & n35579 ;
  assign n35581 = ~x62 & n35580 ;
  assign n35582 = ( x57 & x59 ) | ( x57 & ~n35581 ) | ( x59 & ~n35581 ) ;
  assign n35583 = ~n2096 & n35579 ;
  assign n35584 = x54 & ~n35583 ;
  assign n35585 = n2046 & n35579 ;
  assign n35586 = x87 & n35579 ;
  assign n35587 = n5044 | n5165 ;
  assign n35588 = ~x137 & n35587 ;
  assign n35589 = n5019 & ~n35588 ;
  assign n35590 = x38 & ~x137 ;
  assign n35591 = x39 & n1979 ;
  assign n35592 = n1773 | n10069 ;
  assign n35593 = ( ~n1433 & n1856 ) | ( ~n1433 & n35592 ) | ( n1856 & n35592 ) ;
  assign n35594 = ~n1433 & n35593 ;
  assign n35595 = ( x32 & n1586 ) | ( x32 & ~n35594 ) | ( n1586 & ~n35594 ) ;
  assign n35596 = n35594 | n35595 ;
  assign n35597 = ~n1601 & n35596 ;
  assign n35598 = x95 | n35597 ;
  assign n35599 = ( ~x95 & n1785 ) | ( ~x95 & n35598 ) | ( n1785 & n35598 ) ;
  assign n35600 = n35599 ^ x137 ^ 1'b0 ;
  assign n35601 = ~n1665 & n6442 ;
  assign n35602 = n1288 | n6393 ;
  assign n35603 = n10068 & ~n35602 ;
  assign n35604 = n35601 & n35603 ;
  assign n35605 = ~n1288 & n10069 ;
  assign n35606 = n1654 | n35605 ;
  assign n35607 = ~n1665 & n35606 ;
  assign n35608 = ~n6442 & n35607 ;
  assign n35609 = n35604 | n35608 ;
  assign n35610 = n1666 & ~n6442 ;
  assign n35611 = n1632 & ~n35602 ;
  assign n35612 = ( x32 & n35601 ) | ( x32 & n35611 ) | ( n35601 & n35611 ) ;
  assign n35613 = n35601 & n35612 ;
  assign n35614 = ( x1093 & n35610 ) | ( x1093 & ~n35613 ) | ( n35610 & ~n35613 ) ;
  assign n35615 = ~n35610 & n35614 ;
  assign n35616 = n1407 & ~n35602 ;
  assign n35617 = ( x32 & n35601 ) | ( x32 & n35616 ) | ( n35601 & n35616 ) ;
  assign n35618 = n35601 & n35617 ;
  assign n35619 = x1093 | n35618 ;
  assign n35620 = n35610 | n35619 ;
  assign n35621 = n10151 & ~n35620 ;
  assign n35622 = ( n10151 & n35615 ) | ( n10151 & n35621 ) | ( n35615 & n35621 ) ;
  assign n35623 = ~n35609 & n35622 ;
  assign n35624 = n35609 | n35619 ;
  assign n35625 = x1093 & ~n35607 ;
  assign n35626 = n35624 & ~n35625 ;
  assign n35627 = ( n10196 & ~n35623 ) | ( n10196 & n35626 ) | ( ~n35623 & n35626 ) ;
  assign n35628 = ~n35623 & n35627 ;
  assign n35629 = ( ~x137 & n35599 ) | ( ~x137 & n35600 ) | ( n35599 & n35600 ) ;
  assign n35630 = ( ~n35600 & n35628 ) | ( ~n35600 & n35629 ) | ( n35628 & n35629 ) ;
  assign n35631 = n1785 | n1893 ;
  assign n35632 = x137 & ~n35631 ;
  assign n35633 = x1093 & ~n1666 ;
  assign n35634 = n35620 & ~n35633 ;
  assign n35635 = n10196 | n35634 ;
  assign n35636 = ( n35622 & ~n35632 ) | ( n35622 & n35635 ) | ( ~n35632 & n35635 ) ;
  assign n35637 = ~n35622 & n35636 ;
  assign n35638 = n35630 ^ x332 ^ 1'b0 ;
  assign n35639 = ( n35630 & n35637 ) | ( n35630 & ~n35638 ) | ( n35637 & ~n35638 ) ;
  assign n35640 = ~n1330 & n35639 ;
  assign n35641 = ( n35599 & ~n35600 ) | ( n35599 & n35607 ) | ( ~n35600 & n35607 ) ;
  assign n35642 = n1666 ^ x137 ^ 1'b0 ;
  assign n35643 = ( n1666 & n35631 ) | ( n1666 & n35642 ) | ( n35631 & n35642 ) ;
  assign n35644 = n35641 ^ x332 ^ 1'b0 ;
  assign n35645 = ( n35641 & n35643 ) | ( n35641 & ~n35644 ) | ( n35643 & ~n35644 ) ;
  assign n35646 = n1330 & n35645 ;
  assign n35647 = ( x210 & ~n35640 ) | ( x210 & n35646 ) | ( ~n35640 & n35646 ) ;
  assign n35648 = n35640 | n35647 ;
  assign n35649 = x137 | n1384 ;
  assign n35650 = n35606 & ~n35649 ;
  assign n35651 = ~n1383 & n35596 ;
  assign n35652 = ( x95 & n1426 ) | ( x95 & n35651 ) | ( n1426 & n35651 ) ;
  assign n35653 = n1426 & n35652 ;
  assign n35654 = ( x332 & n35650 ) | ( x332 & ~n35653 ) | ( n35650 & ~n35653 ) ;
  assign n35655 = ~n35650 & n35654 ;
  assign n35656 = ( x137 & n1785 ) | ( x137 & ~n1887 ) | ( n1785 & ~n1887 ) ;
  assign n35657 = ~n1785 & n35656 ;
  assign n35658 = ( x137 & n1655 ) | ( x137 & ~n35657 ) | ( n1655 & ~n35657 ) ;
  assign n35659 = ~n35657 & n35658 ;
  assign n35660 = ( x332 & ~n35655 ) | ( x332 & n35659 ) | ( ~n35655 & n35659 ) ;
  assign n35661 = ~n35655 & n35660 ;
  assign n35662 = ( x299 & n15096 ) | ( x299 & n35661 ) | ( n15096 & n35661 ) ;
  assign n35663 = n35648 & n35662 ;
  assign n35664 = x198 & ~n35661 ;
  assign n35665 = n5412 & n35645 ;
  assign n35666 = ~n5412 & n35639 ;
  assign n35667 = ( x198 & ~n35665 ) | ( x198 & n35666 ) | ( ~n35665 & n35666 ) ;
  assign n35668 = n35665 | n35667 ;
  assign n35669 = ( x299 & ~n35664 ) | ( x299 & n35668 ) | ( ~n35664 & n35668 ) ;
  assign n35670 = ~x299 & n35669 ;
  assign n35671 = ( ~x39 & n35663 ) | ( ~x39 & n35670 ) | ( n35663 & n35670 ) ;
  assign n35672 = ~x39 & n35671 ;
  assign n35673 = ( x38 & ~n35591 ) | ( x38 & n35672 ) | ( ~n35591 & n35672 ) ;
  assign n35674 = n35591 | n35673 ;
  assign n35675 = ( n5054 & ~n35590 ) | ( n5054 & n35674 ) | ( ~n35590 & n35674 ) ;
  assign n35676 = ~n5054 & n35675 ;
  assign n35677 = ( ~x87 & n35589 ) | ( ~x87 & n35676 ) | ( n35589 & n35676 ) ;
  assign n35678 = ~x87 & n35677 ;
  assign n35679 = ( x75 & ~n35586 ) | ( x75 & n35678 ) | ( ~n35586 & n35678 ) ;
  assign n35680 = n35586 | n35679 ;
  assign n35681 = ( x75 & n6256 ) | ( x75 & n35588 ) | ( n6256 & n35588 ) ;
  assign n35682 = ( x92 & n35680 ) | ( x92 & ~n35681 ) | ( n35680 & ~n35681 ) ;
  assign n35683 = ~x92 & n35682 ;
  assign n35684 = ( x54 & ~n35585 ) | ( x54 & n35683 ) | ( ~n35585 & n35683 ) ;
  assign n35685 = n35585 | n35684 ;
  assign n35686 = ( x74 & ~n35584 ) | ( x74 & n35685 ) | ( ~n35584 & n35685 ) ;
  assign n35687 = ~x74 & n35686 ;
  assign n35688 = x74 & ~n5009 ;
  assign n35689 = n35579 & n35688 ;
  assign n35690 = x55 | n35689 ;
  assign n35691 = ( ~n6250 & n35687 ) | ( ~n6250 & n35690 ) | ( n35687 & n35690 ) ;
  assign n35692 = ~n6250 & n35691 ;
  assign n35693 = x56 & ~n2098 ;
  assign n35694 = n35579 & n35693 ;
  assign n35695 = ( ~x62 & n35692 ) | ( ~x62 & n35694 ) | ( n35692 & n35694 ) ;
  assign n35696 = ~x62 & n35695 ;
  assign n35697 = x62 & n35580 ;
  assign n35698 = n2120 | n35697 ;
  assign n35699 = ( ~n35582 & n35696 ) | ( ~n35582 & n35698 ) | ( n35696 & n35698 ) ;
  assign n35700 = ~n35582 & n35699 ;
  assign n35701 = x228 & x231 ;
  assign n35702 = x62 & ~n35701 ;
  assign n35703 = n6352 & n35702 ;
  assign n35704 = x55 & ~n35701 ;
  assign n35705 = n6337 & ~n35701 ;
  assign n35706 = x74 & ~n35705 ;
  assign n35707 = x54 & ~n35701 ;
  assign n35708 = ( ~x70 & n1401 ) | ( ~x70 & n1722 ) | ( n1401 & n1722 ) ;
  assign n35709 = x51 | n35708 ;
  assign n35710 = ~n1435 & n35709 ;
  assign n35711 = ( ~n1433 & n1773 ) | ( ~n1433 & n35710 ) | ( n1773 & n35710 ) ;
  assign n35712 = ~n1433 & n35711 ;
  assign n35713 = ( x32 & n1586 ) | ( x32 & ~n35712 ) | ( n1586 & ~n35712 ) ;
  assign n35714 = n35712 | n35713 ;
  assign n35715 = n35714 ^ n5167 ^ 1'b0 ;
  assign n35716 = ( n5167 & n35714 ) | ( n5167 & n35715 ) | ( n35714 & n35715 ) ;
  assign n35717 = ( x95 & ~n5167 ) | ( x95 & n35716 ) | ( ~n5167 & n35716 ) ;
  assign n35718 = n35717 ^ n1648 ^ 1'b0 ;
  assign n35719 = ( n1648 & n35717 ) | ( n1648 & n35718 ) | ( n35717 & n35718 ) ;
  assign n35720 = ( x39 & ~n1648 ) | ( x39 & n35719 ) | ( ~n1648 & n35719 ) ;
  assign n35721 = ( x38 & ~n2217 ) | ( x38 & n35720 ) | ( ~n2217 & n35720 ) ;
  assign n35722 = ~x38 & n35721 ;
  assign n35723 = ~x228 & n35722 ;
  assign n35724 = ( ~x100 & n35701 ) | ( ~x100 & n35723 ) | ( n35701 & n35723 ) ;
  assign n35725 = ~x100 & n35724 ;
  assign n35726 = n12524 & ~n35701 ;
  assign n35727 = x100 & ~n35726 ;
  assign n35728 = ( x87 & ~n35725 ) | ( x87 & n35727 ) | ( ~n35725 & n35727 ) ;
  assign n35729 = n35725 | n35728 ;
  assign n35730 = x87 & ~n35701 ;
  assign n35731 = n6323 & n35730 ;
  assign n35732 = ( x75 & n35729 ) | ( x75 & ~n35731 ) | ( n35729 & ~n35731 ) ;
  assign n35733 = ~x75 & n35732 ;
  assign n35734 = n12532 & ~n35701 ;
  assign n35735 = x75 & ~n35734 ;
  assign n35736 = ( x92 & ~n35733 ) | ( x92 & n35735 ) | ( ~n35733 & n35735 ) ;
  assign n35737 = n35733 | n35736 ;
  assign n35738 = x92 & ~n35701 ;
  assign n35739 = n6331 & n35738 ;
  assign n35740 = ( x54 & n35737 ) | ( x54 & ~n35739 ) | ( n35737 & ~n35739 ) ;
  assign n35741 = n35740 ^ n35737 ^ 1'b0 ;
  assign n35742 = ( x54 & n35740 ) | ( x54 & ~n35741 ) | ( n35740 & ~n35741 ) ;
  assign n35743 = ( x74 & ~n35707 ) | ( x74 & n35742 ) | ( ~n35707 & n35742 ) ;
  assign n35744 = ~x74 & n35743 ;
  assign n35745 = ( x55 & ~n35706 ) | ( x55 & n35744 ) | ( ~n35706 & n35744 ) ;
  assign n35746 = n35706 | n35745 ;
  assign n35747 = ( x56 & ~n35704 ) | ( x56 & n35746 ) | ( ~n35704 & n35746 ) ;
  assign n35748 = ~x56 & n35747 ;
  assign n35749 = n6347 & ~n35701 ;
  assign n35750 = x56 & ~n35749 ;
  assign n35751 = x62 | n35750 ;
  assign n35752 = ( ~n35703 & n35748 ) | ( ~n35703 & n35751 ) | ( n35748 & n35751 ) ;
  assign n35753 = ~n35703 & n35752 ;
  assign n35754 = n35701 ^ n2120 ^ 1'b0 ;
  assign n35755 = ( n35701 & n35753 ) | ( n35701 & ~n35754 ) | ( n35753 & ~n35754 ) ;
  assign n35756 = x58 | n5261 ;
  assign n35757 = ~n1408 & n9656 ;
  assign n35758 = n9654 & n35757 ;
  assign n35759 = x91 | n1448 ;
  assign n35760 = ~n5020 & n9646 ;
  assign n35761 = ( ~n35758 & n35759 ) | ( ~n35758 & n35760 ) | ( n35759 & n35760 ) ;
  assign n35762 = n35758 | n35761 ;
  assign n35763 = ( n1378 & ~n35756 ) | ( n1378 & n35762 ) | ( ~n35756 & n35762 ) ;
  assign n35764 = ~n1378 & n35763 ;
  assign n35765 = x72 | n35764 ;
  assign n35766 = ~n13121 & n35765 ;
  assign n35767 = ( x829 & n5063 ) | ( x829 & ~n35766 ) | ( n5063 & ~n35766 ) ;
  assign n35768 = ~n5063 & n35767 ;
  assign n35769 = n1378 | n35756 ;
  assign n35770 = n9646 & ~n35769 ;
  assign n35771 = n35759 & ~n35769 ;
  assign n35772 = x72 | n35771 ;
  assign n35773 = n35770 | n35772 ;
  assign n35774 = ~n13121 & n35773 ;
  assign n35775 = n8671 & ~n35774 ;
  assign n35776 = n11569 & n11611 ;
  assign n35777 = ~n13121 & n35776 ;
  assign n35778 = ( x1093 & n5378 ) | ( x1093 & n35777 ) | ( n5378 & n35777 ) ;
  assign n35779 = n35777 ^ n5378 ^ 1'b0 ;
  assign n35780 = ( x1093 & n35778 ) | ( x1093 & n35779 ) | ( n35778 & n35779 ) ;
  assign n35781 = ~n6425 & n35770 ;
  assign n35782 = n7449 | n35772 ;
  assign n35783 = ( ~n13121 & n35781 ) | ( ~n13121 & n35782 ) | ( n35781 & n35782 ) ;
  assign n35784 = ~n13121 & n35783 ;
  assign n35785 = ( ~n35775 & n35780 ) | ( ~n35775 & n35784 ) | ( n35780 & n35784 ) ;
  assign n35786 = ~n35775 & n35785 ;
  assign n35787 = n35786 ^ n35768 ^ 1'b0 ;
  assign n35788 = ( n35768 & n35786 ) | ( n35768 & n35787 ) | ( n35786 & n35787 ) ;
  assign n35789 = ( x39 & ~n35768 ) | ( x39 & n35788 ) | ( ~n35768 & n35788 ) ;
  assign n35790 = ( n9901 & ~n10109 ) | ( n9901 & n35789 ) | ( ~n10109 & n35789 ) ;
  assign n35791 = ~n9901 & n35790 ;
  assign n35792 = x39 | x95 ;
  assign n35793 = x32 | n35792 ;
  assign n35794 = n7450 | n8670 ;
  assign n35795 = ~n35793 & n35794 ;
  assign n35796 = ( n1417 & n10125 ) | ( n1417 & n35795 ) | ( n10125 & n35795 ) ;
  assign n35797 = ~n1417 & n35796 ;
  assign n35798 = n10055 | n10058 ;
  assign n35799 = ( ~x39 & n5371 ) | ( ~x39 & n35798 ) | ( n5371 & n35798 ) ;
  assign n35800 = x39 & n35799 ;
  assign n35801 = ( ~n9901 & n35797 ) | ( ~n9901 & n35800 ) | ( n35797 & n35800 ) ;
  assign n35802 = ~n9901 & n35801 ;
  assign n35803 = ( ~x39 & x228 ) | ( ~x39 & n35802 ) | ( x228 & n35802 ) ;
  assign n35804 = n35802 ^ x39 ^ 1'b0 ;
  assign n35805 = ( n35802 & n35803 ) | ( n35802 & ~n35804 ) | ( n35803 & ~n35804 ) ;
  assign n35816 = n1292 ^ x120 ^ 1'b0 ;
  assign n35817 = n5021 & n6422 ;
  assign n35818 = ~n15409 & n35817 ;
  assign n35819 = n15334 | n35817 ;
  assign n35820 = ( x1091 & n35818 ) | ( x1091 & n35819 ) | ( n35818 & n35819 ) ;
  assign n35821 = ~n35818 & n35820 ;
  assign n35822 = n5365 | n15334 ;
  assign n35823 = n5365 & ~n15409 ;
  assign n35824 = x1091 | n35823 ;
  assign n35825 = ( n35821 & n35822 ) | ( n35821 & ~n35824 ) | ( n35822 & ~n35824 ) ;
  assign n35826 = n35825 ^ n35822 ^ 1'b0 ;
  assign n35827 = ( n35821 & n35825 ) | ( n35821 & ~n35826 ) | ( n35825 & ~n35826 ) ;
  assign n35828 = ( n1292 & ~n35816 ) | ( n1292 & n35827 ) | ( ~n35816 & n35827 ) ;
  assign n35829 = n15336 ^ n5099 ^ 1'b0 ;
  assign n35830 = ( n15336 & n35828 ) | ( n15336 & n35829 ) | ( n35828 & n35829 ) ;
  assign n35841 = ~n5061 & n35830 ;
  assign n35832 = n15336 ^ n5083 ^ 1'b0 ;
  assign n35833 = ( n15336 & n35828 ) | ( n15336 & ~n35832 ) | ( n35828 & ~n35832 ) ;
  assign n35842 = n5061 & n35833 ;
  assign n35843 = ( n2263 & n35841 ) | ( n2263 & ~n35842 ) | ( n35841 & ~n35842 ) ;
  assign n35844 = ~n35841 & n35843 ;
  assign n35845 = ( x215 & n15592 ) | ( x215 & ~n35844 ) | ( n15592 & ~n35844 ) ;
  assign n35846 = ~x215 & n35845 ;
  assign n35806 = x120 & n5074 ;
  assign n35807 = ~n5083 & n35806 ;
  assign n35808 = n15336 | n35807 ;
  assign n35847 = n5061 & ~n35808 ;
  assign n35810 = n5099 & n35806 ;
  assign n35811 = n15336 | n35810 ;
  assign n35848 = n5061 | n35811 ;
  assign n35849 = ( x215 & n35847 ) | ( x215 & n35848 ) | ( n35847 & n35848 ) ;
  assign n35850 = ~n35847 & n35849 ;
  assign n35851 = ( x299 & n35846 ) | ( x299 & ~n35850 ) | ( n35846 & ~n35850 ) ;
  assign n35852 = ~n35846 & n35851 ;
  assign n35809 = n5114 & ~n35808 ;
  assign n35812 = n5114 | n35811 ;
  assign n35813 = ( x223 & n35809 ) | ( x223 & n35812 ) | ( n35809 & n35812 ) ;
  assign n35814 = ~n35809 & n35813 ;
  assign n35815 = n1359 | n15336 ;
  assign n35831 = ~n5114 & n35830 ;
  assign n35834 = n5114 & n35833 ;
  assign n35835 = ( n1359 & n35831 ) | ( n1359 & ~n35834 ) | ( n35831 & ~n35834 ) ;
  assign n35836 = ~n35831 & n35835 ;
  assign n35837 = ( x223 & n35815 ) | ( x223 & ~n35836 ) | ( n35815 & ~n35836 ) ;
  assign n35838 = ~x223 & n35837 ;
  assign n35839 = ( x299 & ~n35814 ) | ( x299 & n35838 ) | ( ~n35814 & n35838 ) ;
  assign n35840 = n35814 | n35839 ;
  assign n35853 = n35852 ^ n35840 ^ 1'b0 ;
  assign n35854 = ( x39 & ~n35840 ) | ( x39 & n35852 ) | ( ~n35840 & n35852 ) ;
  assign n35855 = ( x39 & ~n35853 ) | ( x39 & n35854 ) | ( ~n35853 & n35854 ) ;
  assign n35856 = n5165 | n5367 ;
  assign n35857 = ~n6425 & n15278 ;
  assign n35858 = n15320 | n35857 ;
  assign n35859 = ~n35856 & n35858 ;
  assign n35860 = n5020 & ~n5367 ;
  assign n35861 = x824 & ~n15304 ;
  assign n35862 = x829 & x1091 ;
  assign n35863 = n15308 & n35862 ;
  assign n35864 = x824 | n35863 ;
  assign n35865 = n35862 & ~n35864 ;
  assign n35866 = n35861 | n35865 ;
  assign n35867 = n35860 & n35866 ;
  assign n35868 = ~n5367 & n35864 ;
  assign n35869 = ~n35861 & n35868 ;
  assign n35870 = n15278 | n35869 ;
  assign n35871 = ( n35856 & n35867 ) | ( n35856 & n35870 ) | ( n35867 & n35870 ) ;
  assign n35872 = ~n35867 & n35871 ;
  assign n35873 = ( x1093 & n35859 ) | ( x1093 & ~n35872 ) | ( n35859 & ~n35872 ) ;
  assign n35874 = ~n35859 & n35873 ;
  assign n35875 = n5160 | n15257 ;
  assign n35876 = n15264 & ~n35875 ;
  assign n35877 = x40 | n35876 ;
  assign n35878 = n35877 ^ n8890 ^ 1'b0 ;
  assign n35879 = ( x252 & n8890 ) | ( x252 & ~n35877 ) | ( n8890 & ~n35877 ) ;
  assign n35880 = ( x252 & ~n35878 ) | ( x252 & n35879 ) | ( ~n35878 & n35879 ) ;
  assign n35881 = n15274 ^ n8890 ^ 1'b0 ;
  assign n35882 = ( n8890 & n15274 ) | ( n8890 & n35881 ) | ( n15274 & n35881 ) ;
  assign n35883 = ( x252 & ~n8890 ) | ( x252 & n35882 ) | ( ~n8890 & n35882 ) ;
  assign n35884 = n5022 & n35883 ;
  assign n35885 = n35884 ^ n35880 ^ 1'b0 ;
  assign n35886 = ( n35880 & n35884 ) | ( n35880 & n35885 ) | ( n35884 & n35885 ) ;
  assign n35887 = ( x1093 & ~n35880 ) | ( x1093 & n35886 ) | ( ~n35880 & n35886 ) ;
  assign n35888 = ( ~n5022 & n15278 ) | ( ~n5022 & n35887 ) | ( n15278 & n35887 ) ;
  assign n35889 = n35887 ^ n5022 ^ 1'b0 ;
  assign n35890 = ( n35887 & n35888 ) | ( n35887 & ~n35889 ) | ( n35888 & ~n35889 ) ;
  assign n35891 = ( x39 & ~n35874 ) | ( x39 & n35890 ) | ( ~n35874 & n35890 ) ;
  assign n35892 = ~x39 & n35891 ;
  assign n35893 = ( x38 & ~n35855 ) | ( x38 & n35892 ) | ( ~n35855 & n35892 ) ;
  assign n35894 = n35855 | n35893 ;
  assign n35895 = ( n5053 & ~n8793 ) | ( n5053 & n35894 ) | ( ~n8793 & n35894 ) ;
  assign n35896 = ~n5053 & n35895 ;
  assign n35897 = n5020 & n5065 ;
  assign n35898 = n5363 & n35897 ;
  assign n35899 = ( ~n5083 & n6261 ) | ( ~n5083 & n6263 ) | ( n6261 & n6263 ) ;
  assign n35900 = n35898 & n35899 ;
  assign n35901 = n5070 & n10004 ;
  assign n35902 = n35901 ^ n35900 ^ 1'b0 ;
  assign n35903 = ( n35900 & n35901 ) | ( n35900 & n35902 ) | ( n35901 & n35902 ) ;
  assign n35904 = ( n2217 & ~n35900 ) | ( n2217 & n35903 ) | ( ~n35900 & n35903 ) ;
  assign n35905 = x81 | n1544 ;
  assign n35906 = ~n5208 & n35905 ;
  assign n35907 = n1226 | n35906 ;
  assign n35908 = ~n14213 & n35907 ;
  assign n35909 = ( ~n1469 & n1471 ) | ( ~n1469 & n35908 ) | ( n1471 & n35908 ) ;
  assign n35910 = ~n1469 & n35909 ;
  assign n35911 = ( n1386 & ~n1389 ) | ( n1386 & n35910 ) | ( ~n1389 & n35910 ) ;
  assign n35912 = ~n1389 & n35911 ;
  assign n35913 = x86 | n35912 ;
  assign n35914 = ~n1564 & n35913 ;
  assign n35915 = ( ~n1462 & n1467 ) | ( ~n1462 & n35914 ) | ( n1467 & n35914 ) ;
  assign n35916 = ~n1462 & n35915 ;
  assign n35917 = x108 | n35916 ;
  assign n35918 = ~n1704 & n35917 ;
  assign n35919 = ( ~n1703 & n1841 ) | ( ~n1703 & n35918 ) | ( n1841 & n35918 ) ;
  assign n35920 = ~n1703 & n35919 ;
  assign n35921 = n1452 | n35920 ;
  assign n35922 = ~n1451 & n35921 ;
  assign n35923 = n1444 | n35922 ;
  assign n35924 = ~n1702 & n35923 ;
  assign n35925 = n1268 | n35924 ;
  assign n35926 = ~n14212 & n35925 ;
  assign n35927 = x70 | n35926 ;
  assign n35928 = ~n1693 & n35927 ;
  assign n35929 = x51 | n35928 ;
  assign n35930 = ~n1435 & n35929 ;
  assign n35931 = ( ~n1433 & n1773 ) | ( ~n1433 & n35930 ) | ( n1773 & n35930 ) ;
  assign n35932 = ~n1433 & n35931 ;
  assign n35933 = ~x1082 & n1586 ;
  assign n35934 = x32 | n35933 ;
  assign n35935 = ( ~n1381 & n35932 ) | ( ~n1381 & n35934 ) | ( n35932 & n35934 ) ;
  assign n35936 = ~n1381 & n35935 ;
  assign n35937 = x95 | n35936 ;
  assign n35938 = ( ~x95 & n1785 ) | ( ~x95 & n35937 ) | ( n1785 & n35937 ) ;
  assign n35939 = ( x39 & ~n35904 ) | ( x39 & n35938 ) | ( ~n35904 & n35938 ) ;
  assign n35940 = ~n35904 & n35939 ;
  assign n35941 = x38 | n35940 ;
  assign n35942 = ~n5054 & n35941 ;
  assign n35943 = x87 | n5019 ;
  assign n35944 = ( ~n5013 & n35942 ) | ( ~n5013 & n35943 ) | ( n35942 & n35943 ) ;
  assign n35945 = ~n5013 & n35944 ;
  assign n35946 = ( x75 & x92 ) | ( x75 & ~n35945 ) | ( x92 & ~n35945 ) ;
  assign n35947 = n35945 | n35946 ;
  assign n35948 = ( x54 & ~n6258 ) | ( x54 & n35947 ) | ( ~n6258 & n35947 ) ;
  assign n35949 = ~x54 & n35948 ;
  assign n35950 = n6253 & ~n35949 ;
  assign n35951 = ( x54 & n35949 ) | ( x54 & ~n35950 ) | ( n35949 & ~n35950 ) ;
  assign n35952 = n7447 | n35951 ;
  assign n35953 = ~n14290 & n35952 ;
  assign n35954 = x56 | n35953 ;
  assign n35955 = ~n5008 & n35954 ;
  assign n35956 = x62 | n35955 ;
  assign n35957 = ~n5005 & n35956 ;
  assign n35958 = n2120 | n35957 ;
  assign n35959 = ~n5190 & n35958 ;
  assign n35960 = ~x211 & x1156 ;
  assign n35961 = x211 & x1155 ;
  assign n35962 = n35960 | n35961 ;
  assign n35963 = ~x211 & x1155 ;
  assign n35964 = x211 & x1154 ;
  assign n35965 = n35963 | n35964 ;
  assign n35966 = n35962 ^ x214 ^ 1'b0 ;
  assign n35967 = ( n35962 & n35965 ) | ( n35962 & n35966 ) | ( n35965 & n35966 ) ;
  assign n35968 = x212 & n35967 ;
  assign n35969 = x211 & x1156 ;
  assign n35970 = ~x211 & x1157 ;
  assign n35971 = n35969 | n35970 ;
  assign n35972 = x214 & n35971 ;
  assign n35973 = ~x212 & n35972 ;
  assign n35974 = n35968 | n35973 ;
  assign n35975 = x219 | n35974 ;
  assign n35976 = n35975 ^ x213 ^ 1'b0 ;
  assign n35977 = ~x211 & x214 ;
  assign n35978 = x1155 & n35977 ;
  assign n35979 = x212 | n35978 ;
  assign n35980 = ~x211 & x1153 ;
  assign n35981 = n9344 & ~n35980 ;
  assign n35982 = ~x211 & x1154 ;
  assign n35983 = x214 | n35982 ;
  assign n35984 = ~n35981 & n35983 ;
  assign n35985 = x219 & ~n35984 ;
  assign n35986 = ( x219 & ~n35979 ) | ( x219 & n35985 ) | ( ~n35979 & n35985 ) ;
  assign n35987 = ( x57 & n5193 ) | ( x57 & ~n35986 ) | ( n5193 & ~n35986 ) ;
  assign n35988 = ~n35986 & n35987 ;
  assign n35989 = ( n35975 & ~n35976 ) | ( n35975 & n35988 ) | ( ~n35976 & n35988 ) ;
  assign n35990 = ( x213 & n35976 ) | ( x213 & n35989 ) | ( n35976 & n35989 ) ;
  assign n35991 = x199 & x1142 ;
  assign n35992 = x200 | n35991 ;
  assign n35993 = ~x199 & x1144 ;
  assign n35994 = n35992 | n35993 ;
  assign n35995 = ~x199 & x1143 ;
  assign n35996 = x200 & ~n35995 ;
  assign n35997 = n35994 & ~n35996 ;
  assign n35998 = x299 | n35997 ;
  assign n35999 = ~x207 & n35998 ;
  assign n36000 = x207 & ~x299 ;
  assign n36001 = ~x199 & x1142 ;
  assign n36002 = x200 & ~n36001 ;
  assign n36003 = n36000 & ~n36002 ;
  assign n36004 = n35992 | n35995 ;
  assign n36005 = n36003 & n36004 ;
  assign n36006 = ( x208 & n35999 ) | ( x208 & n36005 ) | ( n35999 & n36005 ) ;
  assign n36007 = n36005 ^ n35999 ^ 1'b0 ;
  assign n36008 = ( x208 & n36006 ) | ( x208 & n36007 ) | ( n36006 & n36007 ) ;
  assign n36009 = x207 & ~x208 ;
  assign n36010 = n36008 ^ n35997 ^ 1'b0 ;
  assign n36011 = ( ~n35997 & n36009 ) | ( ~n35997 & n36010 ) | ( n36009 & n36010 ) ;
  assign n36012 = ( n35997 & n36008 ) | ( n35997 & n36011 ) | ( n36008 & n36011 ) ;
  assign n36013 = ~x299 & n36012 ;
  assign n36014 = ~x212 & x214 ;
  assign n36015 = x299 & x1153 ;
  assign n36016 = x214 & ~n36015 ;
  assign n36017 = x299 & x1154 ;
  assign n36018 = x214 | n36017 ;
  assign n36019 = ( x212 & n36016 ) | ( x212 & n36018 ) | ( n36016 & n36018 ) ;
  assign n36020 = ~n36016 & n36019 ;
  assign n36021 = x299 & x1155 ;
  assign n36022 = ( x299 & n36020 ) | ( x299 & n36021 ) | ( n36020 & n36021 ) ;
  assign n36023 = ( n36014 & n36020 ) | ( n36014 & n36022 ) | ( n36020 & n36022 ) ;
  assign n36024 = ( x211 & x219 ) | ( x211 & n36023 ) | ( x219 & n36023 ) ;
  assign n36025 = ~x211 & n36024 ;
  assign n36026 = ~x219 & x299 ;
  assign n36027 = n36025 ^ n35974 ^ 1'b0 ;
  assign n36028 = ( ~n35974 & n36026 ) | ( ~n35974 & n36027 ) | ( n36026 & n36027 ) ;
  assign n36029 = ( n35974 & n36025 ) | ( n35974 & n36028 ) | ( n36025 & n36028 ) ;
  assign n36030 = ( ~n7318 & n36013 ) | ( ~n7318 & n36029 ) | ( n36013 & n36029 ) ;
  assign n36031 = ~n7318 & n36030 ;
  assign n36032 = ( x209 & n35990 ) | ( x209 & n36031 ) | ( n35990 & n36031 ) ;
  assign n36033 = n36031 ^ n35990 ^ 1'b0 ;
  assign n36034 = ( x209 & n36032 ) | ( x209 & n36033 ) | ( n36032 & n36033 ) ;
  assign n36035 = x212 | x214 ;
  assign n36036 = ~x211 & n36035 ;
  assign n36037 = x219 & ~n36036 ;
  assign n36038 = n7318 & ~n36037 ;
  assign n36039 = x299 | n36012 ;
  assign n36040 = x299 & ~x1142 ;
  assign n36041 = n36036 & ~n36040 ;
  assign n36042 = n36039 & n36041 ;
  assign n36043 = n36013 & ~n36036 ;
  assign n36044 = ( x219 & n36042 ) | ( x219 & ~n36043 ) | ( n36042 & ~n36043 ) ;
  assign n36045 = ~n36042 & n36044 ;
  assign n36046 = ~x211 & x1143 ;
  assign n36047 = x299 & x1142 ;
  assign n36048 = x299 & x1143 ;
  assign n36049 = x211 | n36048 ;
  assign n36050 = ( n36046 & n36047 ) | ( n36046 & n36049 ) | ( n36047 & n36049 ) ;
  assign n36051 = x214 & ~n36050 ;
  assign n36052 = ~n36013 & n36051 ;
  assign n36053 = x211 & x1143 ;
  assign n36054 = ~x211 & x1144 ;
  assign n36055 = n36053 | n36054 ;
  assign n36056 = x299 & n36055 ;
  assign n36057 = x214 | n36013 ;
  assign n36058 = n36056 | n36057 ;
  assign n36059 = ( x212 & n36052 ) | ( x212 & n36058 ) | ( n36052 & n36058 ) ;
  assign n36060 = ~n36052 & n36059 ;
  assign n36061 = n36013 | n36056 ;
  assign n36062 = ~x212 & n36057 ;
  assign n36063 = n36061 & n36062 ;
  assign n36064 = ( x219 & ~n36060 ) | ( x219 & n36063 ) | ( ~n36060 & n36063 ) ;
  assign n36065 = n36060 | n36064 ;
  assign n36066 = ( n7318 & ~n36045 ) | ( n7318 & n36065 ) | ( ~n36045 & n36065 ) ;
  assign n36067 = ~n7318 & n36066 ;
  assign n36068 = n9344 & n36046 ;
  assign n36069 = x214 ^ x212 ^ 1'b0 ;
  assign n36070 = n36055 & n36069 ;
  assign n36071 = ( ~x219 & n36068 ) | ( ~x219 & n36070 ) | ( n36068 & n36070 ) ;
  assign n36072 = ~x219 & n36071 ;
  assign n36073 = n36072 ^ x1142 ^ 1'b0 ;
  assign n36074 = ( ~x1142 & n9275 ) | ( ~x1142 & n36073 ) | ( n9275 & n36073 ) ;
  assign n36075 = ( x1142 & n36072 ) | ( x1142 & n36074 ) | ( n36072 & n36074 ) ;
  assign n36076 = n36067 ^ n36038 ^ 1'b0 ;
  assign n36077 = ( ~n36038 & n36075 ) | ( ~n36038 & n36076 ) | ( n36075 & n36076 ) ;
  assign n36078 = ( n36038 & n36067 ) | ( n36038 & n36077 ) | ( n36067 & n36077 ) ;
  assign n36079 = n36078 ^ n36034 ^ 1'b0 ;
  assign n36080 = ( ~x213 & n36078 ) | ( ~x213 & n36079 ) | ( n36078 & n36079 ) ;
  assign n36081 = ( n36034 & ~n36079 ) | ( n36034 & n36080 ) | ( ~n36079 & n36080 ) ;
  assign n36082 = ~x200 & x1155 ;
  assign n36083 = x199 & n36082 ;
  assign n36084 = ~x299 & n36083 ;
  assign n36085 = x1156 | n36084 ;
  assign n36086 = x200 | x1155 ;
  assign n36087 = x199 & x200 ;
  assign n36088 = n9353 & ~n36087 ;
  assign n36089 = ~x299 & n36088 ;
  assign n36090 = n36086 & n36089 ;
  assign n36091 = n36085 & n36090 ;
  assign n36092 = x207 & n36091 ;
  assign n36093 = ~x208 & n36092 ;
  assign n36106 = x200 | x299 ;
  assign n36107 = x199 & ~x1153 ;
  assign n36108 = n36106 | n36107 ;
  assign n36109 = x199 | x1155 ;
  assign n36110 = ~x1154 & n36109 ;
  assign n36111 = ~n36108 & n36110 ;
  assign n36112 = x299 | n36087 ;
  assign n36113 = x1153 & n36112 ;
  assign n36114 = x1154 & ~n36113 ;
  assign n36115 = ~n10019 & n36082 ;
  assign n36116 = ~x1153 & n10019 ;
  assign n36117 = x1154 & n36088 ;
  assign n36118 = ~n36116 & n36117 ;
  assign n36119 = n36115 | n36118 ;
  assign n36120 = n36114 & n36119 ;
  assign n36121 = n36111 | n36120 ;
  assign n36122 = x207 & ~n36121 ;
  assign n36094 = x200 & ~x299 ;
  assign n36095 = ~x199 & x1155 ;
  assign n36096 = n36094 & n36095 ;
  assign n36097 = x1154 | n36096 ;
  assign n36098 = x200 & ~n36095 ;
  assign n36099 = n9354 & ~n36098 ;
  assign n36100 = n36097 & n36099 ;
  assign n36101 = x200 & ~x1155 ;
  assign n36102 = n10019 | n36101 ;
  assign n36103 = x1156 & ~n36102 ;
  assign n36104 = n36100 | n36103 ;
  assign n36105 = x207 & ~n36104 ;
  assign n36123 = n36122 ^ n36105 ^ n36104 ;
  assign n36124 = x208 & n36123 ;
  assign n36125 = ( x1157 & ~n36093 ) | ( x1157 & n36124 ) | ( ~n36093 & n36124 ) ;
  assign n36126 = n36093 | n36125 ;
  assign n36127 = x199 & ~x1155 ;
  assign n36128 = x1156 & ~n36127 ;
  assign n36129 = ~n36112 & n36128 ;
  assign n36130 = x1156 | n36127 ;
  assign n36131 = n36106 | n36130 ;
  assign n36132 = ~n36129 & n36131 ;
  assign n36133 = x207 & ~n36132 ;
  assign n36134 = ~x208 & n36133 ;
  assign n36135 = ( x1157 & n36124 ) | ( x1157 & ~n36134 ) | ( n36124 & ~n36134 ) ;
  assign n36136 = ~n36124 & n36135 ;
  assign n36137 = n36126 & ~n36136 ;
  assign n36239 = x211 & ~n36137 ;
  assign n36138 = x214 | n36137 ;
  assign n36139 = ~x212 & n36138 ;
  assign n36140 = x211 | x214 ;
  assign n36141 = x207 | x299 ;
  assign n36142 = ~x208 & n36141 ;
  assign n36143 = n10008 & ~n36082 ;
  assign n36144 = ~x1155 & n9354 ;
  assign n36145 = ( n9354 & n36094 ) | ( n9354 & n36144 ) | ( n36094 & n36144 ) ;
  assign n36146 = n36145 ^ x1156 ^ 1'b0 ;
  assign n36147 = ( n36143 & n36145 ) | ( n36143 & n36146 ) | ( n36145 & n36146 ) ;
  assign n36148 = x207 & n36147 ;
  assign n36149 = n36142 & ~n36148 ;
  assign n36150 = x299 & ~x1154 ;
  assign n36151 = x1157 & ~n36150 ;
  assign n36152 = n36149 & n36151 ;
  assign n36153 = n36017 | n36092 ;
  assign n36154 = ~x208 & n36153 ;
  assign n36155 = x1157 | n36154 ;
  assign n36156 = ( ~x1157 & n36152 ) | ( ~x1157 & n36155 ) | ( n36152 & n36155 ) ;
  assign n36157 = x1155 & ~n10008 ;
  assign n36158 = n36089 & ~n36107 ;
  assign n36159 = n36157 | n36158 ;
  assign n36160 = x299 | n36159 ;
  assign n36161 = x1154 & n36160 ;
  assign n36162 = n36111 | n36161 ;
  assign n36163 = x207 & n36162 ;
  assign n36164 = x199 & ~x200 ;
  assign n36165 = x299 | n36164 ;
  assign n36166 = x299 | n36088 ;
  assign n36167 = x1155 & n36166 ;
  assign n36168 = ( n36165 & n36166 ) | ( n36165 & n36167 ) | ( n36166 & n36167 ) ;
  assign n36169 = x1154 & n36168 ;
  assign n36170 = n36104 | n36169 ;
  assign n36171 = ~x207 & n36170 ;
  assign n36172 = n36163 | n36171 ;
  assign n36173 = n36156 ^ x208 ^ 1'b0 ;
  assign n36174 = ( ~x208 & n36172 ) | ( ~x208 & n36173 ) | ( n36172 & n36173 ) ;
  assign n36175 = ( x208 & n36156 ) | ( x208 & n36174 ) | ( n36156 & n36174 ) ;
  assign n36176 = n36140 | n36175 ;
  assign n36177 = ( n9354 & n10008 ) | ( n9354 & n36144 ) | ( n10008 & n36144 ) ;
  assign n36178 = x1156 & ~n36177 ;
  assign n36179 = n36169 | n36178 ;
  assign n36180 = x299 & ~x1155 ;
  assign n36181 = x299 | n10073 ;
  assign n36182 = x1155 & n36181 ;
  assign n36183 = n36180 | n36182 ;
  assign n36184 = n36179 | n36183 ;
  assign n36185 = x299 & ~x1153 ;
  assign n36186 = x207 | n36185 ;
  assign n36187 = n36184 & ~n36186 ;
  assign n36188 = ( ~n36116 & n36119 ) | ( ~n36116 & n36165 ) | ( n36119 & n36165 ) ;
  assign n36189 = x207 & n36188 ;
  assign n36190 = ( x208 & n36187 ) | ( x208 & n36189 ) | ( n36187 & n36189 ) ;
  assign n36191 = n36189 ^ n36187 ^ 1'b0 ;
  assign n36192 = ( x208 & n36190 ) | ( x208 & n36191 ) | ( n36190 & n36191 ) ;
  assign n36193 = x1157 & ~n36149 ;
  assign n36194 = x1156 & ~n36083 ;
  assign n36195 = ~n36181 & n36194 ;
  assign n36196 = n36085 & ~n36195 ;
  assign n36197 = x207 & n36196 ;
  assign n36198 = ( ~x208 & x299 ) | ( ~x208 & n36197 ) | ( x299 & n36197 ) ;
  assign n36199 = ~x208 & n36198 ;
  assign n36200 = x1157 | n36199 ;
  assign n36201 = ~n36185 & n36200 ;
  assign n36202 = ~n36193 & n36201 ;
  assign n36203 = ( n35977 & n36192 ) | ( n35977 & ~n36202 ) | ( n36192 & ~n36202 ) ;
  assign n36204 = ~n36192 & n36203 ;
  assign n36205 = x212 & ~n36204 ;
  assign n36206 = n36176 & n36205 ;
  assign n36207 = x207 | n36021 ;
  assign n36208 = ~x208 & n36207 ;
  assign n36209 = ~x1155 & n10019 ;
  assign n36210 = n36166 & ~n36209 ;
  assign n36211 = x299 | n36085 ;
  assign n36212 = n36210 & n36211 ;
  assign n36213 = n36208 & n36212 ;
  assign n36214 = n36104 | n36207 ;
  assign n36215 = x208 & n36214 ;
  assign n36219 = x1155 & ~n36094 ;
  assign n36216 = x299 | n9353 ;
  assign n36217 = ~x1153 & n36216 ;
  assign n36218 = ( n9354 & n36094 ) | ( n9354 & n36217 ) | ( n36094 & n36217 ) ;
  assign n36220 = n36219 ^ n36218 ^ n36145 ;
  assign n36221 = n36220 ^ x1154 ^ 1'b0 ;
  assign n36222 = ( n36159 & n36220 ) | ( n36159 & n36221 ) | ( n36220 & n36221 ) ;
  assign n36223 = x207 & ~n36222 ;
  assign n36224 = n36215 & ~n36223 ;
  assign n36225 = x1156 & ~n10019 ;
  assign n36226 = ( x1156 & n36219 ) | ( x1156 & n36225 ) | ( n36219 & n36225 ) ;
  assign n36227 = ~x1155 & n36165 ;
  assign n36228 = x1156 | n36094 ;
  assign n36229 = ( ~n36226 & n36227 ) | ( ~n36226 & n36228 ) | ( n36227 & n36228 ) ;
  assign n36230 = ~n36226 & n36229 ;
  assign n36231 = x207 & n36230 ;
  assign n36232 = x1157 & n36208 ;
  assign n36233 = ~n36231 & n36232 ;
  assign n36234 = ( ~n36213 & n36224 ) | ( ~n36213 & n36233 ) | ( n36224 & n36233 ) ;
  assign n36235 = n36213 | n36234 ;
  assign n36236 = n35977 & ~n36235 ;
  assign n36237 = ~n36206 & n36236 ;
  assign n36238 = ( n36139 & n36206 ) | ( n36139 & ~n36237 ) | ( n36206 & ~n36237 ) ;
  assign n36240 = n36239 ^ n36238 ^ 1'b0 ;
  assign n36241 = ( x219 & ~n36238 ) | ( x219 & n36239 ) | ( ~n36238 & n36239 ) ;
  assign n36242 = ( x219 & ~n36240 ) | ( x219 & n36241 ) | ( ~n36240 & n36241 ) ;
  assign n36243 = x207 | n36184 ;
  assign n36244 = n36000 & ~n36188 ;
  assign n36245 = x208 & ~n36244 ;
  assign n36246 = n36193 & ~n36245 ;
  assign n36247 = ( n36193 & ~n36243 ) | ( n36193 & n36246 ) | ( ~n36243 & n36246 ) ;
  assign n36248 = ( x211 & n36126 ) | ( x211 & ~n36247 ) | ( n36126 & ~n36247 ) ;
  assign n36249 = ~x211 & n36248 ;
  assign n36250 = ~x208 & x1157 ;
  assign n36251 = x299 & x1156 ;
  assign n36252 = n36133 | n36251 ;
  assign n36253 = n36250 & n36252 ;
  assign n36254 = x207 & n36121 ;
  assign n36255 = n36100 | n36178 ;
  assign n36256 = n36255 ^ x207 ^ 1'b0 ;
  assign n36257 = ( n36251 & n36255 ) | ( n36251 & n36256 ) | ( n36255 & n36256 ) ;
  assign n36258 = n36254 | n36257 ;
  assign n36259 = x208 & n36258 ;
  assign n36260 = n36085 & n36199 ;
  assign n36261 = ( ~n36253 & n36259 ) | ( ~n36253 & n36260 ) | ( n36259 & n36260 ) ;
  assign n36262 = n36253 | n36261 ;
  assign n36263 = x211 & n36262 ;
  assign n36264 = ( x214 & n36249 ) | ( x214 & ~n36263 ) | ( n36249 & ~n36263 ) ;
  assign n36265 = ~n36249 & n36264 ;
  assign n36266 = ( x212 & n36138 ) | ( x212 & ~n36265 ) | ( n36138 & ~n36265 ) ;
  assign n36267 = ~x212 & n36266 ;
  assign n36268 = x219 ^ x212 ^ 1'b0 ;
  assign n36269 = n9271 & n36175 ;
  assign n36270 = ~n36140 & n36262 ;
  assign n36271 = ~n9271 & n36140 ;
  assign n36272 = n36235 & n36271 ;
  assign n36273 = ( ~n36269 & n36270 ) | ( ~n36269 & n36272 ) | ( n36270 & n36272 ) ;
  assign n36274 = n36269 | n36273 ;
  assign n36275 = ( x212 & ~n36268 ) | ( x212 & n36274 ) | ( ~n36268 & n36274 ) ;
  assign n36276 = ( x219 & n36268 ) | ( x219 & n36275 ) | ( n36268 & n36275 ) ;
  assign n36277 = ( ~n7318 & n36267 ) | ( ~n7318 & n36276 ) | ( n36267 & n36276 ) ;
  assign n36278 = ~n7318 & n36277 ;
  assign n36279 = n36278 ^ n36242 ^ 1'b0 ;
  assign n36280 = ( n36242 & n36278 ) | ( n36242 & n36279 ) | ( n36278 & n36279 ) ;
  assign n36281 = ( n35990 & ~n36242 ) | ( n35990 & n36280 ) | ( ~n36242 & n36280 ) ;
  assign n36282 = n36038 & n36075 ;
  assign n36283 = ~n36040 & n36179 ;
  assign n36284 = n36047 | n36096 ;
  assign n36285 = x1154 | x1156 ;
  assign n36286 = ( x207 & n36284 ) | ( x207 & ~n36285 ) | ( n36284 & ~n36285 ) ;
  assign n36287 = n36286 ^ n36284 ^ 1'b0 ;
  assign n36288 = ( x207 & n36286 ) | ( x207 & ~n36287 ) | ( n36286 & ~n36287 ) ;
  assign n36289 = ( x208 & n36283 ) | ( x208 & n36288 ) | ( n36283 & n36288 ) ;
  assign n36290 = n36288 ^ n36283 ^ 1'b0 ;
  assign n36291 = ( x208 & n36289 ) | ( x208 & n36290 ) | ( n36289 & n36290 ) ;
  assign n36292 = ~x299 & n36222 ;
  assign n36293 = n36292 ^ n36291 ^ 1'b0 ;
  assign n36294 = x207 & ~n36047 ;
  assign n36295 = ( n36292 & n36293 ) | ( n36292 & ~n36294 ) | ( n36293 & ~n36294 ) ;
  assign n36296 = ( n36291 & ~n36293 ) | ( n36291 & n36295 ) | ( ~n36293 & n36295 ) ;
  assign n36297 = ~x219 & n36035 ;
  assign n36298 = n36036 | n36297 ;
  assign n36299 = n9275 & n36298 ;
  assign n36300 = ~n36040 & n36200 ;
  assign n36301 = ~n36193 & n36300 ;
  assign n36302 = ( n36296 & n36299 ) | ( n36296 & ~n36301 ) | ( n36299 & ~n36301 ) ;
  assign n36303 = ~n36296 & n36302 ;
  assign n36304 = ( x57 & n5193 ) | ( x57 & ~n36303 ) | ( n5193 & ~n36303 ) ;
  assign n36305 = n36303 | n36304 ;
  assign n36306 = n36137 | n36298 ;
  assign n36307 = ~x211 & n9344 ;
  assign n36308 = ~n36129 & n36145 ;
  assign n36309 = x299 & ~x1143 ;
  assign n36310 = x207 & ~n36309 ;
  assign n36311 = ~n36308 & n36310 ;
  assign n36312 = ( n36048 & n36250 ) | ( n36048 & n36311 ) | ( n36250 & n36311 ) ;
  assign n36313 = n36311 ^ n36048 ^ 1'b0 ;
  assign n36314 = ( n36250 & n36312 ) | ( n36250 & n36313 ) | ( n36312 & n36313 ) ;
  assign n36315 = ~n36048 & n36122 ;
  assign n36316 = x208 & ~n36315 ;
  assign n36320 = ( ~x1154 & n36177 ) | ( ~x1154 & n36309 ) | ( n36177 & n36309 ) ;
  assign n36317 = x299 | n36098 ;
  assign n36318 = x1154 & n36317 ;
  assign n36319 = ~n36048 & n36318 ;
  assign n36321 = ( x1156 & ~n36319 ) | ( x1156 & n36320 ) | ( ~n36319 & n36320 ) ;
  assign n36322 = ~n36320 & n36321 ;
  assign n36323 = ~x1155 & n36048 ;
  assign n36324 = n36167 & ~n36309 ;
  assign n36325 = x1154 & ~n10008 ;
  assign n36326 = ( x1154 & n36086 ) | ( x1154 & n36325 ) | ( n36086 & n36325 ) ;
  assign n36327 = ( n36323 & ~n36324 ) | ( n36323 & n36326 ) | ( ~n36324 & n36326 ) ;
  assign n36328 = ~n36323 & n36327 ;
  assign n36329 = n36048 | n36097 ;
  assign n36330 = ~x1156 & n36329 ;
  assign n36331 = ( n36322 & ~n36328 ) | ( n36322 & n36330 ) | ( ~n36328 & n36330 ) ;
  assign n36332 = n36328 ^ n36322 ^ 1'b0 ;
  assign n36333 = ( n36322 & n36331 ) | ( n36322 & ~n36332 ) | ( n36331 & ~n36332 ) ;
  assign n36334 = x207 | n36333 ;
  assign n36335 = n36316 & n36334 ;
  assign n36336 = ~x1157 & n36199 ;
  assign n36337 = ~n36309 & n36336 ;
  assign n36338 = ( ~n36314 & n36335 ) | ( ~n36314 & n36337 ) | ( n36335 & n36337 ) ;
  assign n36339 = n36314 | n36338 ;
  assign n36340 = n36307 & ~n36339 ;
  assign n36341 = x299 & x1144 ;
  assign n36342 = n36122 & ~n36341 ;
  assign n36344 = x299 & ~x1144 ;
  assign n36345 = ( ~x1154 & n36177 ) | ( ~x1154 & n36344 ) | ( n36177 & n36344 ) ;
  assign n36343 = n36318 & ~n36341 ;
  assign n36346 = ( x1156 & ~n36343 ) | ( x1156 & n36345 ) | ( ~n36343 & n36345 ) ;
  assign n36347 = ~n36345 & n36346 ;
  assign n36348 = ~x1155 & n36341 ;
  assign n36349 = n36167 & ~n36344 ;
  assign n36350 = ( n36326 & n36348 ) | ( n36326 & ~n36349 ) | ( n36348 & ~n36349 ) ;
  assign n36351 = ~n36348 & n36350 ;
  assign n36352 = n36097 | n36341 ;
  assign n36353 = ~x1156 & n36352 ;
  assign n36354 = ( n36347 & ~n36351 ) | ( n36347 & n36353 ) | ( ~n36351 & n36353 ) ;
  assign n36355 = n36351 ^ n36347 ^ 1'b0 ;
  assign n36356 = ( n36347 & n36354 ) | ( n36347 & ~n36355 ) | ( n36354 & ~n36355 ) ;
  assign n36357 = x207 | n36356 ;
  assign n36358 = ( x208 & n36342 ) | ( x208 & n36357 ) | ( n36342 & n36357 ) ;
  assign n36359 = ~n36342 & n36358 ;
  assign n36360 = x207 & ~n36344 ;
  assign n36361 = n36308 | n36360 ;
  assign n36362 = ( ~n36308 & n36341 ) | ( ~n36308 & n36361 ) | ( n36341 & n36361 ) ;
  assign n36363 = ( x208 & x1157 ) | ( x208 & n36362 ) | ( x1157 & n36362 ) ;
  assign n36364 = ~x208 & n36363 ;
  assign n36365 = n36344 & ~n36364 ;
  assign n36366 = ( n36336 & n36364 ) | ( n36336 & ~n36365 ) | ( n36364 & ~n36365 ) ;
  assign n36367 = ( ~x211 & n36359 ) | ( ~x211 & n36366 ) | ( n36359 & n36366 ) ;
  assign n36368 = ~x211 & n36367 ;
  assign n36369 = ~n9344 & n36035 ;
  assign n36370 = x211 & n36339 ;
  assign n36371 = ( n36368 & n36369 ) | ( n36368 & ~n36370 ) | ( n36369 & ~n36370 ) ;
  assign n36372 = ~n36368 & n36371 ;
  assign n36373 = ( ~x219 & n36340 ) | ( ~x219 & n36372 ) | ( n36340 & n36372 ) ;
  assign n36374 = ~x219 & n36373 ;
  assign n36375 = ( n36305 & n36306 ) | ( n36305 & ~n36374 ) | ( n36306 & ~n36374 ) ;
  assign n36376 = ~n36305 & n36375 ;
  assign n36377 = ( x213 & n36282 ) | ( x213 & ~n36376 ) | ( n36282 & ~n36376 ) ;
  assign n36378 = ~n36282 & n36377 ;
  assign n36379 = ( x209 & n36281 ) | ( x209 & ~n36378 ) | ( n36281 & ~n36378 ) ;
  assign n36380 = ~x209 & n36379 ;
  assign n36381 = ( x230 & n36081 ) | ( x230 & n36380 ) | ( n36081 & n36380 ) ;
  assign n36382 = n36380 ^ n36081 ^ 1'b0 ;
  assign n36383 = ( x230 & n36381 ) | ( x230 & n36382 ) | ( n36381 & n36382 ) ;
  assign n36384 = ( x230 & x233 ) | ( x230 & ~n36383 ) | ( x233 & ~n36383 ) ;
  assign n36385 = ~n36383 & n36384 ;
  assign n36386 = x214 & n35962 ;
  assign n36387 = ~x212 & n36386 ;
  assign n36388 = x219 | n36387 ;
  assign n36389 = n35968 | n36388 ;
  assign n36390 = x219 & ~n35982 ;
  assign n36391 = x213 & ~n36390 ;
  assign n36392 = ( ~n36038 & n36389 ) | ( ~n36038 & n36391 ) | ( n36389 & n36391 ) ;
  assign n36393 = n36038 & n36392 ;
  assign n36394 = x207 | x208 ;
  assign n36395 = ~n9233 & n36394 ;
  assign n36396 = x1154 | n36115 ;
  assign n36397 = x199 | n36086 ;
  assign n36398 = ~n36112 & n36397 ;
  assign n36399 = n36396 & n36398 ;
  assign n36400 = x207 & n36399 ;
  assign n36401 = n36395 | n36400 ;
  assign n36402 = n9233 | n36104 ;
  assign n36403 = n36401 & n36402 ;
  assign n36404 = x219 & ~n36403 ;
  assign n36405 = ( x219 & n36036 ) | ( x219 & n36404 ) | ( n36036 & n36404 ) ;
  assign n36406 = x207 & n36170 ;
  assign n36407 = ~x207 & n36017 ;
  assign n36408 = n36406 | n36407 ;
  assign n36409 = ( n36115 & n36166 ) | ( n36115 & n36396 ) | ( n36166 & n36396 ) ;
  assign n36410 = x207 & n36409 ;
  assign n36411 = n36171 | n36410 ;
  assign n36412 = n36408 ^ x208 ^ 1'b0 ;
  assign n36413 = ( n36408 & n36411 ) | ( n36408 & n36412 ) | ( n36411 & n36412 ) ;
  assign n36414 = x211 & n36413 ;
  assign n36415 = n36413 ^ x211 ^ 1'b0 ;
  assign n36416 = ( n36036 & n36414 ) | ( n36036 & n36415 ) | ( n36414 & n36415 ) ;
  assign n36417 = n36405 & ~n36416 ;
  assign n36418 = n33358 & ~n36417 ;
  assign n36419 = x214 | n36403 ;
  assign n36420 = ~x212 & n36419 ;
  assign n36421 = x207 & n36255 ;
  assign n36422 = n36251 | n36421 ;
  assign n36423 = n36257 | n36400 ;
  assign n36424 = n36422 ^ x208 ^ 1'b0 ;
  assign n36425 = ( n36422 & n36423 ) | ( n36422 & n36424 ) | ( n36423 & n36424 ) ;
  assign n36426 = x207 & ~n36021 ;
  assign n36427 = ~n36399 & n36426 ;
  assign n36428 = ( x208 & n36214 ) | ( x208 & n36427 ) | ( n36214 & n36427 ) ;
  assign n36429 = ~n36427 & n36428 ;
  assign n36430 = n36021 | n36104 ;
  assign n36431 = ( n36214 & n36429 ) | ( n36214 & n36430 ) | ( n36429 & n36430 ) ;
  assign n36432 = ( n36208 & n36429 ) | ( n36208 & n36431 ) | ( n36429 & n36431 ) ;
  assign n36433 = n36425 ^ x211 ^ 1'b0 ;
  assign n36434 = ( n36425 & n36432 ) | ( n36425 & n36433 ) | ( n36432 & n36433 ) ;
  assign n36435 = x214 & ~n36434 ;
  assign n36436 = n36420 & ~n36435 ;
  assign n36437 = ~x211 & n36432 ;
  assign n36438 = ( x214 & n36414 ) | ( x214 & ~n36437 ) | ( n36414 & ~n36437 ) ;
  assign n36439 = ~n36414 & n36438 ;
  assign n36440 = x214 | n36434 ;
  assign n36441 = ( x212 & n36439 ) | ( x212 & n36440 ) | ( n36439 & n36440 ) ;
  assign n36442 = ~n36439 & n36441 ;
  assign n36443 = ( x219 & ~n36436 ) | ( x219 & n36442 ) | ( ~n36436 & n36442 ) ;
  assign n36444 = n36436 | n36443 ;
  assign n36445 = n36418 & n36444 ;
  assign n36446 = x1153 & n36140 ;
  assign n36447 = ( ~x214 & n9271 ) | ( ~x214 & n35983 ) | ( n9271 & n35983 ) ;
  assign n36448 = ( x212 & n36446 ) | ( x212 & n36447 ) | ( n36446 & n36447 ) ;
  assign n36449 = n36447 ^ n36446 ^ 1'b0 ;
  assign n36450 = ( x212 & n36448 ) | ( x212 & n36449 ) | ( n36448 & n36449 ) ;
  assign n36451 = x211 & x1153 ;
  assign n36452 = n35982 | n36451 ;
  assign n36453 = n36014 & n36452 ;
  assign n36454 = x219 | n36453 ;
  assign n36455 = n36450 | n36454 ;
  assign n36456 = n36038 & n36455 ;
  assign n36457 = n36000 & ~n36409 ;
  assign n36458 = ( x208 & n36243 ) | ( x208 & n36457 ) | ( n36243 & n36457 ) ;
  assign n36459 = ~n36457 & n36458 ;
  assign n36460 = x207 & ~n36183 ;
  assign n36461 = ~n36179 & n36460 ;
  assign n36462 = ~n36459 & n36461 ;
  assign n36463 = ( n36142 & n36459 ) | ( n36142 & ~n36462 ) | ( n36459 & ~n36462 ) ;
  assign n36464 = n36036 & n36463 ;
  assign n36465 = n36405 & ~n36464 ;
  assign n36466 = ~n36185 & n36463 ;
  assign n36467 = ( n36413 & n36415 ) | ( n36413 & n36466 ) | ( n36415 & n36466 ) ;
  assign n36468 = ~x214 & n36467 ;
  assign n36469 = x211 | n36466 ;
  assign n36470 = x214 & n36469 ;
  assign n36471 = n36463 & n36470 ;
  assign n36472 = n36468 | n36471 ;
  assign n36473 = x212 & n36472 ;
  assign n36474 = x214 & ~n36467 ;
  assign n36475 = n36420 & ~n36474 ;
  assign n36476 = ( x219 & ~n36473 ) | ( x219 & n36475 ) | ( ~n36473 & n36475 ) ;
  assign n36477 = n36473 | n36476 ;
  assign n36478 = ( n7318 & ~n36465 ) | ( n7318 & n36477 ) | ( ~n36465 & n36477 ) ;
  assign n36479 = ~n7318 & n36478 ;
  assign n36480 = ( x1152 & n36456 ) | ( x1152 & ~n36479 ) | ( n36456 & ~n36479 ) ;
  assign n36481 = ~n36456 & n36480 ;
  assign n36482 = x211 & ~n36403 ;
  assign n36483 = n36470 & ~n36482 ;
  assign n36484 = ( x212 & n36468 ) | ( x212 & n36483 ) | ( n36468 & n36483 ) ;
  assign n36485 = n36483 ^ n36468 ^ 1'b0 ;
  assign n36486 = ( x212 & n36484 ) | ( x212 & n36485 ) | ( n36484 & n36485 ) ;
  assign n36487 = ( x219 & n36475 ) | ( x219 & ~n36486 ) | ( n36475 & ~n36486 ) ;
  assign n36488 = n36486 | n36487 ;
  assign n36489 = ( n7318 & ~n36404 ) | ( n7318 & n36488 ) | ( ~n36404 & n36488 ) ;
  assign n36490 = ~n7318 & n36489 ;
  assign n36491 = n9344 | n36452 ;
  assign n36492 = n36297 & n36491 ;
  assign n36493 = ~n35981 & n36492 ;
  assign n36494 = n7318 & n36493 ;
  assign n36495 = ( x1152 & ~n36490 ) | ( x1152 & n36494 ) | ( ~n36490 & n36494 ) ;
  assign n36496 = n36490 | n36495 ;
  assign n36497 = ( x213 & ~n36481 ) | ( x213 & n36496 ) | ( ~n36481 & n36496 ) ;
  assign n36498 = ~x213 & n36497 ;
  assign n36499 = ( x209 & n36445 ) | ( x209 & ~n36498 ) | ( n36445 & ~n36498 ) ;
  assign n36500 = ~n36445 & n36499 ;
  assign n36501 = x213 ^ x209 ^ 1'b0 ;
  assign n36502 = x199 | x1154 ;
  assign n36503 = x200 | n36502 ;
  assign n36504 = n36141 | n36503 ;
  assign n36505 = x200 | x1153 ;
  assign n36506 = ~x199 & n36505 ;
  assign n36507 = x299 | n36506 ;
  assign n36508 = n36164 | n36507 ;
  assign n36509 = x207 & ~n36508 ;
  assign n36510 = x208 & ~n36509 ;
  assign n36511 = ~x199 & x1153 ;
  assign n36512 = x200 & n36511 ;
  assign n36513 = ~x299 & n36512 ;
  assign n36514 = x1154 | n36513 ;
  assign n36515 = x1154 & n36094 ;
  assign n36516 = ~n36511 & n36515 ;
  assign n36517 = n36514 & ~n36516 ;
  assign n36518 = n36165 | n36517 ;
  assign n36519 = x207 | n36518 ;
  assign n36520 = n36510 & n36519 ;
  assign n36521 = n36208 & n36518 ;
  assign n36522 = n36520 | n36521 ;
  assign n36523 = ( n36180 & n36504 ) | ( n36180 & n36522 ) | ( n36504 & n36522 ) ;
  assign n36524 = ~n36180 & n36523 ;
  assign n36525 = ~x211 & n36524 ;
  assign n36526 = n36114 & ~n36217 ;
  assign n36527 = x199 | x1153 ;
  assign n36528 = n36089 & n36527 ;
  assign n36529 = n36526 | n36528 ;
  assign n36530 = x207 & n36529 ;
  assign n36531 = n36017 | n36530 ;
  assign n36532 = x1154 & ~n9354 ;
  assign n36533 = n36526 | n36532 ;
  assign n36534 = n36528 | n36533 ;
  assign n36535 = ~x207 & n36534 ;
  assign n36536 = x207 & n36508 ;
  assign n36537 = ~n36150 & n36536 ;
  assign n36538 = n36535 | n36537 ;
  assign n36539 = n36531 ^ x208 ^ 1'b0 ;
  assign n36540 = ( n36531 & n36538 ) | ( n36531 & n36539 ) | ( n36538 & n36539 ) ;
  assign n36541 = x211 & n36540 ;
  assign n36542 = ( n9344 & n36525 ) | ( n9344 & ~n36541 ) | ( n36525 & ~n36541 ) ;
  assign n36543 = ~n36525 & n36542 ;
  assign n36544 = x211 & n36524 ;
  assign n36545 = n36251 | n36529 ;
  assign n36546 = ~x207 & n36545 ;
  assign n36547 = x299 & ~x1156 ;
  assign n36548 = n36536 & ~n36547 ;
  assign n36549 = ( x208 & n36546 ) | ( x208 & ~n36548 ) | ( n36546 & ~n36548 ) ;
  assign n36550 = ~n36546 & n36549 ;
  assign n36551 = x208 | n36251 ;
  assign n36552 = n36530 | n36551 ;
  assign n36553 = ( x211 & ~n36550 ) | ( x211 & n36552 ) | ( ~n36550 & n36552 ) ;
  assign n36554 = ~x211 & n36553 ;
  assign n36555 = ( n36069 & n36544 ) | ( n36069 & ~n36554 ) | ( n36544 & ~n36554 ) ;
  assign n36556 = ~n36544 & n36555 ;
  assign n36557 = n9233 | n36529 ;
  assign n36558 = x1153 | n9353 ;
  assign n36559 = ~n36112 & n36558 ;
  assign n36560 = ( n36394 & n36395 ) | ( n36394 & n36559 ) | ( n36395 & n36559 ) ;
  assign n36561 = n36557 & n36560 ;
  assign n36562 = x214 | n36561 ;
  assign n36563 = ~x212 & n36562 ;
  assign n36564 = ( x212 & ~x219 ) | ( x212 & n36563 ) | ( ~x219 & n36563 ) ;
  assign n36565 = ( n36543 & ~n36556 ) | ( n36543 & n36564 ) | ( ~n36556 & n36564 ) ;
  assign n36566 = ~n36543 & n36565 ;
  assign n36567 = ~x211 & n36540 ;
  assign n36568 = n36035 & n36567 ;
  assign n36569 = ~n36036 & n36561 ;
  assign n36570 = n36568 | n36569 ;
  assign n36571 = n36566 ^ x219 ^ 1'b0 ;
  assign n36572 = ( ~x219 & n36570 ) | ( ~x219 & n36571 ) | ( n36570 & n36571 ) ;
  assign n36573 = ( x219 & n36566 ) | ( x219 & n36572 ) | ( n36566 & n36572 ) ;
  assign n36574 = x299 | x1153 ;
  assign n36575 = ~n9354 & n36574 ;
  assign n36576 = ~n36180 & n36575 ;
  assign n36577 = x207 & ~n36576 ;
  assign n36578 = x208 & ~n36577 ;
  assign n36579 = ( x299 & ~x1154 ) | ( x299 & n36513 ) | ( ~x1154 & n36513 ) ;
  assign n36580 = ~n36180 & n36579 ;
  assign n36581 = x1153 & ~n10008 ;
  assign n36582 = ( n36325 & n36532 ) | ( n36325 & n36581 ) | ( n36532 & n36581 ) ;
  assign n36583 = ~n36209 & n36582 ;
  assign n36584 = n36580 | n36583 ;
  assign n36585 = x207 | n36584 ;
  assign n36586 = n36578 & n36585 ;
  assign n36587 = x207 & ~n36584 ;
  assign n36588 = ~n36586 & n36587 ;
  assign n36589 = ( n36208 & n36586 ) | ( n36208 & ~n36588 ) | ( n36586 & ~n36588 ) ;
  assign n36590 = x211 & ~n36589 ;
  assign n36591 = x208 & n36000 ;
  assign n36592 = x1153 & ~n9354 ;
  assign n36593 = n36591 & n36592 ;
  assign n36594 = x200 & ~x1153 ;
  assign n36595 = n10019 | n36594 ;
  assign n36596 = ( n36513 & n36514 ) | ( n36513 & ~n36595 ) | ( n36514 & ~n36595 ) ;
  assign n36597 = n36395 & n36596 ;
  assign n36598 = n36593 | n36597 ;
  assign n36599 = x211 | n36251 ;
  assign n36600 = n36598 | n36599 ;
  assign n36601 = ( n36069 & n36590 ) | ( n36069 & n36600 ) | ( n36590 & n36600 ) ;
  assign n36602 = ~n36590 & n36601 ;
  assign n36603 = x211 | n36589 ;
  assign n36604 = ~n36150 & n36575 ;
  assign n36605 = x207 & ~n36604 ;
  assign n36606 = n36513 | n36582 ;
  assign n36607 = x207 | n36606 ;
  assign n36608 = ( x208 & n36605 ) | ( x208 & n36607 ) | ( n36605 & n36607 ) ;
  assign n36609 = ~n36605 & n36608 ;
  assign n36610 = x207 & n36606 ;
  assign n36611 = ( n36017 & n36606 ) | ( n36017 & n36610 ) | ( n36606 & n36610 ) ;
  assign n36612 = ( ~x208 & n36609 ) | ( ~x208 & n36611 ) | ( n36609 & n36611 ) ;
  assign n36613 = n36609 ^ x208 ^ 1'b0 ;
  assign n36614 = ( n36609 & n36612 ) | ( n36609 & ~n36613 ) | ( n36612 & ~n36613 ) ;
  assign n36615 = ( n9344 & n36307 ) | ( n9344 & n36614 ) | ( n36307 & n36614 ) ;
  assign n36616 = n36603 & n36615 ;
  assign n36617 = ( ~x219 & n36602 ) | ( ~x219 & n36616 ) | ( n36602 & n36616 ) ;
  assign n36618 = ~x219 & n36617 ;
  assign n36619 = ~n36035 & n36598 ;
  assign n36620 = x211 | n36614 ;
  assign n36621 = x219 & n36035 ;
  assign n36622 = x211 & ~n36598 ;
  assign n36623 = n36621 & ~n36622 ;
  assign n36624 = n36620 & n36623 ;
  assign n36625 = ( ~n36618 & n36619 ) | ( ~n36618 & n36624 ) | ( n36619 & n36624 ) ;
  assign n36626 = n36618 | n36625 ;
  assign n36627 = ( x1152 & ~n7318 ) | ( x1152 & n36626 ) | ( ~n7318 & n36626 ) ;
  assign n36628 = ~x1152 & n36627 ;
  assign n36629 = x1152 & ~n7318 ;
  assign n36630 = n36628 ^ n36573 ^ 1'b0 ;
  assign n36631 = ( ~n36573 & n36629 ) | ( ~n36573 & n36630 ) | ( n36629 & n36630 ) ;
  assign n36632 = ( n36573 & n36628 ) | ( n36573 & n36631 ) | ( n36628 & n36631 ) ;
  assign n36633 = ( x213 & ~n36501 ) | ( x213 & n36632 ) | ( ~n36501 & n36632 ) ;
  assign n36634 = ( x209 & n36501 ) | ( x209 & n36633 ) | ( n36501 & n36633 ) ;
  assign n36635 = x219 & ~n36561 ;
  assign n36636 = n36621 | n36635 ;
  assign n36637 = n36142 & n36518 ;
  assign n36638 = n36520 | n36637 ;
  assign n36639 = n36638 ^ x211 ^ 1'b0 ;
  assign n36640 = ( n36561 & n36638 ) | ( n36561 & n36639 ) | ( n36638 & n36639 ) ;
  assign n36641 = n36035 & n36640 ;
  assign n36642 = ( n7318 & n36636 ) | ( n7318 & ~n36641 ) | ( n36636 & ~n36641 ) ;
  assign n36643 = n36642 ^ n36636 ^ 1'b0 ;
  assign n36644 = ( n7318 & n36642 ) | ( n7318 & ~n36643 ) | ( n36642 & ~n36643 ) ;
  assign n36645 = x1153 | n9354 ;
  assign n36646 = ~x299 & n36087 ;
  assign n36647 = x207 & ~n36646 ;
  assign n36648 = n36645 & n36647 ;
  assign n36649 = ~x1153 & n36106 ;
  assign n36650 = n36166 & ~n36649 ;
  assign n36651 = n36325 & ~n36649 ;
  assign n36652 = n36650 | n36651 ;
  assign n36653 = ~x207 & n36652 ;
  assign n36654 = n36648 | n36653 ;
  assign n36655 = x207 | n36015 ;
  assign n36656 = ( n36015 & n36652 ) | ( n36015 & n36655 ) | ( n36652 & n36655 ) ;
  assign n36657 = n36656 ^ x208 ^ 1'b0 ;
  assign n36658 = ( n36654 & n36656 ) | ( n36654 & n36657 ) | ( n36656 & n36657 ) ;
  assign n36659 = ~x211 & n36658 ;
  assign n36660 = n36659 ^ n36658 ^ n36567 ;
  assign n36661 = x214 & ~n36660 ;
  assign n36662 = n36563 & ~n36661 ;
  assign n36664 = x211 & n36638 ;
  assign n36663 = x214 & ~n36659 ;
  assign n36665 = n36664 ^ n36663 ^ 1'b0 ;
  assign n36666 = ( x212 & ~n36663 ) | ( x212 & n36664 ) | ( ~n36663 & n36664 ) ;
  assign n36667 = ( x212 & ~n36665 ) | ( x212 & n36666 ) | ( ~n36665 & n36666 ) ;
  assign n36668 = n36667 ^ x219 ^ 1'b0 ;
  assign n36669 = x214 | n36660 ;
  assign n36670 = ( n36667 & ~n36668 ) | ( n36667 & n36669 ) | ( ~n36668 & n36669 ) ;
  assign n36671 = ( x219 & n36668 ) | ( x219 & n36670 ) | ( n36668 & n36670 ) ;
  assign n36672 = ( ~n36644 & n36662 ) | ( ~n36644 & n36671 ) | ( n36662 & n36671 ) ;
  assign n36673 = ~n36644 & n36672 ;
  assign n36674 = ( x1152 & n36456 ) | ( x1152 & ~n36673 ) | ( n36456 & ~n36673 ) ;
  assign n36675 = ~n36456 & n36674 ;
  assign n36676 = x1152 | n36494 ;
  assign n36677 = x207 & ~n9354 ;
  assign n36678 = x1153 & n36677 ;
  assign n36679 = x1153 & ~x1154 ;
  assign n36680 = n36181 & n36679 ;
  assign n36681 = n36651 | n36680 ;
  assign n36682 = ~x207 & n36681 ;
  assign n36683 = n36678 | n36682 ;
  assign n36684 = ( n36015 & n36655 ) | ( n36015 & n36681 ) | ( n36655 & n36681 ) ;
  assign n36685 = n36684 ^ x208 ^ 1'b0 ;
  assign n36686 = ( n36683 & n36684 ) | ( n36683 & n36685 ) | ( n36684 & n36685 ) ;
  assign n36687 = n36307 & ~n36686 ;
  assign n36688 = n36686 ^ x211 ^ 1'b0 ;
  assign n36689 = ( n36614 & n36686 ) | ( n36614 & ~n36688 ) | ( n36686 & ~n36688 ) ;
  assign n36690 = ( n9344 & n36035 ) | ( n9344 & ~n36689 ) | ( n36035 & ~n36689 ) ;
  assign n36691 = ~n9344 & n36690 ;
  assign n36692 = ( ~x219 & n36687 ) | ( ~x219 & n36691 ) | ( n36687 & n36691 ) ;
  assign n36693 = ~x219 & n36692 ;
  assign n36694 = x219 & ~n36598 ;
  assign n36695 = n7318 | n36694 ;
  assign n36696 = n35977 | n36369 ;
  assign n36697 = n36598 | n36696 ;
  assign n36698 = ( n36693 & ~n36695 ) | ( n36693 & n36697 ) | ( ~n36695 & n36697 ) ;
  assign n36699 = ~n36693 & n36698 ;
  assign n36700 = ( ~n36675 & n36676 ) | ( ~n36675 & n36699 ) | ( n36676 & n36699 ) ;
  assign n36701 = ~n36675 & n36700 ;
  assign n36702 = ( ~x213 & n36634 ) | ( ~x213 & n36701 ) | ( n36634 & n36701 ) ;
  assign n36703 = n36634 ^ x213 ^ 1'b0 ;
  assign n36704 = ( n36634 & n36702 ) | ( n36634 & ~n36703 ) | ( n36702 & ~n36703 ) ;
  assign n36705 = ( n36393 & ~n36500 ) | ( n36393 & n36704 ) | ( ~n36500 & n36704 ) ;
  assign n36706 = n36500 ^ n36393 ^ 1'b0 ;
  assign n36707 = ( n36393 & n36705 ) | ( n36393 & ~n36706 ) | ( n36705 & ~n36706 ) ;
  assign n36708 = x234 ^ x230 ^ 1'b0 ;
  assign n36709 = ( x234 & n36707 ) | ( x234 & n36708 ) | ( n36707 & n36708 ) ;
  assign n36710 = n36103 | n36182 ;
  assign n36711 = x207 & n36710 ;
  assign n36712 = ~x207 & n36212 ;
  assign n36713 = ( x208 & n36711 ) | ( x208 & n36712 ) | ( n36711 & n36712 ) ;
  assign n36714 = ( ~x1157 & n36213 ) | ( ~x1157 & n36713 ) | ( n36213 & n36713 ) ;
  assign n36715 = ~x1157 & n36714 ;
  assign n36716 = x208 & x1157 ;
  assign n36717 = x207 | n36230 ;
  assign n36718 = ~n36711 & n36717 ;
  assign n36719 = n36716 & ~n36718 ;
  assign n36720 = ( n36233 & ~n36715 ) | ( n36233 & n36719 ) | ( ~n36715 & n36719 ) ;
  assign n36721 = n36715 | n36720 ;
  assign n36722 = x211 | n36721 ;
  assign n36723 = ~x1156 & n36096 ;
  assign n36724 = n9233 & ~n36103 ;
  assign n36725 = ~n36723 & n36724 ;
  assign n36726 = ~x207 & n36132 ;
  assign n36727 = n36725 | n36726 ;
  assign n36728 = x208 | n36133 ;
  assign n36729 = x1157 & ~n36728 ;
  assign n36730 = ( x1157 & n36727 ) | ( x1157 & n36729 ) | ( n36727 & n36729 ) ;
  assign n36731 = x208 | n36092 ;
  assign n36732 = x207 | n36091 ;
  assign n36733 = ~n36725 & n36732 ;
  assign n36734 = n36731 & n36733 ;
  assign n36735 = ( x1157 & ~n36730 ) | ( x1157 & n36734 ) | ( ~n36730 & n36734 ) ;
  assign n36736 = ~n36730 & n36735 ;
  assign n36737 = x211 & ~n36736 ;
  assign n36738 = n36069 & ~n36737 ;
  assign n36739 = n36722 & n36738 ;
  assign n36740 = ~n36069 & n36736 ;
  assign n36741 = x219 & ~n36740 ;
  assign n36742 = ~n36739 & n36741 ;
  assign n36743 = ( ~n36085 & n36131 ) | ( ~n36085 & n36143 ) | ( n36131 & n36143 ) ;
  assign n36744 = x207 | n36743 ;
  assign n36745 = ( x207 & n36178 ) | ( x207 & n36723 ) | ( n36178 & n36723 ) ;
  assign n36746 = n36744 & ~n36745 ;
  assign n36747 = n36716 & ~n36746 ;
  assign n36748 = ~x207 & n36196 ;
  assign n36749 = ( x208 & n36745 ) | ( x208 & n36748 ) | ( n36745 & n36748 ) ;
  assign n36750 = ( ~x1157 & n36260 ) | ( ~x1157 & n36749 ) | ( n36260 & n36749 ) ;
  assign n36751 = ~x1157 & n36750 ;
  assign n36752 = ( n36253 & ~n36747 ) | ( n36253 & n36751 ) | ( ~n36747 & n36751 ) ;
  assign n36753 = n36747 | n36752 ;
  assign n36754 = ~x211 & n36753 ;
  assign n36755 = x211 & n36721 ;
  assign n36756 = ( n9344 & n36754 ) | ( n9344 & ~n36755 ) | ( n36754 & ~n36755 ) ;
  assign n36757 = ~n36754 & n36756 ;
  assign n36762 = ~x207 & n36147 ;
  assign n36763 = x208 & ~n36762 ;
  assign n36764 = ~n36178 & n36460 ;
  assign n36765 = n36763 & ~n36764 ;
  assign n36766 = n36149 | n36765 ;
  assign n36767 = x1157 & ~n36766 ;
  assign n36758 = n36731 ^ x1157 ^ 1'b0 ;
  assign n36759 = ( n36731 & n36733 ) | ( n36731 & ~n36758 ) | ( n36733 & ~n36758 ) ;
  assign n36760 = ( x1157 & n36758 ) | ( x1157 & n36759 ) | ( n36758 & n36759 ) ;
  assign n36761 = ~x211 & n36760 ;
  assign n36768 = n36767 ^ n36761 ^ 1'b0 ;
  assign n36769 = ( n36369 & ~n36761 ) | ( n36369 & n36767 ) | ( ~n36761 & n36767 ) ;
  assign n36770 = ( n36369 & ~n36768 ) | ( n36369 & n36769 ) | ( ~n36768 & n36769 ) ;
  assign n36771 = ( x211 & n36753 ) | ( x211 & ~n36770 ) | ( n36753 & ~n36770 ) ;
  assign n36772 = n36771 ^ n36770 ^ 1'b0 ;
  assign n36773 = ( n36770 & ~n36771 ) | ( n36770 & n36772 ) | ( ~n36771 & n36772 ) ;
  assign n36774 = ( n36035 & n36736 ) | ( n36035 & ~n36773 ) | ( n36736 & ~n36773 ) ;
  assign n36775 = ~n36773 & n36774 ;
  assign n36776 = n36775 ^ n36757 ^ 1'b0 ;
  assign n36777 = ( n36757 & n36775 ) | ( n36757 & n36776 ) | ( n36775 & n36776 ) ;
  assign n36778 = ( x219 & ~n36757 ) | ( x219 & n36777 ) | ( ~n36757 & n36777 ) ;
  assign n36779 = ( x209 & n36742 ) | ( x209 & n36778 ) | ( n36742 & n36778 ) ;
  assign n36780 = ~n36742 & n36779 ;
  assign n36781 = n9233 & ~n36596 ;
  assign n36782 = ( x207 & x208 ) | ( x207 & n36121 ) | ( x208 & n36121 ) ;
  assign n36783 = ~n36781 & n36782 ;
  assign n36784 = x211 & ~n36783 ;
  assign n36785 = n36069 & ~n36784 ;
  assign n36786 = n36208 & n36222 ;
  assign n36787 = x207 | n36222 ;
  assign n36788 = x208 & ~n36587 ;
  assign n36789 = n36787 & n36788 ;
  assign n36790 = n36786 | n36789 ;
  assign n36791 = x211 | n36790 ;
  assign n36792 = n36785 & n36791 ;
  assign n36793 = ~n36069 & n36783 ;
  assign n36794 = x219 & ~n36793 ;
  assign n36795 = ~n36792 & n36794 ;
  assign n36796 = n36251 | n36783 ;
  assign n36797 = ~x211 & n36796 ;
  assign n36798 = x211 & n36790 ;
  assign n36799 = ( n9344 & n36797 ) | ( n9344 & ~n36798 ) | ( n36797 & ~n36798 ) ;
  assign n36800 = ~n36797 & n36799 ;
  assign n36801 = ( n36035 & n36783 ) | ( n36035 & ~n36800 ) | ( n36783 & ~n36800 ) ;
  assign n36802 = ~n36800 & n36801 ;
  assign n36803 = x211 & ~n36796 ;
  assign n36804 = ~x1157 & n36783 ;
  assign n36805 = x1157 ^ x211 ^ 1'b0 ;
  assign n36806 = n36579 | n36582 ;
  assign n36807 = x207 & ~n36806 ;
  assign n36808 = n36141 | n36188 ;
  assign n36809 = x208 & n36808 ;
  assign n36810 = ~n36807 & n36809 ;
  assign n36811 = n36142 & ~n36244 ;
  assign n36812 = n36810 | n36811 ;
  assign n36813 = ( x1157 & ~n36805 ) | ( x1157 & n36812 ) | ( ~n36805 & n36812 ) ;
  assign n36814 = ( x211 & n36805 ) | ( x211 & n36813 ) | ( n36805 & n36813 ) ;
  assign n36815 = ( ~n36803 & n36804 ) | ( ~n36803 & n36814 ) | ( n36804 & n36814 ) ;
  assign n36816 = ~n36803 & n36815 ;
  assign n36817 = ( n9344 & n36035 ) | ( n9344 & ~n36816 ) | ( n36035 & ~n36816 ) ;
  assign n36818 = ~n9344 & n36817 ;
  assign n36819 = ( x219 & n36802 ) | ( x219 & ~n36818 ) | ( n36802 & ~n36818 ) ;
  assign n36820 = n36819 ^ n36802 ^ 1'b0 ;
  assign n36821 = ( x219 & n36819 ) | ( x219 & ~n36820 ) | ( n36819 & ~n36820 ) ;
  assign n36822 = ( x209 & ~n36795 ) | ( x209 & n36821 ) | ( ~n36795 & n36821 ) ;
  assign n36823 = ~x209 & n36822 ;
  assign n36824 = ( ~n7318 & n36780 ) | ( ~n7318 & n36823 ) | ( n36780 & n36823 ) ;
  assign n36825 = ~n7318 & n36824 ;
  assign n36830 = x219 & ~n36369 ;
  assign n36831 = x219 & ~n35963 ;
  assign n36832 = ( x219 & n36830 ) | ( x219 & n36831 ) | ( n36830 & n36831 ) ;
  assign n36826 = ( n35962 & ~n35966 ) | ( n35962 & n35971 ) | ( ~n35966 & n35971 ) ;
  assign n36827 = ( x212 & ~n36268 ) | ( x212 & n36826 ) | ( ~n36268 & n36826 ) ;
  assign n36828 = ( x219 & n36268 ) | ( x219 & n36827 ) | ( n36268 & n36827 ) ;
  assign n36829 = n35973 | n36828 ;
  assign n36833 = ( n7318 & n36829 ) | ( n7318 & n36832 ) | ( n36829 & n36832 ) ;
  assign n36834 = ~n36832 & n36833 ;
  assign n36835 = ( x213 & n36825 ) | ( x213 & ~n36834 ) | ( n36825 & ~n36834 ) ;
  assign n36836 = ~n36825 & n36835 ;
  assign n36837 = n36163 | n36407 ;
  assign n36838 = n36837 ^ x208 ^ 1'b0 ;
  assign n36839 = n36162 ^ x207 ^ 1'b0 ;
  assign n36840 = ( n36162 & n36606 ) | ( n36162 & n36839 ) | ( n36606 & n36839 ) ;
  assign n36841 = ( n36837 & n36838 ) | ( n36837 & n36840 ) | ( n36838 & n36840 ) ;
  assign n36842 = ~x211 & n36841 ;
  assign n36843 = n36188 ^ x207 ^ 1'b0 ;
  assign n36844 = ( n36015 & n36188 ) | ( n36015 & ~n36843 ) | ( n36188 & ~n36843 ) ;
  assign n36845 = n36844 ^ x208 ^ 1'b0 ;
  assign n36846 = ( n36188 & n36681 ) | ( n36188 & n36843 ) | ( n36681 & n36843 ) ;
  assign n36847 = ( n36844 & n36845 ) | ( n36844 & n36846 ) | ( n36845 & n36846 ) ;
  assign n36848 = x211 & n36847 ;
  assign n36849 = ( n9344 & n36842 ) | ( n9344 & ~n36848 ) | ( n36842 & ~n36848 ) ;
  assign n36850 = ~n36842 & n36849 ;
  assign n36851 = ( n36035 & n36783 ) | ( n36035 & ~n36850 ) | ( n36783 & ~n36850 ) ;
  assign n36852 = ~n36850 & n36851 ;
  assign n36853 = x211 & ~n36841 ;
  assign n36854 = n36069 & ~n36791 ;
  assign n36855 = ( n36069 & n36853 ) | ( n36069 & n36854 ) | ( n36853 & n36854 ) ;
  assign n36856 = ( x219 & n36852 ) | ( x219 & ~n36855 ) | ( n36852 & ~n36855 ) ;
  assign n36857 = n36856 ^ n36852 ^ 1'b0 ;
  assign n36858 = ( x219 & n36856 ) | ( x219 & ~n36857 ) | ( n36856 & ~n36857 ) ;
  assign n36859 = x211 | n36847 ;
  assign n36860 = n36785 & n36859 ;
  assign n36861 = n36794 & ~n36860 ;
  assign n36862 = ( x209 & n36858 ) | ( x209 & ~n36861 ) | ( n36858 & ~n36861 ) ;
  assign n36863 = n36862 ^ n36858 ^ 1'b0 ;
  assign n36864 = ( x209 & n36862 ) | ( x209 & ~n36863 ) | ( n36862 & ~n36863 ) ;
  assign n36865 = x1157 & n36766 ;
  assign n36866 = ( x299 & ~x1157 ) | ( x299 & n36751 ) | ( ~x1157 & n36751 ) ;
  assign n36867 = ( ~n36185 & n36865 ) | ( ~n36185 & n36866 ) | ( n36865 & n36866 ) ;
  assign n36868 = ~n36185 & n36867 ;
  assign n36869 = x211 | n36868 ;
  assign n36870 = n36738 & n36869 ;
  assign n36871 = n36741 & ~n36870 ;
  assign n36872 = x211 & n36868 ;
  assign n36873 = n36097 & n36183 ;
  assign n36874 = n36103 | n36873 ;
  assign n36875 = x207 & n36874 ;
  assign n36876 = x1154 & ~n36195 ;
  assign n36877 = n36090 | n36876 ;
  assign n36878 = ( x207 & n36211 ) | ( x207 & n36877 ) | ( n36211 & n36877 ) ;
  assign n36879 = ~x207 & n36878 ;
  assign n36880 = ( x208 & n36875 ) | ( x208 & ~n36879 ) | ( n36875 & ~n36879 ) ;
  assign n36881 = ~n36875 & n36880 ;
  assign n36882 = x208 | n36153 ;
  assign n36883 = ( x1157 & ~n36881 ) | ( x1157 & n36882 ) | ( ~n36881 & n36882 ) ;
  assign n36884 = ~x1157 & n36883 ;
  assign n36885 = n36884 ^ n36151 ^ 1'b0 ;
  assign n36886 = ( ~n36151 & n36766 ) | ( ~n36151 & n36885 ) | ( n36766 & n36885 ) ;
  assign n36887 = ( n36151 & n36884 ) | ( n36151 & n36886 ) | ( n36884 & n36886 ) ;
  assign n36888 = ~x211 & n36887 ;
  assign n36889 = ( n9344 & n36872 ) | ( n9344 & ~n36888 ) | ( n36872 & ~n36888 ) ;
  assign n36890 = ~n36872 & n36889 ;
  assign n36891 = x211 & ~n36887 ;
  assign n36892 = n36369 & ~n36722 ;
  assign n36893 = ( n36369 & n36891 ) | ( n36369 & n36892 ) | ( n36891 & n36892 ) ;
  assign n36894 = ( n36035 & n36736 ) | ( n36035 & ~n36893 ) | ( n36736 & ~n36893 ) ;
  assign n36895 = ~n36893 & n36894 ;
  assign n36896 = n36895 ^ n36890 ^ 1'b0 ;
  assign n36897 = ( n36890 & n36895 ) | ( n36890 & n36896 ) | ( n36895 & n36896 ) ;
  assign n36898 = ( x219 & ~n36890 ) | ( x219 & n36897 ) | ( ~n36890 & n36897 ) ;
  assign n36899 = x209 & ~n36898 ;
  assign n36900 = ( x209 & n36871 ) | ( x209 & n36899 ) | ( n36871 & n36899 ) ;
  assign n36901 = ( n7318 & n36864 ) | ( n7318 & ~n36900 ) | ( n36864 & ~n36900 ) ;
  assign n36902 = ~n7318 & n36901 ;
  assign n36903 = n9344 & n36452 ;
  assign n36904 = n35965 & n36369 ;
  assign n36905 = ( x219 & ~n36903 ) | ( x219 & n36904 ) | ( ~n36903 & n36904 ) ;
  assign n36906 = n36903 | n36905 ;
  assign n36907 = n36906 ^ x213 ^ 1'b0 ;
  assign n36908 = x219 & ~n35980 ;
  assign n36909 = n7318 & ~n36908 ;
  assign n36910 = ~n36830 & n36909 ;
  assign n36911 = ( n36906 & ~n36907 ) | ( n36906 & n36910 ) | ( ~n36907 & n36910 ) ;
  assign n36912 = ( x213 & n36907 ) | ( x213 & n36911 ) | ( n36907 & n36911 ) ;
  assign n36913 = ( ~n36836 & n36902 ) | ( ~n36836 & n36912 ) | ( n36902 & n36912 ) ;
  assign n36914 = ~n36836 & n36913 ;
  assign n36915 = x235 ^ x230 ^ 1'b0 ;
  assign n36916 = ( x235 & n36914 ) | ( x235 & n36915 ) | ( n36914 & n36915 ) ;
  assign n36917 = ~x100 & n35722 ;
  assign n36918 = n35943 | n36917 ;
  assign n36919 = ( x75 & ~n5013 ) | ( x75 & n36918 ) | ( ~n5013 & n36918 ) ;
  assign n36920 = ~x75 & n36919 ;
  assign n36921 = x75 & ~n6255 ;
  assign n36922 = ( x92 & ~n36920 ) | ( x92 & n36921 ) | ( ~n36920 & n36921 ) ;
  assign n36923 = n36920 | n36922 ;
  assign n36924 = n36923 ^ n12146 ^ 1'b0 ;
  assign n36925 = ( n12146 & n36923 ) | ( n12146 & n36924 ) | ( n36923 & n36924 ) ;
  assign n36926 = ( x74 & ~n12146 ) | ( x74 & n36925 ) | ( ~n12146 & n36925 ) ;
  assign n36927 = n36926 ^ n5012 ^ 1'b0 ;
  assign n36928 = ( n5012 & n36926 ) | ( n5012 & n36927 ) | ( n36926 & n36927 ) ;
  assign n36929 = ( x56 & ~n5012 ) | ( x56 & n36928 ) | ( ~n5012 & n36928 ) ;
  assign n36930 = n36929 ^ n5008 ^ 1'b0 ;
  assign n36931 = ( n5008 & n36929 ) | ( n5008 & n36930 ) | ( n36929 & n36930 ) ;
  assign n36932 = ( x62 & ~n5008 ) | ( x62 & n36931 ) | ( ~n5008 & n36931 ) ;
  assign n36933 = ( x57 & ~n5006 ) | ( x57 & n36932 ) | ( ~n5006 & n36932 ) ;
  assign n36934 = ~x57 & n36933 ;
  assign n36935 = ( x1157 & x1158 ) | ( x1157 & ~n36805 ) | ( x1158 & ~n36805 ) ;
  assign n36936 = n36014 & n36935 ;
  assign n36937 = n36828 | n36936 ;
  assign n36938 = n36937 ^ x213 ^ 1'b0 ;
  assign n36939 = x1155 & ~n36140 ;
  assign n36940 = x214 & n35982 ;
  assign n36941 = n36939 | n36940 ;
  assign n36942 = ( ~x212 & n7318 ) | ( ~x212 & n36941 ) | ( n7318 & n36941 ) ;
  assign n36943 = x212 & n36942 ;
  assign n36944 = n35960 & n36014 ;
  assign n36945 = x219 & ~n36944 ;
  assign n36946 = ~n36943 & n36945 ;
  assign n36947 = ( n7318 & n36943 ) | ( n7318 & ~n36946 ) | ( n36943 & ~n36946 ) ;
  assign n36948 = ( n36937 & ~n36938 ) | ( n36937 & n36947 ) | ( ~n36938 & n36947 ) ;
  assign n36949 = ( x213 & n36938 ) | ( x213 & n36948 ) | ( n36938 & n36948 ) ;
  assign n36950 = x207 & n36430 ;
  assign n36951 = n36717 & ~n36950 ;
  assign n36952 = n36716 & ~n36951 ;
  assign n36953 = ( x208 & n36712 ) | ( x208 & n36950 ) | ( n36712 & n36950 ) ;
  assign n36954 = n36009 & ~n36106 ;
  assign n36955 = x1158 & ~n36216 ;
  assign n36956 = x199 | x1158 ;
  assign n36957 = x1156 & n36956 ;
  assign n36958 = n36955 | n36957 ;
  assign n36959 = n36954 & n36958 ;
  assign n36960 = ( n36021 & n36208 ) | ( n36021 & n36959 ) | ( n36208 & n36959 ) ;
  assign n36961 = ( ~x1157 & n36953 ) | ( ~x1157 & n36960 ) | ( n36953 & n36960 ) ;
  assign n36962 = ~x1157 & n36961 ;
  assign n36963 = x200 | x1158 ;
  assign n36964 = ~x199 & n36963 ;
  assign n36965 = x1156 & ~n36646 ;
  assign n36966 = x1158 | n36089 ;
  assign n36967 = n36965 & n36966 ;
  assign n36968 = n36964 | n36967 ;
  assign n36969 = n36000 & n36968 ;
  assign n36970 = n36021 | n36969 ;
  assign n36971 = n36250 & n36970 ;
  assign n36972 = ( ~n36952 & n36962 ) | ( ~n36952 & n36971 ) | ( n36962 & n36971 ) ;
  assign n36973 = n36952 | n36972 ;
  assign n36974 = n9271 & n36973 ;
  assign n36975 = ~n36421 & n36744 ;
  assign n36976 = n36716 & ~n36975 ;
  assign n36977 = ~x200 & x207 ;
  assign n36978 = n36958 & n36977 ;
  assign n36979 = n36551 | n36978 ;
  assign n36980 = x208 & ~n36748 ;
  assign n36981 = ~n36421 & n36980 ;
  assign n36982 = ( x1157 & n36979 ) | ( x1157 & ~n36981 ) | ( n36979 & ~n36981 ) ;
  assign n36983 = ~x1157 & n36982 ;
  assign n36984 = x1156 & n36164 ;
  assign n36985 = n36964 | n36984 ;
  assign n36986 = n36000 & n36985 ;
  assign n36987 = ( n36250 & n36251 ) | ( n36250 & n36986 ) | ( n36251 & n36986 ) ;
  assign n36988 = ( ~n36976 & n36983 ) | ( ~n36976 & n36987 ) | ( n36983 & n36987 ) ;
  assign n36989 = n36976 | n36988 ;
  assign n36990 = n36271 & n36989 ;
  assign n36991 = n36974 | n36990 ;
  assign n36992 = x208 & n36732 ;
  assign n36993 = ~n36105 & n36992 ;
  assign n36994 = n36959 | n36993 ;
  assign n36995 = n36994 ^ x1157 ^ 1'b0 ;
  assign n36996 = x299 | n36985 ;
  assign n36997 = n36142 & n36996 ;
  assign n36998 = ~n36461 & n36763 ;
  assign n36999 = n36997 | n36998 ;
  assign n37000 = ( n36994 & n36995 ) | ( n36994 & n36999 ) | ( n36995 & n36999 ) ;
  assign n37001 = ~n36140 & n37000 ;
  assign n37002 = ( x212 & n36991 ) | ( x212 & n37001 ) | ( n36991 & n37001 ) ;
  assign n37003 = n37001 ^ n36991 ^ 1'b0 ;
  assign n37004 = ( x212 & n37002 ) | ( x212 & n37003 ) | ( n37002 & n37003 ) ;
  assign n37005 = ~x208 & n36986 ;
  assign n37006 = x208 & ~n36726 ;
  assign n37007 = ~n36105 & n37006 ;
  assign n37008 = n37005 | n37007 ;
  assign n37009 = ( n36994 & n36995 ) | ( n36994 & n37008 ) | ( n36995 & n37008 ) ;
  assign n37010 = x214 | n37009 ;
  assign n37011 = x211 & ~n37000 ;
  assign n37012 = n36089 & n36228 ;
  assign n37013 = x1157 & ~n36955 ;
  assign n37014 = ~n37012 & n37013 ;
  assign n37015 = x207 & ~n37014 ;
  assign n37016 = x299 & x1158 ;
  assign n37017 = ( x1158 & n36677 ) | ( x1158 & n37016 ) | ( n36677 & n37016 ) ;
  assign n37018 = n37015 | n37017 ;
  assign n37019 = n36250 & n37018 ;
  assign n37020 = n36000 & n36984 ;
  assign n37021 = x208 | n37020 ;
  assign n37022 = n37017 | n37021 ;
  assign n37023 = x1158 | n36104 ;
  assign n37024 = x1158 & ~n36184 ;
  assign n37025 = x207 & ~n37024 ;
  assign n37026 = n37023 & n37025 ;
  assign n37027 = x299 | n36196 ;
  assign n37028 = x299 & ~x1158 ;
  assign n37029 = x207 | n37028 ;
  assign n37030 = n37027 & ~n37029 ;
  assign n37031 = ( x208 & n37026 ) | ( x208 & ~n37030 ) | ( n37026 & ~n37030 ) ;
  assign n37032 = ~n37026 & n37031 ;
  assign n37033 = ( x1157 & n37022 ) | ( x1157 & ~n37032 ) | ( n37022 & ~n37032 ) ;
  assign n37034 = ~x1157 & n37033 ;
  assign n37035 = ( x211 & ~n37019 ) | ( x211 & n37034 ) | ( ~n37019 & n37034 ) ;
  assign n37036 = n37019 | n37035 ;
  assign n37037 = ( n36762 & ~n37026 ) | ( n36762 & n37029 ) | ( ~n37026 & n37029 ) ;
  assign n37038 = ~n37036 & n37037 ;
  assign n37039 = ( n36716 & n37036 ) | ( n36716 & ~n37038 ) | ( n37036 & ~n37038 ) ;
  assign n37040 = x214 & ~n37039 ;
  assign n37041 = ( x214 & n37011 ) | ( x214 & n37040 ) | ( n37011 & n37040 ) ;
  assign n37042 = ( x212 & n37010 ) | ( x212 & ~n37041 ) | ( n37010 & ~n37041 ) ;
  assign n37043 = ~x212 & n37042 ;
  assign n37044 = ( x219 & ~n37004 ) | ( x219 & n37043 ) | ( ~n37004 & n37043 ) ;
  assign n37045 = n37004 | n37044 ;
  assign n37046 = ~x214 & n36973 ;
  assign n37047 = x207 | n36147 ;
  assign n37048 = n36150 | n37047 ;
  assign n37049 = x1157 & n37048 ;
  assign n37050 = x1157 | n36959 ;
  assign n37051 = n36879 | n37050 ;
  assign n37052 = ~n37049 & n37051 ;
  assign n37053 = ( x208 & n36406 ) | ( x208 & ~n37052 ) | ( n36406 & ~n37052 ) ;
  assign n37054 = ~n36406 & n37053 ;
  assign n37055 = n36969 & n37050 ;
  assign n37056 = x208 | n36017 ;
  assign n37057 = n37055 | n37056 ;
  assign n37058 = ( x214 & n37054 ) | ( x214 & n37057 ) | ( n37054 & n37057 ) ;
  assign n37059 = ~n37054 & n37058 ;
  assign n37060 = ( x212 & n37046 ) | ( x212 & ~n37059 ) | ( n37046 & ~n37059 ) ;
  assign n37061 = ~n37046 & n37060 ;
  assign n37062 = n36014 & ~n36989 ;
  assign n37063 = ( ~x211 & n37061 ) | ( ~x211 & n37062 ) | ( n37061 & n37062 ) ;
  assign n37064 = ~x211 & n37063 ;
  assign n37065 = n36036 | n37009 ;
  assign n37066 = x219 & ~n37065 ;
  assign n37067 = ( x219 & n37064 ) | ( x219 & n37066 ) | ( n37064 & n37066 ) ;
  assign n37068 = ( x57 & n5193 ) | ( x57 & ~n37067 ) | ( n5193 & ~n37067 ) ;
  assign n37069 = n37067 | n37068 ;
  assign n37070 = ( n36949 & n37045 ) | ( n36949 & ~n37069 ) | ( n37045 & ~n37069 ) ;
  assign n37071 = n37070 ^ n37045 ^ 1'b0 ;
  assign n37072 = ( n36949 & n37070 ) | ( n36949 & ~n37071 ) | ( n37070 & ~n37071 ) ;
  assign n37073 = x219 & ~n36046 ;
  assign n37074 = n36038 & ~n37073 ;
  assign n37075 = ~x211 & x1145 ;
  assign n37076 = x211 & x1144 ;
  assign n37077 = n37075 | n37076 ;
  assign n37078 = n9344 | n37077 ;
  assign n37079 = ( n36035 & n36055 ) | ( n36035 & n36369 ) | ( n36055 & n36369 ) ;
  assign n37080 = n37078 & n37079 ;
  assign n37081 = x219 | n37080 ;
  assign n37082 = n37074 & n37081 ;
  assign n37083 = x207 & n36333 ;
  assign n37084 = ~x200 & x1157 ;
  assign n37085 = ~x199 & n37084 ;
  assign n37086 = n37027 | n37085 ;
  assign n37087 = x207 | n36309 ;
  assign n37088 = n37086 & ~n37087 ;
  assign n37089 = ( x208 & n37083 ) | ( x208 & ~n37088 ) | ( n37083 & ~n37088 ) ;
  assign n37090 = ~n37083 & n37089 ;
  assign n37091 = x1157 | n36978 ;
  assign n37092 = ( x208 & n36969 ) | ( x208 & n37091 ) | ( n36969 & n37091 ) ;
  assign n37093 = ~x208 & n37092 ;
  assign n37094 = x208 | n37093 ;
  assign n37095 = ( n36048 & ~n37090 ) | ( n36048 & n37094 ) | ( ~n37090 & n37094 ) ;
  assign n37096 = ~n37090 & n37095 ;
  assign n37097 = n36036 & ~n37096 ;
  assign n37098 = ( x219 & n37066 ) | ( x219 & n37097 ) | ( n37066 & n37097 ) ;
  assign n37099 = ~x212 & n37010 ;
  assign n37102 = x299 & ~x1145 ;
  assign n37103 = ( ~x1154 & n36177 ) | ( ~x1154 & n37102 ) | ( n36177 & n37102 ) ;
  assign n37100 = x299 & x1145 ;
  assign n37101 = n36318 & ~n37100 ;
  assign n37104 = ( x1156 & ~n37101 ) | ( x1156 & n37103 ) | ( ~n37101 & n37103 ) ;
  assign n37105 = ~n37103 & n37104 ;
  assign n37106 = n36168 & ~n37102 ;
  assign n37107 = x1154 & ~n37106 ;
  assign n37108 = n36097 | n37100 ;
  assign n37109 = ( x1156 & ~n37107 ) | ( x1156 & n37108 ) | ( ~n37107 & n37108 ) ;
  assign n37110 = ~x1156 & n37109 ;
  assign n37111 = ( x207 & n37105 ) | ( x207 & n37110 ) | ( n37105 & n37110 ) ;
  assign n37112 = n37110 ^ n37105 ^ 1'b0 ;
  assign n37113 = ( x207 & n37111 ) | ( x207 & n37112 ) | ( n37111 & n37112 ) ;
  assign n37114 = x207 | n37102 ;
  assign n37115 = n37086 & ~n37114 ;
  assign n37116 = ( x208 & n37113 ) | ( x208 & ~n37115 ) | ( n37113 & ~n37115 ) ;
  assign n37117 = ~n37113 & n37116 ;
  assign n37118 = x208 | n37100 ;
  assign n37119 = x1157 | n36955 ;
  assign n37120 = ~x299 & n36984 ;
  assign n37121 = n37119 | n37120 ;
  assign n37122 = n37015 & n37121 ;
  assign n37123 = ( ~n37117 & n37118 ) | ( ~n37117 & n37122 ) | ( n37118 & n37122 ) ;
  assign n37124 = ~n37117 & n37123 ;
  assign n37125 = x207 & n36356 ;
  assign n37126 = x207 | n36344 ;
  assign n37127 = n37086 & ~n37126 ;
  assign n37128 = ( x208 & n37125 ) | ( x208 & ~n37127 ) | ( n37125 & ~n37127 ) ;
  assign n37129 = ~n37125 & n37128 ;
  assign n37130 = ( n36341 & n37094 ) | ( n36341 & ~n37129 ) | ( n37094 & ~n37129 ) ;
  assign n37131 = ~n37129 & n37130 ;
  assign n37132 = n37124 ^ x211 ^ 1'b0 ;
  assign n37133 = ( n37124 & n37131 ) | ( n37124 & n37132 ) | ( n37131 & n37132 ) ;
  assign n37134 = x214 & ~n37133 ;
  assign n37135 = n37099 & ~n37134 ;
  assign n37138 = x211 & n37096 ;
  assign n37136 = ~x211 & n37131 ;
  assign n37137 = x214 & ~n37136 ;
  assign n37139 = n37138 ^ n37137 ^ 1'b0 ;
  assign n37140 = ( x212 & ~n37137 ) | ( x212 & n37138 ) | ( ~n37137 & n37138 ) ;
  assign n37141 = ( x212 & ~n37139 ) | ( x212 & n37140 ) | ( ~n37139 & n37140 ) ;
  assign n37142 = n37133 ^ x214 ^ 1'b0 ;
  assign n37143 = ( x214 & n37133 ) | ( x214 & ~n37142 ) | ( n37133 & ~n37142 ) ;
  assign n37144 = ( n37141 & n37142 ) | ( n37141 & n37143 ) | ( n37142 & n37143 ) ;
  assign n37145 = ( x219 & ~n37135 ) | ( x219 & n37144 ) | ( ~n37135 & n37144 ) ;
  assign n37146 = n37135 | n37145 ;
  assign n37147 = ( n7318 & ~n37098 ) | ( n7318 & n37146 ) | ( ~n37098 & n37146 ) ;
  assign n37148 = ~n7318 & n37147 ;
  assign n37149 = ( x213 & n37082 ) | ( x213 & ~n37148 ) | ( n37082 & ~n37148 ) ;
  assign n37150 = ~n37082 & n37149 ;
  assign n37151 = ( x209 & n37072 ) | ( x209 & ~n37150 ) | ( n37072 & ~n37150 ) ;
  assign n37152 = ~x209 & n37151 ;
  assign n37153 = x214 & ~n36017 ;
  assign n37154 = x214 | n36021 ;
  assign n37155 = ( x212 & n37153 ) | ( x212 & n37154 ) | ( n37153 & n37154 ) ;
  assign n37156 = ~n37153 & n37155 ;
  assign n37157 = ( x299 & n36251 ) | ( x299 & n37156 ) | ( n36251 & n37156 ) ;
  assign n37158 = ( n36014 & n37156 ) | ( n36014 & n37157 ) | ( n37156 & n37157 ) ;
  assign n37159 = ( x211 & x219 ) | ( x211 & n37158 ) | ( x219 & n37158 ) ;
  assign n37160 = ~x211 & n37159 ;
  assign n37161 = x199 & x1143 ;
  assign n37162 = x200 | n37161 ;
  assign n37163 = ~x199 & x1145 ;
  assign n37164 = n37162 | n37163 ;
  assign n37165 = x200 & ~n35993 ;
  assign n37166 = n36395 & ~n37165 ;
  assign n37167 = n37164 & n37166 ;
  assign n37168 = n35993 | n37162 ;
  assign n37169 = ~n35996 & n36591 ;
  assign n37170 = n37168 & n37169 ;
  assign n37171 = ( ~x299 & n37167 ) | ( ~x299 & n37170 ) | ( n37167 & n37170 ) ;
  assign n37172 = ~x299 & n37171 ;
  assign n37173 = n36026 & n36937 ;
  assign n37174 = ( ~n37160 & n37172 ) | ( ~n37160 & n37173 ) | ( n37172 & n37173 ) ;
  assign n37175 = n37160 | n37174 ;
  assign n37176 = n7318 | n37175 ;
  assign n37177 = ( ~n7318 & n36949 ) | ( ~n7318 & n37176 ) | ( n36949 & n37176 ) ;
  assign n37178 = n36026 & n37080 ;
  assign n37179 = x299 & n36621 ;
  assign n37180 = n36046 & n37179 ;
  assign n37181 = ( n37172 & ~n37178 ) | ( n37172 & n37180 ) | ( ~n37178 & n37180 ) ;
  assign n37182 = n37178 | n37181 ;
  assign n37183 = n7318 | n37182 ;
  assign n37184 = ( ~n7318 & n37082 ) | ( ~n7318 & n37183 ) | ( n37082 & n37183 ) ;
  assign n37185 = x213 & ~n37184 ;
  assign n37186 = x209 & ~n37185 ;
  assign n37187 = n37177 & n37186 ;
  assign n37188 = ( x230 & n37152 ) | ( x230 & n37187 ) | ( n37152 & n37187 ) ;
  assign n37189 = n37187 ^ n37152 ^ 1'b0 ;
  assign n37190 = ( x230 & n37188 ) | ( x230 & n37189 ) | ( n37188 & n37189 ) ;
  assign n37191 = ( x230 & x237 ) | ( x230 & ~n37190 ) | ( x237 & ~n37190 ) ;
  assign n37192 = ~n37190 & n37191 ;
  assign n37193 = n36089 & n36679 ;
  assign n37194 = n9233 & ~n37193 ;
  assign n37195 = ~n36526 & n37194 ;
  assign n37196 = n36782 & ~n37195 ;
  assign n37197 = ~x219 & n36369 ;
  assign n37198 = n37196 | n37197 ;
  assign n37199 = x211 & ~n37196 ;
  assign n37200 = x1153 & n36166 ;
  assign n37201 = n36526 | n37200 ;
  assign n37202 = ( n36188 & n36843 ) | ( n36188 & n37201 ) | ( n36843 & n37201 ) ;
  assign n37203 = ( n36844 & n36845 ) | ( n36844 & n37202 ) | ( n36845 & n37202 ) ;
  assign n37204 = x211 | n37203 ;
  assign n37205 = ~n37199 & n37204 ;
  assign n37206 = n37197 & ~n37205 ;
  assign n37207 = ( n7318 & n37198 ) | ( n7318 & ~n37206 ) | ( n37198 & ~n37206 ) ;
  assign n37208 = ~n7318 & n37207 ;
  assign n37209 = ~x211 & n36369 ;
  assign n37210 = x1153 & n37209 ;
  assign n37211 = ~x219 & n7318 ;
  assign n37212 = n37210 & n37211 ;
  assign n37213 = ( x1151 & ~n37208 ) | ( x1151 & n37212 ) | ( ~n37208 & n37212 ) ;
  assign n37214 = n37208 | n37213 ;
  assign n37215 = n9275 | n37210 ;
  assign n37216 = n36038 & n37215 ;
  assign n37217 = ~x1154 & n36574 ;
  assign n37218 = x207 & ~n37217 ;
  assign n37219 = ( x207 & ~n36166 ) | ( x207 & n37218 ) | ( ~n36166 & n37218 ) ;
  assign n37220 = n37219 ^ n36533 ^ 1'b0 ;
  assign n37221 = ( x208 & n36533 ) | ( x208 & ~n37219 ) | ( n36533 & ~n37219 ) ;
  assign n37222 = ( x208 & ~n37220 ) | ( x208 & n37221 ) | ( ~n37220 & n37221 ) ;
  assign n37223 = ( n36808 & n36811 ) | ( n36808 & n37222 ) | ( n36811 & n37222 ) ;
  assign n37224 = x211 & ~n37223 ;
  assign n37225 = n37224 ^ n37223 ^ n37199 ;
  assign n37226 = n36035 & ~n37225 ;
  assign n37227 = x214 | n37196 ;
  assign n37228 = x212 | n37227 ;
  assign n37229 = x219 & ~n37228 ;
  assign n37230 = ( x219 & n37226 ) | ( x219 & n37229 ) | ( n37226 & n37229 ) ;
  assign n37231 = n37225 ^ n37223 ^ n37196 ;
  assign n37232 = x214 & n37231 ;
  assign n37233 = ~x214 & n37205 ;
  assign n37234 = ( x212 & n37232 ) | ( x212 & ~n37233 ) | ( n37232 & ~n37233 ) ;
  assign n37235 = ~n37232 & n37234 ;
  assign n37236 = x214 & ~n37205 ;
  assign n37237 = n37227 & ~n37236 ;
  assign n37238 = x212 | n37237 ;
  assign n37239 = n37238 ^ n37235 ^ 1'b0 ;
  assign n37240 = ( n37235 & n37238 ) | ( n37235 & n37239 ) | ( n37238 & n37239 ) ;
  assign n37241 = ( x219 & ~n37235 ) | ( x219 & n37240 ) | ( ~n37235 & n37240 ) ;
  assign n37242 = ( n7318 & ~n37230 ) | ( n7318 & n37241 ) | ( ~n37230 & n37241 ) ;
  assign n37243 = ~n7318 & n37242 ;
  assign n37244 = ( x1151 & n37216 ) | ( x1151 & ~n37243 ) | ( n37216 & ~n37243 ) ;
  assign n37245 = ~n37216 & n37244 ;
  assign n37246 = ( x1152 & n37214 ) | ( x1152 & ~n37245 ) | ( n37214 & ~n37245 ) ;
  assign n37247 = ~x1152 & n37246 ;
  assign n37248 = x219 & ~n37196 ;
  assign n37249 = n37204 & ~n37224 ;
  assign n37250 = x214 & ~n37249 ;
  assign n37251 = ( ~x212 & n37227 ) | ( ~x212 & n37250 ) | ( n37227 & n37250 ) ;
  assign n37252 = ( x219 & ~n37250 ) | ( x219 & n37251 ) | ( ~n37250 & n37251 ) ;
  assign n37253 = n37252 ^ x212 ^ 1'b0 ;
  assign n37254 = n37223 ^ x214 ^ 1'b0 ;
  assign n37255 = ( n37223 & n37249 ) | ( n37223 & ~n37254 ) | ( n37249 & ~n37254 ) ;
  assign n37256 = n37255 ^ n37250 ^ n37236 ;
  assign n37257 = ( x212 & ~n37253 ) | ( x212 & n37256 ) | ( ~n37253 & n37256 ) ;
  assign n37258 = ( n37252 & n37253 ) | ( n37252 & n37257 ) | ( n37253 & n37257 ) ;
  assign n37259 = ( n7318 & ~n37248 ) | ( n7318 & n37258 ) | ( ~n37248 & n37258 ) ;
  assign n37260 = ~n7318 & n37259 ;
  assign n37261 = ~n9272 & n36297 ;
  assign n37262 = n7318 & n37261 ;
  assign n37263 = n9344 ^ x211 ^ 1'b0 ;
  assign n37264 = x211 | x1153 ;
  assign n37265 = ( ~x211 & n37263 ) | ( ~x211 & n37264 ) | ( n37263 & n37264 ) ;
  assign n37266 = n37262 & n37265 ;
  assign n37267 = ( x1151 & ~n37260 ) | ( x1151 & n37266 ) | ( ~n37260 & n37266 ) ;
  assign n37268 = n37260 | n37267 ;
  assign n37269 = n9275 & n36038 ;
  assign n37270 = x1151 & ~n37269 ;
  assign n37271 = ( n37241 & n37255 ) | ( n37241 & n37258 ) | ( n37255 & n37258 ) ;
  assign n37272 = ( n7318 & ~n37230 ) | ( n7318 & n37271 ) | ( ~n37230 & n37271 ) ;
  assign n37273 = ~n7318 & n37272 ;
  assign n37274 = ( n37266 & n37270 ) | ( n37266 & ~n37273 ) | ( n37270 & ~n37273 ) ;
  assign n37275 = ~n37266 & n37274 ;
  assign n37276 = x1152 & ~n37275 ;
  assign n37277 = n37268 & n37276 ;
  assign n37278 = ( x209 & n37247 ) | ( x209 & ~n37277 ) | ( n37247 & ~n37277 ) ;
  assign n37279 = ~n37247 & n37278 ;
  assign n37285 = x299 | n36977 ;
  assign n37286 = ~x208 & n37285 ;
  assign n37287 = x200 & ~n36141 ;
  assign n37282 = n36088 & n36591 ;
  assign n37288 = n37282 ^ n36591 ^ x208 ;
  assign n37289 = ~n37287 & n37288 ;
  assign n37290 = n37286 | n37289 ;
  assign n37291 = x211 & n37290 ;
  assign n37280 = n9233 | n36106 ;
  assign n37281 = n36394 & ~n37280 ;
  assign n37283 = n37281 | n37282 ;
  assign n37284 = x211 & n37283 ;
  assign n37292 = n37291 ^ n37290 ^ n37284 ;
  assign n37293 = n36645 & n37292 ;
  assign n37294 = ~x214 & n37293 ;
  assign n37295 = n36558 & n37283 ;
  assign n37296 = ~n36216 & n36395 ;
  assign n37297 = x1153 & n37296 ;
  assign n37298 = n11549 | n37297 ;
  assign n37299 = n37295 | n37298 ;
  assign n37300 = ( x212 & n36069 ) | ( x212 & ~n37299 ) | ( n36069 & ~n37299 ) ;
  assign n37301 = ( x212 & ~x214 ) | ( x212 & n37300 ) | ( ~x214 & n37300 ) ;
  assign n37302 = ~n37294 & n37301 ;
  assign n37303 = n36035 | n37295 ;
  assign n37304 = n37293 & n37303 ;
  assign n37305 = x212 | n37304 ;
  assign n37306 = n37305 ^ n37302 ^ 1'b0 ;
  assign n37307 = ( n37302 & n37305 ) | ( n37302 & n37306 ) | ( n37305 & n37306 ) ;
  assign n37308 = ( x219 & ~n37302 ) | ( x219 & n37307 ) | ( ~n37302 & n37307 ) ;
  assign n37309 = ~x211 & x299 ;
  assign n37310 = n37297 | n37309 ;
  assign n37311 = n37295 | n37310 ;
  assign n37312 = n37303 & n37311 ;
  assign n37313 = x219 & ~n37312 ;
  assign n37314 = ( n7318 & n37308 ) | ( n7318 & ~n37313 ) | ( n37308 & ~n37313 ) ;
  assign n37315 = ~n7318 & n37314 ;
  assign n37316 = ( x1151 & n37216 ) | ( x1151 & ~n37315 ) | ( n37216 & ~n37315 ) ;
  assign n37317 = ~n37216 & n37316 ;
  assign n37318 = x1151 | n37212 ;
  assign n37319 = x214 | n37296 ;
  assign n37320 = ~n9353 & n36395 ;
  assign n37321 = x299 | n37320 ;
  assign n37322 = ~n11549 & n37321 ;
  assign n37323 = x212 | n37319 ;
  assign n37324 = n37322 & n37323 ;
  assign n37325 = x1153 & n37324 ;
  assign n37326 = ~n37319 & n37325 ;
  assign n37327 = x212 & n37319 ;
  assign n37328 = n37298 & n37327 ;
  assign n37329 = x219 | n37328 ;
  assign n37330 = ~x211 & n36015 ;
  assign n37331 = n36014 & n37330 ;
  assign n37332 = n37296 | n37331 ;
  assign n37333 = ( ~n37326 & n37329 ) | ( ~n37326 & n37332 ) | ( n37329 & n37332 ) ;
  assign n37334 = n37326 | n37333 ;
  assign n37335 = x219 & ~n37296 ;
  assign n37336 = n7318 | n37335 ;
  assign n37337 = n37325 & ~n37336 ;
  assign n37338 = n37334 & n37337 ;
  assign n37339 = n37318 | n37338 ;
  assign n37340 = ( x1152 & ~n37317 ) | ( x1152 & n37339 ) | ( ~n37317 & n37339 ) ;
  assign n37341 = ~x1152 & n37340 ;
  assign n37342 = x208 & ~n36112 ;
  assign n37343 = ( n36141 & n36508 ) | ( n36141 & n37342 ) | ( n36508 & n37342 ) ;
  assign n37344 = ~x211 & n37343 ;
  assign n37345 = ( n36000 & n36089 ) | ( n36000 & n37342 ) | ( n36089 & n37342 ) ;
  assign n37346 = n37297 | n37345 ;
  assign n37347 = n37344 | n37346 ;
  assign n37350 = x214 | n37345 ;
  assign n37351 = n37297 | n37350 ;
  assign n37352 = ~x212 & n37351 ;
  assign n37348 = x214 & ~n37347 ;
  assign n37349 = x212 & ~n37348 ;
  assign n37353 = n37352 ^ n37349 ^ n37348 ;
  assign n37354 = n37347 & n37353 ;
  assign n37355 = x219 & ~n37354 ;
  assign n37356 = x211 & n37343 ;
  assign n37357 = x1153 & n37321 ;
  assign n37358 = n37356 | n37357 ;
  assign n37359 = x214 & ~n37345 ;
  assign n37360 = ~n37358 & n37359 ;
  assign n37361 = n37352 & ~n37360 ;
  assign n37362 = x214 & ~n37343 ;
  assign n37363 = x212 & ~n37362 ;
  assign n37364 = n37350 | n37358 ;
  assign n37365 = n37363 & n37364 ;
  assign n37366 = ( x219 & ~n37361 ) | ( x219 & n37365 ) | ( ~n37361 & n37365 ) ;
  assign n37367 = n37361 | n37366 ;
  assign n37368 = ( n7318 & ~n37355 ) | ( n7318 & n37367 ) | ( ~n37355 & n37367 ) ;
  assign n37369 = ~n7318 & n37368 ;
  assign n37370 = ( n37266 & n37270 ) | ( n37266 & ~n37369 ) | ( n37270 & ~n37369 ) ;
  assign n37371 = ~n37266 & n37370 ;
  assign n37372 = x1151 | n37266 ;
  assign n37373 = n9233 | n36505 ;
  assign n37374 = n36395 | n36977 ;
  assign n37375 = ~n10019 & n37374 ;
  assign n37376 = n37373 & n37375 ;
  assign n37377 = x219 & ~n37376 ;
  assign n37378 = ~n36369 & n37376 ;
  assign n37379 = n36507 ^ x207 ^ 1'b0 ;
  assign n37380 = ( ~n9354 & n36507 ) | ( ~n9354 & n37379 ) | ( n36507 & n37379 ) ;
  assign n37381 = x208 & n37380 ;
  assign n37382 = n37381 ^ n36142 ^ 1'b0 ;
  assign n37383 = ( ~n36142 & n36507 ) | ( ~n36142 & n37382 ) | ( n36507 & n37382 ) ;
  assign n37384 = ( n36142 & n37381 ) | ( n36142 & n37383 ) | ( n37381 & n37383 ) ;
  assign n37385 = n36069 & n37384 ;
  assign n37386 = x200 & x207 ;
  assign n37387 = x199 | n37386 ;
  assign n37388 = ~x299 & n37387 ;
  assign n37389 = x208 & ~n37388 ;
  assign n37390 = n10074 | n36581 ;
  assign n37391 = x207 & ~n37390 ;
  assign n37392 = ( x208 & n36655 ) | ( x208 & ~n37391 ) | ( n36655 & ~n37391 ) ;
  assign n37393 = ~x208 & n37392 ;
  assign n37394 = ( x207 & ~x299 ) | ( x207 & n9354 ) | ( ~x299 & n9354 ) ;
  assign n37395 = x1153 | n37394 ;
  assign n37396 = n37393 ^ n37389 ^ 1'b0 ;
  assign n37397 = ( ~n37389 & n37395 ) | ( ~n37389 & n37396 ) | ( n37395 & n37396 ) ;
  assign n37398 = ( n37389 & n37393 ) | ( n37389 & n37397 ) | ( n37393 & n37397 ) ;
  assign n37399 = x211 | n37398 ;
  assign n37400 = n37385 & n37399 ;
  assign n37401 = x299 & n36307 ;
  assign n37402 = x219 | n37401 ;
  assign n37403 = ( ~n37378 & n37400 ) | ( ~n37378 & n37402 ) | ( n37400 & n37402 ) ;
  assign n37404 = n37378 | n37403 ;
  assign n37405 = ( n7318 & ~n37377 ) | ( n7318 & n37404 ) | ( ~n37377 & n37404 ) ;
  assign n37406 = ~n7318 & n37405 ;
  assign n37407 = ( x1152 & n37372 ) | ( x1152 & n37406 ) | ( n37372 & n37406 ) ;
  assign n37408 = n37406 ^ n37372 ^ 1'b0 ;
  assign n37409 = ( x1152 & n37407 ) | ( x1152 & n37408 ) | ( n37407 & n37408 ) ;
  assign n37410 = n37409 ^ n37371 ^ 1'b0 ;
  assign n37411 = ( n37371 & n37409 ) | ( n37371 & n37410 ) | ( n37409 & n37410 ) ;
  assign n37412 = ( n37341 & ~n37371 ) | ( n37341 & n37411 ) | ( ~n37371 & n37411 ) ;
  assign n37413 = x209 | n37412 ;
  assign n37414 = ( x213 & ~n37279 ) | ( x213 & n37413 ) | ( ~n37279 & n37413 ) ;
  assign n37415 = ~x213 & n37414 ;
  assign n37416 = x219 & ~n37304 ;
  assign n37417 = x214 | n37295 ;
  assign n37418 = ~x212 & n37417 ;
  assign n37419 = n36208 | n37288 ;
  assign n37420 = n37419 ^ n37282 ^ 1'b0 ;
  assign n37421 = ~n36106 & n36527 ;
  assign n37422 = x1153 & n36094 ;
  assign n37423 = x1153 | n36165 ;
  assign n37424 = ~n37422 & n37423 ;
  assign n37425 = x1155 & n37424 ;
  assign n37426 = n37421 | n37425 ;
  assign n37427 = ( n37419 & ~n37420 ) | ( n37419 & n37426 ) | ( ~n37420 & n37426 ) ;
  assign n37428 = ( n37282 & n37420 ) | ( n37282 & n37427 ) | ( n37420 & n37427 ) ;
  assign n37429 = n36140 | n37428 ;
  assign n37430 = n37429 ^ x219 ^ 1'b0 ;
  assign n37431 = ~n36017 & n36271 ;
  assign n37432 = ~n37295 & n37431 ;
  assign n37433 = n36645 & n37290 ;
  assign n37434 = n9271 & ~n37433 ;
  assign n37435 = ( x212 & n37432 ) | ( x212 & ~n37434 ) | ( n37432 & ~n37434 ) ;
  assign n37436 = ~n37432 & n37435 ;
  assign n37437 = ( n37429 & ~n37430 ) | ( n37429 & n37436 ) | ( ~n37430 & n37436 ) ;
  assign n37438 = ( x219 & n37430 ) | ( x219 & n37437 ) | ( n37430 & n37437 ) ;
  assign n37439 = x299 & n35965 ;
  assign n37440 = x214 & ~n37439 ;
  assign n37441 = ~x299 & n37428 ;
  assign n37442 = n37440 & ~n37441 ;
  assign n37443 = ~n37438 & n37442 ;
  assign n37444 = ( n37418 & n37438 ) | ( n37418 & ~n37443 ) | ( n37438 & ~n37443 ) ;
  assign n37445 = x1151 & ~n7318 ;
  assign n37446 = ( n37416 & n37444 ) | ( n37416 & n37445 ) | ( n37444 & n37445 ) ;
  assign n37447 = ~n37416 & n37446 ;
  assign n37448 = n36451 & n37321 ;
  assign n37449 = n36017 | n37297 ;
  assign n37450 = ~x211 & n37449 ;
  assign n37451 = ( n9344 & n37448 ) | ( n9344 & ~n37450 ) | ( n37448 & ~n37450 ) ;
  assign n37452 = ~n37448 & n37451 ;
  assign n37453 = n36069 & ~n37439 ;
  assign n37454 = ~n37297 & n37453 ;
  assign n37455 = ( ~x219 & n37452 ) | ( ~x219 & n37454 ) | ( n37452 & n37454 ) ;
  assign n37456 = ~x219 & n37455 ;
  assign n37457 = x1151 | n7318 ;
  assign n37458 = n36297 | n37325 ;
  assign n37459 = ( n37456 & ~n37457 ) | ( n37456 & n37458 ) | ( ~n37457 & n37458 ) ;
  assign n37460 = ~n37456 & n37459 ;
  assign n37461 = ( x1152 & ~n37447 ) | ( x1152 & n37460 ) | ( ~n37447 & n37460 ) ;
  assign n37462 = n37447 | n37461 ;
  assign n37463 = x211 & n37398 ;
  assign n37464 = x211 | n36150 ;
  assign n37465 = n37384 & ~n37464 ;
  assign n37466 = n37463 | n37465 ;
  assign n37467 = n9344 & n37466 ;
  assign n37468 = x299 & ~n35965 ;
  assign n37469 = n37385 & ~n37468 ;
  assign n37470 = ( ~x219 & n37467 ) | ( ~x219 & n37469 ) | ( n37467 & n37469 ) ;
  assign n37471 = ~x219 & n37470 ;
  assign n37472 = n36035 & n37330 ;
  assign n37473 = ( ~n36297 & n37376 ) | ( ~n36297 & n37472 ) | ( n37376 & n37472 ) ;
  assign n37474 = ~n36297 & n37473 ;
  assign n37475 = ( ~n37457 & n37471 ) | ( ~n37457 & n37474 ) | ( n37471 & n37474 ) ;
  assign n37476 = ~n37457 & n37475 ;
  assign n37477 = x219 & ~n37345 ;
  assign n37478 = ~n37325 & n37477 ;
  assign n37479 = ~n36150 & n37356 ;
  assign n37480 = ~n36180 & n37344 ;
  assign n37481 = ( n36069 & n37479 ) | ( n36069 & n37480 ) | ( n37479 & n37480 ) ;
  assign n37482 = n37480 ^ n37479 ^ 1'b0 ;
  assign n37483 = ( n36069 & n37481 ) | ( n36069 & n37482 ) | ( n37481 & n37482 ) ;
  assign n37484 = n37345 | n37448 ;
  assign n37485 = n37465 | n37484 ;
  assign n37486 = n9344 & n37485 ;
  assign n37487 = ~x214 & n37352 ;
  assign n37488 = x219 | n37487 ;
  assign n37489 = ( ~n37483 & n37486 ) | ( ~n37483 & n37488 ) | ( n37486 & n37488 ) ;
  assign n37490 = n37483 | n37489 ;
  assign n37491 = ( n37445 & n37478 ) | ( n37445 & n37490 ) | ( n37478 & n37490 ) ;
  assign n37492 = ~n37478 & n37491 ;
  assign n37493 = ( x1152 & n37476 ) | ( x1152 & ~n37492 ) | ( n37476 & ~n37492 ) ;
  assign n37494 = ~n37476 & n37493 ;
  assign n37495 = ( x209 & n37462 ) | ( x209 & ~n37494 ) | ( n37462 & ~n37494 ) ;
  assign n37496 = n37495 ^ n37462 ^ 1'b0 ;
  assign n37497 = ( x209 & n37495 ) | ( x209 & ~n37496 ) | ( n37495 & ~n37496 ) ;
  assign n37498 = x219 & ~n37264 ;
  assign n37499 = ( n36038 & n36906 ) | ( n36038 & n37498 ) | ( n36906 & n37498 ) ;
  assign n37500 = ~n37498 & n37499 ;
  assign n37504 = n36112 & n36577 ;
  assign n37505 = n36787 & ~n37504 ;
  assign n37506 = n37222 & n37505 ;
  assign n37507 = n36786 | n37506 ;
  assign n37508 = ~x211 & n37507 ;
  assign n37509 = n36533 | n37193 ;
  assign n37510 = ( n36162 & n36839 ) | ( n36162 & n37509 ) | ( n36839 & n37509 ) ;
  assign n37511 = ( n36837 & n36838 ) | ( n36837 & n37510 ) | ( n36838 & n37510 ) ;
  assign n37512 = x211 & n37511 ;
  assign n37513 = ( n36014 & n37508 ) | ( n36014 & ~n37512 ) | ( n37508 & ~n37512 ) ;
  assign n37514 = ~n37508 & n37513 ;
  assign n37515 = n9271 & n37203 ;
  assign n37516 = ~n36140 & n37507 ;
  assign n37517 = ( x212 & n37515 ) | ( x212 & ~n37516 ) | ( n37515 & ~n37516 ) ;
  assign n37518 = ~n37515 & n37517 ;
  assign n37519 = ( n36271 & n37511 ) | ( n36271 & ~n37518 ) | ( n37511 & ~n37518 ) ;
  assign n37520 = n37519 ^ n37518 ^ 1'b0 ;
  assign n37521 = ( n37518 & ~n37519 ) | ( n37518 & n37520 ) | ( ~n37519 & n37520 ) ;
  assign n37522 = ( ~x219 & n37514 ) | ( ~x219 & n37521 ) | ( n37514 & n37521 ) ;
  assign n37523 = ~x219 & n37522 ;
  assign n37501 = ~n7318 & n37228 ;
  assign n37502 = n36621 & ~n37205 ;
  assign n37503 = n37501 & ~n37502 ;
  assign n37524 = n37523 ^ n37503 ^ 1'b0 ;
  assign n37525 = ( x209 & ~n37503 ) | ( x209 & n37523 ) | ( ~n37503 & n37523 ) ;
  assign n37526 = ( x209 & ~n37524 ) | ( x209 & n37525 ) | ( ~n37524 & n37525 ) ;
  assign n37527 = ~n37500 & n37526 ;
  assign n37528 = ( n37497 & n37500 ) | ( n37497 & ~n37527 ) | ( n37500 & ~n37527 ) ;
  assign n37529 = ( ~x213 & n37414 ) | ( ~x213 & n37528 ) | ( n37414 & n37528 ) ;
  assign n37530 = ( x213 & n37415 ) | ( x213 & n37529 ) | ( n37415 & n37529 ) ;
  assign n37531 = x238 ^ x230 ^ 1'b0 ;
  assign n37532 = ( x238 & n37530 ) | ( x238 & n37531 ) | ( n37530 & n37531 ) ;
  assign n37533 = n37005 & n37050 ;
  assign n37534 = ~x214 & n37533 ;
  assign n37535 = x212 | n37534 ;
  assign n37536 = x219 & ~n37535 ;
  assign n37537 = x211 & ~n37533 ;
  assign n37538 = n36599 | n37533 ;
  assign n37539 = x214 & n37538 ;
  assign n37540 = ~n37537 & n37539 ;
  assign n37541 = n37536 & ~n37540 ;
  assign n37542 = x208 & x299 ;
  assign n37543 = x1157 & ~n37542 ;
  assign n37544 = ~n36997 & n37543 ;
  assign n37545 = x211 & ~n37050 ;
  assign n37546 = ( x211 & n37544 ) | ( x211 & n37545 ) | ( n37544 & n37545 ) ;
  assign n37547 = x208 & ~n37016 ;
  assign n37548 = ( n36250 & n37022 ) | ( n36250 & ~n37547 ) | ( n37022 & ~n37547 ) ;
  assign n37549 = ~n36250 & n37548 ;
  assign n37550 = ( x211 & n37019 ) | ( x211 & ~n37549 ) | ( n37019 & ~n37549 ) ;
  assign n37551 = n37549 | n37550 ;
  assign n37552 = ( x214 & n37546 ) | ( x214 & n37551 ) | ( n37546 & n37551 ) ;
  assign n37553 = ~n37546 & n37552 ;
  assign n37554 = ( x219 & n37535 ) | ( x219 & ~n37553 ) | ( n37535 & ~n37553 ) ;
  assign n37555 = n37553 | n37554 ;
  assign n37556 = x212 & ~n37533 ;
  assign n37557 = n7318 | n37556 ;
  assign n37558 = x209 & ~n37557 ;
  assign n37559 = ( n37541 & n37555 ) | ( n37541 & n37558 ) | ( n37555 & n37558 ) ;
  assign n37560 = ~n37541 & n37559 ;
  assign n37561 = n7318 & ~n36945 ;
  assign n37562 = x219 | n36936 ;
  assign n37563 = x213 & ~n37562 ;
  assign n37564 = ( x213 & ~n37561 ) | ( x213 & n37563 ) | ( ~n37561 & n37563 ) ;
  assign n37565 = n36009 & n36104 ;
  assign n37566 = x212 & ~n37565 ;
  assign n37567 = n7318 | n37566 ;
  assign n37568 = x209 | n37567 ;
  assign n37569 = n36142 & ~n36461 ;
  assign n37570 = n37543 & ~n37569 ;
  assign n37571 = x1157 | n37565 ;
  assign n37572 = ( x211 & n37570 ) | ( x211 & n37571 ) | ( n37570 & n37571 ) ;
  assign n37573 = ~n37570 & n37572 ;
  assign n37574 = ~n36009 & n37016 ;
  assign n37575 = ~x208 & n37026 ;
  assign n37576 = ( ~x211 & n37574 ) | ( ~x211 & n37575 ) | ( n37574 & n37575 ) ;
  assign n37577 = ~x211 & n37576 ;
  assign n37578 = ( x214 & n37573 ) | ( x214 & n37577 ) | ( n37573 & n37577 ) ;
  assign n37579 = n37577 ^ n37573 ^ 1'b0 ;
  assign n37580 = ( x214 & n37578 ) | ( x214 & n37579 ) | ( n37578 & n37579 ) ;
  assign n37581 = ~x214 & n37565 ;
  assign n37582 = x212 | n37581 ;
  assign n37583 = ( x219 & ~n37580 ) | ( x219 & n37582 ) | ( ~n37580 & n37582 ) ;
  assign n37584 = n37580 | n37583 ;
  assign n37585 = x219 & ~n37582 ;
  assign n37586 = x211 & ~n37565 ;
  assign n37587 = x214 & ~n37586 ;
  assign n37588 = ~x208 & n36422 ;
  assign n37589 = n36599 | n37588 ;
  assign n37590 = n37587 & n37589 ;
  assign n37591 = n37585 & ~n37590 ;
  assign n37592 = ( n37568 & n37584 ) | ( n37568 & ~n37591 ) | ( n37584 & ~n37591 ) ;
  assign n37593 = ~n37568 & n37592 ;
  assign n37594 = ( n37560 & n37564 ) | ( n37560 & ~n37593 ) | ( n37564 & ~n37593 ) ;
  assign n37595 = ~n37560 & n37594 ;
  assign n37596 = x211 | n36017 ;
  assign n37597 = n37093 | n37596 ;
  assign n37598 = x214 & ~n37537 ;
  assign n37599 = n37536 & ~n37598 ;
  assign n37600 = ( n37536 & ~n37597 ) | ( n37536 & n37599 ) | ( ~n37597 & n37599 ) ;
  assign n37601 = x219 | n37535 ;
  assign n37602 = x211 & ~n36021 ;
  assign n37603 = ~n37093 & n37602 ;
  assign n37604 = n37539 & ~n37603 ;
  assign n37605 = n37601 | n37604 ;
  assign n37606 = ~n37557 & n37605 ;
  assign n37607 = x209 & ~n37606 ;
  assign n37608 = ( x209 & n37600 ) | ( x209 & n37607 ) | ( n37600 & n37607 ) ;
  assign n37609 = ~x208 & n36408 ;
  assign n37610 = n36017 | n37609 ;
  assign n37611 = n37585 & ~n37610 ;
  assign n37612 = ( n37585 & ~n37587 ) | ( n37585 & n37611 ) | ( ~n37587 & n37611 ) ;
  assign n37613 = n36208 & n36430 ;
  assign n37614 = n37602 & ~n37613 ;
  assign n37615 = ( x214 & n37589 ) | ( x214 & n37614 ) | ( n37589 & n37614 ) ;
  assign n37616 = ~n37614 & n37615 ;
  assign n37617 = ( x219 & n37582 ) | ( x219 & ~n37616 ) | ( n37582 & ~n37616 ) ;
  assign n37618 = n37616 | n37617 ;
  assign n37619 = ( n37567 & ~n37612 ) | ( n37567 & n37618 ) | ( ~n37612 & n37618 ) ;
  assign n37620 = ~n37567 & n37619 ;
  assign n37621 = ( x209 & ~n37608 ) | ( x209 & n37620 ) | ( ~n37608 & n37620 ) ;
  assign n37622 = ~n37608 & n37621 ;
  assign n37623 = n7318 & ~n36390 ;
  assign n37624 = n36014 & n36388 ;
  assign n37625 = n37623 & n37624 ;
  assign n37626 = x213 | n37625 ;
  assign n37627 = ( ~n37595 & n37622 ) | ( ~n37595 & n37626 ) | ( n37622 & n37626 ) ;
  assign n37628 = ~n37595 & n37627 ;
  assign n37629 = x239 ^ x230 ^ 1'b0 ;
  assign n37630 = ( x239 & n37628 ) | ( x239 & n37629 ) | ( n37628 & n37629 ) ;
  assign n37631 = ~n15098 & n37320 ;
  assign n37633 = x211 & x1145 ;
  assign n37632 = x211 & x1146 ;
  assign n37634 = n37633 ^ n37632 ^ x1146 ;
  assign n37635 = x214 & n37634 ;
  assign n37636 = ~x214 & n37632 ;
  assign n37637 = n37635 | n37636 ;
  assign n37638 = x212 & n37637 ;
  assign n37639 = n36014 & n37632 ;
  assign n37640 = n37638 | n37639 ;
  assign n37641 = n36621 | n37640 ;
  assign n37642 = x219 & ~n37075 ;
  assign n37643 = n7318 & ~n37642 ;
  assign n37644 = n37641 & n37643 ;
  assign n37645 = x1147 | n37644 ;
  assign n37650 = x219 | n7318 ;
  assign n37651 = x299 & n37640 ;
  assign n37652 = ~n37650 & n37651 ;
  assign n37646 = n7318 | n36037 ;
  assign n37647 = ~x211 & n37100 ;
  assign n37648 = x219 & ~n37647 ;
  assign n37649 = n37646 | n37648 ;
  assign n37653 = n37652 ^ n37650 ^ n37649 ;
  assign n37654 = n37645 | n37653 ;
  assign n37655 = n37631 | n37654 ;
  assign n37656 = ~n9741 & n36297 ;
  assign n37657 = n7318 & n37656 ;
  assign n37658 = x1147 & ~n37657 ;
  assign n37659 = ~n37644 & n37658 ;
  assign n37660 = x219 & ~n37283 ;
  assign n37661 = n7318 | n37660 ;
  assign n37662 = n37649 & n37661 ;
  assign n37663 = x214 | n37283 ;
  assign n37664 = ~x212 & n37663 ;
  assign n37665 = ~x211 & n37290 ;
  assign n37666 = x299 & x1146 ;
  assign n37667 = x211 & n37666 ;
  assign n37668 = ( ~n36112 & n36954 ) | ( ~n36112 & n37289 ) | ( n36954 & n37289 ) ;
  assign n37669 = ( x211 & n37667 ) | ( x211 & n37668 ) | ( n37667 & n37668 ) ;
  assign n37670 = n37665 | n37669 ;
  assign n37671 = x214 & ~n37670 ;
  assign n37672 = n37664 & ~n37671 ;
  assign n37673 = x299 & n37634 ;
  assign n37674 = x214 & ~n37673 ;
  assign n37675 = ~n37668 & n37674 ;
  assign n37676 = x212 & ~n37675 ;
  assign n37677 = x214 | n37670 ;
  assign n37678 = n37676 & n37677 ;
  assign n37679 = ( x219 & ~n37672 ) | ( x219 & n37678 ) | ( ~n37672 & n37678 ) ;
  assign n37680 = n37672 | n37679 ;
  assign n37681 = n37659 & ~n37680 ;
  assign n37682 = ( n37659 & n37662 ) | ( n37659 & n37681 ) | ( n37662 & n37681 ) ;
  assign n37683 = ( x1148 & n37655 ) | ( x1148 & ~n37682 ) | ( n37655 & ~n37682 ) ;
  assign n37684 = ~x1148 & n37683 ;
  assign n37685 = ~n36112 & n36394 ;
  assign n37686 = x219 & ~n37685 ;
  assign n37687 = x211 & ~n37685 ;
  assign n37688 = x214 & x299 ;
  assign n37689 = ( ~x212 & n37685 ) | ( ~x212 & n37688 ) | ( n37685 & n37688 ) ;
  assign n37690 = ~n37687 & n37689 ;
  assign n37691 = x212 & n36140 ;
  assign n37692 = x299 & n37691 ;
  assign n37693 = ( x212 & x299 ) | ( x212 & n37685 ) | ( x299 & n37685 ) ;
  assign n37694 = ~n37692 & n37693 ;
  assign n37695 = ( x219 & ~n37690 ) | ( x219 & n37694 ) | ( ~n37690 & n37694 ) ;
  assign n37696 = n37690 | n37695 ;
  assign n37697 = ( n7318 & ~n37686 ) | ( n7318 & n37696 ) | ( ~n37686 & n37696 ) ;
  assign n37698 = ~n7318 & n37697 ;
  assign n37699 = ~n37653 & n37659 ;
  assign n37700 = ~n37698 & n37699 ;
  assign n37701 = x1148 & ~n37700 ;
  assign n37702 = ~x199 & n36009 ;
  assign n37703 = ( x299 & n37389 ) | ( x299 & ~n37702 ) | ( n37389 & ~n37702 ) ;
  assign n37704 = n37702 | n37703 ;
  assign n37705 = x212 & n37704 ;
  assign n37706 = n37375 | n37637 ;
  assign n37707 = n37705 & n37706 ;
  assign n37708 = x214 | n37375 ;
  assign n37709 = ~x212 & n37708 ;
  assign n37710 = ~x212 & n37375 ;
  assign n37711 = ( n37667 & n37709 ) | ( n37667 & n37710 ) | ( n37709 & n37710 ) ;
  assign n37712 = ( x219 & ~n37707 ) | ( x219 & n37711 ) | ( ~n37707 & n37711 ) ;
  assign n37713 = n37707 | n37712 ;
  assign n37714 = ~n36036 & n37375 ;
  assign n37715 = ~x211 & n37704 ;
  assign n37716 = n36035 & n37715 ;
  assign n37717 = ( x219 & n37714 ) | ( x219 & ~n37716 ) | ( n37714 & ~n37716 ) ;
  assign n37718 = ~n37714 & n37717 ;
  assign n37719 = n7318 | n37718 ;
  assign n37720 = n10019 | n37719 ;
  assign n37721 = ( n37649 & ~n37713 ) | ( n37649 & n37720 ) | ( ~n37713 & n37720 ) ;
  assign n37722 = n37721 ^ n37713 ^ 1'b0 ;
  assign n37723 = ( n37713 & ~n37721 ) | ( n37713 & n37722 ) | ( ~n37721 & n37722 ) ;
  assign n37724 = ( x1147 & n37644 ) | ( x1147 & ~n37723 ) | ( n37644 & ~n37723 ) ;
  assign n37725 = n37723 | n37724 ;
  assign n37726 = n37701 & n37725 ;
  assign n37727 = ( x1149 & n37684 ) | ( x1149 & ~n37726 ) | ( n37684 & ~n37726 ) ;
  assign n37728 = ~n37684 & n37727 ;
  assign n37731 = ( n9344 & n37345 ) | ( n9344 & n37673 ) | ( n37345 & n37673 ) ;
  assign n37729 = ~n36035 & n37345 ;
  assign n37730 = x219 | n37729 ;
  assign n37732 = n37309 | n37345 ;
  assign n37733 = ( n36369 & n37667 ) | ( n36369 & n37732 ) | ( n37667 & n37732 ) ;
  assign n37734 = ( n37730 & ~n37731 ) | ( n37730 & n37733 ) | ( ~n37731 & n37733 ) ;
  assign n37735 = n37731 | n37734 ;
  assign n37736 = ~n7318 & n37345 ;
  assign n37737 = n37736 ^ n37735 ^ 1'b0 ;
  assign n37738 = ( ~n37649 & n37736 ) | ( ~n37649 & n37737 ) | ( n37736 & n37737 ) ;
  assign n37739 = ( n37735 & ~n37737 ) | ( n37735 & n37738 ) | ( ~n37737 & n37738 ) ;
  assign n37740 = x1148 & ~n37659 ;
  assign n37741 = ( x1148 & n37739 ) | ( x1148 & n37740 ) | ( n37739 & n37740 ) ;
  assign n37742 = n36395 | n36677 ;
  assign n37743 = n9233 | n36181 ;
  assign n37744 = n37742 & n37743 ;
  assign n37745 = n37394 & n37744 ;
  assign n37746 = ~n7318 & n37745 ;
  assign n37747 = n37746 ^ n37654 ^ 1'b0 ;
  assign n37748 = ( n37654 & n37746 ) | ( n37654 & ~n37747 ) | ( n37746 & ~n37747 ) ;
  assign n37749 = ( n37741 & n37747 ) | ( n37741 & n37748 ) | ( n37747 & n37748 ) ;
  assign n37750 = n37075 & n37179 ;
  assign n37751 = n36165 | n37386 ;
  assign n37752 = x208 & n37751 ;
  assign n37753 = x199 | n37752 ;
  assign n37754 = n37345 & n37753 ;
  assign n37755 = ~n36297 & n37754 ;
  assign n37756 = n37750 | n37755 ;
  assign n37757 = x299 | n37754 ;
  assign n37758 = ~x1146 & n11549 ;
  assign n37759 = n36369 & ~n37758 ;
  assign n37760 = n37731 | n37759 ;
  assign n37761 = ( x219 & n37757 ) | ( x219 & n37760 ) | ( n37757 & n37760 ) ;
  assign n37762 = ~x219 & n37761 ;
  assign n37763 = ( ~n7318 & n37756 ) | ( ~n7318 & n37762 ) | ( n37756 & n37762 ) ;
  assign n37764 = ~n7318 & n37763 ;
  assign n37765 = ( n37644 & n37658 ) | ( n37644 & ~n37764 ) | ( n37658 & ~n37764 ) ;
  assign n37766 = ~n37644 & n37765 ;
  assign n37767 = ~x1148 & n37654 ;
  assign n37768 = n37767 ^ n37766 ^ 1'b0 ;
  assign n37769 = ( n37766 & n37767 ) | ( n37766 & n37768 ) | ( n37767 & n37768 ) ;
  assign n37770 = ( n37749 & ~n37766 ) | ( n37749 & n37769 ) | ( ~n37766 & n37769 ) ;
  assign n37771 = ( x1149 & ~n37728 ) | ( x1149 & n37770 ) | ( ~n37728 & n37770 ) ;
  assign n37772 = ~n37728 & n37771 ;
  assign n37773 = ( x209 & x213 ) | ( x209 & ~n37772 ) | ( x213 & ~n37772 ) ;
  assign n37774 = ( x209 & ~n36501 ) | ( x209 & n37773 ) | ( ~n36501 & n37773 ) ;
  assign n37775 = ~x211 & n7318 ;
  assign n37776 = n37211 | n37775 ;
  assign n37777 = n36035 & n37776 ;
  assign n37778 = x299 & n36035 ;
  assign n37779 = ~n37646 & n37778 ;
  assign n37780 = ~n7318 & n37685 ;
  assign n37781 = n37779 | n37780 ;
  assign n37782 = n37777 | n37781 ;
  assign n37783 = x1147 & ~n37782 ;
  assign n37784 = x1149 & ~n37783 ;
  assign n37785 = x211 & n36014 ;
  assign n37786 = x219 | n37785 ;
  assign n37787 = n37691 | n37786 ;
  assign n37788 = n37779 & n37787 ;
  assign n37789 = n36038 & n37787 ;
  assign n37790 = n37736 | n37789 ;
  assign n37791 = n37788 | n37790 ;
  assign n37792 = x1147 & ~n37791 ;
  assign n37793 = x1149 | n37792 ;
  assign n37794 = n37691 ^ n36271 ^ n36140 ;
  assign n37795 = n37211 & n37794 ;
  assign n37796 = x219 & ~n37745 ;
  assign n37797 = n7318 | n37796 ;
  assign n37798 = x299 & n9271 ;
  assign n37799 = n37745 | n37798 ;
  assign n37800 = ~x212 & n37799 ;
  assign n37801 = x219 | n37800 ;
  assign n37802 = x299 | n37744 ;
  assign n37803 = x214 & n37802 ;
  assign n37804 = ~x214 & n37745 ;
  assign n37805 = x212 | n37804 ;
  assign n37806 = n37803 | n37805 ;
  assign n37807 = ~x214 & n37802 ;
  assign n37808 = ~x211 & n37802 ;
  assign n37809 = n37745 | n37808 ;
  assign n37810 = x214 & n37809 ;
  assign n37811 = x212 & ~n37810 ;
  assign n37812 = n37806 & ~n37811 ;
  assign n37813 = ( n37806 & n37807 ) | ( n37806 & n37812 ) | ( n37807 & n37812 ) ;
  assign n37814 = ~x214 & n11549 ;
  assign n37815 = n37814 ^ n37804 ^ n37803 ;
  assign n37816 = x212 & n37815 ;
  assign n37817 = n37801 | n37816 ;
  assign n37818 = ( n37801 & n37813 ) | ( n37801 & n37817 ) | ( n37813 & n37817 ) ;
  assign n37819 = ~n37797 & n37818 ;
  assign n37820 = n37795 | n37819 ;
  assign n37821 = ( x1147 & ~n37793 ) | ( x1147 & n37820 ) | ( ~n37793 & n37820 ) ;
  assign n37822 = ~n37793 & n37821 ;
  assign n37823 = ~n7318 & n37375 ;
  assign n37824 = n37336 & ~n37823 ;
  assign n37825 = x211 & n37375 ;
  assign n37826 = x214 & ~n37825 ;
  assign n37827 = ~n37715 & n37826 ;
  assign n37828 = x212 & ~n37827 ;
  assign n37829 = x211 & n37704 ;
  assign n37830 = n37375 | n37829 ;
  assign n37831 = x214 | n37830 ;
  assign n37832 = n37828 & n37831 ;
  assign n37833 = x219 | n37832 ;
  assign n37834 = n37708 & n37830 ;
  assign n37835 = ~x212 & n37834 ;
  assign n37836 = n37833 | n37835 ;
  assign n37837 = x214 & ~n37704 ;
  assign n37838 = n37709 & ~n37837 ;
  assign n37839 = x219 | n37838 ;
  assign n37840 = n37705 | n37839 ;
  assign n37841 = ( n37715 & n37836 ) | ( n37715 & n37840 ) | ( n37836 & n37840 ) ;
  assign n37842 = ~n37824 & n37841 ;
  assign n37843 = n37262 | n37842 ;
  assign n37844 = x1147 | n37843 ;
  assign n37845 = n37822 ^ n37784 ^ 1'b0 ;
  assign n37846 = ( ~n37784 & n37844 ) | ( ~n37784 & n37845 ) | ( n37844 & n37845 ) ;
  assign n37847 = ( n37784 & n37822 ) | ( n37784 & n37846 ) | ( n37822 & n37846 ) ;
  assign n37848 = n9275 | n37209 ;
  assign n37849 = n36038 & n37848 ;
  assign n37850 = ~x211 & n37283 ;
  assign n37851 = x214 & ~n37291 ;
  assign n37852 = ~n37850 & n37851 ;
  assign n37853 = n9344 & ~n37852 ;
  assign n37854 = x214 & ~n37292 ;
  assign n37855 = n37664 & ~n37854 ;
  assign n37856 = x219 | n37855 ;
  assign n37857 = x212 & ~n37852 ;
  assign n37858 = n37292 & n37857 ;
  assign n37859 = n37856 | n37858 ;
  assign n37860 = n37853 | n37859 ;
  assign n37861 = x212 & n37292 ;
  assign n37862 = ( x219 & n37855 ) | ( x219 & ~n37861 ) | ( n37855 & ~n37861 ) ;
  assign n37863 = ~n37855 & n37862 ;
  assign n37864 = ( x57 & n5193 ) | ( x57 & ~n37863 ) | ( n5193 & ~n37863 ) ;
  assign n37865 = n37863 | n37864 ;
  assign n37866 = n37860 & ~n37865 ;
  assign n37867 = n37849 | n37866 ;
  assign n37868 = x1147 & ~n37867 ;
  assign n37869 = ~x219 & n15098 ;
  assign n37870 = n37209 & n37869 ;
  assign n37871 = n37631 | n37870 ;
  assign n37872 = x1147 | n37871 ;
  assign n37873 = ( x1149 & n37868 ) | ( x1149 & n37872 ) | ( n37868 & n37872 ) ;
  assign n37874 = ~n37868 & n37873 ;
  assign n37875 = n37350 & n37732 ;
  assign n37876 = x212 & ~n37814 ;
  assign n37877 = ~n37875 & n37876 ;
  assign n37878 = x212 | n37798 ;
  assign n37879 = ( n37345 & ~n37877 ) | ( n37345 & n37878 ) | ( ~n37877 & n37878 ) ;
  assign n37880 = ~n37877 & n37879 ;
  assign n37881 = x219 | n37880 ;
  assign n37882 = x219 | n37757 ;
  assign n37883 = n37881 & n37882 ;
  assign n37884 = x211 | n37883 ;
  assign n37885 = x214 | n37732 ;
  assign n37886 = x212 & n37885 ;
  assign n37887 = ~n11549 & n37359 ;
  assign n37888 = n37886 & ~n37887 ;
  assign n37889 = ~x212 & n37875 ;
  assign n37890 = x219 | n37889 ;
  assign n37891 = n37888 | n37890 ;
  assign n37892 = x219 & ~n37309 ;
  assign n37893 = n37646 | n37892 ;
  assign n37894 = ~n37736 & n37893 ;
  assign n37895 = n37891 & ~n37894 ;
  assign n37896 = n37757 & n37895 ;
  assign n37897 = n37884 & n37896 ;
  assign n37898 = n37269 | n37897 ;
  assign n37899 = n37898 ^ n37874 ^ 1'b0 ;
  assign n37900 = x1147 & ~x1149 ;
  assign n37901 = ( n37898 & ~n37899 ) | ( n37898 & n37900 ) | ( ~n37899 & n37900 ) ;
  assign n37902 = ( n37874 & n37899 ) | ( n37874 & n37901 ) | ( n37899 & n37901 ) ;
  assign n37903 = n37847 ^ x1148 ^ 1'b0 ;
  assign n37904 = ( n37847 & n37902 ) | ( n37847 & ~n37903 ) | ( n37902 & ~n37903 ) ;
  assign n37905 = ( x213 & ~n37774 ) | ( x213 & n37904 ) | ( ~n37774 & n37904 ) ;
  assign n37906 = n37905 ^ n37774 ^ 1'b0 ;
  assign n37907 = ( n37774 & ~n37905 ) | ( n37774 & n37906 ) | ( ~n37905 & n37906 ) ;
  assign n37908 = x200 & ~n37163 ;
  assign n37909 = n36000 & ~n37908 ;
  assign n37910 = x199 & x1145 ;
  assign n37911 = x200 | n37910 ;
  assign n37912 = ~x199 & x1146 ;
  assign n37913 = n37911 | n37912 ;
  assign n37914 = n37909 & n37913 ;
  assign n37915 = n37666 | n37914 ;
  assign n37916 = x200 & ~n37912 ;
  assign n37917 = x299 | n37916 ;
  assign n37923 = n37911 & ~n37917 ;
  assign n37918 = x199 & x1146 ;
  assign n37921 = n36164 & ~n37918 ;
  assign n37922 = n37917 | n37921 ;
  assign n37919 = x200 | n37918 ;
  assign n37920 = ~n37917 & n37919 ;
  assign n37924 = n37923 ^ n37922 ^ n37920 ;
  assign n37925 = x207 | n37924 ;
  assign n37926 = x208 & ~n37925 ;
  assign n37927 = ( x208 & n37915 ) | ( x208 & n37926 ) | ( n37915 & n37926 ) ;
  assign n37928 = n36009 & ~n37924 ;
  assign n37929 = n37927 | n37928 ;
  assign n37930 = x299 | n37929 ;
  assign n37931 = x211 & n37930 ;
  assign n37932 = ~n37102 & n37931 ;
  assign n37933 = n9271 & n37930 ;
  assign n37934 = n37674 & ~n37929 ;
  assign n37935 = n37933 | n37934 ;
  assign n37936 = ~n37932 & n37935 ;
  assign n37937 = n37309 | n37667 ;
  assign n37938 = x214 | n37937 ;
  assign n37939 = n37929 | n37938 ;
  assign n37940 = ( x212 & n37936 ) | ( x212 & n37939 ) | ( n37936 & n37939 ) ;
  assign n37941 = ~n37936 & n37940 ;
  assign n37942 = n36395 | n37914 ;
  assign n37943 = ~n9233 & n37924 ;
  assign n37944 = n37942 & ~n37943 ;
  assign n37945 = ~x211 & n37930 ;
  assign n37946 = n37944 | n37945 ;
  assign n37947 = x214 | n37944 ;
  assign n37948 = ~x212 & n37947 ;
  assign n37949 = n37946 & n37948 ;
  assign n37950 = n9233 | n37923 ;
  assign n37951 = n37942 & n37950 ;
  assign n37952 = n37667 | n37951 ;
  assign n37953 = ~x214 & n37951 ;
  assign n37954 = ( ~x212 & x214 ) | ( ~x212 & n37953 ) | ( x214 & n37953 ) ;
  assign n37955 = n37952 & n37954 ;
  assign n37956 = x219 | n37955 ;
  assign n37957 = ( ~n37941 & n37949 ) | ( ~n37941 & n37956 ) | ( n37949 & n37956 ) ;
  assign n37958 = n37941 | n37957 ;
  assign n37959 = ~n36036 & n37944 ;
  assign n37960 = x219 & ~n37959 ;
  assign n37961 = n36035 & n37945 ;
  assign n37962 = n37960 & ~n37961 ;
  assign n37963 = ( n37102 & n37960 ) | ( n37102 & n37962 ) | ( n37960 & n37962 ) ;
  assign n37964 = ( n7318 & n37958 ) | ( n7318 & ~n37963 ) | ( n37958 & ~n37963 ) ;
  assign n37965 = ~n7318 & n37964 ;
  assign n37966 = ( n37644 & n37658 ) | ( n37644 & ~n37965 ) | ( n37658 & ~n37965 ) ;
  assign n37967 = ~n37644 & n37966 ;
  assign n37968 = ~n36035 & n37951 ;
  assign n37969 = x219 & ~n37968 ;
  assign n37970 = n37911 | n37925 ;
  assign n37971 = n37927 & n37970 ;
  assign n37972 = n36009 & n37923 ;
  assign n37973 = n37971 | n37972 ;
  assign n37974 = ~x299 & n37973 ;
  assign n37975 = x211 | n37100 ;
  assign n37976 = n37974 | n37975 ;
  assign n37977 = n37969 & ~n37976 ;
  assign n37978 = ( n36035 & n36036 ) | ( n36035 & n37951 ) | ( n36036 & n37951 ) ;
  assign n37979 = ( n37969 & n37977 ) | ( n37969 & ~n37978 ) | ( n37977 & ~n37978 ) ;
  assign n37980 = n37674 & ~n37974 ;
  assign n37981 = x214 | n37952 ;
  assign n37982 = ( x212 & n37980 ) | ( x212 & n37981 ) | ( n37980 & n37981 ) ;
  assign n37983 = ~n37980 & n37982 ;
  assign n37984 = ( x219 & n37955 ) | ( x219 & ~n37983 ) | ( n37955 & ~n37983 ) ;
  assign n37985 = n37983 | n37984 ;
  assign n37986 = ( n7318 & ~n37979 ) | ( n7318 & n37985 ) | ( ~n37979 & n37985 ) ;
  assign n37987 = ~n7318 & n37986 ;
  assign n37988 = ( n37645 & ~n37967 ) | ( n37645 & n37987 ) | ( ~n37967 & n37987 ) ;
  assign n37989 = ~n37967 & n37988 ;
  assign n37990 = ~x213 & n37989 ;
  assign n37991 = x209 | n37990 ;
  assign n37992 = n7318 | n37962 ;
  assign n37993 = x219 | n37944 ;
  assign n37994 = x299 | n37973 ;
  assign n37995 = x214 & n37994 ;
  assign n37996 = n37931 | n37995 ;
  assign n37997 = x212 & n37996 ;
  assign n37998 = ( n37933 & ~n37993 ) | ( n37933 & n37997 ) | ( ~n37993 & n37997 ) ;
  assign n37999 = n37993 | n37998 ;
  assign n38000 = ~n37992 & n37999 ;
  assign n38001 = x1147 & ~n37789 ;
  assign n38002 = ~n38000 & n38001 ;
  assign n38003 = x219 & ~n37951 ;
  assign n38004 = ( x212 & ~n37953 ) | ( x212 & n37995 ) | ( ~n37953 & n37995 ) ;
  assign n38005 = n37953 | n38004 ;
  assign n38006 = x214 & ~n37946 ;
  assign n38007 = x212 & ~n37994 ;
  assign n38008 = ( x212 & n38006 ) | ( x212 & n38007 ) | ( n38006 & n38007 ) ;
  assign n38009 = ( x219 & n38005 ) | ( x219 & ~n38008 ) | ( n38005 & ~n38008 ) ;
  assign n38010 = n38009 ^ n38005 ^ 1'b0 ;
  assign n38011 = ( x219 & n38009 ) | ( x219 & ~n38010 ) | ( n38009 & ~n38010 ) ;
  assign n38012 = ( n7318 & ~n38003 ) | ( n7318 & n38011 ) | ( ~n38003 & n38011 ) ;
  assign n38013 = ~n7318 & n38012 ;
  assign n38014 = n37968 | n37999 ;
  assign n38015 = n38013 & n38014 ;
  assign n38016 = ( x1147 & n37795 ) | ( x1147 & ~n38015 ) | ( n37795 & ~n38015 ) ;
  assign n38017 = n38015 | n38016 ;
  assign n38018 = ( x1149 & ~n38002 ) | ( x1149 & n38017 ) | ( ~n38002 & n38017 ) ;
  assign n38019 = ~x1149 & n38018 ;
  assign n38021 = n37778 | n37993 ;
  assign n38022 = ~n37992 & n38021 ;
  assign n38020 = x1147 & ~n37777 ;
  assign n38023 = n38022 ^ n38020 ^ 1'b0 ;
  assign n38024 = ( x1149 & ~n38020 ) | ( x1149 & n38022 ) | ( ~n38020 & n38022 ) ;
  assign n38025 = ( x1149 & ~n38023 ) | ( x1149 & n38024 ) | ( ~n38023 & n38024 ) ;
  assign n38026 = x1147 | n37262 ;
  assign n38027 = n38026 ^ n38013 ^ 1'b0 ;
  assign n38028 = ( n38013 & n38026 ) | ( n38013 & ~n38027 ) | ( n38026 & ~n38027 ) ;
  assign n38029 = ( n38025 & n38027 ) | ( n38025 & n38028 ) | ( n38027 & n38028 ) ;
  assign n38030 = ( x1148 & n38019 ) | ( x1148 & ~n38029 ) | ( n38019 & ~n38029 ) ;
  assign n38031 = ~n38019 & n38030 ;
  assign n38032 = x1147 | n7318 ;
  assign n38033 = n37951 & ~n38032 ;
  assign n38034 = x214 & ~n37944 ;
  assign n38035 = ~n37931 & n38034 ;
  assign n38036 = n37945 | n37947 ;
  assign n38037 = ( x212 & n38035 ) | ( x212 & n38036 ) | ( n38035 & n38036 ) ;
  assign n38038 = ~n38035 & n38037 ;
  assign n38039 = ( x219 & ~n37949 ) | ( x219 & n38038 ) | ( ~n37949 & n38038 ) ;
  assign n38040 = n37949 | n38039 ;
  assign n38041 = n38000 & n38040 ;
  assign n38042 = n37269 | n38041 ;
  assign n38043 = x1147 & n38042 ;
  assign n38044 = ( ~x1149 & n38033 ) | ( ~x1149 & n38043 ) | ( n38033 & n38043 ) ;
  assign n38045 = ~x1149 & n38044 ;
  assign n38046 = ~n15098 & n37656 ;
  assign n38047 = ~n37973 & n38046 ;
  assign n38048 = ~x1147 & n37656 ;
  assign n38049 = ( n38033 & ~n38047 ) | ( n38033 & n38048 ) | ( ~n38047 & n38048 ) ;
  assign n38050 = ~n38047 & n38049 ;
  assign n38051 = ~n37992 & n38040 ;
  assign n38052 = n37849 | n38051 ;
  assign n38053 = x1147 & n38052 ;
  assign n38054 = ( x1149 & n38050 ) | ( x1149 & n38053 ) | ( n38050 & n38053 ) ;
  assign n38055 = n38053 ^ n38050 ^ 1'b0 ;
  assign n38056 = ( x1149 & n38054 ) | ( x1149 & n38055 ) | ( n38054 & n38055 ) ;
  assign n38057 = ( x1148 & ~n38045 ) | ( x1148 & n38056 ) | ( ~n38045 & n38056 ) ;
  assign n38058 = n38045 | n38057 ;
  assign n38059 = ( x213 & n38031 ) | ( x213 & n38058 ) | ( n38031 & n38058 ) ;
  assign n38060 = ~n38031 & n38059 ;
  assign n38061 = ( ~n37907 & n37991 ) | ( ~n37907 & n38060 ) | ( n37991 & n38060 ) ;
  assign n38062 = ~n37907 & n38061 ;
  assign n38063 = x240 ^ x230 ^ 1'b0 ;
  assign n38064 = ( x240 & n38062 ) | ( x240 & n38063 ) | ( n38062 & n38063 ) ;
  assign n38065 = x213 & n37412 ;
  assign n38073 = n7318 | n37377 ;
  assign n38074 = x219 & ~n37297 ;
  assign n38075 = n7318 | n38074 ;
  assign n38076 = n37893 & n38075 ;
  assign n38077 = n38073 & n38076 ;
  assign n38066 = n9344 & ~n37384 ;
  assign n38067 = n37298 & n37323 ;
  assign n38068 = n9344 | n37376 ;
  assign n38069 = n38067 | n38068 ;
  assign n38070 = n38069 ^ n38066 ^ 1'b0 ;
  assign n38071 = ( n38066 & n38069 ) | ( n38066 & n38070 ) | ( n38069 & n38070 ) ;
  assign n38072 = ( x219 & ~n38066 ) | ( x219 & n38071 ) | ( ~n38066 & n38071 ) ;
  assign n38078 = n38077 ^ n38072 ^ 1'b0 ;
  assign n38079 = ( x1152 & ~n38072 ) | ( x1152 & n38077 ) | ( ~n38072 & n38077 ) ;
  assign n38080 = ( x1152 & ~n38078 ) | ( x1152 & n38079 ) | ( ~n38078 & n38079 ) ;
  assign n38081 = ~x212 & n37321 ;
  assign n38082 = n37319 & n38081 ;
  assign n38083 = ~n37309 & n38082 ;
  assign n38084 = x219 | n38083 ;
  assign n38085 = x212 & n37321 ;
  assign n38086 = x211 | n37319 ;
  assign n38087 = n38085 & n38086 ;
  assign n38088 = ( n37324 & n37814 ) | ( n37324 & n38087 ) | ( n37814 & n38087 ) ;
  assign n38089 = n38084 | n38088 ;
  assign n38090 = n37297 | n37329 ;
  assign n38091 = x299 | n38090 ;
  assign n38092 = n38089 & n38091 ;
  assign n38093 = ~n38075 & n38092 ;
  assign n38094 = x1152 | n38093 ;
  assign n38095 = ~n38076 & n38090 ;
  assign n38096 = ( ~n38080 & n38094 ) | ( ~n38080 & n38095 ) | ( n38094 & n38095 ) ;
  assign n38097 = ~n38080 & n38096 ;
  assign n38098 = ( x1151 & n37789 ) | ( x1151 & ~n38097 ) | ( n37789 & ~n38097 ) ;
  assign n38099 = n38097 | n38098 ;
  assign n38100 = n7318 | n37313 ;
  assign n38101 = x1152 | n38100 ;
  assign n38102 = x299 | n37433 ;
  assign n38103 = n37303 & n38102 ;
  assign n38104 = x219 | n38103 ;
  assign n38105 = ~n38101 & n38104 ;
  assign n38106 = x1151 & ~n37777 ;
  assign n38107 = n7318 | n37355 ;
  assign n38108 = x1152 & ~n38107 ;
  assign n38109 = n37352 & ~n37362 ;
  assign n38110 = x219 | n38109 ;
  assign n38111 = x212 & n37343 ;
  assign n38112 = n38110 | n38111 ;
  assign n38113 = n38108 & n38112 ;
  assign n38114 = ( n38105 & n38106 ) | ( n38105 & ~n38113 ) | ( n38106 & ~n38113 ) ;
  assign n38115 = ~n38105 & n38114 ;
  assign n38116 = x1150 & ~n38115 ;
  assign n38117 = n38099 & n38116 ;
  assign n38118 = ~x214 & n37311 ;
  assign n38119 = n37301 & ~n38118 ;
  assign n38120 = ( x212 & n37303 ) | ( x212 & n37312 ) | ( n37303 & n37312 ) ;
  assign n38121 = ( x219 & ~n38119 ) | ( x219 & n38120 ) | ( ~n38119 & n38120 ) ;
  assign n38122 = ( x1152 & ~n38100 ) | ( x1152 & n38121 ) | ( ~n38100 & n38121 ) ;
  assign n38123 = ~x1152 & n38122 ;
  assign n38124 = x1151 & ~n37849 ;
  assign n38125 = ~n36271 & n37343 ;
  assign n38126 = ( n37346 & n37352 ) | ( n37346 & n37354 ) | ( n37352 & n37354 ) ;
  assign n38127 = ( n37353 & n38125 ) | ( n37353 & n38126 ) | ( n38125 & n38126 ) ;
  assign n38128 = ( x219 & x1152 ) | ( x219 & n38127 ) | ( x1152 & n38127 ) ;
  assign n38129 = x1152 & n38128 ;
  assign n38130 = ( n7318 & ~n37355 ) | ( n7318 & n38129 ) | ( ~n37355 & n38129 ) ;
  assign n38131 = ~n7318 & n38130 ;
  assign n38132 = ( n38123 & n38124 ) | ( n38123 & ~n38131 ) | ( n38124 & ~n38131 ) ;
  assign n38133 = ~n38123 & n38132 ;
  assign n38134 = ~x1152 & n38095 ;
  assign n38135 = x1152 & ~n38077 ;
  assign n38136 = n37329 | n37376 ;
  assign n38137 = n38135 & n38136 ;
  assign n38138 = x1151 | n37269 ;
  assign n38139 = ( ~n38134 & n38137 ) | ( ~n38134 & n38138 ) | ( n38137 & n38138 ) ;
  assign n38140 = n38134 | n38139 ;
  assign n38141 = ( x1150 & ~n38133 ) | ( x1150 & n38140 ) | ( ~n38133 & n38140 ) ;
  assign n38142 = ~x1150 & n38141 ;
  assign n38143 = ( x1149 & n38117 ) | ( x1149 & n38142 ) | ( n38117 & n38142 ) ;
  assign n38144 = n38142 ^ n38117 ^ 1'b0 ;
  assign n38145 = ( x1149 & n38143 ) | ( x1149 & n38144 ) | ( n38143 & n38144 ) ;
  assign n38146 = n37376 | n38092 ;
  assign n38147 = ~n38073 & n38146 ;
  assign n38148 = n38093 ^ x1152 ^ 1'b0 ;
  assign n38149 = ( n38093 & n38147 ) | ( n38093 & n38148 ) | ( n38147 & n38148 ) ;
  assign n38150 = ( x1151 & n37795 ) | ( x1151 & ~n38149 ) | ( n37795 & ~n38149 ) ;
  assign n38151 = n38149 | n38150 ;
  assign n38152 = n38111 ^ n37363 ^ n37349 ;
  assign n38153 = ( x1152 & n38110 ) | ( x1152 & n38152 ) | ( n38110 & n38152 ) ;
  assign n38154 = n38152 ^ n38110 ^ 1'b0 ;
  assign n38155 = ( x1152 & n38153 ) | ( x1152 & n38154 ) | ( n38153 & n38154 ) ;
  assign n38156 = x1152 | n37660 ;
  assign n38157 = x212 & n37290 ;
  assign n38158 = ( x212 & x214 ) | ( x212 & n38157 ) | ( x214 & n38157 ) ;
  assign n38159 = ~n37854 & n38158 ;
  assign n38160 = ( n37418 & n38102 ) | ( n37418 & n38159 ) | ( n38102 & n38159 ) ;
  assign n38161 = x219 | n38160 ;
  assign n38162 = n38161 ^ n38156 ^ 1'b0 ;
  assign n38163 = ( n38156 & n38161 ) | ( n38156 & n38162 ) | ( n38161 & n38162 ) ;
  assign n38164 = ( n38155 & ~n38156 ) | ( n38155 & n38163 ) | ( ~n38156 & n38163 ) ;
  assign n38165 = n38164 ^ n37736 ^ 1'b0 ;
  assign n38166 = ( n37736 & ~n38075 ) | ( n37736 & n38165 ) | ( ~n38075 & n38165 ) ;
  assign n38167 = ( n38164 & ~n38165 ) | ( n38164 & n38166 ) | ( ~n38165 & n38166 ) ;
  assign n38168 = ( x1151 & n37262 ) | ( x1151 & ~n38167 ) | ( n37262 & ~n38167 ) ;
  assign n38169 = ~n37262 & n38168 ;
  assign n38170 = x1150 & ~n38169 ;
  assign n38171 = n38151 & n38170 ;
  assign n38172 = n7318 & ~n37656 ;
  assign n38173 = x1151 & ~n38172 ;
  assign n38174 = n36026 & n37209 ;
  assign n38175 = n37295 | n38174 ;
  assign n38176 = n38173 & n38175 ;
  assign n38177 = n37297 & ~n37457 ;
  assign n38178 = ( ~x1152 & n38176 ) | ( ~x1152 & n38177 ) | ( n38176 & n38177 ) ;
  assign n38179 = ~x1152 & n38178 ;
  assign n38180 = x1152 & ~n37457 ;
  assign n38181 = n38179 ^ n37376 ^ 1'b0 ;
  assign n38182 = ( ~n37376 & n38180 ) | ( ~n37376 & n38181 ) | ( n38180 & n38181 ) ;
  assign n38183 = ( n37376 & n38179 ) | ( n37376 & n38182 ) | ( n38179 & n38182 ) ;
  assign n38184 = n7318 ^ x1152 ^ 1'b0 ;
  assign n38185 = n37343 & n37656 ;
  assign n38186 = n37346 | n38185 ;
  assign n38187 = ( x1152 & ~n38184 ) | ( x1152 & n38186 ) | ( ~n38184 & n38186 ) ;
  assign n38188 = ( n7318 & n38184 ) | ( n7318 & n38187 ) | ( n38184 & n38187 ) ;
  assign n38189 = n38173 & n38188 ;
  assign n38190 = ( ~x1150 & n38183 ) | ( ~x1150 & n38189 ) | ( n38183 & n38189 ) ;
  assign n38191 = ~x1150 & n38190 ;
  assign n38192 = ( ~x1149 & n38171 ) | ( ~x1149 & n38191 ) | ( n38171 & n38191 ) ;
  assign n38193 = ~x1149 & n38192 ;
  assign n38194 = ( ~x213 & n38145 ) | ( ~x213 & n38193 ) | ( n38145 & n38193 ) ;
  assign n38195 = ~x213 & n38194 ;
  assign n38196 = ( x209 & n38065 ) | ( x209 & ~n38195 ) | ( n38065 & ~n38195 ) ;
  assign n38197 = ~n38065 & n38196 ;
  assign n38198 = x211 | n36185 ;
  assign n38199 = ~n10008 & n36142 ;
  assign n38200 = ( n37389 & ~n38198 ) | ( n37389 & n38199 ) | ( ~n38198 & n38199 ) ;
  assign n38201 = ~n38198 & n38200 ;
  assign n38202 = n37829 | n38201 ;
  assign n38203 = x214 & ~n37830 ;
  assign n38204 = n37708 | n37715 ;
  assign n38205 = ( x212 & n38203 ) | ( x212 & n38204 ) | ( n38203 & n38204 ) ;
  assign n38206 = ~n38203 & n38205 ;
  assign n38207 = n38202 & n38206 ;
  assign n38208 = ( n37709 & n37825 ) | ( n37709 & n38201 ) | ( n37825 & n38201 ) ;
  assign n38209 = x219 | n38208 ;
  assign n38210 = ( ~n37719 & n38207 ) | ( ~n37719 & n38209 ) | ( n38207 & n38209 ) ;
  assign n38211 = ~n37719 & n38210 ;
  assign n38212 = ( x1151 & n37216 ) | ( x1151 & ~n38211 ) | ( n37216 & ~n38211 ) ;
  assign n38213 = ~n37216 & n38212 ;
  assign n38214 = ( ~x299 & n36015 ) | ( ~x299 & n37802 ) | ( n36015 & n37802 ) ;
  assign n38215 = n37197 & n37809 ;
  assign n38216 = ( n37745 & n38214 ) | ( n37745 & n38215 ) | ( n38214 & n38215 ) ;
  assign n38217 = n7318 | n38216 ;
  assign n38218 = ( ~n7318 & n37318 ) | ( ~n7318 & n38217 ) | ( n37318 & n38217 ) ;
  assign n38219 = ( x1152 & ~n38213 ) | ( x1152 & n38218 ) | ( ~n38213 & n38218 ) ;
  assign n38220 = ~x1152 & n38219 ;
  assign n38221 = x214 & ~n38202 ;
  assign n38222 = n37709 & ~n38221 ;
  assign n38223 = x219 | n38222 ;
  assign n38224 = ( n37705 & n38202 ) | ( n37705 & n38221 ) | ( n38202 & n38221 ) ;
  assign n38225 = ( ~n37719 & n38223 ) | ( ~n37719 & n38224 ) | ( n38223 & n38224 ) ;
  assign n38226 = ~n37719 & n38225 ;
  assign n38227 = ( n37266 & n37270 ) | ( n37266 & ~n38226 ) | ( n37270 & ~n38226 ) ;
  assign n38228 = ~n37266 & n38227 ;
  assign n38229 = x299 & ~n37264 ;
  assign n38230 = n37802 & ~n38229 ;
  assign n38231 = ~x214 & n38230 ;
  assign n38232 = n37811 & ~n38231 ;
  assign n38233 = ( n37805 & n37812 ) | ( n37805 & n38230 ) | ( n37812 & n38230 ) ;
  assign n38234 = ~n38232 & n38233 ;
  assign n38235 = x219 | n38234 ;
  assign n38236 = ~n37797 & n38235 ;
  assign n38237 = ( x1151 & n37266 ) | ( x1151 & ~n38236 ) | ( n37266 & ~n38236 ) ;
  assign n38238 = n38236 | n38237 ;
  assign n38239 = ( x1152 & n38228 ) | ( x1152 & n38238 ) | ( n38228 & n38238 ) ;
  assign n38240 = ~n38228 & n38239 ;
  assign n38241 = ( x1150 & n38220 ) | ( x1150 & ~n38240 ) | ( n38220 & ~n38240 ) ;
  assign n38242 = ~n38220 & n38241 ;
  assign n38243 = x1153 & n38174 ;
  assign n38244 = ( ~x1152 & n37318 ) | ( ~x1152 & n38243 ) | ( n37318 & n38243 ) ;
  assign n38245 = ~x1152 & n38244 ;
  assign n38246 = x1151 & ~n37215 ;
  assign n38247 = ( x1151 & ~n36038 ) | ( x1151 & n38246 ) | ( ~n36038 & n38246 ) ;
  assign n38248 = x219 & ~n37324 ;
  assign n38249 = n7318 | n38248 ;
  assign n38250 = n37334 & ~n38249 ;
  assign n38251 = n38247 & ~n38250 ;
  assign n38252 = n38245 & ~n38251 ;
  assign n38253 = n38084 | n38087 ;
  assign n38254 = ~n38249 & n38253 ;
  assign n38255 = ~n37266 & n37270 ;
  assign n38256 = ~n38250 & n38255 ;
  assign n38257 = ~n38254 & n38256 ;
  assign n38258 = x299 & n37261 ;
  assign n38259 = n37265 & n38258 ;
  assign n38260 = n37372 | n38259 ;
  assign n38261 = ( x1152 & n38257 ) | ( x1152 & n38260 ) | ( n38257 & n38260 ) ;
  assign n38262 = ~n38257 & n38261 ;
  assign n38263 = ( x1150 & ~n38252 ) | ( x1150 & n38262 ) | ( ~n38252 & n38262 ) ;
  assign n38264 = n38252 | n38263 ;
  assign n38265 = ( x1149 & ~n38242 ) | ( x1149 & n38264 ) | ( ~n38242 & n38264 ) ;
  assign n38266 = ~x1149 & n38265 ;
  assign n38267 = n9344 & n37732 ;
  assign n38268 = n36069 & ~n38229 ;
  assign n38269 = x299 | n37345 ;
  assign n38270 = n38268 & n38269 ;
  assign n38271 = ( n37730 & ~n38267 ) | ( n37730 & n38270 ) | ( ~n38267 & n38270 ) ;
  assign n38272 = n38267 | n38271 ;
  assign n38273 = ( n7318 & ~n37477 ) | ( n7318 & n38272 ) | ( ~n37477 & n38272 ) ;
  assign n38274 = ~n7318 & n38273 ;
  assign n38275 = ( x1151 & n37266 ) | ( x1151 & ~n38274 ) | ( n37266 & ~n38274 ) ;
  assign n38276 = n38274 | n38275 ;
  assign n38277 = x219 | n37685 ;
  assign n38278 = n37692 | n38277 ;
  assign n38279 = x1153 | n38278 ;
  assign n38280 = x299 & n9272 ;
  assign n38281 = x219 | n38280 ;
  assign n38282 = ~n37893 & n38281 ;
  assign n38283 = n37698 | n38282 ;
  assign n38284 = n38279 & n38283 ;
  assign n38285 = x211 | n38278 ;
  assign n38286 = n37781 & n38285 ;
  assign n38287 = n38255 & ~n38286 ;
  assign n38288 = ~n38284 & n38287 ;
  assign n38289 = x1152 & ~n38288 ;
  assign n38290 = n38276 & n38289 ;
  assign n38291 = n38247 & ~n38284 ;
  assign n38292 = x1151 | n37736 ;
  assign n38293 = ~x1152 & n38292 ;
  assign n38294 = n38245 | n38293 ;
  assign n38295 = ~n38291 & n38294 ;
  assign n38296 = ( x1150 & n38290 ) | ( x1150 & ~n38295 ) | ( n38290 & ~n38295 ) ;
  assign n38297 = ~n38290 & n38296 ;
  assign n38298 = n37664 | n37857 ;
  assign n38299 = ~n36185 & n37665 ;
  assign n38300 = n37284 | n38299 ;
  assign n38301 = ( n37853 & n38298 ) | ( n37853 & n38300 ) | ( n38298 & n38300 ) ;
  assign n38302 = n38298 & n38301 ;
  assign n38303 = x219 | n38302 ;
  assign n38304 = ~n37865 & n38303 ;
  assign n38305 = ( x1151 & n37216 ) | ( x1151 & ~n38304 ) | ( n37216 & ~n38304 ) ;
  assign n38306 = ~n37216 & n38305 ;
  assign n38307 = n37736 & n37753 ;
  assign n38308 = ( ~n7318 & n38174 ) | ( ~n7318 & n38307 ) | ( n38174 & n38307 ) ;
  assign n38309 = ~n38229 & n38308 ;
  assign n38310 = n37318 | n38309 ;
  assign n38311 = ( x1152 & ~n38306 ) | ( x1152 & n38310 ) | ( ~n38306 & n38310 ) ;
  assign n38312 = ~x1152 & n38311 ;
  assign n38313 = n37663 & ~n37852 ;
  assign n38314 = x219 | n37692 ;
  assign n38315 = n37304 | n38314 ;
  assign n38316 = ( ~n37865 & n38313 ) | ( ~n37865 & n38315 ) | ( n38313 & n38315 ) ;
  assign n38317 = ~n37865 & n38316 ;
  assign n38318 = ( n37266 & n37270 ) | ( n37266 & ~n38317 ) | ( n37270 & ~n38317 ) ;
  assign n38319 = ~n37266 & n38318 ;
  assign n38320 = x219 & ~n37754 ;
  assign n38321 = n7318 | n38320 ;
  assign n38322 = n37754 | n37778 ;
  assign n38323 = n36089 | n37265 ;
  assign n38324 = n38322 & n38323 ;
  assign n38325 = ( x219 & ~n38321 ) | ( x219 & n38324 ) | ( ~n38321 & n38324 ) ;
  assign n38326 = ~n38321 & n38325 ;
  assign n38327 = ( x1151 & n37266 ) | ( x1151 & ~n38326 ) | ( n37266 & ~n38326 ) ;
  assign n38328 = n38326 | n38327 ;
  assign n38329 = ( x1152 & n38319 ) | ( x1152 & n38328 ) | ( n38319 & n38328 ) ;
  assign n38330 = ~n38319 & n38329 ;
  assign n38331 = ( x1150 & ~n38312 ) | ( x1150 & n38330 ) | ( ~n38312 & n38330 ) ;
  assign n38332 = n38312 | n38331 ;
  assign n38333 = ( x1149 & n38297 ) | ( x1149 & n38332 ) | ( n38297 & n38332 ) ;
  assign n38334 = ~n38297 & n38333 ;
  assign n38335 = ( x213 & n38266 ) | ( x213 & n38334 ) | ( n38266 & n38334 ) ;
  assign n38336 = n38334 ^ n38266 ^ 1'b0 ;
  assign n38337 = ( x213 & n38335 ) | ( x213 & n38336 ) | ( n38335 & n38336 ) ;
  assign n38338 = ~n37866 & n38124 ;
  assign n38339 = n37897 | n38138 ;
  assign n38340 = ~x1150 & n38339 ;
  assign n38341 = ~n38338 & n38340 ;
  assign n38342 = x1151 | n37791 ;
  assign n38343 = ~n37781 & n38106 ;
  assign n38344 = x1150 & ~n38343 ;
  assign n38345 = n38342 & n38344 ;
  assign n38346 = ( x1149 & n38341 ) | ( x1149 & ~n38345 ) | ( n38341 & ~n38345 ) ;
  assign n38347 = ~n38341 & n38346 ;
  assign n38348 = x1151 | n37795 ;
  assign n38349 = n37819 | n38348 ;
  assign n38350 = x1151 & ~n37262 ;
  assign n38351 = ~n37842 & n38350 ;
  assign n38352 = x1150 & ~n38351 ;
  assign n38353 = n38349 & n38352 ;
  assign n38354 = ~x1150 & x1151 ;
  assign n38355 = n37871 & n38354 ;
  assign n38356 = x1149 | n38355 ;
  assign n38357 = ( ~n38347 & n38353 ) | ( ~n38347 & n38356 ) | ( n38353 & n38356 ) ;
  assign n38358 = ~n38347 & n38357 ;
  assign n38359 = ~x213 & n38358 ;
  assign n38360 = x209 | n38359 ;
  assign n38361 = ( ~n38197 & n38337 ) | ( ~n38197 & n38360 ) | ( n38337 & n38360 ) ;
  assign n38362 = ~n38197 & n38361 ;
  assign n38363 = x241 ^ x230 ^ 1'b0 ;
  assign n38364 = ( x241 & n38362 ) | ( x241 & n38363 ) | ( n38362 & n38363 ) ;
  assign n38397 = n37077 ^ x214 ^ 1'b0 ;
  assign n38398 = ( n37077 & n37634 ) | ( n37077 & ~n38397 ) | ( n37634 & ~n38397 ) ;
  assign n38399 = x212 & n38398 ;
  assign n38400 = ~x212 & n37635 ;
  assign n38401 = ( x219 & ~n38399 ) | ( x219 & n38400 ) | ( ~n38399 & n38400 ) ;
  assign n38402 = n38399 | n38401 ;
  assign n38365 = x199 & x1144 ;
  assign n38366 = x200 | n38365 ;
  assign n38367 = n37912 | n38366 ;
  assign n38368 = x299 | n37908 ;
  assign n38369 = n38367 & ~n38368 ;
  assign n38370 = x207 | n38369 ;
  assign n38371 = x299 | n37165 ;
  assign n38372 = n37163 | n38366 ;
  assign n38373 = ~n38371 & n38372 ;
  assign n38374 = x207 & ~n38373 ;
  assign n38375 = x208 & ~n38374 ;
  assign n38376 = n38370 & n38375 ;
  assign n38383 = n36395 & n38369 ;
  assign n38403 = n38376 | n38383 ;
  assign n38404 = ~n36036 & n38403 ;
  assign n38405 = x219 & ~n38404 ;
  assign n38377 = n36009 & n38369 ;
  assign n38406 = n36341 | n38377 ;
  assign n38407 = n38376 | n38406 ;
  assign n38408 = n36036 & n38407 ;
  assign n38409 = n38405 & ~n38408 ;
  assign n38410 = x214 | n38403 ;
  assign n38411 = ~x212 & n38410 ;
  assign n38412 = n37666 | n38377 ;
  assign n38413 = n38376 | n38412 ;
  assign n38414 = ~x211 & n38413 ;
  assign n38415 = n37100 | n38377 ;
  assign n38416 = n38376 | n38415 ;
  assign n38417 = x211 | n37666 ;
  assign n38418 = ( n38414 & n38416 ) | ( n38414 & n38417 ) | ( n38416 & n38417 ) ;
  assign n38419 = x214 & ~n38418 ;
  assign n38420 = n38411 & ~n38419 ;
  assign n38423 = x211 & n38407 ;
  assign n38421 = ~x211 & n38416 ;
  assign n38422 = x214 & ~n38421 ;
  assign n38424 = n38423 ^ n38422 ^ 1'b0 ;
  assign n38425 = ( x212 & ~n38422 ) | ( x212 & n38423 ) | ( ~n38422 & n38423 ) ;
  assign n38426 = ( x212 & ~n38424 ) | ( x212 & n38425 ) | ( ~n38424 & n38425 ) ;
  assign n38427 = n38418 ^ x214 ^ 1'b0 ;
  assign n38428 = ( x214 & n38418 ) | ( x214 & ~n38427 ) | ( n38418 & ~n38427 ) ;
  assign n38429 = ( n38426 & n38427 ) | ( n38426 & n38428 ) | ( n38427 & n38428 ) ;
  assign n38430 = ( x219 & ~n38420 ) | ( x219 & n38429 ) | ( ~n38420 & n38429 ) ;
  assign n38431 = n38420 | n38430 ;
  assign n38432 = ( n7318 & ~n38409 ) | ( n7318 & n38431 ) | ( ~n38409 & n38431 ) ;
  assign n38433 = ~n7318 & n38432 ;
  assign n38434 = x219 & ~n36054 ;
  assign n38435 = n36038 & ~n38434 ;
  assign n38436 = n38433 ^ n38402 ^ 1'b0 ;
  assign n38437 = ( ~n38402 & n38435 ) | ( ~n38402 & n38436 ) | ( n38435 & n38436 ) ;
  assign n38438 = ( n38402 & n38433 ) | ( n38402 & n38437 ) | ( n38433 & n38437 ) ;
  assign n38439 = x213 & ~n38438 ;
  assign n38378 = ~n36056 & n36369 ;
  assign n38379 = n9344 & ~n36050 ;
  assign n38380 = n38378 | n38379 ;
  assign n38381 = ( x219 & ~n38377 ) | ( x219 & n38380 ) | ( ~n38377 & n38380 ) ;
  assign n38382 = ~x219 & n38381 ;
  assign n38384 = n36035 | n38383 ;
  assign n38385 = n36036 & ~n36047 ;
  assign n38386 = ~n38377 & n38385 ;
  assign n38387 = x211 & ~n38383 ;
  assign n38388 = ( x219 & n38386 ) | ( x219 & n38387 ) | ( n38386 & n38387 ) ;
  assign n38389 = n38387 ^ n38386 ^ 1'b0 ;
  assign n38390 = ( x219 & n38388 ) | ( x219 & n38389 ) | ( n38388 & n38389 ) ;
  assign n38391 = ( n38382 & n38384 ) | ( n38382 & ~n38390 ) | ( n38384 & ~n38390 ) ;
  assign n38392 = ~n38382 & n38391 ;
  assign n38393 = ( ~n7318 & n38376 ) | ( ~n7318 & n38392 ) | ( n38376 & n38392 ) ;
  assign n38394 = ~n7318 & n38393 ;
  assign n38395 = ( x213 & n36282 ) | ( x213 & ~n38394 ) | ( n36282 & ~n38394 ) ;
  assign n38396 = n38394 | n38395 ;
  assign n38440 = n38439 ^ n38396 ^ 1'b0 ;
  assign n38441 = ( x209 & ~n38396 ) | ( x209 & n38439 ) | ( ~n38396 & n38439 ) ;
  assign n38442 = ( x209 & ~n38440 ) | ( x209 & n38441 ) | ( ~n38440 & n38441 ) ;
  assign n38443 = ( x219 & ~n36035 ) | ( x219 & n38434 ) | ( ~n36035 & n38434 ) ;
  assign n38444 = x299 & ~n38402 ;
  assign n38445 = ( x299 & n38443 ) | ( x299 & n38444 ) | ( n38443 & n38444 ) ;
  assign n38446 = ( n7318 & n36039 ) | ( n7318 & ~n38445 ) | ( n36039 & ~n38445 ) ;
  assign n38447 = ~n7318 & n38446 ;
  assign n38448 = n38447 ^ n38402 ^ 1'b0 ;
  assign n38449 = ( ~n38402 & n38435 ) | ( ~n38402 & n38448 ) | ( n38435 & n38448 ) ;
  assign n38450 = ( n38402 & n38447 ) | ( n38402 & n38449 ) | ( n38447 & n38449 ) ;
  assign n38451 = ( x213 & ~n36501 ) | ( x213 & n38450 ) | ( ~n36501 & n38450 ) ;
  assign n38452 = ( x209 & n36501 ) | ( x209 & n38451 ) | ( n36501 & n38451 ) ;
  assign n38453 = ~x213 & n36078 ;
  assign n38454 = ( ~n38442 & n38452 ) | ( ~n38442 & n38453 ) | ( n38452 & n38453 ) ;
  assign n38455 = ~n38442 & n38454 ;
  assign n38456 = x242 ^ x230 ^ 1'b0 ;
  assign n38457 = ( x242 & n38455 ) | ( x242 & n38456 ) | ( n38455 & n38456 ) ;
  assign n38458 = x253 & x254 ;
  assign n38459 = x267 & n38458 ;
  assign n38460 = ~x263 & n38459 ;
  assign n38461 = x83 | x85 ;
  assign n38462 = x314 & n38461 ;
  assign n38463 = x802 & n38462 ;
  assign n38464 = x276 & n38463 ;
  assign n38465 = ~x1091 & n38464 ;
  assign n38470 = x243 & ~x1091 ;
  assign n38471 = n35970 & ~n38470 ;
  assign n38472 = ~n38465 & n38471 ;
  assign n38466 = x271 & n38465 ;
  assign n38473 = x273 & n38466 ;
  assign n38474 = x243 & n38473 ;
  assign n38475 = n38472 | n38474 ;
  assign n38467 = ( x273 & x1091 ) | ( x273 & n38466 ) | ( x1091 & n38466 ) ;
  assign n38468 = x1091 | n38467 ;
  assign n38469 = x243 | n38468 ;
  assign n38476 = n38475 ^ n38469 ^ 1'b0 ;
  assign n38477 = ( x219 & ~n38469 ) | ( x219 & n38475 ) | ( ~n38469 & n38475 ) ;
  assign n38478 = ( x219 & ~n38476 ) | ( x219 & n38477 ) | ( ~n38476 & n38477 ) ;
  assign n38479 = ( x81 & x314 ) | ( x81 & n38462 ) | ( x314 & n38462 ) ;
  assign n38480 = x802 & n38479 ;
  assign n38481 = x276 & n38480 ;
  assign n38482 = ~x1091 & n38481 ;
  assign n38483 = x271 & n38482 ;
  assign n38484 = x273 & n38483 ;
  assign n38485 = ~x243 & n38484 ;
  assign n38486 = n35963 | n35969 ;
  assign n38487 = x1091 & ~n38486 ;
  assign n38488 = ( x219 & ~n38485 ) | ( x219 & n38487 ) | ( ~n38485 & n38487 ) ;
  assign n38489 = n38485 | n38488 ;
  assign n38490 = n38467 | n38484 ;
  assign n38491 = ~n38489 & n38490 ;
  assign n38492 = ( n38470 & n38489 ) | ( n38470 & ~n38491 ) | ( n38489 & ~n38491 ) ;
  assign n38493 = n38460 & ~n38492 ;
  assign n38494 = ( n38460 & n38478 ) | ( n38460 & n38493 ) | ( n38478 & n38493 ) ;
  assign n38495 = ~x219 & n38486 ;
  assign n38496 = ~x211 & x219 ;
  assign n38497 = x1157 & n38496 ;
  assign n38498 = n38495 | n38497 ;
  assign n38499 = x243 | x1091 ;
  assign n38500 = ( n38470 & ~n38498 ) | ( n38470 & n38499 ) | ( ~n38498 & n38499 ) ;
  assign n38501 = n38460 | n38500 ;
  assign n38502 = ( n7318 & n38494 ) | ( n7318 & n38501 ) | ( n38494 & n38501 ) ;
  assign n38503 = ~n38494 & n38502 ;
  assign n38504 = x272 & x283 ;
  assign n38505 = x275 & n38504 ;
  assign n38506 = x268 & n38505 ;
  assign n38507 = x1091 | n38490 ;
  assign n38508 = ~x199 & n38507 ;
  assign n38509 = ( n38468 & n38507 ) | ( n38468 & n38508 ) | ( n38507 & n38508 ) ;
  assign n38510 = n38482 & n38509 ;
  assign n38511 = x299 | n38510 ;
  assign n38512 = n38508 | n38511 ;
  assign n38513 = x299 & ~n38473 ;
  assign n38514 = ~x200 & n38468 ;
  assign n38515 = n38511 | n38514 ;
  assign n38516 = ~n38513 & n38515 ;
  assign n38517 = x243 & n38516 ;
  assign n38518 = n38512 & n38517 ;
  assign n38519 = x199 & n38468 ;
  assign n38520 = x200 | n38482 ;
  assign n38521 = n38509 & n38520 ;
  assign n38522 = x299 | n38521 ;
  assign n38523 = n38519 | n38522 ;
  assign n38524 = x299 & ~n38468 ;
  assign n38525 = n38523 & ~n38524 ;
  assign n38526 = x243 | n38525 ;
  assign n38527 = ( x1155 & n38518 ) | ( x1155 & n38526 ) | ( n38518 & n38526 ) ;
  assign n38528 = ~n38518 & n38527 ;
  assign n38529 = n38511 & ~n38513 ;
  assign n38530 = n38499 | n38529 ;
  assign n38531 = ~x1155 & n38530 ;
  assign n38532 = x243 & n38529 ;
  assign n38533 = n38531 & ~n38532 ;
  assign n38534 = x1156 | n38533 ;
  assign n38535 = ( ~x1157 & n38528 ) | ( ~x1157 & n38534 ) | ( n38528 & n38534 ) ;
  assign n38536 = ~x1157 & n38535 ;
  assign n38537 = n38508 | n38522 ;
  assign n38538 = ~n38524 & n38537 ;
  assign n38539 = x243 | n38538 ;
  assign n38540 = n38511 | n38519 ;
  assign n38541 = n38516 & n38540 ;
  assign n38542 = x243 & n38541 ;
  assign n38543 = n38539 & ~n38542 ;
  assign n38544 = ~n38484 & n38524 ;
  assign n38545 = n38522 & ~n38544 ;
  assign n38546 = x243 | n38545 ;
  assign n38547 = ~n38517 & n38546 ;
  assign n38548 = x1155 & ~n38547 ;
  assign n38549 = ( x1156 & n38543 ) | ( x1156 & ~n38548 ) | ( n38543 & ~n38548 ) ;
  assign n38550 = n38549 ^ n38543 ^ 1'b0 ;
  assign n38551 = ( x1156 & n38549 ) | ( x1156 & ~n38550 ) | ( n38549 & ~n38550 ) ;
  assign n38552 = x211 & x1157 ;
  assign n38553 = n38514 | n38540 ;
  assign n38554 = ~n38524 & n38553 ;
  assign n38555 = ~x243 & n38554 ;
  assign n38556 = n38508 | n38515 ;
  assign n38557 = ~n38513 & n38556 ;
  assign n38558 = n38523 & n38557 ;
  assign n38559 = x243 & ~n38558 ;
  assign n38560 = n38555 | n38559 ;
  assign n38561 = ~x1155 & n38539 ;
  assign n38562 = x1155 & n38546 ;
  assign n38563 = x243 & n38557 ;
  assign n38564 = n38562 & ~n38563 ;
  assign n38565 = n38561 | n38564 ;
  assign n38566 = x1156 & ~n38565 ;
  assign n38567 = ( x1156 & ~n38560 ) | ( x1156 & n38566 ) | ( ~n38560 & n38566 ) ;
  assign n38568 = n38552 & ~n38567 ;
  assign n38569 = n38551 & n38568 ;
  assign n38577 = n38512 & ~n38513 ;
  assign n38578 = x1155 & n38577 ;
  assign n38579 = n38522 & n38577 ;
  assign n38580 = n38578 | n38579 ;
  assign n38581 = x243 & n38580 ;
  assign n38570 = x299 & ~n38484 ;
  assign n38571 = n38515 & ~n38570 ;
  assign n38572 = ~x1155 & n38571 ;
  assign n38573 = ~n38482 & n38572 ;
  assign n38574 = ~n38524 & n38540 ;
  assign n38575 = x243 | n38574 ;
  assign n38576 = n38573 | n38575 ;
  assign n38582 = n38581 ^ n38576 ^ 1'b0 ;
  assign n38583 = ( x1156 & ~n38576 ) | ( x1156 & n38581 ) | ( ~n38576 & n38581 ) ;
  assign n38584 = ( x1156 & ~n38582 ) | ( x1156 & n38583 ) | ( ~n38582 & n38583 ) ;
  assign n38585 = ~n38569 & n38584 ;
  assign n38586 = ( n38536 & n38569 ) | ( n38536 & ~n38585 ) | ( n38569 & ~n38585 ) ;
  assign n38587 = ~n38513 & n38522 ;
  assign n38588 = ~x243 & x1155 ;
  assign n38589 = n38587 & n38588 ;
  assign n38590 = x1156 | n38589 ;
  assign n38591 = n38515 & ~n38524 ;
  assign n38592 = x243 & ~n38591 ;
  assign n38593 = x243 & n38540 ;
  assign n38594 = x1155 | n38593 ;
  assign n38595 = ~n38513 & n38537 ;
  assign n38596 = ( x243 & ~n38594 ) | ( x243 & n38595 ) | ( ~n38594 & n38595 ) ;
  assign n38597 = ~n38594 & n38596 ;
  assign n38598 = ( ~n38590 & n38592 ) | ( ~n38590 & n38597 ) | ( n38592 & n38597 ) ;
  assign n38599 = n38590 | n38598 ;
  assign n38605 = ~n38558 & n38592 ;
  assign n38606 = x1155 & ~n38605 ;
  assign n38607 = n38555 & n38587 ;
  assign n38608 = n38606 & ~n38607 ;
  assign n38600 = n38553 & ~n38570 ;
  assign n38601 = n38470 | n38600 ;
  assign n38602 = n38539 & n38601 ;
  assign n38603 = n38560 & n38602 ;
  assign n38604 = x1155 | n38603 ;
  assign n38609 = n38608 ^ n38604 ^ 1'b0 ;
  assign n38610 = ( x1156 & ~n38604 ) | ( x1156 & n38608 ) | ( ~n38604 & n38608 ) ;
  assign n38611 = ( x1156 & ~n38609 ) | ( x1156 & n38610 ) | ( ~n38609 & n38610 ) ;
  assign n38612 = n35970 & ~n38611 ;
  assign n38613 = n38599 & n38612 ;
  assign n38614 = ( x219 & n38586 ) | ( x219 & n38613 ) | ( n38586 & n38613 ) ;
  assign n38615 = n38613 ^ n38586 ^ 1'b0 ;
  assign n38616 = ( x219 & n38614 ) | ( x219 & n38615 ) | ( n38614 & n38615 ) ;
  assign n38617 = n38511 & ~n38570 ;
  assign n38618 = x243 & n38617 ;
  assign n38619 = ~x1155 & n38617 ;
  assign n38620 = n38531 | n38619 ;
  assign n38621 = n38620 ^ n38618 ^ 1'b0 ;
  assign n38622 = ( n38618 & n38620 ) | ( n38618 & n38621 ) | ( n38620 & n38621 ) ;
  assign n38623 = ( x1156 & ~n38618 ) | ( x1156 & n38622 ) | ( ~n38618 & n38622 ) ;
  assign n38624 = x243 & n38571 ;
  assign n38625 = n38562 & ~n38624 ;
  assign n38626 = x1155 & ~n38470 ;
  assign n38627 = n38519 & n38626 ;
  assign n38628 = n38625 | n38627 ;
  assign n38629 = n38623 | n38628 ;
  assign n38630 = n38512 & ~n38544 ;
  assign n38631 = n38540 & ~n38570 ;
  assign n38632 = n38631 ^ x243 ^ 1'b0 ;
  assign n38633 = ( ~n38630 & n38631 ) | ( ~n38630 & n38632 ) | ( n38631 & n38632 ) ;
  assign n38634 = x1156 & ~n38573 ;
  assign n38635 = ~n38633 & n38634 ;
  assign n38636 = ( x1157 & n38629 ) | ( x1157 & ~n38635 ) | ( n38629 & ~n38635 ) ;
  assign n38637 = ~x1157 & n38636 ;
  assign n38638 = n38540 & n38624 ;
  assign n38639 = n38561 | n38619 ;
  assign n38640 = n38639 ^ n38638 ^ 1'b0 ;
  assign n38641 = ( n38638 & n38639 ) | ( n38638 & n38640 ) | ( n38639 & n38640 ) ;
  assign n38642 = ( x1156 & ~n38638 ) | ( x1156 & n38641 ) | ( ~n38638 & n38641 ) ;
  assign n38643 = n38625 | n38642 ;
  assign n38644 = n38522 & ~n38570 ;
  assign n38645 = ~x243 & n38644 ;
  assign n38646 = n38553 & n38645 ;
  assign n38647 = ~n38544 & n38556 ;
  assign n38648 = x1155 & n38647 ;
  assign n38649 = ( n38606 & ~n38646 ) | ( n38606 & n38648 ) | ( ~n38646 & n38648 ) ;
  assign n38650 = ~n38646 & n38649 ;
  assign n38651 = n38523 & ~n38570 ;
  assign n38652 = x243 & n38556 ;
  assign n38653 = n38651 & n38652 ;
  assign n38654 = n38537 & n38553 ;
  assign n38655 = ~n38544 & n38654 ;
  assign n38656 = ( x243 & ~n38653 ) | ( x243 & n38655 ) | ( ~n38653 & n38655 ) ;
  assign n38657 = ~n38653 & n38656 ;
  assign n38658 = ( x1155 & ~n38650 ) | ( x1155 & n38657 ) | ( ~n38650 & n38657 ) ;
  assign n38659 = ~n38650 & n38658 ;
  assign n38660 = n38601 & n38659 ;
  assign n38661 = x1156 & ~n38660 ;
  assign n38662 = x1157 & ~n38661 ;
  assign n38663 = n38643 & n38662 ;
  assign n38664 = ( x211 & n38637 ) | ( x211 & ~n38663 ) | ( n38637 & ~n38663 ) ;
  assign n38665 = ~n38637 & n38664 ;
  assign n38666 = n38515 & ~n38544 ;
  assign n38667 = n38644 ^ x243 ^ 1'b0 ;
  assign n38668 = ( n38644 & ~n38666 ) | ( n38644 & n38667 ) | ( ~n38666 & n38667 ) ;
  assign n38669 = n38633 | n38668 ;
  assign n38670 = x1155 & n38669 ;
  assign n38671 = n38623 | n38670 ;
  assign n38672 = ~x1155 & n38666 ;
  assign n38673 = ~n38644 & n38672 ;
  assign n38674 = n38635 & ~n38673 ;
  assign n38675 = ( x1157 & n38671 ) | ( x1157 & ~n38674 ) | ( n38671 & ~n38674 ) ;
  assign n38676 = ~x1157 & n38675 ;
  assign n38677 = x1156 & ~n38659 ;
  assign n38678 = n38642 | n38668 ;
  assign n38679 = ( x1157 & n38677 ) | ( x1157 & n38678 ) | ( n38677 & n38678 ) ;
  assign n38680 = ~n38677 & n38679 ;
  assign n38681 = ( x211 & ~n38676 ) | ( x211 & n38680 ) | ( ~n38676 & n38680 ) ;
  assign n38682 = n38676 | n38681 ;
  assign n38683 = ( x219 & ~n38665 ) | ( x219 & n38682 ) | ( ~n38665 & n38682 ) ;
  assign n38684 = ~x219 & n38683 ;
  assign n38685 = ( n38460 & n38616 ) | ( n38460 & ~n38684 ) | ( n38616 & ~n38684 ) ;
  assign n38686 = ~n38616 & n38685 ;
  assign n38713 = x299 & x1091 ;
  assign n38714 = ~x299 & x1091 ;
  assign n38715 = x200 & ~x1156 ;
  assign n38716 = n38714 & n38715 ;
  assign n38717 = x199 & x1091 ;
  assign n38718 = ~x299 & n38717 ;
  assign n38719 = n38626 & ~n38718 ;
  assign n38720 = x1091 & ~n10074 ;
  assign n38721 = ( n38470 & ~n38719 ) | ( n38470 & n38720 ) | ( ~n38719 & n38720 ) ;
  assign n38722 = n38716 | n38721 ;
  assign n38723 = ~x1157 & n38722 ;
  assign n38724 = ( ~x1157 & n38713 ) | ( ~x1157 & n38723 ) | ( n38713 & n38723 ) ;
  assign n38687 = ~x299 & n36164 ;
  assign n38688 = x1091 & ~n38687 ;
  assign n38689 = n38688 ^ n38499 ^ x1091 ;
  assign n38690 = ( n38470 & n38499 ) | ( n38470 & ~n38626 ) | ( n38499 & ~n38626 ) ;
  assign n38691 = ( n36106 & n38689 ) | ( n36106 & n38690 ) | ( n38689 & n38690 ) ;
  assign n38692 = x1156 | n38691 ;
  assign n38694 = x1091 & n36216 ;
  assign n38695 = n38690 | n38694 ;
  assign n38693 = x1091 & ~n36089 ;
  assign n38696 = n38695 ^ n38693 ^ x1091 ;
  assign n38697 = x1156 & ~n38696 ;
  assign n38698 = n38552 & ~n38697 ;
  assign n38699 = x219 & ~n38698 ;
  assign n38700 = ( x219 & ~n38692 ) | ( x219 & n38699 ) | ( ~n38692 & n38699 ) ;
  assign n38701 = x200 & x1091 ;
  assign n38702 = ~x299 & n38701 ;
  assign n38703 = n38626 & ~n38702 ;
  assign n38704 = x1155 | n38470 ;
  assign n38705 = x1091 & ~n36165 ;
  assign n38706 = n38704 | n38705 ;
  assign n38707 = ~n38703 & n38706 ;
  assign n38708 = x1156 | n38707 ;
  assign n38709 = n36965 & n38694 ;
  assign n38710 = n38697 | n38709 ;
  assign n38711 = n35970 & ~n38710 ;
  assign n38712 = n38708 & n38711 ;
  assign n38725 = ( n38700 & ~n38712 ) | ( n38700 & n38724 ) | ( ~n38712 & n38724 ) ;
  assign n38726 = ~n38724 & n38725 ;
  assign n38733 = n38692 & ~n38710 ;
  assign n38734 = x1157 & ~n38733 ;
  assign n38727 = ~x1156 & n38695 ;
  assign n38728 = x1156 & ~n38719 ;
  assign n38729 = ~n10073 & n38714 ;
  assign n38730 = ( n38470 & n38728 ) | ( n38470 & n38729 ) | ( n38728 & n38729 ) ;
  assign n38731 = ( x1157 & ~n38727 ) | ( x1157 & n38730 ) | ( ~n38727 & n38730 ) ;
  assign n38732 = n38727 | n38731 ;
  assign n38735 = n38734 ^ n38732 ^ 1'b0 ;
  assign n38736 = ( x211 & ~n38732 ) | ( x211 & n38734 ) | ( ~n38732 & n38734 ) ;
  assign n38737 = ( x211 & ~n38735 ) | ( x211 & n38736 ) | ( ~n38735 & n38736 ) ;
  assign n38738 = x211 | n38723 ;
  assign n38739 = x1155 | n38689 ;
  assign n38740 = x1156 | n38703 ;
  assign n38741 = n38739 & ~n38740 ;
  assign n38742 = n38696 & n38728 ;
  assign n38743 = ( x1157 & n38741 ) | ( x1157 & n38742 ) | ( n38741 & n38742 ) ;
  assign n38744 = n38742 ^ n38741 ^ 1'b0 ;
  assign n38745 = ( x1157 & n38743 ) | ( x1157 & n38744 ) | ( n38743 & n38744 ) ;
  assign n38746 = ( ~n38737 & n38738 ) | ( ~n38737 & n38745 ) | ( n38738 & n38745 ) ;
  assign n38747 = ~n38737 & n38746 ;
  assign n38748 = ( x219 & ~n38726 ) | ( x219 & n38747 ) | ( ~n38726 & n38747 ) ;
  assign n38749 = ~n38726 & n38748 ;
  assign n38750 = n38460 | n38749 ;
  assign n38751 = ( n7318 & ~n38686 ) | ( n7318 & n38750 ) | ( ~n38686 & n38750 ) ;
  assign n38752 = ~n7318 & n38751 ;
  assign n38753 = ( n38503 & n38506 ) | ( n38503 & ~n38752 ) | ( n38506 & ~n38752 ) ;
  assign n38754 = ~n38503 & n38753 ;
  assign n38755 = n7318 & n38500 ;
  assign n38756 = ~n7318 & n38749 ;
  assign n38757 = ( n38506 & ~n38755 ) | ( n38506 & n38756 ) | ( ~n38755 & n38756 ) ;
  assign n38758 = n38755 | n38757 ;
  assign n38759 = ( x230 & ~n38754 ) | ( x230 & n38758 ) | ( ~n38754 & n38758 ) ;
  assign n38760 = ~x230 & n38759 ;
  assign n38761 = x199 & ~n37084 ;
  assign n38762 = x1155 | n9353 ;
  assign n38763 = ~n38715 & n38762 ;
  assign n38764 = ( n15098 & ~n38761 ) | ( n15098 & n38763 ) | ( ~n38761 & n38763 ) ;
  assign n38765 = ~n15098 & n38764 ;
  assign n38766 = ~n38760 & n38765 ;
  assign n38767 = x230 & ~n15098 ;
  assign n38768 = ( x230 & ~n38498 ) | ( x230 & n38767 ) | ( ~n38498 & n38767 ) ;
  assign n38769 = ( n38760 & ~n38766 ) | ( n38760 & n38768 ) | ( ~n38766 & n38768 ) ;
  assign n38770 = x213 & ~n37989 ;
  assign n38771 = x213 | n37082 ;
  assign n38772 = n36049 | n37974 ;
  assign n38773 = n37969 & ~n38772 ;
  assign n38774 = ( n37969 & ~n37978 ) | ( n37969 & n38773 ) | ( ~n37978 & n38773 ) ;
  assign n38775 = ~n37102 & n37945 ;
  assign n38776 = ~n36344 & n37931 ;
  assign n38777 = n38775 | n38776 ;
  assign n38778 = n37994 & n38777 ;
  assign n38779 = x214 & ~n38778 ;
  assign n38780 = n37954 & ~n38779 ;
  assign n38781 = ~n36055 & n37688 ;
  assign n38782 = x214 | n38777 ;
  assign n38783 = ( x212 & n38781 ) | ( x212 & n38782 ) | ( n38781 & n38782 ) ;
  assign n38784 = ~n38781 & n38783 ;
  assign n38785 = n37994 & n38784 ;
  assign n38786 = ( x219 & ~n38780 ) | ( x219 & n38785 ) | ( ~n38780 & n38785 ) ;
  assign n38787 = n38780 | n38786 ;
  assign n38788 = ( n38032 & ~n38774 ) | ( n38032 & n38787 ) | ( ~n38774 & n38787 ) ;
  assign n38789 = ~n38032 & n38788 ;
  assign n38790 = x299 & n37073 ;
  assign n38791 = x1147 & ~n38790 ;
  assign n38792 = x214 & ~n38777 ;
  assign n38793 = n37948 & ~n38792 ;
  assign n38794 = n37930 & n38784 ;
  assign n38795 = ( x219 & ~n38793 ) | ( x219 & n38794 ) | ( ~n38793 & n38794 ) ;
  assign n38796 = n38793 | n38795 ;
  assign n38797 = ( n37992 & n38791 ) | ( n37992 & n38796 ) | ( n38791 & n38796 ) ;
  assign n38798 = ~n37992 & n38797 ;
  assign n38799 = ( ~n38771 & n38789 ) | ( ~n38771 & n38798 ) | ( n38789 & n38798 ) ;
  assign n38800 = n38771 | n38799 ;
  assign n38801 = x209 & ~n38800 ;
  assign n38802 = ( x209 & n38770 ) | ( x209 & n38801 ) | ( n38770 & n38801 ) ;
  assign n38803 = n37645 | n37652 ;
  assign n38804 = ~n37659 & n38803 ;
  assign n38805 = n9344 & ~n37673 ;
  assign n38806 = n37645 | n37651 ;
  assign n38807 = n9344 | n37937 ;
  assign n38808 = n36297 & n38807 ;
  assign n38809 = ( n38805 & n38806 ) | ( n38805 & n38808 ) | ( n38806 & n38808 ) ;
  assign n38810 = ~n38805 & n38809 ;
  assign n38811 = n37172 | n37750 ;
  assign n38812 = ( ~n7318 & n38810 ) | ( ~n7318 & n38811 ) | ( n38810 & n38811 ) ;
  assign n38813 = ~n7318 & n38812 ;
  assign n38814 = ( x213 & n38804 ) | ( x213 & n38813 ) | ( n38804 & n38813 ) ;
  assign n38815 = n38813 ^ n38804 ^ 1'b0 ;
  assign n38816 = ( x213 & n38814 ) | ( x213 & n38815 ) | ( n38814 & n38815 ) ;
  assign n38817 = ~x213 & n37184 ;
  assign n38818 = x209 | n38817 ;
  assign n38819 = ( ~n38802 & n38816 ) | ( ~n38802 & n38818 ) | ( n38816 & n38818 ) ;
  assign n38820 = ~n38802 & n38819 ;
  assign n38821 = x244 ^ x230 ^ 1'b0 ;
  assign n38822 = ( x244 & n38820 ) | ( x244 & n38821 ) | ( n38820 & n38821 ) ;
  assign n38823 = x207 & ~n37922 ;
  assign n38824 = n36395 | n38823 ;
  assign n38825 = n36112 | n37921 ;
  assign n38826 = ~n9233 & n38825 ;
  assign n38827 = n38824 & ~n38826 ;
  assign n38828 = ~n36036 & n38827 ;
  assign n38829 = x219 & ~n38828 ;
  assign n38830 = n36009 & ~n38825 ;
  assign n38831 = x208 & ~n37922 ;
  assign n38832 = ~n36112 & n37919 ;
  assign n38833 = ~x207 & n38832 ;
  assign n38834 = ( n37666 & n38823 ) | ( n37666 & ~n38833 ) | ( n38823 & ~n38833 ) ;
  assign n38835 = n38833 | n38834 ;
  assign n38836 = x208 & n38835 ;
  assign n38837 = ~x299 & n38836 ;
  assign n38838 = ( ~n38830 & n38831 ) | ( ~n38830 & n38837 ) | ( n38831 & n38837 ) ;
  assign n38839 = n38830 | n38838 ;
  assign n38840 = n37666 | n38839 ;
  assign n38841 = n36036 & n38840 ;
  assign n38842 = n38829 & ~n38841 ;
  assign n38843 = n7318 | n38842 ;
  assign n38844 = x214 | n38827 ;
  assign n38845 = ~x212 & n38844 ;
  assign n38846 = x299 | n38839 ;
  assign n38847 = n38845 & n38846 ;
  assign n38848 = x219 | n38847 ;
  assign n38849 = x212 & n38846 ;
  assign n38850 = n9271 & ~n38840 ;
  assign n38851 = n38849 & ~n38850 ;
  assign n38852 = ( ~n38843 & n38848 ) | ( ~n38843 & n38851 ) | ( n38848 & n38851 ) ;
  assign n38853 = ~n38843 & n38852 ;
  assign n38854 = x1147 & ~n37262 ;
  assign n38855 = x1146 & n37269 ;
  assign n38856 = n38854 & ~n38855 ;
  assign n38857 = x1148 & ~n38856 ;
  assign n38858 = ( x1148 & n38853 ) | ( x1148 & n38857 ) | ( n38853 & n38857 ) ;
  assign n38891 = x1147 | n38855 ;
  assign n38892 = n37262 & n37848 ;
  assign n38893 = n38891 | n38892 ;
  assign n38859 = x207 | n38831 ;
  assign n38861 = x207 & n37920 ;
  assign n38862 = x1146 & n36165 ;
  assign n38863 = n38861 | n38862 ;
  assign n38864 = ( x208 & n37666 ) | ( x208 & n38863 ) | ( n37666 & n38863 ) ;
  assign n38860 = n37280 | n37921 ;
  assign n38865 = n38860 & ~n38864 ;
  assign n38866 = ( n38859 & n38864 ) | ( n38859 & ~n38865 ) | ( n38864 & ~n38865 ) ;
  assign n38867 = ~x299 & n38866 ;
  assign n38868 = ~n36036 & n38867 ;
  assign n38869 = x219 & ~n38868 ;
  assign n38870 = n36036 & n38866 ;
  assign n38871 = n38869 & ~n38870 ;
  assign n38872 = n7318 | n38871 ;
  assign n38873 = x214 | n38867 ;
  assign n38874 = ~x212 & n38873 ;
  assign n38875 = x299 | n37920 ;
  assign n38876 = n38866 & n38875 ;
  assign n38877 = x299 | n38876 ;
  assign n38878 = ( n9233 & n37281 ) | ( n9233 & n37920 ) | ( n37281 & n37920 ) ;
  assign n38879 = n38878 ^ x211 ^ 1'b0 ;
  assign n38880 = ( n38877 & n38878 ) | ( n38877 & ~n38879 ) | ( n38878 & ~n38879 ) ;
  assign n38881 = n38867 | n38880 ;
  assign n38882 = n38874 & n38881 ;
  assign n38883 = x219 | n38882 ;
  assign n38884 = x214 | n38881 ;
  assign n38885 = x212 & n38884 ;
  assign n38886 = x214 & ~n37667 ;
  assign n38887 = x212 & ~n38886 ;
  assign n38888 = ( n38867 & n38885 ) | ( n38867 & n38887 ) | ( n38885 & n38887 ) ;
  assign n38889 = ( ~n38872 & n38883 ) | ( ~n38872 & n38888 ) | ( n38883 & n38888 ) ;
  assign n38890 = ~n38872 & n38889 ;
  assign n38894 = n38893 ^ n38890 ^ 1'b0 ;
  assign n38895 = ( n38890 & n38893 ) | ( n38890 & ~n38894 ) | ( n38893 & ~n38894 ) ;
  assign n38896 = ( n38858 & n38894 ) | ( n38858 & n38895 ) | ( n38894 & n38895 ) ;
  assign n38897 = x219 & ~n38878 ;
  assign n38898 = n36621 | n38897 ;
  assign n38899 = ( n36035 & n36036 ) | ( n36035 & n38878 ) | ( n36036 & n38878 ) ;
  assign n38900 = n38876 & n38899 ;
  assign n38901 = n38898 & ~n38900 ;
  assign n38902 = n38280 | n38867 ;
  assign n38903 = x219 | n38902 ;
  assign n38904 = ( x219 & n38863 ) | ( x219 & n38903 ) | ( n38863 & n38903 ) ;
  assign n38905 = ( n7318 & ~n38901 ) | ( n7318 & n38904 ) | ( ~n38901 & n38904 ) ;
  assign n38906 = ~n7318 & n38905 ;
  assign n38907 = ( ~x1148 & n38891 ) | ( ~x1148 & n38906 ) | ( n38891 & n38906 ) ;
  assign n38908 = ~x1148 & n38907 ;
  assign n38909 = ~x208 & n37666 ;
  assign n38910 = n36009 & n38832 ;
  assign n38911 = ( n38836 & ~n38909 ) | ( n38836 & n38910 ) | ( ~n38909 & n38910 ) ;
  assign n38912 = n38909 | n38911 ;
  assign n38913 = n9233 | n38832 ;
  assign n38914 = n38824 & n38913 ;
  assign n38915 = ( n36035 & n36036 ) | ( n36035 & n38914 ) | ( n36036 & n38914 ) ;
  assign n38916 = n38912 & n38915 ;
  assign n38917 = ~x214 & n38914 ;
  assign n38918 = ~x212 & n38917 ;
  assign n38919 = x219 & ~n38918 ;
  assign n38920 = ~n38916 & n38919 ;
  assign n38921 = n7318 | n38920 ;
  assign n38922 = n11549 | n38914 ;
  assign n38923 = ~x214 & n38922 ;
  assign n38924 = x299 | n38912 ;
  assign n38925 = x214 & n38924 ;
  assign n38926 = ~x211 & n38846 ;
  assign n38927 = n38827 | n38926 ;
  assign n38928 = n38925 & n38927 ;
  assign n38929 = x212 & ~n38928 ;
  assign n38930 = ~n38923 & n38929 ;
  assign n38931 = x214 & n38922 ;
  assign n38932 = x212 | n38917 ;
  assign n38933 = n38931 | n38932 ;
  assign n38934 = n38933 ^ n38930 ^ 1'b0 ;
  assign n38935 = ( n38930 & n38933 ) | ( n38930 & n38934 ) | ( n38933 & n38934 ) ;
  assign n38936 = ( x219 & ~n38930 ) | ( x219 & n38935 ) | ( ~n38930 & n38935 ) ;
  assign n38937 = x1146 | n36271 ;
  assign n38938 = n37692 & n38937 ;
  assign n38939 = ( ~n38921 & n38936 ) | ( ~n38921 & n38938 ) | ( n38936 & n38938 ) ;
  assign n38940 = ~n38921 & n38939 ;
  assign n38941 = ( n38001 & n38856 ) | ( n38001 & ~n38940 ) | ( n38856 & ~n38940 ) ;
  assign n38942 = ~n38940 & n38941 ;
  assign n38943 = ( n38896 & n38908 ) | ( n38896 & ~n38942 ) | ( n38908 & ~n38942 ) ;
  assign n38944 = n38943 ^ n38908 ^ 1'b0 ;
  assign n38945 = ( n38896 & n38943 ) | ( n38896 & ~n38944 ) | ( n38943 & ~n38944 ) ;
  assign n38946 = x213 & n38945 ;
  assign n38947 = ~x214 & n38878 ;
  assign n38948 = n37673 | n38867 ;
  assign n38949 = x214 & n38877 ;
  assign n38950 = n38948 & n38949 ;
  assign n38951 = ( ~x212 & n38947 ) | ( ~x212 & n38950 ) | ( n38947 & n38950 ) ;
  assign n38952 = ~x212 & n38951 ;
  assign n38953 = x299 & n38398 ;
  assign n38954 = ( x212 & n38867 ) | ( x212 & n38953 ) | ( n38867 & n38953 ) ;
  assign n38955 = n38875 & n38954 ;
  assign n38956 = ( x219 & ~n38952 ) | ( x219 & n38955 ) | ( ~n38952 & n38955 ) ;
  assign n38957 = n38952 | n38956 ;
  assign n38958 = n36341 | n38839 ;
  assign n38959 = n38924 & n38958 ;
  assign n38960 = ( x211 & n38915 ) | ( x211 & n38959 ) | ( n38915 & n38959 ) ;
  assign n38961 = n38915 & n38960 ;
  assign n38962 = ( x219 & n38918 ) | ( x219 & ~n38961 ) | ( n38918 & ~n38961 ) ;
  assign n38963 = ~n38918 & n38962 ;
  assign n38964 = x1147 & ~n7318 ;
  assign n38965 = ( n38399 & n38839 ) | ( n38399 & n38849 ) | ( n38839 & n38849 ) ;
  assign n38966 = n38924 & n38965 ;
  assign n38967 = n37673 | n38839 ;
  assign n38968 = n38925 & n38967 ;
  assign n38969 = ( ~x212 & n38917 ) | ( ~x212 & n38968 ) | ( n38917 & n38968 ) ;
  assign n38970 = ~x212 & n38969 ;
  assign n38971 = ( x219 & ~n38966 ) | ( x219 & n38970 ) | ( ~n38966 & n38970 ) ;
  assign n38972 = n38966 | n38971 ;
  assign n38973 = ( n38963 & n38964 ) | ( n38963 & n38972 ) | ( n38964 & n38972 ) ;
  assign n38974 = ~n38963 & n38973 ;
  assign n38975 = n38402 & n38435 ;
  assign n38976 = ( x1148 & ~n38974 ) | ( x1148 & n38975 ) | ( ~n38974 & n38975 ) ;
  assign n38977 = n38974 | n38976 ;
  assign n38978 = ~n36344 & n38877 ;
  assign n38979 = x211 | n38978 ;
  assign n38980 = n38898 & ~n38979 ;
  assign n38981 = ( n38898 & ~n38899 ) | ( n38898 & n38980 ) | ( ~n38899 & n38980 ) ;
  assign n38982 = ( x1147 & n7318 ) | ( x1147 & ~n38981 ) | ( n7318 & ~n38981 ) ;
  assign n38983 = n38981 | n38982 ;
  assign n38984 = ~n38977 & n38983 ;
  assign n38985 = ( n38957 & n38977 ) | ( n38957 & ~n38984 ) | ( n38977 & ~n38984 ) ;
  assign n38986 = x299 | n38866 ;
  assign n38987 = n36036 & n38986 ;
  assign n38988 = n38869 & ~n38987 ;
  assign n38989 = ( n36344 & n38869 ) | ( n36344 & n38988 ) | ( n38869 & n38988 ) ;
  assign n38990 = n38032 | n38989 ;
  assign n38991 = n38874 & n38948 ;
  assign n38992 = x219 | n38954 ;
  assign n38993 = ( ~n38990 & n38991 ) | ( ~n38990 & n38992 ) | ( n38991 & n38992 ) ;
  assign n38994 = ~n38990 & n38993 ;
  assign n38995 = x1148 & ~n38975 ;
  assign n38996 = n36036 & n38958 ;
  assign n38997 = n38829 & ~n38996 ;
  assign n38998 = x214 & ~n38967 ;
  assign n38999 = n38845 & ~n38998 ;
  assign n39000 = ( x219 & n38965 ) | ( x219 & ~n38999 ) | ( n38965 & ~n38999 ) ;
  assign n39001 = n38999 | n39000 ;
  assign n39002 = ( n38964 & n38997 ) | ( n38964 & n39001 ) | ( n38997 & n39001 ) ;
  assign n39003 = ~n38997 & n39002 ;
  assign n39004 = ( n38994 & n38995 ) | ( n38994 & ~n39003 ) | ( n38995 & ~n39003 ) ;
  assign n39005 = ~n38994 & n39004 ;
  assign n39006 = ( x213 & n38985 ) | ( x213 & ~n39005 ) | ( n38985 & ~n39005 ) ;
  assign n39007 = ~x213 & n39006 ;
  assign n39008 = ( x209 & n38946 ) | ( x209 & ~n39007 ) | ( n38946 & ~n39007 ) ;
  assign n39009 = ~n38946 & n39008 ;
  assign n39010 = ~x213 & n38438 ;
  assign n39011 = x209 | n39010 ;
  assign n39012 = n36035 & n38414 ;
  assign n39013 = n38405 & ~n39012 ;
  assign n39014 = n7318 | n39013 ;
  assign n39015 = ~x212 & n38403 ;
  assign n39016 = ~x299 & n38418 ;
  assign n39017 = ( x212 & n38887 ) | ( x212 & n39016 ) | ( n38887 & n39016 ) ;
  assign n39018 = n38410 & n39017 ;
  assign n39019 = ( x219 & ~n39015 ) | ( x219 & n39018 ) | ( ~n39015 & n39018 ) ;
  assign n39020 = n39015 | n39019 ;
  assign n39021 = n39014 | n39020 ;
  assign n39022 = ( n38891 & ~n39014 ) | ( n38891 & n39021 ) | ( ~n39014 & n39021 ) ;
  assign n39023 = x299 | n38416 ;
  assign n39024 = ~x211 & n39023 ;
  assign n39025 = ( n38413 & n39023 ) | ( n38413 & n39024 ) | ( n39023 & n39024 ) ;
  assign n39026 = x214 & n39025 ;
  assign n39027 = n11549 | n38403 ;
  assign n39028 = ~x214 & n39027 ;
  assign n39029 = n39026 | n39028 ;
  assign n39030 = x212 & n39029 ;
  assign n39031 = n38411 & n39027 ;
  assign n39032 = x219 | n39031 ;
  assign n39033 = ( ~n39014 & n39030 ) | ( ~n39014 & n39032 ) | ( n39030 & n39032 ) ;
  assign n39034 = ~n39014 & n39033 ;
  assign n39035 = ( n38001 & n38856 ) | ( n38001 & ~n39034 ) | ( n38856 & ~n39034 ) ;
  assign n39036 = ~n39034 & n39035 ;
  assign n39037 = ( x1148 & n39022 ) | ( x1148 & ~n39036 ) | ( n39022 & ~n39036 ) ;
  assign n39038 = ~x1148 & n39037 ;
  assign n39039 = n38403 | n39024 ;
  assign n39040 = n38411 & n39039 ;
  assign n39041 = ( n39017 & n39018 ) | ( n39017 & n39024 ) | ( n39018 & n39024 ) ;
  assign n39042 = ( x219 & ~n39040 ) | ( x219 & n39041 ) | ( ~n39040 & n39041 ) ;
  assign n39043 = n39040 | n39042 ;
  assign n39044 = ( n7318 & ~n39013 ) | ( n7318 & n39043 ) | ( ~n39013 & n39043 ) ;
  assign n39045 = ~n7318 & n39044 ;
  assign n39046 = ( n38891 & n38892 ) | ( n38891 & ~n39045 ) | ( n38892 & ~n39045 ) ;
  assign n39047 = n39045 | n39046 ;
  assign n39048 = ~x214 & n39023 ;
  assign n39049 = n39026 | n39048 ;
  assign n39050 = x212 & n39049 ;
  assign n39051 = n38411 & n39023 ;
  assign n39052 = ( x219 & ~n39050 ) | ( x219 & n39051 ) | ( ~n39050 & n39051 ) ;
  assign n39053 = n39050 | n39052 ;
  assign n39054 = ( n7318 & ~n39013 ) | ( n7318 & n39053 ) | ( ~n39013 & n39053 ) ;
  assign n39055 = ~n7318 & n39054 ;
  assign n39056 = ( n38854 & n38855 ) | ( n38854 & ~n39055 ) | ( n38855 & ~n39055 ) ;
  assign n39057 = ~n38855 & n39056 ;
  assign n39058 = x1148 & ~n39057 ;
  assign n39059 = n39047 & n39058 ;
  assign n39060 = ( x213 & n39038 ) | ( x213 & n39059 ) | ( n39038 & n39059 ) ;
  assign n39061 = n39059 ^ n39038 ^ 1'b0 ;
  assign n39062 = ( x213 & n39060 ) | ( x213 & n39061 ) | ( n39060 & n39061 ) ;
  assign n39063 = ( ~n39009 & n39011 ) | ( ~n39009 & n39062 ) | ( n39011 & n39062 ) ;
  assign n39064 = ~n39009 & n39063 ;
  assign n39065 = x245 ^ x230 ^ 1'b0 ;
  assign n39066 = ( x245 & n39064 ) | ( x245 & n39065 ) | ( n39064 & n39065 ) ;
  assign n39067 = x1150 & ~n37782 ;
  assign n39068 = x1150 | n37791 ;
  assign n39069 = ( x1149 & n39067 ) | ( x1149 & n39068 ) | ( n39067 & n39068 ) ;
  assign n39070 = ~n39067 & n39069 ;
  assign n39071 = x1150 & ~n37867 ;
  assign n39072 = x1150 | n37898 ;
  assign n39073 = ( x1149 & ~n39071 ) | ( x1149 & n39072 ) | ( ~n39071 & n39072 ) ;
  assign n39074 = ~x1149 & n39073 ;
  assign n39075 = ( x1148 & n39070 ) | ( x1148 & ~n39074 ) | ( n39070 & ~n39074 ) ;
  assign n39076 = ~n39070 & n39075 ;
  assign n39077 = x1150 & ~n37843 ;
  assign n39078 = x1149 & ~n39077 ;
  assign n39079 = x1150 | n37820 ;
  assign n39080 = n39078 & n39079 ;
  assign n39081 = n39080 ^ n37871 ^ 1'b0 ;
  assign n39082 = ~x1149 & x1150 ;
  assign n39083 = ( n37871 & ~n39081 ) | ( n37871 & n39082 ) | ( ~n39081 & n39082 ) ;
  assign n39084 = ( n39080 & n39081 ) | ( n39080 & n39083 ) | ( n39081 & n39083 ) ;
  assign n39085 = ( x1148 & ~n39076 ) | ( x1148 & n39084 ) | ( ~n39076 & n39084 ) ;
  assign n39086 = ~n39076 & n39085 ;
  assign n39087 = x213 & n39086 ;
  assign n39088 = ~n38856 & n38893 ;
  assign n39092 = ( n37345 & n37886 ) | ( n37345 & n38887 ) | ( n37886 & n38887 ) ;
  assign n39089 = n37732 & n37888 ;
  assign n39090 = n37880 | n39089 ;
  assign n39091 = n38893 & n39090 ;
  assign n39093 = ( n37890 & n39091 ) | ( n37890 & ~n39092 ) | ( n39091 & ~n39092 ) ;
  assign n39094 = n39092 | n39093 ;
  assign n39095 = n39094 ^ n37736 ^ 1'b0 ;
  assign n39096 = x219 & ~n37666 ;
  assign n39097 = n37646 | n39096 ;
  assign n39098 = ( n37736 & n39095 ) | ( n37736 & ~n39097 ) | ( n39095 & ~n39097 ) ;
  assign n39099 = ( n39094 & ~n39095 ) | ( n39094 & n39098 ) | ( ~n39095 & n39098 ) ;
  assign n39100 = ( ~x1150 & n39088 ) | ( ~x1150 & n39099 ) | ( n39088 & n39099 ) ;
  assign n39101 = ~x1150 & n39100 ;
  assign n39102 = x214 & n37687 ;
  assign n39103 = n37693 & ~n39102 ;
  assign n39104 = ( x219 & n37689 ) | ( x219 & ~n39103 ) | ( n37689 & ~n39103 ) ;
  assign n39105 = n39103 | n39104 ;
  assign n39106 = ( n7318 & ~n37686 ) | ( n7318 & n39105 ) | ( ~n37686 & n39105 ) ;
  assign n39107 = ~n7318 & n39106 ;
  assign n39108 = x1146 & n37779 ;
  assign n39109 = n38856 & ~n39108 ;
  assign n39110 = ~n39107 & n39109 ;
  assign n39111 = x219 | n37632 ;
  assign n39112 = n38281 & n39111 ;
  assign n39113 = ~n39097 & n39112 ;
  assign n39114 = n37698 | n39113 ;
  assign n39115 = n38893 | n39114 ;
  assign n39116 = ( x1150 & n39110 ) | ( x1150 & n39115 ) | ( n39110 & n39115 ) ;
  assign n39117 = ~n39110 & n39116 ;
  assign n39118 = ( x1148 & n39101 ) | ( x1148 & ~n39117 ) | ( n39101 & ~n39117 ) ;
  assign n39119 = ~n39101 & n39118 ;
  assign n39120 = n38001 | n38856 ;
  assign n39121 = n37720 & n39097 ;
  assign n39122 = n37833 | n37834 ;
  assign n39123 = n37704 ^ n37666 ^ x299 ;
  assign n39124 = ( n37833 & n37835 ) | ( n37833 & ~n39123 ) | ( n37835 & ~n39123 ) ;
  assign n39125 = n39123 | n39124 ;
  assign n39126 = ( n39121 & n39122 ) | ( n39121 & n39125 ) | ( n39122 & n39125 ) ;
  assign n39127 = ~n39121 & n39126 ;
  assign n39128 = n39120 & ~n39127 ;
  assign n39129 = x1150 & ~n39128 ;
  assign n39130 = n37709 & ~n37827 ;
  assign n39131 = ( x219 & n38206 ) | ( x219 & ~n39130 ) | ( n38206 & ~n39130 ) ;
  assign n39132 = n39130 | n39131 ;
  assign n39133 = ~n37719 & n39132 ;
  assign n39134 = n37823 | n39127 ;
  assign n39135 = n39133 & n39134 ;
  assign n39136 = n38891 | n39135 ;
  assign n39137 = n39129 & n39136 ;
  assign n39138 = ~n37646 & n37802 ;
  assign n39139 = n37797 & ~n39138 ;
  assign n39140 = n37799 & ~n38081 ;
  assign n39141 = x219 | n39140 ;
  assign n39142 = ~n39139 & n39141 ;
  assign n39143 = x1146 | n37745 ;
  assign n39144 = n39142 & n39143 ;
  assign n39145 = ( ~x1150 & n38891 ) | ( ~x1150 & n39144 ) | ( n38891 & n39144 ) ;
  assign n39146 = ~x1150 & n39145 ;
  assign n39147 = ~x1146 & n37796 ;
  assign n39148 = n37632 & n37688 ;
  assign n39149 = ( n37745 & n37818 ) | ( n37745 & ~n39148 ) | ( n37818 & ~n39148 ) ;
  assign n39150 = n39148 | n39149 ;
  assign n39151 = ( n39139 & ~n39147 ) | ( n39139 & n39150 ) | ( ~n39147 & n39150 ) ;
  assign n39152 = ~n39139 & n39151 ;
  assign n39153 = n39152 ^ n39146 ^ 1'b0 ;
  assign n39154 = ( ~n39120 & n39152 ) | ( ~n39120 & n39153 ) | ( n39152 & n39153 ) ;
  assign n39155 = ( n39146 & ~n39153 ) | ( n39146 & n39154 ) | ( ~n39153 & n39154 ) ;
  assign n39156 = ( x1148 & ~n39137 ) | ( x1148 & n39155 ) | ( ~n39137 & n39155 ) ;
  assign n39157 = n39137 | n39156 ;
  assign n39158 = ( x1149 & n39119 ) | ( x1149 & n39157 ) | ( n39119 & n39157 ) ;
  assign n39159 = ~n39119 & n39158 ;
  assign n39160 = x299 & n37785 ;
  assign n39161 = ( x219 & n38938 ) | ( x219 & ~n39160 ) | ( n38938 & ~n39160 ) ;
  assign n39162 = n39160 | n39161 ;
  assign n39163 = n39162 ^ x1150 ^ 1'b0 ;
  assign n39164 = ( ~x1150 & n37296 ) | ( ~x1150 & n39163 ) | ( n37296 & n39163 ) ;
  assign n39165 = ( x1150 & n39162 ) | ( x1150 & n39164 ) | ( n39162 & n39164 ) ;
  assign n39166 = ( x1148 & n39120 ) | ( x1148 & ~n39165 ) | ( n39120 & ~n39165 ) ;
  assign n39167 = n39166 ^ n39120 ^ 1'b0 ;
  assign n39168 = ( x1148 & n39166 ) | ( x1148 & ~n39167 ) | ( n39166 & ~n39167 ) ;
  assign n39169 = n38891 | n39113 ;
  assign n39170 = n39097 & n39120 ;
  assign n39171 = n39169 & ~n39170 ;
  assign n39172 = x1150 & n37631 ;
  assign n39173 = ( ~n39168 & n39171 ) | ( ~n39168 & n39172 ) | ( n39171 & n39172 ) ;
  assign n39174 = ~n39168 & n39173 ;
  assign n39175 = n37661 & n39097 ;
  assign n39176 = x214 & ~n37850 ;
  assign n39177 = ~n37669 & n39176 ;
  assign n39178 = x214 | n37292 ;
  assign n39179 = ( x212 & n39177 ) | ( x212 & n39178 ) | ( n39177 & n39178 ) ;
  assign n39180 = ~n39177 & n39179 ;
  assign n39181 = n37856 | n39180 ;
  assign n39182 = ~n39175 & n39181 ;
  assign n39183 = ( n38891 & n38892 ) | ( n38891 & ~n39182 ) | ( n38892 & ~n39182 ) ;
  assign n39184 = n39182 | n39183 ;
  assign n39185 = ~x212 & n37283 ;
  assign n39186 = x219 | n39185 ;
  assign n39187 = n38082 | n39186 ;
  assign n39188 = ~n37671 & n38158 ;
  assign n39189 = n39187 | n39188 ;
  assign n39190 = n39189 ^ n39175 ^ 1'b0 ;
  assign n39191 = ( n38856 & n39175 ) | ( n38856 & ~n39189 ) | ( n39175 & ~n39189 ) ;
  assign n39192 = ( n38856 & ~n39190 ) | ( n38856 & n39191 ) | ( ~n39190 & n39191 ) ;
  assign n39193 = x1150 & ~n39192 ;
  assign n39194 = n39184 & n39193 ;
  assign n39195 = ~n38307 & n39097 ;
  assign n39196 = n37757 & ~n37758 ;
  assign n39197 = ( n36069 & n38322 ) | ( n36069 & n39196 ) | ( n38322 & n39196 ) ;
  assign n39198 = n38322 & n39197 ;
  assign n39199 = ( x219 & ~n39195 ) | ( x219 & n39198 ) | ( ~n39195 & n39198 ) ;
  assign n39200 = ~n39195 & n39199 ;
  assign n39201 = ( ~n38856 & n38893 ) | ( ~n38856 & n39200 ) | ( n38893 & n39200 ) ;
  assign n39202 = n39200 ^ n38856 ^ 1'b0 ;
  assign n39203 = ( n39200 & n39201 ) | ( n39200 & ~n39202 ) | ( n39201 & ~n39202 ) ;
  assign n39204 = n37882 & n37891 ;
  assign n39205 = n38893 | n39204 ;
  assign n39206 = ( x1150 & n39203 ) | ( x1150 & n39205 ) | ( n39203 & n39205 ) ;
  assign n39207 = ~x1150 & n39206 ;
  assign n39208 = ( x1148 & n39194 ) | ( x1148 & n39207 ) | ( n39194 & n39207 ) ;
  assign n39209 = n39207 ^ n39194 ^ 1'b0 ;
  assign n39210 = ( x1148 & n39208 ) | ( x1148 & n39209 ) | ( n39208 & n39209 ) ;
  assign n39211 = ( ~x1149 & n39174 ) | ( ~x1149 & n39210 ) | ( n39174 & n39210 ) ;
  assign n39212 = ~x1149 & n39211 ;
  assign n39213 = ( ~x213 & n39159 ) | ( ~x213 & n39212 ) | ( n39159 & n39212 ) ;
  assign n39214 = ~x213 & n39213 ;
  assign n39215 = ( x209 & n39087 ) | ( x209 & ~n39214 ) | ( n39087 & ~n39214 ) ;
  assign n39216 = ~n39087 & n39215 ;
  assign n39217 = x1150 & n37656 ;
  assign n39218 = ~x1147 & n38876 ;
  assign n39219 = ( n15098 & n39217 ) | ( n15098 & n39218 ) | ( n39217 & n39218 ) ;
  assign n39220 = n39217 & n39219 ;
  assign n39221 = x1147 & ~n38914 ;
  assign n39222 = n38878 & ~n39217 ;
  assign n39223 = x1147 | n39222 ;
  assign n39224 = ( n7318 & ~n39221 ) | ( n7318 & n39223 ) | ( ~n39221 & n39223 ) ;
  assign n39225 = ~n7318 & n39224 ;
  assign n39226 = ( x1149 & ~n39220 ) | ( x1149 & n39225 ) | ( ~n39220 & n39225 ) ;
  assign n39227 = n39220 | n39226 ;
  assign n39236 = x212 | n38947 ;
  assign n39247 = n38949 | n39236 ;
  assign n39231 = x214 & n38880 ;
  assign n39232 = x212 & ~n39231 ;
  assign n39248 = ~x214 & n38877 ;
  assign n39249 = n39232 & ~n39248 ;
  assign n39250 = ( x219 & n39247 ) | ( x219 & ~n39249 ) | ( n39247 & ~n39249 ) ;
  assign n39251 = n39250 ^ n39247 ^ 1'b0 ;
  assign n39252 = ( x219 & n39250 ) | ( x219 & ~n39251 ) | ( n39250 & ~n39251 ) ;
  assign n39253 = n39252 ^ n38897 ^ 1'b0 ;
  assign n39254 = ( n38897 & n39252 ) | ( n38897 & n39253 ) | ( n39252 & n39253 ) ;
  assign n39255 = ( x1147 & ~n38897 ) | ( x1147 & n39254 ) | ( ~n38897 & n39254 ) ;
  assign n39256 = x219 & n38914 ;
  assign n39257 = n38925 | n38932 ;
  assign n39258 = ~x214 & n38924 ;
  assign n39259 = n38929 & ~n39258 ;
  assign n39260 = ( x219 & n39257 ) | ( x219 & ~n39259 ) | ( n39257 & ~n39259 ) ;
  assign n39261 = ~x219 & n39260 ;
  assign n39262 = ( x1147 & n39256 ) | ( x1147 & ~n39261 ) | ( n39256 & ~n39261 ) ;
  assign n39263 = ~n39256 & n39262 ;
  assign n39264 = ( n7318 & n39255 ) | ( n7318 & ~n39263 ) | ( n39255 & ~n39263 ) ;
  assign n39265 = ~n7318 & n39264 ;
  assign n39266 = ( x1150 & n37262 ) | ( x1150 & ~n39265 ) | ( n37262 & ~n39265 ) ;
  assign n39267 = ~n37262 & n39266 ;
  assign n39228 = x219 & ~n38914 ;
  assign n39229 = ( n38936 & n38964 ) | ( n38936 & n39228 ) | ( n38964 & n39228 ) ;
  assign n39230 = ~n39228 & n39229 ;
  assign n39233 = n11549 | n38878 ;
  assign n39234 = ~x214 & n39233 ;
  assign n39235 = n39232 & ~n39234 ;
  assign n39237 = x214 & n39233 ;
  assign n39238 = n39236 | n39237 ;
  assign n39239 = n39238 ^ n39235 ^ 1'b0 ;
  assign n39240 = ( n39235 & n39238 ) | ( n39235 & n39239 ) | ( n39238 & n39239 ) ;
  assign n39241 = ( x219 & ~n39235 ) | ( x219 & n39240 ) | ( ~n39235 & n39240 ) ;
  assign n39242 = ( n38032 & ~n38897 ) | ( n38032 & n39241 ) | ( ~n38897 & n39241 ) ;
  assign n39243 = ~n38032 & n39242 ;
  assign n39244 = x1150 | n37795 ;
  assign n39245 = ( ~n39230 & n39243 ) | ( ~n39230 & n39244 ) | ( n39243 & n39244 ) ;
  assign n39246 = n39230 | n39245 ;
  assign n39268 = n39267 ^ n39246 ^ 1'b0 ;
  assign n39269 = ( x1149 & ~n39246 ) | ( x1149 & n39267 ) | ( ~n39246 & n39267 ) ;
  assign n39270 = ( x1149 & ~n39268 ) | ( x1149 & n39269 ) | ( ~n39268 & n39269 ) ;
  assign n39271 = ( x1148 & n39227 ) | ( x1148 & ~n39270 ) | ( n39227 & ~n39270 ) ;
  assign n39272 = n39271 ^ n39227 ^ 1'b0 ;
  assign n39273 = ( x1148 & n39271 ) | ( x1148 & ~n39272 ) | ( n39271 & ~n39272 ) ;
  assign n39274 = n36035 & n38926 ;
  assign n39275 = n38829 & ~n39274 ;
  assign n39276 = n38964 & ~n39275 ;
  assign n39278 = x214 & ~n11549 ;
  assign n39279 = ~n38839 & n39278 ;
  assign n39280 = x212 & ~n39279 ;
  assign n39281 = n38844 & n39280 ;
  assign n39282 = ( n38926 & n39280 ) | ( n38926 & n39281 ) | ( n39280 & n39281 ) ;
  assign n39277 = n38845 & n38927 ;
  assign n39283 = ( x219 & n39277 ) | ( x219 & ~n39282 ) | ( n39277 & ~n39282 ) ;
  assign n39284 = n39282 | n39283 ;
  assign n39285 = n39276 & n39284 ;
  assign n39286 = ( x1150 & n37849 ) | ( x1150 & ~n39285 ) | ( n37849 & ~n39285 ) ;
  assign n39287 = ~n37849 & n39286 ;
  assign n39288 = n38032 | n38988 ;
  assign n39289 = n39288 ^ n39287 ^ 1'b0 ;
  assign n39290 = n38867 | n39233 ;
  assign n39291 = x214 & ~n39290 ;
  assign n39292 = n38885 & ~n39291 ;
  assign n39293 = n38883 | n39292 ;
  assign n39294 = ( n39288 & n39289 ) | ( n39288 & ~n39293 ) | ( n39289 & ~n39293 ) ;
  assign n39295 = ( n39287 & ~n39289 ) | ( n39287 & n39294 ) | ( ~n39289 & n39294 ) ;
  assign n39296 = x1150 | n37269 ;
  assign n39297 = n38903 & ~n39288 ;
  assign n39298 = ~x212 & n38827 ;
  assign n39299 = ( x219 & ~n39281 ) | ( x219 & n39298 ) | ( ~n39281 & n39298 ) ;
  assign n39300 = n39281 | n39299 ;
  assign n39301 = n39276 & n39300 ;
  assign n39302 = ( ~n39296 & n39297 ) | ( ~n39296 & n39301 ) | ( n39297 & n39301 ) ;
  assign n39303 = n39296 | n39302 ;
  assign n39304 = ( x1149 & ~n39295 ) | ( x1149 & n39303 ) | ( ~n39295 & n39303 ) ;
  assign n39305 = ~x1149 & n39304 ;
  assign n39306 = n38848 | n38849 ;
  assign n39307 = ~n39275 & n39306 ;
  assign n39308 = n38285 & n38964 ;
  assign n39309 = n39307 & n39308 ;
  assign n39310 = n38949 | n39290 ;
  assign n39311 = x212 & n39310 ;
  assign n39312 = n38874 & ~n39291 ;
  assign n39313 = x219 | n39312 ;
  assign n39314 = ( ~n39288 & n39311 ) | ( ~n39288 & n39313 ) | ( n39311 & n39313 ) ;
  assign n39315 = ~n39288 & n39314 ;
  assign n39316 = x1150 | n37789 ;
  assign n39317 = ( ~n39309 & n39315 ) | ( ~n39309 & n39316 ) | ( n39315 & n39316 ) ;
  assign n39318 = n39309 | n39317 ;
  assign n39320 = n5193 & n36298 ;
  assign n39330 = ~x57 & x1147 ;
  assign n39331 = ~n5193 & n39307 ;
  assign n39332 = ( n39320 & n39330 ) | ( n39320 & ~n39331 ) | ( n39330 & ~n39331 ) ;
  assign n39333 = ~n39320 & n39332 ;
  assign n39319 = n36298 & n38986 ;
  assign n39321 = x57 | x1147 ;
  assign n39322 = ( ~n39319 & n39320 ) | ( ~n39319 & n39321 ) | ( n39320 & n39321 ) ;
  assign n39323 = n39319 | n39322 ;
  assign n39324 = n5193 | n36297 ;
  assign n39325 = ~n39323 & n39324 ;
  assign n39326 = ( n38868 & n39323 ) | ( n38868 & ~n39325 ) | ( n39323 & ~n39325 ) ;
  assign n39327 = n39326 ^ n36298 ^ 1'b0 ;
  assign n39328 = ( ~x57 & n36298 ) | ( ~x57 & n39327 ) | ( n36298 & n39327 ) ;
  assign n39329 = ( n39326 & ~n39327 ) | ( n39326 & n39328 ) | ( ~n39327 & n39328 ) ;
  assign n39334 = n39333 ^ n39329 ^ 1'b0 ;
  assign n39335 = ( x1150 & ~n39329 ) | ( x1150 & n39333 ) | ( ~n39329 & n39333 ) ;
  assign n39336 = ( x1150 & ~n39334 ) | ( x1150 & n39335 ) | ( ~n39334 & n39335 ) ;
  assign n39337 = x1149 & ~n39336 ;
  assign n39338 = n39318 & n39337 ;
  assign n39339 = ( x1148 & n39305 ) | ( x1148 & ~n39338 ) | ( n39305 & ~n39338 ) ;
  assign n39340 = ~n39305 & n39339 ;
  assign n39341 = x213 & ~n39340 ;
  assign n39342 = n39273 & n39341 ;
  assign n39343 = ~x213 & n38945 ;
  assign n39344 = x209 | n39343 ;
  assign n39345 = ( ~n39216 & n39342 ) | ( ~n39216 & n39344 ) | ( n39342 & n39344 ) ;
  assign n39346 = ~n39216 & n39345 ;
  assign n39347 = x246 ^ x230 ^ 1'b0 ;
  assign n39348 = ( x246 & n39346 ) | ( x246 & n39347 ) | ( n39346 & n39347 ) ;
  assign n39349 = x213 & n38358 ;
  assign n39350 = ~x1147 & x1151 ;
  assign n39351 = n37631 & n39350 ;
  assign n39352 = n38138 | n38282 ;
  assign n39353 = x1147 & n39352 ;
  assign n39354 = n37296 | n38281 ;
  assign n39355 = ~n38249 & n39354 ;
  assign n39356 = n37270 & ~n39355 ;
  assign n39357 = n39353 & ~n39356 ;
  assign n39358 = ( x1150 & ~n39351 ) | ( x1150 & n39357 ) | ( ~n39351 & n39357 ) ;
  assign n39359 = n39351 | n39358 ;
  assign n39360 = ~n37719 & n39122 ;
  assign n39361 = n39132 & n39360 ;
  assign n39362 = n37270 & ~n39361 ;
  assign n39363 = n37269 | n39142 ;
  assign n39364 = x1151 & ~n39363 ;
  assign n39365 = ( x1147 & n39363 ) | ( x1147 & n39364 ) | ( n39363 & n39364 ) ;
  assign n39366 = ~n39362 & n39365 ;
  assign n39367 = x1151 | n37746 ;
  assign n39368 = ~x1147 & n39367 ;
  assign n39369 = x1151 & ~n37823 ;
  assign n39370 = n39368 & ~n39369 ;
  assign n39371 = ( x1150 & n39366 ) | ( x1150 & ~n39370 ) | ( n39366 & ~n39370 ) ;
  assign n39372 = ~n39366 & n39371 ;
  assign n39373 = ( x1149 & n39359 ) | ( x1149 & ~n39372 ) | ( n39359 & ~n39372 ) ;
  assign n39374 = n39373 ^ n39359 ^ 1'b0 ;
  assign n39375 = ( x1149 & n39373 ) | ( x1149 & ~n39374 ) | ( n39373 & ~n39374 ) ;
  assign n39376 = x1151 | n37657 ;
  assign n39389 = n7318 | n37477 ;
  assign n39390 = n37890 | n39089 ;
  assign n39391 = ~n39389 & n39390 ;
  assign n39392 = n39376 | n39391 ;
  assign n39393 = x1151 & ~n37657 ;
  assign n39394 = ~n37698 & n39393 ;
  assign n39395 = x1147 | n39394 ;
  assign n39396 = n39392 & ~n39395 ;
  assign n39397 = n38124 & ~n38283 ;
  assign n39398 = x1147 & ~n39397 ;
  assign n39399 = n37849 | n37895 ;
  assign n39400 = x1151 & ~n39399 ;
  assign n39401 = ( n39398 & n39399 ) | ( n39398 & n39400 ) | ( n39399 & n39400 ) ;
  assign n39402 = ( x1150 & n39396 ) | ( x1150 & ~n39401 ) | ( n39396 & ~n39401 ) ;
  assign n39403 = ~n39396 & n39402 ;
  assign n39377 = n38308 | n39376 ;
  assign n39378 = ~x1147 & n39377 ;
  assign n39379 = ~n37661 & n37859 ;
  assign n39380 = n37657 | n39379 ;
  assign n39381 = x1151 & ~n39380 ;
  assign n39382 = n39378 & ~n39381 ;
  assign n39383 = x1147 & ~n38338 ;
  assign n39384 = x1151 | n37849 ;
  assign n39385 = n37896 | n39384 ;
  assign n39386 = n39383 & n39385 ;
  assign n39387 = ( x1150 & ~n39382 ) | ( x1150 & n39386 ) | ( ~n39382 & n39386 ) ;
  assign n39388 = n39382 | n39387 ;
  assign n39404 = n39403 ^ n39388 ^ 1'b0 ;
  assign n39405 = ( x1149 & ~n39388 ) | ( x1149 & n39403 ) | ( ~n39388 & n39403 ) ;
  assign n39406 = ( x1149 & ~n39404 ) | ( x1149 & n39405 ) | ( ~n39404 & n39405 ) ;
  assign n39407 = ( x1148 & n39375 ) | ( x1148 & ~n39406 ) | ( n39375 & ~n39406 ) ;
  assign n39408 = ~x1148 & n39407 ;
  assign n39415 = n38159 | n39187 ;
  assign n39416 = ~n37661 & n39415 ;
  assign n39417 = n37262 | n39416 ;
  assign n39418 = x1151 & ~n39417 ;
  assign n39409 = x1151 | n37262 ;
  assign n39410 = n37757 & ~n38321 ;
  assign n39411 = n36069 | n37875 ;
  assign n39412 = n39410 & n39411 ;
  assign n39413 = n39409 | n39412 ;
  assign n39414 = ~x1147 & n39413 ;
  assign n39419 = n39418 ^ n39414 ^ 1'b0 ;
  assign n39420 = ( x1149 & ~n39414 ) | ( x1149 & n39418 ) | ( ~n39414 & n39418 ) ;
  assign n39421 = ( x1149 & ~n39419 ) | ( x1149 & n39420 ) | ( ~n39419 & n39420 ) ;
  assign n39422 = ( ~n37865 & n38157 ) | ( ~n37865 & n39187 ) | ( n38157 & n39187 ) ;
  assign n39423 = ~n37865 & n39422 ;
  assign n39424 = n38106 & ~n39423 ;
  assign n39425 = x1147 & ~n39424 ;
  assign n39426 = x1151 | n37777 ;
  assign n39427 = n39412 | n39426 ;
  assign n39428 = n37896 | n39427 ;
  assign n39429 = ( ~n39421 & n39425 ) | ( ~n39421 & n39428 ) | ( n39425 & n39428 ) ;
  assign n39430 = n39429 ^ n39421 ^ 1'b0 ;
  assign n39431 = ( n39421 & ~n39429 ) | ( n39421 & n39430 ) | ( ~n39429 & n39430 ) ;
  assign n39432 = x1151 & ~n37789 ;
  assign n39433 = ~n38254 & n39432 ;
  assign n39434 = x1151 | n37789 ;
  assign n39435 = n37788 | n39434 ;
  assign n39436 = x1147 & n39435 ;
  assign n39437 = ~n39433 & n39436 ;
  assign n39438 = n37794 & n37869 ;
  assign n39439 = x1151 | n39438 ;
  assign n39440 = ~x1147 & n39439 ;
  assign n39441 = x1151 & ~n37795 ;
  assign n39442 = ~n37336 & n38089 ;
  assign n39443 = n39441 & ~n39442 ;
  assign n39444 = n39440 & ~n39443 ;
  assign n39445 = ( x1149 & ~n39437 ) | ( x1149 & n39444 ) | ( ~n39437 & n39444 ) ;
  assign n39446 = n39437 | n39445 ;
  assign n39447 = ( x1150 & ~n39431 ) | ( x1150 & n39446 ) | ( ~n39431 & n39446 ) ;
  assign n39448 = ~x1150 & n39447 ;
  assign n39449 = n38350 & ~n39107 ;
  assign n39450 = x1147 | n39449 ;
  assign n39451 = n37881 & ~n39389 ;
  assign n39452 = n39391 | n39451 ;
  assign n39453 = n39409 | n39452 ;
  assign n39454 = ~n39450 & n39453 ;
  assign n39455 = x1147 & ~n38343 ;
  assign n39456 = n37777 | n37779 ;
  assign n39457 = x1147 & n38292 ;
  assign n39458 = ( n39455 & n39456 ) | ( n39455 & n39457 ) | ( n39456 & n39457 ) ;
  assign n39459 = ( x1149 & n39454 ) | ( x1149 & ~n39458 ) | ( n39454 & ~n39458 ) ;
  assign n39460 = ~n39454 & n39459 ;
  assign n39461 = ~x1147 & n38349 ;
  assign n39462 = n37817 & ~n39139 ;
  assign n39463 = n37789 | n39462 ;
  assign n39464 = x1151 | n39463 ;
  assign n39465 = n39464 ^ x1149 ^ 1'b0 ;
  assign n39466 = ~n39360 & n39432 ;
  assign n39467 = x1147 & ~n39466 ;
  assign n39468 = ( n39464 & ~n39465 ) | ( n39464 & n39467 ) | ( ~n39465 & n39467 ) ;
  assign n39469 = ( x1149 & n39465 ) | ( x1149 & n39468 ) | ( n39465 & n39468 ) ;
  assign n39470 = ~n37824 & n37836 ;
  assign n39471 = n39441 & ~n39470 ;
  assign n39472 = ~n39469 & n39471 ;
  assign n39473 = ( n39461 & n39469 ) | ( n39461 & ~n39472 ) | ( n39469 & ~n39472 ) ;
  assign n39474 = ( x1150 & n39460 ) | ( x1150 & n39473 ) | ( n39460 & n39473 ) ;
  assign n39475 = ~n39460 & n39474 ;
  assign n39476 = ( x1148 & n39448 ) | ( x1148 & n39475 ) | ( n39448 & n39475 ) ;
  assign n39477 = n39475 ^ n39448 ^ 1'b0 ;
  assign n39478 = ( x1148 & n39476 ) | ( x1148 & n39477 ) | ( n39476 & n39477 ) ;
  assign n39479 = ( ~x213 & n39408 ) | ( ~x213 & n39478 ) | ( n39408 & n39478 ) ;
  assign n39480 = ~x213 & n39479 ;
  assign n39481 = ( x209 & n39349 ) | ( x209 & ~n39480 ) | ( n39349 & ~n39480 ) ;
  assign n39482 = ~n39349 & n39481 ;
  assign n39485 = n38350 & ~n39452 ;
  assign n39483 = n38348 | n39451 ;
  assign n39484 = x1147 & n39483 ;
  assign n39486 = n39485 ^ n39484 ^ 1'b0 ;
  assign n39487 = ( x1150 & ~n39484 ) | ( x1150 & n39485 ) | ( ~n39484 & n39485 ) ;
  assign n39488 = ( x1150 & ~n39486 ) | ( x1150 & n39487 ) | ( ~n39486 & n39487 ) ;
  assign n39489 = ~n37797 & n37813 ;
  assign n39490 = n38350 & ~n39489 ;
  assign n39491 = n39490 ^ n39488 ^ 1'b0 ;
  assign n39492 = ( ~n39461 & n39490 ) | ( ~n39461 & n39491 ) | ( n39490 & n39491 ) ;
  assign n39493 = ( n39488 & ~n39491 ) | ( n39488 & n39492 ) | ( ~n39491 & n39492 ) ;
  assign n39494 = ~n37197 & n37745 ;
  assign n39495 = n7318 | n39494 ;
  assign n39496 = ( ~n38172 & n38215 ) | ( ~n38172 & n39495 ) | ( n38215 & n39495 ) ;
  assign n39497 = ~n38172 & n39496 ;
  assign n39498 = n39368 & n39497 ;
  assign n39499 = ~n39391 & n39393 ;
  assign n39500 = n39457 & ~n39499 ;
  assign n39501 = ( x1150 & ~n39498 ) | ( x1150 & n39500 ) | ( ~n39498 & n39500 ) ;
  assign n39502 = n39498 | n39501 ;
  assign n39503 = n39502 ^ n39493 ^ 1'b0 ;
  assign n39504 = ( n39493 & n39502 ) | ( n39493 & n39503 ) | ( n39502 & n39503 ) ;
  assign n39505 = ( x1149 & ~n39493 ) | ( x1149 & n39504 ) | ( ~n39493 & n39504 ) ;
  assign n39515 = ~n37719 & n37840 ;
  assign n39516 = n38106 & ~n39515 ;
  assign n39517 = x1147 | n39516 ;
  assign n39518 = n39360 | n39434 ;
  assign n39519 = ~n39517 & n39518 ;
  assign n39520 = n37789 | n38286 ;
  assign n39521 = x1151 & ~n39520 ;
  assign n39522 = ( n39455 & n39520 ) | ( n39455 & n39521 ) | ( n39520 & n39521 ) ;
  assign n39523 = ( x1150 & n39519 ) | ( x1150 & ~n39522 ) | ( n39519 & ~n39522 ) ;
  assign n39524 = ~n39519 & n39523 ;
  assign n39506 = n37780 | n39352 ;
  assign n39507 = n39398 & n39506 ;
  assign n39508 = n38138 | n39361 ;
  assign n39509 = n37849 | n39133 ;
  assign n39510 = x1151 & ~n39509 ;
  assign n39511 = x1147 | n39510 ;
  assign n39512 = n39508 & ~n39511 ;
  assign n39513 = ( x1150 & ~n39507 ) | ( x1150 & n39512 ) | ( ~n39507 & n39512 ) ;
  assign n39514 = n39507 | n39513 ;
  assign n39525 = n39524 ^ n39514 ^ 1'b0 ;
  assign n39526 = ( x1149 & ~n39514 ) | ( x1149 & n39524 ) | ( ~n39514 & n39524 ) ;
  assign n39527 = ( x1149 & ~n39525 ) | ( x1149 & n39526 ) | ( ~n39525 & n39526 ) ;
  assign n39528 = x1148 & ~n39527 ;
  assign n39529 = n39505 & n39528 ;
  assign n39530 = n37870 & n39350 ;
  assign n39531 = x1151 | n38307 ;
  assign n39532 = x1147 & n39531 ;
  assign n39533 = n37657 | n38308 ;
  assign n39534 = n39532 & n39533 ;
  assign n39535 = ( x1150 & ~n39530 ) | ( x1150 & n39534 ) | ( ~n39530 & n39534 ) ;
  assign n39536 = n39530 | n39535 ;
  assign n39537 = n37883 & ~n38321 ;
  assign n39538 = n37795 | n39537 ;
  assign n39539 = x1151 | n39538 ;
  assign n39540 = n38350 & ~n39412 ;
  assign n39541 = x1147 & ~n39540 ;
  assign n39542 = n39539 & n39541 ;
  assign n39543 = n15098 & n37261 ;
  assign n39544 = x1151 & ~n39543 ;
  assign n39545 = n39440 & ~n39544 ;
  assign n39546 = ( x1150 & n39542 ) | ( x1150 & ~n39545 ) | ( n39542 & ~n39545 ) ;
  assign n39547 = ~n39542 & n39546 ;
  assign n39548 = ( x1149 & n39536 ) | ( x1149 & ~n39547 ) | ( n39536 & ~n39547 ) ;
  assign n39549 = n39548 ^ n39536 ^ 1'b0 ;
  assign n39550 = ( x1149 & n39548 ) | ( x1149 & ~n39549 ) | ( n39548 & ~n39549 ) ;
  assign n39557 = x219 | n38087 ;
  assign n39558 = ( ~n37865 & n38313 ) | ( ~n37865 & n39557 ) | ( n38313 & n39557 ) ;
  assign n39559 = ~n37865 & n39558 ;
  assign n39560 = n37789 | n39559 ;
  assign n39561 = x1151 & ~n39560 ;
  assign n39562 = ( n39425 & n39560 ) | ( n39425 & n39561 ) | ( n39560 & n39561 ) ;
  assign n39551 = n38254 | n39434 ;
  assign n39552 = n37324 & ~n37336 ;
  assign n39553 = n38106 & ~n39552 ;
  assign n39554 = ~n38254 & n39553 ;
  assign n39555 = x1147 | n39554 ;
  assign n39556 = n39551 & ~n39555 ;
  assign n39563 = ( x1150 & ~n39556 ) | ( x1150 & n39562 ) | ( ~n39556 & n39562 ) ;
  assign n39564 = ~n39562 & n39563 ;
  assign n39565 = ~n9344 & n39552 ;
  assign n39566 = n39355 | n39565 ;
  assign n39567 = n38124 & ~n39566 ;
  assign n39568 = n38138 | n39355 ;
  assign n39569 = ~x1147 & n39568 ;
  assign n39570 = n39569 ^ n39567 ^ 1'b0 ;
  assign n39571 = ( n39567 & n39569 ) | ( n39567 & n39570 ) | ( n39569 & n39570 ) ;
  assign n39572 = ( x1150 & ~n39567 ) | ( x1150 & n39571 ) | ( ~n39567 & n39571 ) ;
  assign n39573 = n37860 & n39559 ;
  assign n39574 = n38138 | n39573 ;
  assign n39575 = n39572 ^ n39383 ^ 1'b0 ;
  assign n39576 = ( ~n39383 & n39574 ) | ( ~n39383 & n39575 ) | ( n39574 & n39575 ) ;
  assign n39577 = ( n39383 & n39572 ) | ( n39383 & n39576 ) | ( n39572 & n39576 ) ;
  assign n39578 = x1149 & ~n39577 ;
  assign n39579 = ( x1149 & n39564 ) | ( x1149 & n39578 ) | ( n39564 & n39578 ) ;
  assign n39580 = ( x1148 & n39550 ) | ( x1148 & ~n39579 ) | ( n39550 & ~n39579 ) ;
  assign n39581 = ~x1148 & n39580 ;
  assign n39582 = ( x213 & n39529 ) | ( x213 & n39581 ) | ( n39529 & n39581 ) ;
  assign n39583 = n39581 ^ n39529 ^ 1'b0 ;
  assign n39584 = ( x213 & n39582 ) | ( x213 & n39583 ) | ( n39582 & n39583 ) ;
  assign n39585 = ~x213 & n37904 ;
  assign n39586 = x209 | n39585 ;
  assign n39587 = ( ~n39482 & n39584 ) | ( ~n39482 & n39586 ) | ( n39584 & n39586 ) ;
  assign n39588 = ~n39482 & n39587 ;
  assign n39589 = x247 ^ x230 ^ 1'b0 ;
  assign n39590 = ( x247 & n39588 ) | ( x247 & n39589 ) | ( n39588 & n39589 ) ;
  assign n39591 = ~n39362 & n39568 ;
  assign n39592 = x1152 & ~n39591 ;
  assign n39593 = n39352 & ~n39364 ;
  assign n39594 = x1152 | n39593 ;
  assign n39595 = ( x1150 & ~n39592 ) | ( x1150 & n39594 ) | ( ~n39592 & n39594 ) ;
  assign n39596 = ~x1150 & n39595 ;
  assign n39597 = n37866 | n39384 ;
  assign n39598 = x1152 & n39597 ;
  assign n39599 = ~n39397 & n39598 ;
  assign n39600 = ~x1152 & n39385 ;
  assign n39601 = ~n39400 & n39600 ;
  assign n39602 = ( x1150 & n39599 ) | ( x1150 & n39601 ) | ( n39599 & n39601 ) ;
  assign n39603 = n39601 ^ n39599 ^ 1'b0 ;
  assign n39604 = ( x1150 & n39602 ) | ( x1150 & n39603 ) | ( n39602 & n39603 ) ;
  assign n39605 = ( x1148 & n39596 ) | ( x1148 & ~n39604 ) | ( n39596 & ~n39604 ) ;
  assign n39606 = ~n39596 & n39605 ;
  assign n39607 = x1151 & ~x1152 ;
  assign n39608 = n37746 & n39607 ;
  assign n39609 = x1152 & ~n39369 ;
  assign n39610 = x1151 | n37631 ;
  assign n39611 = n39609 & n39610 ;
  assign n39612 = ( x1150 & ~n39608 ) | ( x1150 & n39611 ) | ( ~n39608 & n39611 ) ;
  assign n39613 = n39608 | n39612 ;
  assign n39614 = x1151 | n39380 ;
  assign n39615 = x1152 & ~n39394 ;
  assign n39616 = n39614 & n39615 ;
  assign n39617 = ~x1152 & n39377 ;
  assign n39618 = ~n39499 & n39617 ;
  assign n39619 = ( x1150 & n39616 ) | ( x1150 & ~n39618 ) | ( n39616 & ~n39618 ) ;
  assign n39620 = ~n39616 & n39619 ;
  assign n39621 = ( x1148 & n39613 ) | ( x1148 & ~n39620 ) | ( n39613 & ~n39620 ) ;
  assign n39622 = n39621 ^ n39613 ^ 1'b0 ;
  assign n39623 = ( x1148 & n39621 ) | ( x1148 & ~n39622 ) | ( n39621 & ~n39622 ) ;
  assign n39624 = ( x1149 & ~n39606 ) | ( x1149 & n39623 ) | ( ~n39606 & n39623 ) ;
  assign n39625 = ~x1149 & n39624 ;
  assign n39626 = x1152 & ~n38343 ;
  assign n39627 = n39423 | n39426 ;
  assign n39628 = n39626 & n39627 ;
  assign n39629 = x1151 & ~n37736 ;
  assign n39630 = ~n39456 & n39629 ;
  assign n39631 = ( x1152 & n39428 ) | ( x1152 & ~n39630 ) | ( n39428 & ~n39630 ) ;
  assign n39632 = ~x1152 & n39631 ;
  assign n39633 = ( x1150 & n39628 ) | ( x1150 & ~n39632 ) | ( n39628 & ~n39632 ) ;
  assign n39634 = ~n39628 & n39633 ;
  assign n39635 = x1152 & n39551 ;
  assign n39636 = ~n39466 & n39635 ;
  assign n39637 = ~x1152 & n39435 ;
  assign n39638 = x1151 & ~n39463 ;
  assign n39639 = n39637 & ~n39638 ;
  assign n39640 = ( x1150 & ~n39636 ) | ( x1150 & n39639 ) | ( ~n39636 & n39639 ) ;
  assign n39641 = n39636 | n39640 ;
  assign n39642 = ( x1148 & n39634 ) | ( x1148 & n39641 ) | ( n39634 & n39641 ) ;
  assign n39643 = ~n39634 & n39642 ;
  assign n39644 = n38348 | n39442 ;
  assign n39645 = x1152 & ~n39471 ;
  assign n39646 = n39644 & n39645 ;
  assign n39647 = x1150 | n39646 ;
  assign n39648 = ~n37819 & n39441 ;
  assign n39649 = x1152 | n39648 ;
  assign n39650 = ~n39647 & n39649 ;
  assign n39651 = ( n39439 & n39647 ) | ( n39439 & ~n39650 ) | ( n39647 & ~n39650 ) ;
  assign n39652 = ~x1152 & n39413 ;
  assign n39653 = ~n39485 & n39652 ;
  assign n39654 = x1152 & ~n39449 ;
  assign n39655 = x1151 | n39417 ;
  assign n39656 = n39654 & n39655 ;
  assign n39657 = ( x1150 & n39653 ) | ( x1150 & ~n39656 ) | ( n39653 & ~n39656 ) ;
  assign n39658 = ~n39653 & n39657 ;
  assign n39659 = ( x1148 & n39651 ) | ( x1148 & ~n39658 ) | ( n39651 & ~n39658 ) ;
  assign n39660 = ~x1148 & n39659 ;
  assign n39661 = ( x1149 & n39643 ) | ( x1149 & n39660 ) | ( n39643 & n39660 ) ;
  assign n39662 = n39660 ^ n39643 ^ 1'b0 ;
  assign n39663 = ( x1149 & n39661 ) | ( x1149 & n39662 ) | ( n39661 & n39662 ) ;
  assign n39664 = ( ~x213 & n39625 ) | ( ~x213 & n39663 ) | ( n39625 & n39663 ) ;
  assign n39665 = ~x213 & n39664 ;
  assign n39666 = n39597 & n39626 ;
  assign n39667 = x1151 & ~n37791 ;
  assign n39668 = ( x1152 & n38339 ) | ( x1152 & ~n39667 ) | ( n38339 & ~n39667 ) ;
  assign n39669 = ~x1152 & n39668 ;
  assign n39670 = ( x1150 & n39666 ) | ( x1150 & ~n39669 ) | ( n39666 & ~n39669 ) ;
  assign n39671 = ~n39666 & n39670 ;
  assign n39672 = x1151 | n37870 ;
  assign n39673 = n37631 | n39672 ;
  assign n39674 = x1152 & ~n38351 ;
  assign n39675 = n39673 & n39674 ;
  assign n39676 = x1150 | n39675 ;
  assign n39677 = n37820 & n39607 ;
  assign n39678 = ( ~n39671 & n39676 ) | ( ~n39671 & n39677 ) | ( n39676 & n39677 ) ;
  assign n39679 = ~n39671 & n39678 ;
  assign n39680 = x213 & n39679 ;
  assign n39681 = ( x209 & n39665 ) | ( x209 & ~n39680 ) | ( n39665 & ~n39680 ) ;
  assign n39682 = ~n39665 & n39681 ;
  assign n39683 = x1152 & n39377 ;
  assign n39684 = ~n39540 & n39683 ;
  assign n39685 = ~x1152 & n39531 ;
  assign n39686 = x1151 & ~n39538 ;
  assign n39687 = n39685 & ~n39686 ;
  assign n39688 = ( x1150 & ~n39684 ) | ( x1150 & n39687 ) | ( ~n39684 & n39687 ) ;
  assign n39689 = n39684 | n39688 ;
  assign n39690 = ~x1152 & n39574 ;
  assign n39691 = ~n39561 & n39690 ;
  assign n39692 = ~n39424 & n39598 ;
  assign n39693 = ( x1150 & n39691 ) | ( x1150 & ~n39692 ) | ( n39691 & ~n39692 ) ;
  assign n39694 = ~n39691 & n39693 ;
  assign n39695 = ( x1149 & n39689 ) | ( x1149 & ~n39694 ) | ( n39689 & ~n39694 ) ;
  assign n39696 = ~x1149 & n39695 ;
  assign n39697 = n38283 | n39384 ;
  assign n39698 = n39626 & n39697 ;
  assign n39699 = ~x1152 & n39506 ;
  assign n39700 = ~n39521 & n39699 ;
  assign n39701 = ( x1150 & n39698 ) | ( x1150 & ~n39700 ) | ( n39698 & ~n39700 ) ;
  assign n39702 = ~n39698 & n39701 ;
  assign n39703 = x1152 & n39392 ;
  assign n39704 = ~n39485 & n39703 ;
  assign n39705 = n39441 & ~n39451 ;
  assign n39706 = n38293 & ~n39705 ;
  assign n39707 = ( x1150 & ~n39704 ) | ( x1150 & n39706 ) | ( ~n39704 & n39706 ) ;
  assign n39708 = n39704 | n39707 ;
  assign n39709 = ( x1149 & n39702 ) | ( x1149 & n39708 ) | ( n39702 & n39708 ) ;
  assign n39710 = ~n39702 & n39709 ;
  assign n39711 = ( x1148 & n39696 ) | ( x1148 & ~n39710 ) | ( n39696 & ~n39710 ) ;
  assign n39712 = ~n39696 & n39711 ;
  assign n39713 = x1152 | n39466 ;
  assign n39714 = n39508 & ~n39713 ;
  assign n39715 = x1152 & ~n39516 ;
  assign n39716 = x1151 | n39509 ;
  assign n39717 = n39715 & n39716 ;
  assign n39718 = ( x1150 & n39714 ) | ( x1150 & ~n39717 ) | ( n39714 & ~n39717 ) ;
  assign n39719 = ~n39714 & n39718 ;
  assign n39720 = x1151 | n39497 ;
  assign n39721 = x1152 & ~n39490 ;
  assign n39722 = n39720 & n39721 ;
  assign n39723 = x1150 | n39722 ;
  assign n39724 = n39649 & ~n39723 ;
  assign n39725 = ( n39367 & n39723 ) | ( n39367 & ~n39724 ) | ( n39723 & ~n39724 ) ;
  assign n39726 = ( x1149 & n39719 ) | ( x1149 & n39725 ) | ( n39719 & n39725 ) ;
  assign n39727 = ~n39719 & n39726 ;
  assign n39728 = n39438 & n39607 ;
  assign n39729 = x1152 & ~n39544 ;
  assign n39730 = n39672 & n39729 ;
  assign n39731 = ( x1150 & ~n39728 ) | ( x1150 & n39730 ) | ( ~n39728 & n39730 ) ;
  assign n39732 = n39728 | n39731 ;
  assign n39733 = n39384 | n39566 ;
  assign n39734 = x1152 & ~n39554 ;
  assign n39735 = n39733 & n39734 ;
  assign n39736 = ~x1152 & n39568 ;
  assign n39737 = ~n39433 & n39736 ;
  assign n39738 = ( x1150 & n39735 ) | ( x1150 & ~n39737 ) | ( n39735 & ~n39737 ) ;
  assign n39739 = ~n39735 & n39738 ;
  assign n39740 = ( x1149 & n39732 ) | ( x1149 & ~n39739 ) | ( n39732 & ~n39739 ) ;
  assign n39741 = ~x1149 & n39740 ;
  assign n39742 = ( x1148 & ~n39727 ) | ( x1148 & n39741 ) | ( ~n39727 & n39741 ) ;
  assign n39743 = n39727 | n39742 ;
  assign n39744 = ( x213 & n39712 ) | ( x213 & n39743 ) | ( n39712 & n39743 ) ;
  assign n39745 = ~n39712 & n39744 ;
  assign n39746 = ~x213 & n39086 ;
  assign n39747 = x209 | n39746 ;
  assign n39748 = ( ~n39682 & n39745 ) | ( ~n39682 & n39747 ) | ( n39745 & n39747 ) ;
  assign n39749 = ~n39682 & n39748 ;
  assign n39750 = x248 ^ x230 ^ 1'b0 ;
  assign n39751 = ( x248 & n39749 ) | ( x248 & n39750 ) | ( n39749 & n39750 ) ;
  assign n39752 = x214 & ~n36638 ;
  assign n39753 = n36563 & ~n39752 ;
  assign n39754 = x219 | n39753 ;
  assign n39755 = x212 & n36638 ;
  assign n39756 = ( ~n36644 & n39754 ) | ( ~n36644 & n39755 ) | ( n39754 & n39755 ) ;
  assign n39757 = ~n36644 & n39756 ;
  assign n39758 = ( x1151 & n37777 ) | ( x1151 & ~n39757 ) | ( n37777 & ~n39757 ) ;
  assign n39759 = ~n37777 & n39758 ;
  assign n39760 = x214 & ~n36640 ;
  assign n39761 = n36562 & ~n39760 ;
  assign n39762 = x212 | n39761 ;
  assign n39763 = ( n36561 & n36638 ) | ( n36561 & ~n36639 ) | ( n36638 & ~n36639 ) ;
  assign n39764 = ( x212 & n36069 ) | ( x212 & ~n39763 ) | ( n36069 & ~n39763 ) ;
  assign n39765 = ( x212 & ~x214 ) | ( x212 & n39764 ) | ( ~x214 & n39764 ) ;
  assign n39766 = n39765 ^ x214 ^ 1'b0 ;
  assign n39767 = ( x214 & ~n36640 ) | ( x214 & n39766 ) | ( ~n36640 & n39766 ) ;
  assign n39768 = ( n39765 & ~n39766 ) | ( n39765 & n39767 ) | ( ~n39766 & n39767 ) ;
  assign n39769 = ( x219 & n39762 ) | ( x219 & ~n39768 ) | ( n39762 & ~n39768 ) ;
  assign n39770 = n39769 ^ n39762 ^ 1'b0 ;
  assign n39771 = ( x219 & n39769 ) | ( x219 & ~n39770 ) | ( n39769 & ~n39770 ) ;
  assign n39772 = n36644 | n39771 ;
  assign n39773 = ( ~n36644 & n39384 ) | ( ~n36644 & n39772 ) | ( n39384 & n39772 ) ;
  assign n39774 = ( x1152 & n39759 ) | ( x1152 & n39773 ) | ( n39759 & n39773 ) ;
  assign n39775 = ~n39759 & n39774 ;
  assign n39777 = n36678 ^ n36186 ^ n36185 ;
  assign n39776 = x207 | n36806 ;
  assign n39778 = ( x208 & n39776 ) | ( x208 & n39777 ) | ( n39776 & n39777 ) ;
  assign n39779 = ~n39777 & n39778 ;
  assign n39780 = n36807 & ~n39779 ;
  assign n39781 = ( n36142 & n39779 ) | ( n36142 & ~n39780 ) | ( n39779 & ~n39780 ) ;
  assign n39782 = x211 | n39781 ;
  assign n39783 = ~n36622 & n39782 ;
  assign n39796 = n36035 & n39783 ;
  assign n39797 = x219 & ~n36619 ;
  assign n39798 = n39797 ^ n39796 ^ 1'b0 ;
  assign n39799 = ( n39796 & n39797 ) | ( n39796 & n39798 ) | ( n39797 & n39798 ) ;
  assign n39800 = ( n7318 & ~n39796 ) | ( n7318 & n39799 ) | ( ~n39796 & n39799 ) ;
  assign n39785 = x214 & ~n39781 ;
  assign n39784 = x214 & ~n39783 ;
  assign n39786 = n39785 ^ n39784 ^ n36598 ;
  assign n39787 = ~x212 & n39786 ;
  assign n39788 = x219 | n39787 ;
  assign n39789 = ~x211 & n36598 ;
  assign n39790 = x211 & n39781 ;
  assign n39791 = ( x214 & ~n39789 ) | ( x214 & n39790 ) | ( ~n39789 & n39790 ) ;
  assign n39792 = n39789 | n39791 ;
  assign n39793 = x212 & n39792 ;
  assign n39794 = ~n39785 & n39793 ;
  assign n39795 = n39788 | n39794 ;
  assign n39801 = n39800 ^ n39795 ^ 1'b0 ;
  assign n39802 = ( n39432 & ~n39795 ) | ( n39432 & n39800 ) | ( ~n39795 & n39800 ) ;
  assign n39803 = ( n39432 & ~n39801 ) | ( n39432 & n39802 ) | ( ~n39801 & n39802 ) ;
  assign n39804 = ~x212 & n36598 ;
  assign n39805 = x219 | n39804 ;
  assign n39806 = x212 & n39786 ;
  assign n39807 = ( ~n39800 & n39805 ) | ( ~n39800 & n39806 ) | ( n39805 & n39806 ) ;
  assign n39808 = ~n39800 & n39807 ;
  assign n39809 = ( x1151 & n37269 ) | ( x1151 & ~n39808 ) | ( n37269 & ~n39808 ) ;
  assign n39810 = n39808 | n39809 ;
  assign n39811 = ( x1152 & ~n39803 ) | ( x1152 & n39810 ) | ( ~n39803 & n39810 ) ;
  assign n39812 = ~x1152 & n39811 ;
  assign n39813 = ( x1150 & n39775 ) | ( x1150 & ~n39812 ) | ( n39775 & ~n39812 ) ;
  assign n39814 = ~n39775 & n39813 ;
  assign n39815 = n36561 | n37197 ;
  assign n39816 = ~n36640 & n37197 ;
  assign n39817 = ( n7318 & n39815 ) | ( n7318 & ~n39816 ) | ( n39815 & ~n39816 ) ;
  assign n39818 = ~n7318 & n39817 ;
  assign n39819 = ( x1151 & n37657 ) | ( x1151 & ~n39818 ) | ( n37657 & ~n39818 ) ;
  assign n39820 = n39818 | n39819 ;
  assign n39821 = n7318 | n36635 ;
  assign n39822 = ( x212 & x214 ) | ( x212 & n39755 ) | ( x214 & n39755 ) ;
  assign n39823 = ~n39760 & n39822 ;
  assign n39824 = ( x219 & n39753 ) | ( x219 & ~n39823 ) | ( n39753 & ~n39823 ) ;
  assign n39825 = n39823 | n39824 ;
  assign n39826 = n38350 & ~n39825 ;
  assign n39827 = ( n38350 & n39821 ) | ( n38350 & n39826 ) | ( n39821 & n39826 ) ;
  assign n39828 = x1152 & ~n39827 ;
  assign n39829 = n39820 & n39828 ;
  assign n39830 = ~n39784 & n39793 ;
  assign n39831 = ( ~n36695 & n39788 ) | ( ~n36695 & n39830 ) | ( n39788 & n39830 ) ;
  assign n39832 = ~n36695 & n39831 ;
  assign n39833 = ( x1151 & n37795 ) | ( x1151 & ~n39832 ) | ( n37795 & ~n39832 ) ;
  assign n39834 = ~n37795 & n39833 ;
  assign n39835 = x1152 | n7318 ;
  assign n39836 = n36598 & ~n39835 ;
  assign n39837 = ( n39607 & ~n39834 ) | ( n39607 & n39836 ) | ( ~n39834 & n39836 ) ;
  assign n39838 = ~n39834 & n39837 ;
  assign n39839 = ( x1150 & ~n39829 ) | ( x1150 & n39838 ) | ( ~n39829 & n39838 ) ;
  assign n39840 = n39829 | n39839 ;
  assign n39841 = ( x213 & ~n39814 ) | ( x213 & n39840 ) | ( ~n39814 & n39840 ) ;
  assign n39842 = ~x213 & n39841 ;
  assign n39843 = x213 & n36701 ;
  assign n39844 = ( x209 & n39842 ) | ( x209 & ~n39843 ) | ( n39842 & ~n39843 ) ;
  assign n39845 = ~n39842 & n39844 ;
  assign n39846 = ~x213 & n39679 ;
  assign n39847 = ~n36150 & n37808 ;
  assign n39848 = x211 & n38214 ;
  assign n39849 = ( n36369 & n39847 ) | ( n36369 & ~n39848 ) | ( n39847 & ~n39848 ) ;
  assign n39850 = ~n39847 & n39849 ;
  assign n39851 = x211 | n38214 ;
  assign n39852 = n9344 & ~n39851 ;
  assign n39853 = n36696 | n37745 ;
  assign n39854 = ~n39852 & n39853 ;
  assign n39855 = n39854 ^ n39850 ^ 1'b0 ;
  assign n39856 = ( n39850 & n39854 ) | ( n39850 & n39855 ) | ( n39854 & n39855 ) ;
  assign n39857 = ( x219 & ~n39850 ) | ( x219 & n39856 ) | ( ~n39850 & n39856 ) ;
  assign n39858 = x1151 & ~n37797 ;
  assign n39859 = n39857 & n39858 ;
  assign n39860 = n36492 & ~n37457 ;
  assign n39861 = x299 & n36452 ;
  assign n39862 = ~n9344 & n39861 ;
  assign n39863 = n37330 | n39862 ;
  assign n39864 = n39860 & n39863 ;
  assign n39865 = ( n36676 & ~n39859 ) | ( n36676 & n39864 ) | ( ~n39859 & n39864 ) ;
  assign n39866 = n39859 | n39865 ;
  assign n39867 = x299 & ~n36452 ;
  assign n39868 = n38082 & ~n39867 ;
  assign n39869 = n37290 & ~n39867 ;
  assign n39870 = ( x212 & x214 ) | ( x212 & n39869 ) | ( x214 & n39869 ) ;
  assign n39871 = ( x212 & ~n36069 ) | ( x212 & n39870 ) | ( ~n36069 & n39870 ) ;
  assign n39872 = n39871 ^ n38299 ^ 1'b0 ;
  assign n39873 = ( ~n37851 & n38299 ) | ( ~n37851 & n39872 ) | ( n38299 & n39872 ) ;
  assign n39874 = ( n39871 & ~n39872 ) | ( n39871 & n39873 ) | ( ~n39872 & n39873 ) ;
  assign n39875 = ( n39186 & ~n39868 ) | ( n39186 & n39874 ) | ( ~n39868 & n39874 ) ;
  assign n39876 = n39868 | n39875 ;
  assign n39877 = ( x1151 & ~n37865 ) | ( x1151 & n39876 ) | ( ~n37865 & n39876 ) ;
  assign n39878 = ~x1151 & n39877 ;
  assign n39879 = x1152 & ~n36455 ;
  assign n39880 = ( x1152 & ~n36038 ) | ( x1152 & n39879 ) | ( ~n36038 & n39879 ) ;
  assign n39884 = ( n7318 & n37686 ) | ( n7318 & n37893 ) | ( n37686 & n37893 ) ;
  assign n39881 = n36450 | n39862 ;
  assign n39882 = n37778 & n39881 ;
  assign n39883 = n38277 | n39882 ;
  assign n39885 = ( x1151 & n39883 ) | ( x1151 & n39884 ) | ( n39883 & n39884 ) ;
  assign n39886 = ~n39884 & n39885 ;
  assign n39887 = ( n39878 & n39880 ) | ( n39878 & ~n39886 ) | ( n39880 & ~n39886 ) ;
  assign n39888 = ~n39878 & n39887 ;
  assign n39889 = n37757 & ~n39867 ;
  assign n39890 = n37350 & n39889 ;
  assign n39891 = x212 | n39890 ;
  assign n39892 = n37309 | n37754 ;
  assign n39893 = x214 & ~n38229 ;
  assign n39894 = x212 & ~n39893 ;
  assign n39895 = ( x212 & ~n39892 ) | ( x212 & n39894 ) | ( ~n39892 & n39894 ) ;
  assign n39896 = n39895 ^ x214 ^ 1'b0 ;
  assign n39897 = ( x214 & ~n39889 ) | ( x214 & n39896 ) | ( ~n39889 & n39896 ) ;
  assign n39898 = ( n39895 & ~n39896 ) | ( n39895 & n39897 ) | ( ~n39896 & n39897 ) ;
  assign n39899 = ( x219 & n39891 ) | ( x219 & ~n39898 ) | ( n39891 & ~n39898 ) ;
  assign n39900 = n39899 ^ n39891 ^ 1'b0 ;
  assign n39901 = ( x219 & n39899 ) | ( x219 & ~n39900 ) | ( n39899 & ~n39900 ) ;
  assign n39902 = ( n5193 & ~n38320 ) | ( n5193 & n39901 ) | ( ~n38320 & n39901 ) ;
  assign n39903 = ~n5193 & n39902 ;
  assign n39904 = n5193 & n36493 ;
  assign n39905 = x57 | x1151 ;
  assign n39906 = ( ~n39903 & n39904 ) | ( ~n39903 & n39905 ) | ( n39904 & n39905 ) ;
  assign n39907 = n39903 | n39906 ;
  assign n39908 = ~n37330 & n37359 ;
  assign n39909 = n37345 | n39861 ;
  assign n39910 = x214 | n39909 ;
  assign n39911 = ( x212 & n39908 ) | ( x212 & n39910 ) | ( n39908 & n39910 ) ;
  assign n39912 = ~n39908 & n39911 ;
  assign n39913 = x214 & ~n39909 ;
  assign n39914 = ~x212 & n37350 ;
  assign n39915 = ~n39913 & n39914 ;
  assign n39916 = ( x219 & ~n39912 ) | ( x219 & n39915 ) | ( ~n39912 & n39915 ) ;
  assign n39917 = n39912 | n39916 ;
  assign n39918 = ( n5193 & ~n37477 ) | ( n5193 & n39917 ) | ( ~n37477 & n39917 ) ;
  assign n39919 = ~n5193 & n39918 ;
  assign n39920 = ~x57 & x1151 ;
  assign n39921 = ( n39904 & ~n39919 ) | ( n39904 & n39920 ) | ( ~n39919 & n39920 ) ;
  assign n39922 = ~n39904 & n39921 ;
  assign n39923 = n36493 & ~n39922 ;
  assign n39924 = ( x57 & n39922 ) | ( x57 & ~n39923 ) | ( n39922 & ~n39923 ) ;
  assign n39925 = ( x1152 & n39907 ) | ( x1152 & ~n39924 ) | ( n39907 & ~n39924 ) ;
  assign n39926 = n39925 ^ n39907 ^ 1'b0 ;
  assign n39927 = ( x1152 & n39925 ) | ( x1152 & ~n39926 ) | ( n39925 & ~n39926 ) ;
  assign n39928 = ( x1150 & n39888 ) | ( x1150 & n39927 ) | ( n39888 & n39927 ) ;
  assign n39929 = ~n39888 & n39928 ;
  assign n39930 = n37445 & ~n37718 ;
  assign n39931 = x219 | n37710 ;
  assign n39932 = n37708 | n39861 ;
  assign n39933 = x212 & ~n38221 ;
  assign n39934 = n39932 & n39933 ;
  assign n39935 = ( n39868 & ~n39931 ) | ( n39868 & n39934 ) | ( ~n39931 & n39934 ) ;
  assign n39936 = n39931 | n39935 ;
  assign n39937 = n39930 & n39936 ;
  assign n39938 = ~n39864 & n39880 ;
  assign n39939 = ~x1151 & n39355 ;
  assign n39940 = n39938 & ~n39939 ;
  assign n39941 = n39940 ^ n39937 ^ 1'b0 ;
  assign n39942 = ( n39937 & n39940 ) | ( n39937 & n39941 ) | ( n39940 & n39941 ) ;
  assign n39943 = ( x1150 & ~n39937 ) | ( x1150 & n39942 ) | ( ~n39937 & n39942 ) ;
  assign n39944 = ~n39929 & n39943 ;
  assign n39945 = ( n39866 & n39929 ) | ( n39866 & ~n39944 ) | ( n39929 & ~n39944 ) ;
  assign n39946 = ( x213 & ~n36501 ) | ( x213 & n39945 ) | ( ~n36501 & n39945 ) ;
  assign n39947 = ( x209 & n36501 ) | ( x209 & n39946 ) | ( n36501 & n39946 ) ;
  assign n39948 = ( ~n39845 & n39846 ) | ( ~n39845 & n39947 ) | ( n39846 & n39947 ) ;
  assign n39949 = ~n39845 & n39948 ;
  assign n39950 = x249 ^ x230 ^ 1'b0 ;
  assign n39951 = ( x249 & n39949 ) | ( x249 & n39950 ) | ( n39949 & n39950 ) ;
  assign n39952 = ~n2095 & n10164 ;
  assign n39953 = ( ~x75 & n5019 ) | ( ~x75 & n39952 ) | ( n5019 & n39952 ) ;
  assign n39954 = ~x75 & n39953 ;
  assign n39955 = ( ~n6259 & n7460 ) | ( ~n6259 & n39954 ) | ( n7460 & n39954 ) ;
  assign n39956 = n39954 ^ n6259 ^ 1'b0 ;
  assign n39957 = ( n39954 & n39955 ) | ( n39954 & ~n39956 ) | ( n39955 & ~n39956 ) ;
  assign n39958 = x87 | x250 ;
  assign n39959 = ( n10138 & n39957 ) | ( n10138 & ~n39958 ) | ( n39957 & ~n39958 ) ;
  assign n39960 = ~n10138 & n39959 ;
  assign n39961 = ~x200 & x1053 ;
  assign n39962 = x200 & x1039 ;
  assign n39963 = ( x199 & ~n39961 ) | ( x199 & n39962 ) | ( ~n39961 & n39962 ) ;
  assign n39964 = n39961 | n39963 ;
  assign n39965 = ~x476 & n10073 ;
  assign n39966 = x897 & ~n9353 ;
  assign n39967 = n39965 | n39966 ;
  assign n39968 = n39967 ^ x251 ^ 1'b0 ;
  assign n39969 = ( x251 & n39964 ) | ( x251 & n39968 ) | ( n39964 & n39968 ) ;
  assign n39970 = ~n9605 & n10184 ;
  assign n39971 = x979 | x984 ;
  assign n39972 = x1001 & ~n39971 ;
  assign n39973 = n5071 & n39972 ;
  assign n39974 = n5021 & n39973 ;
  assign n39975 = ~n5362 & n39974 ;
  assign n39976 = x252 | n39975 ;
  assign n39977 = x1092 & ~x1093 ;
  assign n39978 = n39976 & n39977 ;
  assign n39979 = n39978 ^ n5371 ^ 1'b0 ;
  assign n39980 = ( ~n5371 & n5374 ) | ( ~n5371 & n39979 ) | ( n5374 & n39979 ) ;
  assign n39981 = n10184 ^ n5083 ^ 1'b0 ;
  assign n39982 = ( n10184 & n39980 ) | ( n10184 & ~n39981 ) | ( n39980 & ~n39981 ) ;
  assign n39983 = n5061 & n39982 ;
  assign n39984 = n10184 ^ n5099 ^ 1'b0 ;
  assign n39985 = ( n10184 & n39980 ) | ( n10184 & n39984 ) | ( n39980 & n39984 ) ;
  assign n39986 = ~n5061 & n39985 ;
  assign n39987 = ( x299 & n39983 ) | ( x299 & ~n39986 ) | ( n39983 & ~n39986 ) ;
  assign n39988 = ~n39983 & n39987 ;
  assign n39989 = ~n5114 & n39985 ;
  assign n39990 = n5114 & n39982 ;
  assign n39991 = ( x299 & ~n39989 ) | ( x299 & n39990 ) | ( ~n39989 & n39990 ) ;
  assign n39992 = n39989 | n39991 ;
  assign n39993 = ( n9605 & n39988 ) | ( n9605 & n39992 ) | ( n39988 & n39992 ) ;
  assign n39994 = ~n39988 & n39993 ;
  assign n39995 = ( n10841 & n39970 ) | ( n10841 & ~n39994 ) | ( n39970 & ~n39994 ) ;
  assign n39996 = ~n39970 & n39995 ;
  assign n39997 = x57 & n10183 ;
  assign n39998 = n10841 | n39997 ;
  assign n39999 = n9604 & n39973 ;
  assign n40000 = ~n19509 & n39999 ;
  assign n40001 = ( ~n5065 & n35899 ) | ( ~n5065 & n40000 ) | ( n35899 & n40000 ) ;
  assign n40002 = n5065 & n40001 ;
  assign n40003 = n40002 ^ n5362 ^ 1'b0 ;
  assign n40004 = ( n5362 & n40002 ) | ( n5362 & n40003 ) | ( n40002 & n40003 ) ;
  assign n40005 = ( x252 & ~n5362 ) | ( x252 & n40004 ) | ( ~n5362 & n40004 ) ;
  assign n40006 = ( x57 & x1092 ) | ( x57 & n40005 ) | ( x1092 & n40005 ) ;
  assign n40007 = ~x57 & n40006 ;
  assign n40008 = ( ~n39996 & n39998 ) | ( ~n39996 & n40007 ) | ( n39998 & n40007 ) ;
  assign n40009 = ~n39996 & n40008 ;
  assign n40010 = x1151 | n9343 ;
  assign n40011 = n36909 & n40010 ;
  assign n40012 = n37200 & n38496 ;
  assign n40013 = x1151 | n10076 ;
  assign n40014 = ( n36158 & ~n40012 ) | ( n36158 & n40013 ) | ( ~n40012 & n40013 ) ;
  assign n40015 = n40012 | n40014 ;
  assign n40016 = n11549 | n36094 ;
  assign n40017 = x1153 & ~n40016 ;
  assign n40018 = n10008 | n11550 ;
  assign n40019 = x1151 & n40018 ;
  assign n40020 = ~n40017 & n40019 ;
  assign n40021 = ( n7318 & n40015 ) | ( n7318 & ~n40020 ) | ( n40015 & ~n40020 ) ;
  assign n40022 = ~n7318 & n40021 ;
  assign n40023 = ( x1152 & n40011 ) | ( x1152 & ~n40022 ) | ( n40011 & ~n40022 ) ;
  assign n40024 = ~n40011 & n40023 ;
  assign n40025 = ~n10075 & n36909 ;
  assign n40026 = n36094 | n36116 ;
  assign n40027 = n38496 & n40026 ;
  assign n40028 = ~n9343 & n36218 ;
  assign n40029 = x211 & n36108 ;
  assign n40030 = n40028 | n40029 ;
  assign n40031 = ( n7318 & ~n40027 ) | ( n7318 & n40030 ) | ( ~n40027 & n40030 ) ;
  assign n40032 = n40027 | n40031 ;
  assign n40033 = ( x1151 & n40025 ) | ( x1151 & n40032 ) | ( n40025 & n40032 ) ;
  assign n40034 = ~n40025 & n40033 ;
  assign n40035 = n11549 | n36026 ;
  assign n40036 = n36165 & ~n40035 ;
  assign n40037 = ~n7318 & n40036 ;
  assign n40038 = x219 & n37775 ;
  assign n40039 = n40037 | n40038 ;
  assign n40040 = x1151 | n40039 ;
  assign n40041 = ( x1151 & x1153 ) | ( x1151 & n40040 ) | ( x1153 & n40040 ) ;
  assign n40042 = ( x1152 & ~n40034 ) | ( x1152 & n40041 ) | ( ~n40034 & n40041 ) ;
  assign n40043 = n40042 ^ n40041 ^ 1'b0 ;
  assign n40044 = ( x1152 & n40042 ) | ( x1152 & ~n40043 ) | ( n40042 & ~n40043 ) ;
  assign n40045 = x230 & ~n40044 ;
  assign n40046 = ( x230 & n40024 ) | ( x230 & n40045 ) | ( n40024 & n40045 ) ;
  assign n40047 = ~x219 & n38507 ;
  assign n40048 = x219 & x1091 ;
  assign n40049 = ~n35980 & n40048 ;
  assign n40050 = n38473 | n40049 ;
  assign n40051 = n40047 | n40050 ;
  assign n40052 = x253 & n40051 ;
  assign n40053 = ~x211 & n38468 ;
  assign n40054 = x211 & n38473 ;
  assign n40055 = x219 & ~n40054 ;
  assign n40056 = ~n40053 & n40055 ;
  assign n40057 = x219 | n38484 ;
  assign n40058 = ~n40049 & n40057 ;
  assign n40059 = ~n40056 & n40058 ;
  assign n40060 = x253 | n40059 ;
  assign n40061 = ( n7318 & n40052 ) | ( n7318 & n40060 ) | ( n40052 & n40060 ) ;
  assign n40062 = ~n40052 & n40061 ;
  assign n40063 = n40053 | n40057 ;
  assign n40064 = n40047 & n40063 ;
  assign n40065 = x219 & n38468 ;
  assign n40066 = n7318 & ~n40065 ;
  assign n40067 = ~n40064 & n40066 ;
  assign n40068 = n38468 & n40067 ;
  assign n40069 = n40062 | n40068 ;
  assign n40070 = n40063 ^ n40057 ^ n40047 ;
  assign n40071 = x219 | n40070 ;
  assign n40072 = n7318 & ~n40071 ;
  assign n40073 = n38468 & n40072 ;
  assign n40074 = x1151 & ~n40073 ;
  assign n40075 = n38523 & ~n38544 ;
  assign n40076 = ~x211 & n38570 ;
  assign n40077 = n40075 & ~n40076 ;
  assign n40078 = n38538 & n38553 ;
  assign n40079 = n40077 & n40078 ;
  assign n40080 = x1153 & ~n40079 ;
  assign n40081 = x1153 | n38574 ;
  assign n40082 = x219 & n40081 ;
  assign n40083 = ~n40080 & n40082 ;
  assign n40084 = n38545 & n38600 ;
  assign n40085 = x1153 & ~n40084 ;
  assign n40086 = x1153 | n38631 ;
  assign n40087 = ~x219 & n40086 ;
  assign n40088 = ~n40085 & n40087 ;
  assign n40089 = ( x253 & n40083 ) | ( x253 & ~n40088 ) | ( n40083 & ~n40088 ) ;
  assign n40090 = ~n40083 & n40089 ;
  assign n40091 = n38515 & n38574 ;
  assign n40092 = ~x211 & n40091 ;
  assign n40093 = n38557 | n40092 ;
  assign n40094 = x1153 | n38529 ;
  assign n40095 = ( n38577 & n40093 ) | ( n38577 & n40094 ) | ( n40093 & n40094 ) ;
  assign n40096 = x219 & ~n40095 ;
  assign n40097 = ~x1153 & n38630 ;
  assign n40098 = x219 | n40097 ;
  assign n40099 = x1153 & n38647 ;
  assign n40100 = n40098 | n40099 ;
  assign n40101 = ~x253 & n40100 ;
  assign n40102 = ~n40096 & n40101 ;
  assign n40103 = ( ~n7318 & n40090 ) | ( ~n7318 & n40102 ) | ( n40090 & n40102 ) ;
  assign n40104 = ~n7318 & n40103 ;
  assign n40105 = ( n40062 & n40074 ) | ( n40062 & ~n40104 ) | ( n40074 & ~n40104 ) ;
  assign n40106 = ~n40062 & n40105 ;
  assign n40107 = n38537 & ~n38544 ;
  assign n40108 = x1153 | n40107 ;
  assign n40109 = n38556 & n40077 ;
  assign n40110 = n40108 & n40109 ;
  assign n40111 = ( x219 & n38523 ) | ( x219 & n40110 ) | ( n38523 & n40110 ) ;
  assign n40112 = n40111 ^ n40096 ^ 1'b0 ;
  assign n40113 = ( n40096 & n40111 ) | ( n40096 & n40112 ) | ( n40111 & n40112 ) ;
  assign n40114 = ( x253 & ~n40096 ) | ( x253 & n40113 ) | ( ~n40096 & n40113 ) ;
  assign n40115 = x219 & n38554 ;
  assign n40116 = ~n38595 & n40080 ;
  assign n40117 = n40115 & ~n40116 ;
  assign n40118 = n38600 | n40092 ;
  assign n40119 = n40047 & n40118 ;
  assign n40120 = ~n38654 & n40108 ;
  assign n40121 = n40119 & ~n40120 ;
  assign n40122 = ( x253 & n40117 ) | ( x253 & n40121 ) | ( n40117 & n40121 ) ;
  assign n40123 = n40121 ^ n40117 ^ 1'b0 ;
  assign n40124 = ( x253 & n40122 ) | ( x253 & n40123 ) | ( n40122 & n40123 ) ;
  assign n40125 = ( n7318 & n40114 ) | ( n7318 & ~n40124 ) | ( n40114 & ~n40124 ) ;
  assign n40126 = ~n7318 & n40125 ;
  assign n40127 = x1151 | n40126 ;
  assign n40128 = ~n40106 & n40127 ;
  assign n40129 = ( x1152 & n40069 ) | ( x1152 & n40128 ) | ( n40069 & n40128 ) ;
  assign n40130 = n40128 ^ n40069 ^ 1'b0 ;
  assign n40131 = ( x1152 & n40129 ) | ( x1152 & n40130 ) | ( n40129 & n40130 ) ;
  assign n40132 = x1151 | n40062 ;
  assign n40133 = x219 & n40095 ;
  assign n40134 = n38540 & n40133 ;
  assign n40135 = x1153 | n38617 ;
  assign n40136 = n38515 & n40135 ;
  assign n40137 = ~x219 & n38631 ;
  assign n40138 = n40136 & n40137 ;
  assign n40139 = ( x253 & ~n40134 ) | ( x253 & n40138 ) | ( ~n40134 & n40138 ) ;
  assign n40140 = n40134 | n40139 ;
  assign n40141 = n38595 | n40079 ;
  assign n40142 = x1091 | n38577 ;
  assign n40143 = ~x1153 & n40142 ;
  assign n40144 = ~x219 & n40107 ;
  assign n40145 = n40143 | n40144 ;
  assign n40146 = n40141 | n40145 ;
  assign n40147 = x253 & n40146 ;
  assign n40148 = ( n7318 & n40140 ) | ( n7318 & ~n40147 ) | ( n40140 & ~n40147 ) ;
  assign n40149 = ~n7318 & n40148 ;
  assign n40150 = ( ~x1152 & n40132 ) | ( ~x1152 & n40149 ) | ( n40132 & n40149 ) ;
  assign n40151 = ~x1152 & n40150 ;
  assign n40152 = n7318 ^ x253 ^ 1'b0 ;
  assign n40153 = x1153 & ~n38545 ;
  assign n40154 = n40047 & n40077 ;
  assign n40155 = ~n40153 & n40154 ;
  assign n40156 = n38587 | n40079 ;
  assign n40157 = x1153 & ~n40156 ;
  assign n40158 = x1153 | n38525 ;
  assign n40159 = ( x219 & n40157 ) | ( x219 & n40158 ) | ( n40157 & n40158 ) ;
  assign n40160 = ( n40155 & ~n40157 ) | ( n40155 & n40159 ) | ( ~n40157 & n40159 ) ;
  assign n40161 = ( x253 & ~n40152 ) | ( x253 & n40160 ) | ( ~n40152 & n40160 ) ;
  assign n40162 = ( n7318 & n40152 ) | ( n7318 & n40161 ) | ( n40152 & n40161 ) ;
  assign n40163 = n40100 & n40119 ;
  assign n40164 = n40133 | n40163 ;
  assign n40165 = n38515 & n40164 ;
  assign n40166 = ( x253 & ~n40162 ) | ( x253 & n40165 ) | ( ~n40162 & n40165 ) ;
  assign n40167 = ~n40162 & n40166 ;
  assign n40168 = ( n40062 & n40074 ) | ( n40062 & ~n40167 ) | ( n40074 & ~n40167 ) ;
  assign n40169 = ~n40062 & n40168 ;
  assign n40170 = ( n40131 & n40151 ) | ( n40131 & ~n40169 ) | ( n40151 & ~n40169 ) ;
  assign n40171 = n40170 ^ n40151 ^ 1'b0 ;
  assign n40172 = ( n40131 & n40170 ) | ( n40131 & ~n40171 ) | ( n40170 & ~n40171 ) ;
  assign n40173 = ( ~x268 & n38505 ) | ( ~x268 & n40172 ) | ( n38505 & n40172 ) ;
  assign n40174 = x268 & n40173 ;
  assign n40175 = x1091 & x1153 ;
  assign n40176 = n40037 & n40175 ;
  assign n40177 = x253 | x1091 ;
  assign n40178 = n7318 & n40177 ;
  assign n40179 = ~n40049 & n40178 ;
  assign n40180 = x219 & n40179 ;
  assign n40181 = x253 & ~x1091 ;
  assign n40182 = x1151 | n40181 ;
  assign n40183 = ( ~n40176 & n40180 ) | ( ~n40176 & n40182 ) | ( n40180 & n40182 ) ;
  assign n40184 = n40176 | n40183 ;
  assign n40185 = n11552 & ~n40017 ;
  assign n40186 = x1091 & ~n40185 ;
  assign n40187 = x253 | n40186 ;
  assign n40188 = x1153 | n38694 ;
  assign n40189 = x1153 & ~n38702 ;
  assign n40190 = n38496 & ~n40189 ;
  assign n40191 = n40188 & n40190 ;
  assign n40192 = x1091 & n40030 ;
  assign n40193 = ( x253 & n40191 ) | ( x253 & n40192 ) | ( n40191 & n40192 ) ;
  assign n40194 = n40192 ^ n40191 ^ 1'b0 ;
  assign n40195 = ( x253 & n40193 ) | ( x253 & n40194 ) | ( n40193 & n40194 ) ;
  assign n40196 = ( n7318 & n40187 ) | ( n7318 & ~n40195 ) | ( n40187 & ~n40195 ) ;
  assign n40197 = ~n7318 & n40196 ;
  assign n40198 = x211 & x1091 ;
  assign n40199 = x1091 & ~x1153 ;
  assign n40200 = x219 & n40199 ;
  assign n40201 = n40198 | n40200 ;
  assign n40202 = n40178 & ~n40201 ;
  assign n40203 = ( x1151 & n40197 ) | ( x1151 & ~n40202 ) | ( n40197 & ~n40202 ) ;
  assign n40204 = ~n40197 & n40203 ;
  assign n40205 = ( x1152 & n40184 ) | ( x1152 & ~n40204 ) | ( n40184 & ~n40204 ) ;
  assign n40206 = n40205 ^ n40184 ^ 1'b0 ;
  assign n40207 = ( x1152 & n40205 ) | ( x1152 & ~n40206 ) | ( n40205 & ~n40206 ) ;
  assign n40208 = x1091 & n36158 ;
  assign n40209 = n10075 | n38496 ;
  assign n40210 = n40181 | n40209 ;
  assign n40211 = n40208 | n40210 ;
  assign n40212 = n10075 & n38714 ;
  assign n40213 = ~n36158 & n40212 ;
  assign n40214 = x1153 | n38720 ;
  assign n40215 = x1091 & n37200 ;
  assign n40216 = ( ~x1091 & n40188 ) | ( ~x1091 & n40215 ) | ( n40188 & n40215 ) ;
  assign n40217 = n38496 & ~n40216 ;
  assign n40218 = n40214 & n40217 ;
  assign n40219 = ( x253 & n40213 ) | ( x253 & ~n40218 ) | ( n40213 & ~n40218 ) ;
  assign n40220 = ~n40213 & n40219 ;
  assign n40221 = x1091 & n36094 ;
  assign n40222 = ~n36527 & n40221 ;
  assign n40223 = n38496 & ~n40222 ;
  assign n40224 = n40223 ^ n40215 ^ 1'b0 ;
  assign n40225 = ( n40215 & n40223 ) | ( n40215 & n40224 ) | ( n40223 & n40224 ) ;
  assign n40226 = ( x253 & ~n40215 ) | ( x253 & n40225 ) | ( ~n40215 & n40225 ) ;
  assign n40227 = x211 & ~n38713 ;
  assign n40228 = ~n40208 & n40227 ;
  assign n40229 = ( ~n40220 & n40226 ) | ( ~n40220 & n40228 ) | ( n40226 & n40228 ) ;
  assign n40230 = ~n40220 & n40229 ;
  assign n40231 = ( n37457 & n40211 ) | ( n37457 & ~n40230 ) | ( n40211 & ~n40230 ) ;
  assign n40232 = ~n37457 & n40231 ;
  assign n40233 = ~x211 & x1091 ;
  assign n40234 = ~x219 & n40233 ;
  assign n40235 = n40179 & ~n40234 ;
  assign n40236 = n40016 & ~n40181 ;
  assign n40237 = n40199 | n40236 ;
  assign n40238 = n40018 & n40237 ;
  assign n40239 = ( n7318 & n40177 ) | ( n7318 & ~n40238 ) | ( n40177 & ~n40238 ) ;
  assign n40240 = ~n7318 & n40239 ;
  assign n40241 = ( x1151 & n40179 ) | ( x1151 & n40240 ) | ( n40179 & n40240 ) ;
  assign n40242 = n40240 ^ n40179 ^ 1'b0 ;
  assign n40243 = ( x1151 & n40241 ) | ( x1151 & n40242 ) | ( n40241 & n40242 ) ;
  assign n40244 = ( x1152 & n40235 ) | ( x1152 & ~n40243 ) | ( n40235 & ~n40243 ) ;
  assign n40245 = ~n40235 & n40244 ;
  assign n40246 = n40245 ^ n40232 ^ 1'b0 ;
  assign n40247 = ( n40232 & n40245 ) | ( n40232 & n40246 ) | ( n40245 & n40246 ) ;
  assign n40248 = ( n38506 & ~n40232 ) | ( n38506 & n40247 ) | ( ~n40232 & n40247 ) ;
  assign n40249 = ( x230 & n40207 ) | ( x230 & ~n40248 ) | ( n40207 & ~n40248 ) ;
  assign n40250 = n40249 ^ n40207 ^ 1'b0 ;
  assign n40251 = ( x230 & n40249 ) | ( x230 & ~n40250 ) | ( n40249 & ~n40250 ) ;
  assign n40252 = ( ~n40046 & n40174 ) | ( ~n40046 & n40251 ) | ( n40174 & n40251 ) ;
  assign n40253 = ~n40046 & n40252 ;
  assign n40268 = n35982 ^ x219 ^ 1'b0 ;
  assign n40269 = ( n35982 & n36451 ) | ( n35982 & ~n40268 ) | ( n36451 & ~n40268 ) ;
  assign n40270 = n7318 & n40269 ;
  assign n40271 = n10075 ^ n7318 ^ 1'b0 ;
  assign n40272 = ( n37623 & n40270 ) | ( n37623 & n40271 ) | ( n40270 & n40271 ) ;
  assign n40254 = ~x1154 & n36595 ;
  assign n40255 = ( n36106 & n36112 ) | ( n36106 & n36649 ) | ( n36112 & n36649 ) ;
  assign n40256 = ( ~x211 & x1154 ) | ( ~x211 & n40255 ) | ( x1154 & n40255 ) ;
  assign n40257 = x211 & n40256 ;
  assign n40258 = ( n36516 & ~n40254 ) | ( n36516 & n40257 ) | ( ~n40254 & n40257 ) ;
  assign n40259 = n40254 | n40258 ;
  assign n40260 = x219 & n40259 ;
  assign n40261 = ~x200 & x1154 ;
  assign n40262 = n10008 & ~n40261 ;
  assign n40263 = n36649 & ~n37309 ;
  assign n40264 = ( ~x219 & n40262 ) | ( ~x219 & n40263 ) | ( n40262 & n40263 ) ;
  assign n40265 = ~x219 & n40264 ;
  assign n40266 = n7318 | n40265 ;
  assign n40267 = n40260 | n40266 ;
  assign n40273 = ( x1152 & n40267 ) | ( x1152 & n40272 ) | ( n40267 & n40272 ) ;
  assign n40274 = ~n40272 & n40273 ;
  assign n40275 = ~n10075 & n36528 ;
  assign n40276 = x299 & n38496 ;
  assign n40277 = n40275 | n40276 ;
  assign n40278 = n36514 & n40277 ;
  assign n40279 = ( x1154 & n36650 ) | ( x1154 & n36680 ) | ( n36650 & n36680 ) ;
  assign n40280 = n10075 & n40279 ;
  assign n40281 = ( ~n7318 & n40278 ) | ( ~n7318 & n40280 ) | ( n40278 & n40280 ) ;
  assign n40282 = ~n7318 & n40281 ;
  assign n40283 = ( x1152 & n40270 ) | ( x1152 & ~n40282 ) | ( n40270 & ~n40282 ) ;
  assign n40284 = n40282 | n40283 ;
  assign n40285 = x230 & ~n40284 ;
  assign n40286 = ( x230 & n40274 ) | ( x230 & n40285 ) | ( n40274 & n40285 ) ;
  assign n40287 = x1154 & n40233 ;
  assign n40288 = n40048 | n40287 ;
  assign n40289 = n40259 & n40288 ;
  assign n40290 = x1091 & n35964 ;
  assign n40291 = n36106 & ~n36581 ;
  assign n40292 = n40290 & n40291 ;
  assign n40293 = x211 | n36645 ;
  assign n40294 = x1153 & ~n38718 ;
  assign n40295 = x1154 | n40294 ;
  assign n40296 = n40188 & ~n40295 ;
  assign n40297 = n40293 & n40296 ;
  assign n40298 = ( ~x219 & n40292 ) | ( ~x219 & n40297 ) | ( n40292 & n40297 ) ;
  assign n40299 = ~x219 & n40298 ;
  assign n40300 = ( x254 & n40289 ) | ( x254 & n40299 ) | ( n40289 & n40299 ) ;
  assign n40301 = n40299 ^ n40289 ^ 1'b0 ;
  assign n40302 = ( x254 & n40300 ) | ( x254 & n40301 ) | ( n40300 & n40301 ) ;
  assign n40303 = x1154 & ~n40016 ;
  assign n40304 = x219 & n36595 ;
  assign n40305 = ~n40303 & n40304 ;
  assign n40306 = ( x1091 & n40265 ) | ( x1091 & ~n40305 ) | ( n40265 & ~n40305 ) ;
  assign n40307 = ~n40265 & n40306 ;
  assign n40308 = ( x254 & ~n40302 ) | ( x254 & n40307 ) | ( ~n40302 & n40307 ) ;
  assign n40309 = ~n40302 & n40308 ;
  assign n40310 = x253 | n40309 ;
  assign n40311 = x1154 & n38522 ;
  assign n40312 = n40077 & n40311 ;
  assign n40313 = ~n40085 & n40312 ;
  assign n40314 = ~x1153 & n40110 ;
  assign n40315 = ( ~x1154 & n38631 ) | ( ~x1154 & n40314 ) | ( n38631 & n40314 ) ;
  assign n40316 = ~x1154 & n40315 ;
  assign n40317 = ( x254 & n40313 ) | ( x254 & ~n40316 ) | ( n40313 & ~n40316 ) ;
  assign n40318 = ~n40313 & n40317 ;
  assign n40319 = x211 & n38570 ;
  assign n40320 = n38515 & ~n40319 ;
  assign n40321 = ( ~x254 & x1153 ) | ( ~x254 & n40320 ) | ( x1153 & n40320 ) ;
  assign n40322 = ~x254 & n40321 ;
  assign n40323 = n38525 & n38556 ;
  assign n40324 = x1154 & n40323 ;
  assign n40325 = n40324 ^ n38630 ^ 1'b0 ;
  assign n40326 = ( n38630 & n40324 ) | ( n38630 & ~n40325 ) | ( n40324 & ~n40325 ) ;
  assign n40327 = ( n40322 & n40325 ) | ( n40322 & n40326 ) | ( n40325 & n40326 ) ;
  assign n40328 = ( ~x219 & n40318 ) | ( ~x219 & n40327 ) | ( n40318 & n40327 ) ;
  assign n40329 = ~x219 & n40328 ;
  assign n40331 = x1153 & ~n38574 ;
  assign n40330 = ~x1154 & n40158 ;
  assign n40332 = n40331 ^ n40330 ^ 1'b0 ;
  assign n40333 = ( x254 & ~n40330 ) | ( x254 & n40331 ) | ( ~n40330 & n40331 ) ;
  assign n40334 = ( x254 & ~n40332 ) | ( x254 & n40333 ) | ( ~n40332 & n40333 ) ;
  assign n40335 = x1154 & ~n40080 ;
  assign n40336 = ( n40156 & ~n40334 ) | ( n40156 & n40335 ) | ( ~n40334 & n40335 ) ;
  assign n40337 = n40336 ^ n40334 ^ 1'b0 ;
  assign n40338 = ( n40334 & ~n40336 ) | ( n40334 & n40337 ) | ( ~n40336 & n40337 ) ;
  assign n40339 = n40081 & n40323 ;
  assign n40340 = n35982 & ~n40339 ;
  assign n40341 = ~n38514 & n40340 ;
  assign n40342 = x1153 & n38557 ;
  assign n40343 = n35964 & ~n38516 ;
  assign n40344 = ~n40342 & n40343 ;
  assign n40345 = ( x254 & ~n40341 ) | ( x254 & n40344 ) | ( ~n40341 & n40344 ) ;
  assign n40346 = n40341 | n40345 ;
  assign n40347 = n38579 & n40094 ;
  assign n40348 = x1154 | n40347 ;
  assign n40349 = n38515 & n38577 ;
  assign n40350 = ( ~n40346 & n40348 ) | ( ~n40346 & n40349 ) | ( n40348 & n40349 ) ;
  assign n40351 = ~n40346 & n40350 ;
  assign n40352 = ( x219 & n40338 ) | ( x219 & n40351 ) | ( n40338 & n40351 ) ;
  assign n40353 = n40351 ^ n40338 ^ 1'b0 ;
  assign n40354 = ( x219 & n40352 ) | ( x219 & n40353 ) | ( n40352 & n40353 ) ;
  assign n40355 = ( x253 & n40329 ) | ( x253 & ~n40354 ) | ( n40329 & ~n40354 ) ;
  assign n40356 = ~n40329 & n40355 ;
  assign n40357 = ( n7318 & n40310 ) | ( n7318 & ~n40356 ) | ( n40310 & ~n40356 ) ;
  assign n40358 = ~n7318 & n40357 ;
  assign n40359 = n40063 | n40175 ;
  assign n40360 = x1091 & n36390 ;
  assign n40361 = x254 | n40360 ;
  assign n40362 = ( n40056 & n40359 ) | ( n40056 & ~n40361 ) | ( n40359 & ~n40361 ) ;
  assign n40363 = ~n40056 & n40362 ;
  assign n40368 = ( n38473 & n40056 ) | ( n38473 & n40065 ) | ( n40056 & n40065 ) ;
  assign n40364 = ~x219 & n38484 ;
  assign n40365 = n10075 & n40199 ;
  assign n40366 = ( x254 & n40360 ) | ( x254 & ~n40365 ) | ( n40360 & ~n40365 ) ;
  assign n40367 = ~n40360 & n40366 ;
  assign n40369 = ( ~n40364 & n40367 ) | ( ~n40364 & n40368 ) | ( n40367 & n40368 ) ;
  assign n40370 = ~n40368 & n40369 ;
  assign n40371 = x253 & ~n40370 ;
  assign n40372 = ~n40363 & n40371 ;
  assign n40373 = x253 & n7318 ;
  assign n40374 = x254 | x1091 ;
  assign n40375 = x1091 & ~n40269 ;
  assign n40376 = n7318 & ~n40375 ;
  assign n40377 = n40374 & n40376 ;
  assign n40378 = ( n7318 & n40234 ) | ( n7318 & n40377 ) | ( n40234 & n40377 ) ;
  assign n40379 = ( ~n40372 & n40373 ) | ( ~n40372 & n40378 ) | ( n40373 & n40378 ) ;
  assign n40380 = ~n40372 & n40379 ;
  assign n40381 = ( x1152 & n40358 ) | ( x1152 & ~n40380 ) | ( n40358 & ~n40380 ) ;
  assign n40382 = ~n40358 & n40381 ;
  assign n40383 = n40071 & n40363 ;
  assign n40384 = ~n40064 & n40370 ;
  assign n40385 = ( x253 & n40383 ) | ( x253 & ~n40384 ) | ( n40383 & ~n40384 ) ;
  assign n40386 = ~n40383 & n40385 ;
  assign n40387 = ( n40373 & n40377 ) | ( n40373 & ~n40386 ) | ( n40377 & ~n40386 ) ;
  assign n40388 = ~n40386 & n40387 ;
  assign n40389 = x1153 | n38688 ;
  assign n40390 = ~n40216 & n40389 ;
  assign n40391 = n38693 | n40390 ;
  assign n40392 = ~n40209 & n40391 ;
  assign n40393 = n38705 & n40217 ;
  assign n40394 = ( x1154 & n40392 ) | ( x1154 & ~n40393 ) | ( n40392 & ~n40393 ) ;
  assign n40395 = ~n40392 & n40394 ;
  assign n40396 = x1091 & ~n10075 ;
  assign n40397 = ~n36513 & n40396 ;
  assign n40398 = ( x1154 & ~n40395 ) | ( x1154 & n40397 ) | ( ~n40395 & n40397 ) ;
  assign n40399 = ~n40395 & n40398 ;
  assign n40400 = x1091 & ~x1154 ;
  assign n40401 = ~n36181 & n40400 ;
  assign n40402 = n40390 | n40401 ;
  assign n40403 = n10075 & n40402 ;
  assign n40404 = ( x254 & n40399 ) | ( x254 & ~n40403 ) | ( n40399 & ~n40403 ) ;
  assign n40405 = ~n40399 & n40404 ;
  assign n40406 = x1091 & n36528 ;
  assign n40407 = x1154 & ~n40406 ;
  assign n40408 = x211 & n40407 ;
  assign n40409 = n10074 & n40175 ;
  assign n40410 = x1154 | n40409 ;
  assign n40411 = x219 & n40410 ;
  assign n40412 = n36165 & n40199 ;
  assign n40413 = ( n35982 & n40215 ) | ( n35982 & ~n40412 ) | ( n40215 & ~n40412 ) ;
  assign n40414 = ~n40215 & n40413 ;
  assign n40415 = ( n40408 & n40411 ) | ( n40408 & ~n40414 ) | ( n40411 & ~n40414 ) ;
  assign n40416 = ~n40408 & n40415 ;
  assign n40417 = n38687 & n40199 ;
  assign n40418 = n40215 | n40417 ;
  assign n40419 = ~x211 & n40410 ;
  assign n40420 = ~n40407 & n40419 ;
  assign n40421 = x211 & n40295 ;
  assign n40422 = n40420 ^ n40418 ^ 1'b0 ;
  assign n40423 = ( ~n40418 & n40421 ) | ( ~n40418 & n40422 ) | ( n40421 & n40422 ) ;
  assign n40424 = ( n40418 & n40420 ) | ( n40418 & n40423 ) | ( n40420 & n40423 ) ;
  assign n40425 = ( ~x219 & n40416 ) | ( ~x219 & n40424 ) | ( n40416 & n40424 ) ;
  assign n40426 = n40416 ^ x219 ^ 1'b0 ;
  assign n40427 = ( n40416 & n40425 ) | ( n40416 & ~n40426 ) | ( n40425 & ~n40426 ) ;
  assign n40428 = ( ~x254 & n40405 ) | ( ~x254 & n40427 ) | ( n40405 & n40427 ) ;
  assign n40429 = n40405 ^ x254 ^ 1'b0 ;
  assign n40430 = ( n40405 & n40428 ) | ( n40405 & ~n40429 ) | ( n40428 & ~n40429 ) ;
  assign n40431 = x253 | n40430 ;
  assign n40432 = ~x1153 & n38538 ;
  assign n40433 = n40118 | n40432 ;
  assign n40434 = x1154 & ~n38537 ;
  assign n40435 = x219 | n40434 ;
  assign n40436 = n40433 & ~n40435 ;
  assign n40437 = n35982 & ~n38595 ;
  assign n40438 = n40078 | n40432 ;
  assign n40439 = ~x1154 & n38541 ;
  assign n40440 = n40438 | n40439 ;
  assign n40441 = ( x219 & n40437 ) | ( x219 & n40440 ) | ( n40437 & n40440 ) ;
  assign n40442 = ~n40437 & n40441 ;
  assign n40443 = ( x254 & n40436 ) | ( x254 & n40442 ) | ( n40436 & n40442 ) ;
  assign n40444 = n40442 ^ n40436 ^ 1'b0 ;
  assign n40445 = ( x254 & n40443 ) | ( x254 & n40444 ) | ( n40443 & n40444 ) ;
  assign n40446 = x219 & ~n40340 ;
  assign n40447 = n38558 & n40081 ;
  assign n40448 = n35964 & ~n40447 ;
  assign n40449 = n40348 & ~n40448 ;
  assign n40450 = n40446 & n40449 ;
  assign n40451 = n38522 & n38630 ;
  assign n40452 = n40135 & n40451 ;
  assign n40453 = n38515 & n38631 ;
  assign n40454 = x1154 & ~n40453 ;
  assign n40455 = ~n40452 & n40454 ;
  assign n40456 = n38523 ^ x1154 ^ 1'b0 ;
  assign n40457 = ( n38570 & ~n38651 ) | ( n38570 & n40456 ) | ( ~n38651 & n40456 ) ;
  assign n40458 = x211 | n40457 ;
  assign n40459 = ( ~x211 & x219 ) | ( ~x211 & n40458 ) | ( x219 & n40458 ) ;
  assign n40460 = x1154 | n40452 ;
  assign n40461 = ( n40455 & ~n40459 ) | ( n40455 & n40460 ) | ( ~n40459 & n40460 ) ;
  assign n40462 = ~n40455 & n40461 ;
  assign n40463 = ( x254 & ~n40450 ) | ( x254 & n40462 ) | ( ~n40450 & n40462 ) ;
  assign n40464 = n40450 | n40463 ;
  assign n40465 = x253 & ~n40464 ;
  assign n40466 = ( x253 & n40445 ) | ( x253 & n40465 ) | ( n40445 & n40465 ) ;
  assign n40467 = ( n7318 & n40431 ) | ( n7318 & ~n40466 ) | ( n40431 & ~n40466 ) ;
  assign n40468 = ~n7318 & n40467 ;
  assign n40469 = ( x1152 & ~n40388 ) | ( x1152 & n40468 ) | ( ~n40388 & n40468 ) ;
  assign n40470 = n40388 | n40469 ;
  assign n40471 = ( n38506 & n40382 ) | ( n38506 & n40470 ) | ( n40382 & n40470 ) ;
  assign n40472 = ~n40382 & n40471 ;
  assign n40473 = x1152 | n40377 ;
  assign n40474 = ~n7318 & n40430 ;
  assign n40475 = n40473 | n40474 ;
  assign n40476 = x1152 & ~n40378 ;
  assign n40477 = ~n7318 & n40309 ;
  assign n40478 = ( n38506 & n40476 ) | ( n38506 & ~n40477 ) | ( n40476 & ~n40477 ) ;
  assign n40479 = n40478 ^ n40476 ^ 1'b0 ;
  assign n40480 = ( n38506 & n40478 ) | ( n38506 & ~n40479 ) | ( n40478 & ~n40479 ) ;
  assign n40481 = ( x230 & n40475 ) | ( x230 & ~n40480 ) | ( n40475 & ~n40480 ) ;
  assign n40482 = n40481 ^ n40475 ^ 1'b0 ;
  assign n40483 = ( x230 & n40481 ) | ( x230 & ~n40482 ) | ( n40481 & ~n40482 ) ;
  assign n40484 = ( ~n40286 & n40472 ) | ( ~n40286 & n40483 ) | ( n40472 & n40483 ) ;
  assign n40485 = ~n40286 & n40484 ;
  assign n40486 = x1036 ^ x200 ^ 1'b0 ;
  assign n40487 = ( x1036 & x1049 ) | ( x1036 & ~n40486 ) | ( x1049 & ~n40486 ) ;
  assign n40488 = n39967 ^ x255 ^ 1'b0 ;
  assign n40489 = ( x255 & n40487 ) | ( x255 & n40488 ) | ( n40487 & n40488 ) ;
  assign n40490 = x1048 ^ x200 ^ 1'b0 ;
  assign n40491 = ( x1048 & x1070 ) | ( x1048 & n40490 ) | ( x1070 & n40490 ) ;
  assign n40492 = n39967 ^ x256 ^ 1'b0 ;
  assign n40493 = ( x256 & n40491 ) | ( x256 & n40492 ) | ( n40491 & n40492 ) ;
  assign n40494 = x1065 ^ x200 ^ 1'b0 ;
  assign n40495 = ( x1065 & x1084 ) | ( x1065 & ~n40494 ) | ( x1084 & ~n40494 ) ;
  assign n40496 = n39967 ^ x257 ^ 1'b0 ;
  assign n40497 = ( x257 & n40495 ) | ( x257 & n40496 ) | ( n40495 & n40496 ) ;
  assign n40498 = x1062 ^ x200 ^ 1'b0 ;
  assign n40499 = ( x1062 & x1072 ) | ( x1062 & ~n40498 ) | ( x1072 & ~n40498 ) ;
  assign n40500 = n39967 ^ x258 ^ 1'b0 ;
  assign n40501 = ( x258 & n40499 ) | ( x258 & n40500 ) | ( n40499 & n40500 ) ;
  assign n40502 = x1059 ^ x200 ^ 1'b0 ;
  assign n40503 = ( x1059 & x1069 ) | ( x1059 & n40502 ) | ( x1069 & n40502 ) ;
  assign n40504 = n39967 ^ x259 ^ 1'b0 ;
  assign n40505 = ( x259 & n40503 ) | ( x259 & n40504 ) | ( n40503 & n40504 ) ;
  assign n40506 = ~x200 & x1044 ;
  assign n40507 = x200 & x1067 ;
  assign n40508 = ( x199 & ~n40506 ) | ( x199 & n40507 ) | ( ~n40506 & n40507 ) ;
  assign n40509 = n40506 | n40508 ;
  assign n40510 = n39967 ^ x260 ^ 1'b0 ;
  assign n40511 = ( x260 & n40509 ) | ( x260 & n40510 ) | ( n40509 & n40510 ) ;
  assign n40512 = ~x200 & x1037 ;
  assign n40513 = x200 & x1040 ;
  assign n40514 = ( x199 & ~n40512 ) | ( x199 & n40513 ) | ( ~n40512 & n40513 ) ;
  assign n40515 = n40512 | n40514 ;
  assign n40516 = n39967 ^ x261 ^ 1'b0 ;
  assign n40517 = ( x261 & n40515 ) | ( x261 & n40516 ) | ( n40515 & n40516 ) ;
  assign n40518 = x123 & x262 ;
  assign n40519 = x123 | x1142 ;
  assign n40520 = ( x228 & n40518 ) | ( x228 & n40519 ) | ( n40518 & n40519 ) ;
  assign n40521 = ~n40518 & n40520 ;
  assign n40522 = x1093 & x1142 ;
  assign n40523 = x262 | x1093 ;
  assign n40524 = ~n40522 & n40523 ;
  assign n40525 = ( x228 & ~n40521 ) | ( x228 & n40524 ) | ( ~n40521 & n40524 ) ;
  assign n40526 = ~n40521 & n40525 ;
  assign n40527 = n7318 & ~n40526 ;
  assign n40528 = x228 ^ x123 ^ 1'b0 ;
  assign n40529 = ( ~x123 & x1093 ) | ( ~x123 & n40528 ) | ( x1093 & n40528 ) ;
  assign n40530 = ~n37261 & n40529 ;
  assign n40531 = n40527 & ~n40530 ;
  assign n40532 = x262 | n40529 ;
  assign n40533 = ~n38258 & n40532 ;
  assign n40534 = x199 & n40529 ;
  assign n40535 = n36000 & ~n40534 ;
  assign n40536 = n40533 & ~n40535 ;
  assign n40537 = n40526 | n40536 ;
  assign n40538 = x207 | n40532 ;
  assign n40539 = ~x208 & n40538 ;
  assign n40540 = ( n38258 & n40537 ) | ( n38258 & n40539 ) | ( n40537 & n40539 ) ;
  assign n40541 = n40537 & n40540 ;
  assign n40542 = n37387 & n40529 ;
  assign n40543 = ( x299 & n40526 ) | ( x299 & ~n40542 ) | ( n40526 & ~n40542 ) ;
  assign n40544 = n40542 | n40543 ;
  assign n40545 = x299 & ~n40533 ;
  assign n40546 = x208 & ~n40545 ;
  assign n40547 = n40544 & n40546 ;
  assign n40548 = ( x57 & n5193 ) | ( x57 & ~n40547 ) | ( n5193 & ~n40547 ) ;
  assign n40549 = n40547 | n40548 ;
  assign n40550 = ( ~n40531 & n40541 ) | ( ~n40531 & n40549 ) | ( n40541 & n40549 ) ;
  assign n40551 = ~n40531 & n40550 ;
  assign n40552 = n36097 & ~n36102 ;
  assign n40553 = x1156 | n40552 ;
  assign n40554 = ( n36317 & n36503 ) | ( n36317 & n40553 ) | ( n36503 & n40553 ) ;
  assign n40555 = ~n36317 & n40554 ;
  assign n40556 = ( x219 & ~x1156 ) | ( x219 & n37892 ) | ( ~x1156 & n37892 ) ;
  assign n40557 = n40556 ^ n40555 ^ 1'b0 ;
  assign n40558 = ( n40555 & n40556 ) | ( n40555 & n40557 ) | ( n40556 & n40557 ) ;
  assign n40559 = ( n7318 & ~n40555 ) | ( n7318 & n40558 ) | ( ~n40555 & n40558 ) ;
  assign n40560 = ~n36101 & n37012 ;
  assign n40561 = n36532 | n40560 ;
  assign n40562 = x211 | n40561 ;
  assign n40563 = ( ~x211 & x219 ) | ( ~x211 & n40562 ) | ( x219 & n40562 ) ;
  assign n40564 = n36021 | n40555 ;
  assign n40565 = x211 & n40564 ;
  assign n40566 = ( ~n40559 & n40563 ) | ( ~n40559 & n40565 ) | ( n40563 & n40565 ) ;
  assign n40567 = ~n40559 & n40566 ;
  assign n40568 = x219 & ~n35960 ;
  assign n40569 = x219 | n35961 ;
  assign n40570 = n35982 | n40569 ;
  assign n40571 = ~n40568 & n40570 ;
  assign n40572 = n7318 & n40571 ;
  assign n40573 = ( x230 & n40567 ) | ( x230 & ~n40572 ) | ( n40567 & ~n40572 ) ;
  assign n40574 = ~n40567 & n40573 ;
  assign n40575 = x211 & ~n38468 ;
  assign n40576 = n35961 | n40287 ;
  assign n40577 = ~n40575 & n40576 ;
  assign n40578 = n40057 | n40577 ;
  assign n40579 = x263 & ~n40056 ;
  assign n40580 = n40578 & n40579 ;
  assign n40581 = n40400 ^ x211 ^ 1'b0 ;
  assign n40582 = ( ~x1155 & n40400 ) | ( ~x1155 & n40581 ) | ( n40400 & n40581 ) ;
  assign n40583 = ~n40575 & n40582 ;
  assign n40584 = ( ~x219 & n38484 ) | ( ~x219 & n40583 ) | ( n38484 & n40583 ) ;
  assign n40585 = ~x219 & n40584 ;
  assign n40586 = x263 | n40368 ;
  assign n40587 = ( ~n40580 & n40585 ) | ( ~n40580 & n40586 ) | ( n40585 & n40586 ) ;
  assign n40588 = ~n40580 & n40587 ;
  assign n40589 = x1091 & n40568 ;
  assign n40590 = ( n38459 & n40588 ) | ( n38459 & ~n40589 ) | ( n40588 & ~n40589 ) ;
  assign n40591 = ~n40588 & n40590 ;
  assign n40592 = n40571 ^ x1091 ^ 1'b0 ;
  assign n40593 = ( x263 & ~n40571 ) | ( x263 & n40592 ) | ( ~n40571 & n40592 ) ;
  assign n40594 = n38459 | n40593 ;
  assign n40595 = ( n7318 & n40591 ) | ( n7318 & n40594 ) | ( n40591 & n40594 ) ;
  assign n40596 = ~n40591 & n40595 ;
  assign n40597 = ~n38570 & n38654 ;
  assign n40598 = x1155 & ~n38600 ;
  assign n40599 = x1154 | n40598 ;
  assign n40600 = x1155 & ~n38554 ;
  assign n40601 = x1154 | n40600 ;
  assign n40602 = n38538 & ~n40601 ;
  assign n40603 = ( n40597 & ~n40599 ) | ( n40597 & n40602 ) | ( ~n40599 & n40602 ) ;
  assign n40604 = x1156 & ~n40603 ;
  assign n40605 = x1155 & ~n38631 ;
  assign n40606 = x1154 & ~n40605 ;
  assign n40607 = n38545 & n40606 ;
  assign n40608 = n40604 & ~n40607 ;
  assign n40609 = x1155 | n40142 ;
  assign n40610 = n38630 | n40609 ;
  assign n40611 = n40610 ^ n40599 ^ 1'b0 ;
  assign n40612 = ( n40599 & n40610 ) | ( n40599 & n40611 ) | ( n40610 & n40611 ) ;
  assign n40613 = ( x1156 & ~n40599 ) | ( x1156 & n40612 ) | ( ~n40599 & n40612 ) ;
  assign n40614 = n40075 & n40606 ;
  assign n40615 = n40613 | n40614 ;
  assign n40616 = ( x211 & n40608 ) | ( x211 & n40615 ) | ( n40608 & n40615 ) ;
  assign n40617 = ~n40608 & n40616 ;
  assign n40618 = n38651 & n40606 ;
  assign n40619 = n38520 & n40618 ;
  assign n40620 = ( ~n40602 & n40604 ) | ( ~n40602 & n40619 ) | ( n40604 & n40619 ) ;
  assign n40621 = ~n40619 & n40620 ;
  assign n40622 = ~n40601 & n40609 ;
  assign n40623 = n40618 | n40622 ;
  assign n40624 = n40613 | n40623 ;
  assign n40625 = ( x211 & ~n40621 ) | ( x211 & n40624 ) | ( ~n40621 & n40624 ) ;
  assign n40626 = ~x211 & n40625 ;
  assign n40627 = ( x219 & ~n40617 ) | ( x219 & n40626 ) | ( ~n40617 & n40626 ) ;
  assign n40628 = n40617 | n40627 ;
  assign n40629 = x1154 & n38525 ;
  assign n40630 = x1155 & ~n38553 ;
  assign n40631 = n40629 & ~n40630 ;
  assign n40632 = n40622 | n40631 ;
  assign n40633 = ~x1156 & n40632 ;
  assign n40634 = ~x1154 & n38577 ;
  assign n40635 = n38587 | n40634 ;
  assign n40636 = ( x219 & n40568 ) | ( x219 & n40630 ) | ( n40568 & n40630 ) ;
  assign n40637 = ( x219 & ~n40635 ) | ( x219 & n40636 ) | ( ~n40635 & n40636 ) ;
  assign n40638 = n38522 & n40631 ;
  assign n40639 = n40602 | n40638 ;
  assign n40640 = n35969 & n40639 ;
  assign n40641 = ( n40633 & n40637 ) | ( n40633 & ~n40640 ) | ( n40637 & ~n40640 ) ;
  assign n40642 = ~n40633 & n40641 ;
  assign n40643 = ( x263 & n40628 ) | ( x263 & ~n40642 ) | ( n40628 & ~n40642 ) ;
  assign n40644 = ~x263 & n40643 ;
  assign n40645 = x1154 | n38619 ;
  assign n40646 = n38512 & n38644 ;
  assign n40647 = x1155 & n40646 ;
  assign n40648 = n40645 | n40647 ;
  assign n40649 = n40453 | n40648 ;
  assign n40650 = x1154 & ~n38648 ;
  assign n40651 = ~n38672 & n40650 ;
  assign n40652 = x1156 & ~n40651 ;
  assign n40653 = n40649 & n40652 ;
  assign n40654 = x1156 | n40434 ;
  assign n40655 = n40651 | n40654 ;
  assign n40656 = n40648 & ~n40655 ;
  assign n40657 = ( x211 & ~n40653 ) | ( x211 & n40656 ) | ( ~n40653 & n40656 ) ;
  assign n40658 = n40653 | n40657 ;
  assign n40659 = ~n38572 & n40650 ;
  assign n40660 = ~x1156 & n40655 ;
  assign n40661 = x1155 & n40451 ;
  assign n40662 = ( n40645 & ~n40660 ) | ( n40645 & n40661 ) | ( ~n40660 & n40661 ) ;
  assign n40663 = ~n40660 & n40662 ;
  assign n40664 = n40663 ^ x1156 ^ 1'b0 ;
  assign n40665 = ( ~x1156 & n40453 ) | ( ~x1156 & n40664 ) | ( n40453 & n40664 ) ;
  assign n40666 = ( x1156 & n40663 ) | ( x1156 & n40665 ) | ( n40663 & n40665 ) ;
  assign n40667 = x211 & ~n40666 ;
  assign n40668 = ( x211 & n40659 ) | ( x211 & n40667 ) | ( n40659 & n40667 ) ;
  assign n40669 = ( x219 & n40658 ) | ( x219 & ~n40668 ) | ( n40658 & ~n40668 ) ;
  assign n40670 = ~x219 & n40669 ;
  assign n40671 = n38578 | n38591 ;
  assign n40672 = ( x1154 & n38557 ) | ( x1154 & n40456 ) | ( n38557 & n40456 ) ;
  assign n40673 = n40671 & n40672 ;
  assign n40674 = n35969 & ~n40673 ;
  assign n40675 = n38512 & n40673 ;
  assign n40676 = x1156 | n40675 ;
  assign n40679 = x1155 & ~n40323 ;
  assign n40680 = x1154 | n40679 ;
  assign n40681 = x1155 | n40091 ;
  assign n40682 = ~n40680 & n40681 ;
  assign n40677 = x1154 & n40671 ;
  assign n40678 = n35960 & ~n40677 ;
  assign n40683 = n40682 ^ n40678 ^ 1'b0 ;
  assign n40684 = ( x219 & ~n40678 ) | ( x219 & n40682 ) | ( ~n40678 & n40682 ) ;
  assign n40685 = ( x219 & ~n40683 ) | ( x219 & n40684 ) | ( ~n40683 & n40684 ) ;
  assign n40686 = ( n40674 & n40676 ) | ( n40674 & n40685 ) | ( n40676 & n40685 ) ;
  assign n40687 = ~n40674 & n40686 ;
  assign n40688 = ( x263 & n40670 ) | ( x263 & ~n40687 ) | ( n40670 & ~n40687 ) ;
  assign n40689 = ~n40670 & n40688 ;
  assign n40690 = ( n38459 & n40644 ) | ( n38459 & ~n40689 ) | ( n40644 & ~n40689 ) ;
  assign n40691 = ~n40644 & n40690 ;
  assign n40692 = ~x1154 & n36099 ;
  assign n40693 = n37309 | n40692 ;
  assign n40694 = x1154 & ~n36098 ;
  assign n40695 = x1156 & ~n40694 ;
  assign n40696 = x299 | n40695 ;
  assign n40697 = x1156 & ~n40696 ;
  assign n40698 = ( x1156 & n40693 ) | ( x1156 & n40697 ) | ( n40693 & n40697 ) ;
  assign n40699 = n36096 | n36532 ;
  assign n40700 = ~n40696 & n40699 ;
  assign n40701 = ( x219 & n40698 ) | ( x219 & ~n40700 ) | ( n40698 & ~n40700 ) ;
  assign n40702 = ~n40698 & n40701 ;
  assign n40703 = n36106 & ~n36157 ;
  assign n40704 = x1154 & ~n40703 ;
  assign n40705 = ~x1154 & n36168 ;
  assign n40706 = ( n36144 & n36167 ) | ( n36144 & n40705 ) | ( n36167 & n40705 ) ;
  assign n40707 = ( x1156 & n40704 ) | ( x1156 & ~n40706 ) | ( n40704 & ~n40706 ) ;
  assign n40708 = ~n40704 & n40707 ;
  assign n40709 = n38694 | n40400 ;
  assign n40710 = ~n36182 & n40709 ;
  assign n40711 = ~x1156 & n40710 ;
  assign n40712 = ( x211 & n40708 ) | ( x211 & ~n40711 ) | ( n40708 & ~n40711 ) ;
  assign n40713 = ~n40708 & n40712 ;
  assign n40714 = ( ~x211 & n36532 ) | ( ~x211 & n40560 ) | ( n36532 & n40560 ) ;
  assign n40715 = ~x211 & n40714 ;
  assign n40716 = ( x219 & ~n40713 ) | ( x219 & n40715 ) | ( ~n40713 & n40715 ) ;
  assign n40717 = n40713 | n40716 ;
  assign n40718 = x263 & x1091 ;
  assign n40719 = ( n40702 & n40717 ) | ( n40702 & n40718 ) | ( n40717 & n40718 ) ;
  assign n40720 = ~n40702 & n40719 ;
  assign n40721 = x1155 & ~n36646 ;
  assign n40722 = n38702 & ~n40721 ;
  assign n40723 = ~x1154 & n38693 ;
  assign n40724 = n40722 | n40723 ;
  assign n40725 = n38713 | n40724 ;
  assign n40726 = n35969 & n40725 ;
  assign n40727 = x1156 | n36096 ;
  assign n40728 = x219 & ~n40709 ;
  assign n40729 = ( x219 & n40727 ) | ( x219 & n40728 ) | ( n40727 & n40728 ) ;
  assign n40730 = x1091 & n35960 ;
  assign n40731 = ( x299 & x1154 ) | ( x299 & n40694 ) | ( x1154 & n40694 ) ;
  assign n40732 = ( n40705 & n40730 ) | ( n40705 & ~n40731 ) | ( n40730 & ~n40731 ) ;
  assign n40733 = ~n40705 & n40732 ;
  assign n40734 = ( n40726 & n40729 ) | ( n40726 & ~n40733 ) | ( n40729 & ~n40733 ) ;
  assign n40735 = ~n40726 & n40734 ;
  assign n40736 = ~n36106 & n36502 ;
  assign n40737 = ( n36182 & n40198 ) | ( n36182 & ~n40736 ) | ( n40198 & ~n40736 ) ;
  assign n40738 = ~n36182 & n40737 ;
  assign n40739 = ~x211 & n40724 ;
  assign n40740 = ( x1156 & n40738 ) | ( x1156 & n40739 ) | ( n40738 & n40739 ) ;
  assign n40741 = n40739 ^ n40738 ^ 1'b0 ;
  assign n40742 = ( x1156 & n40740 ) | ( x1156 & n40741 ) | ( n40740 & n40741 ) ;
  assign n40743 = n40233 & ~n40699 ;
  assign n40744 = x211 & n40710 ;
  assign n40745 = n40743 | n40744 ;
  assign n40746 = n40745 ^ x1156 ^ 1'b0 ;
  assign n40747 = ( x1156 & n40745 ) | ( x1156 & n40746 ) | ( n40745 & n40746 ) ;
  assign n40748 = ( x219 & ~x1156 ) | ( x219 & n40747 ) | ( ~x1156 & n40747 ) ;
  assign n40749 = ( ~n40735 & n40742 ) | ( ~n40735 & n40748 ) | ( n40742 & n40748 ) ;
  assign n40750 = ~n40735 & n40749 ;
  assign n40751 = ( x263 & ~n40720 ) | ( x263 & n40750 ) | ( ~n40720 & n40750 ) ;
  assign n40752 = ~n40720 & n40751 ;
  assign n40753 = n38459 | n40752 ;
  assign n40754 = ( n7318 & ~n40691 ) | ( n7318 & n40753 ) | ( ~n40691 & n40753 ) ;
  assign n40755 = ~n7318 & n40754 ;
  assign n40756 = ( n38506 & n40596 ) | ( n38506 & ~n40755 ) | ( n40596 & ~n40755 ) ;
  assign n40757 = ~n40596 & n40756 ;
  assign n40758 = n7318 & n40593 ;
  assign n40759 = n38506 | n40758 ;
  assign n40760 = ~n7318 & n40752 ;
  assign n40761 = ( ~x230 & n40759 ) | ( ~x230 & n40760 ) | ( n40759 & n40760 ) ;
  assign n40762 = ~x230 & n40761 ;
  assign n40763 = ( n40574 & ~n40757 ) | ( n40574 & n40762 ) | ( ~n40757 & n40762 ) ;
  assign n40764 = n40757 ^ n40574 ^ 1'b0 ;
  assign n40765 = ( n40574 & n40763 ) | ( n40574 & ~n40764 ) | ( n40763 & ~n40764 ) ;
  assign n40766 = ~x211 & x1141 ;
  assign n40767 = x211 & x1142 ;
  assign n40768 = x219 | n40767 ;
  assign n40769 = ( ~n37073 & n40766 ) | ( ~n37073 & n40768 ) | ( n40766 & n40768 ) ;
  assign n40770 = ~n37073 & n40769 ;
  assign n40771 = ( x230 & n38767 ) | ( x230 & n40770 ) | ( n38767 & n40770 ) ;
  assign n40772 = ~x199 & x1141 ;
  assign n40773 = n37162 | n40772 ;
  assign n40774 = ~n36002 & n40773 ;
  assign n40775 = n40774 ^ n15098 ^ 1'b0 ;
  assign n40776 = ( n15098 & n40774 ) | ( n15098 & ~n40775 ) | ( n40774 & ~n40775 ) ;
  assign n40777 = ( n40771 & n40775 ) | ( n40771 & n40776 ) | ( n40775 & n40776 ) ;
  assign n40778 = ~x796 & n38479 ;
  assign n40779 = x1091 | n40778 ;
  assign n40780 = n38479 & ~n40779 ;
  assign n40781 = ( x264 & n40779 ) | ( x264 & ~n40780 ) | ( n40779 & ~n40780 ) ;
  assign n40782 = x1091 & x1141 ;
  assign n40783 = n40781 & ~n40782 ;
  assign n40784 = x211 | n40783 ;
  assign n40785 = x1091 & x1142 ;
  assign n40786 = n40781 & ~n40785 ;
  assign n40787 = x211 & ~n40786 ;
  assign n40788 = ( x219 & n40784 ) | ( x219 & ~n40787 ) | ( n40784 & ~n40787 ) ;
  assign n40789 = ~x219 & n40788 ;
  assign n40790 = ~x796 & n38462 ;
  assign n40791 = x1091 | n40790 ;
  assign n40792 = n38462 & ~n40791 ;
  assign n40793 = ( x264 & n40791 ) | ( x264 & ~n40792 ) | ( n40791 & ~n40792 ) ;
  assign n40794 = x219 & ~n40233 ;
  assign n40795 = n37073 | n40794 ;
  assign n40796 = n40793 & n40795 ;
  assign n40797 = ( n15098 & n40789 ) | ( n15098 & ~n40796 ) | ( n40789 & ~n40796 ) ;
  assign n40798 = ~n40789 & n40797 ;
  assign n40799 = x200 | n40783 ;
  assign n40800 = x200 & ~n40786 ;
  assign n40801 = ( x199 & n40799 ) | ( x199 & ~n40800 ) | ( n40799 & ~n40800 ) ;
  assign n40802 = ~x199 & n40801 ;
  assign n40803 = n40793 ^ n15098 ^ 1'b0 ;
  assign n40804 = x1091 & x1143 ;
  assign n40805 = ~x200 & n40804 ;
  assign n40806 = x199 & ~n40805 ;
  assign n40807 = ( n40793 & ~n40803 ) | ( n40793 & n40806 ) | ( ~n40803 & n40806 ) ;
  assign n40808 = ( n15098 & n40803 ) | ( n15098 & n40807 ) | ( n40803 & n40807 ) ;
  assign n40809 = ( ~n40798 & n40802 ) | ( ~n40798 & n40808 ) | ( n40802 & n40808 ) ;
  assign n40810 = ~n40798 & n40809 ;
  assign n40811 = ( x230 & ~n40777 ) | ( x230 & n40810 ) | ( ~n40777 & n40810 ) ;
  assign n40812 = ~n40777 & n40811 ;
  assign n40813 = ~x211 & x1142 ;
  assign n40814 = x219 | n36053 ;
  assign n40815 = ( ~n38434 & n40813 ) | ( ~n38434 & n40814 ) | ( n40813 & n40814 ) ;
  assign n40816 = ~n38434 & n40815 ;
  assign n40817 = ( x230 & n38767 ) | ( x230 & n40816 ) | ( n38767 & n40816 ) ;
  assign n40818 = n36001 | n38366 ;
  assign n40819 = ~n35996 & n40818 ;
  assign n40820 = n40819 ^ n15098 ^ 1'b0 ;
  assign n40821 = ( n15098 & n40819 ) | ( n15098 & ~n40820 ) | ( n40819 & ~n40820 ) ;
  assign n40822 = ( n40817 & n40820 ) | ( n40817 & n40821 ) | ( n40820 & n40821 ) ;
  assign n40823 = ~x819 & n38479 ;
  assign n40824 = x1091 | n40823 ;
  assign n40825 = n38479 & ~n40824 ;
  assign n40826 = ( x265 & n40824 ) | ( x265 & ~n40825 ) | ( n40824 & ~n40825 ) ;
  assign n40827 = ~n40785 & n40826 ;
  assign n40828 = x211 | n40827 ;
  assign n40829 = ~n40804 & n40826 ;
  assign n40830 = x211 & ~n40829 ;
  assign n40831 = ( x219 & n40828 ) | ( x219 & ~n40830 ) | ( n40828 & ~n40830 ) ;
  assign n40832 = ~x219 & n40831 ;
  assign n40833 = ~x819 & n38462 ;
  assign n40834 = x1091 | n40833 ;
  assign n40835 = n38462 & ~n40834 ;
  assign n40836 = ( x265 & n40834 ) | ( x265 & ~n40835 ) | ( n40834 & ~n40835 ) ;
  assign n40837 = n38434 | n40794 ;
  assign n40838 = n40836 & n40837 ;
  assign n40839 = ( n15098 & n40832 ) | ( n15098 & ~n40838 ) | ( n40832 & ~n40838 ) ;
  assign n40840 = ~n40832 & n40839 ;
  assign n40841 = x200 | n40827 ;
  assign n40842 = x200 & ~n40829 ;
  assign n40843 = ( x199 & n40841 ) | ( x199 & ~n40842 ) | ( n40841 & ~n40842 ) ;
  assign n40844 = ~x199 & n40843 ;
  assign n40845 = x1091 & x1144 ;
  assign n40846 = ~x200 & n40845 ;
  assign n40847 = x199 & ~n40846 ;
  assign n40848 = n40836 & n40847 ;
  assign n40849 = n15098 | n40848 ;
  assign n40850 = ( ~n40840 & n40844 ) | ( ~n40840 & n40849 ) | ( n40844 & n40849 ) ;
  assign n40851 = ~n40840 & n40850 ;
  assign n40852 = ( x230 & ~n40822 ) | ( x230 & n40851 ) | ( ~n40822 & n40851 ) ;
  assign n40853 = ~n40822 & n40852 ;
  assign n40854 = ~x211 & x1136 ;
  assign n40855 = x219 & ~n40854 ;
  assign n40856 = x211 & ~x1135 ;
  assign n40857 = n40855 | n40856 ;
  assign n40858 = n9343 & ~n40857 ;
  assign n40859 = n7318 & n40858 ;
  assign n40860 = x199 & x1136 ;
  assign n40861 = x200 | n40860 ;
  assign n40862 = ~x199 & x1135 ;
  assign n40863 = x200 & ~n40862 ;
  assign n40864 = x299 | n40863 ;
  assign n40865 = n40861 & ~n40864 ;
  assign n40866 = x299 & n40858 ;
  assign n40867 = ( ~n7318 & n40865 ) | ( ~n7318 & n40866 ) | ( n40865 & n40866 ) ;
  assign n40868 = ~n7318 & n40867 ;
  assign n40869 = ( x230 & n40859 ) | ( x230 & ~n40868 ) | ( n40859 & ~n40868 ) ;
  assign n40870 = ~n40859 & n40869 ;
  assign n40871 = x266 | n38462 ;
  assign n40872 = ~x948 & n38462 ;
  assign n40873 = ( x1091 & n40871 ) | ( x1091 & ~n40872 ) | ( n40871 & ~n40872 ) ;
  assign n40874 = ~x1091 & n40873 ;
  assign n40875 = n40794 | n40855 ;
  assign n40876 = ~n40874 & n40875 ;
  assign n40877 = n15098 & ~n40876 ;
  assign n40878 = n40877 ^ x230 ^ 1'b0 ;
  assign n40879 = ~x948 & n38479 ;
  assign n40880 = x266 | n38479 ;
  assign n40881 = ( x1091 & ~n40879 ) | ( x1091 & n40880 ) | ( ~n40879 & n40880 ) ;
  assign n40882 = ~x1091 & n40881 ;
  assign n40883 = x219 | n40882 ;
  assign n40884 = x1135 & n40198 ;
  assign n40885 = n40883 | n40884 ;
  assign n40886 = ( n40877 & ~n40878 ) | ( n40877 & n40885 ) | ( ~n40878 & n40885 ) ;
  assign n40887 = ( x230 & n40878 ) | ( x230 & n40886 ) | ( n40878 & n40886 ) ;
  assign n40888 = x199 | n40882 ;
  assign n40889 = x1091 & x1136 ;
  assign n40890 = x199 & ~n40874 ;
  assign n40891 = ~n40889 & n40890 ;
  assign n40892 = n40888 & ~n40891 ;
  assign n40893 = ~x200 & n40892 ;
  assign n40894 = x1091 & x1135 ;
  assign n40895 = n40888 | n40894 ;
  assign n40896 = x200 & ~n40890 ;
  assign n40897 = n40895 & n40896 ;
  assign n40898 = ( ~n15098 & n40893 ) | ( ~n15098 & n40897 ) | ( n40893 & n40897 ) ;
  assign n40899 = ~n15098 & n40898 ;
  assign n40900 = ( ~n40870 & n40887 ) | ( ~n40870 & n40899 ) | ( n40887 & n40899 ) ;
  assign n40901 = ~n40870 & n40900 ;
  assign n40902 = n15098 & ~n40857 ;
  assign n40903 = n36164 & ~n40860 ;
  assign n40904 = ( n15098 & n40863 ) | ( n15098 & ~n40903 ) | ( n40863 & ~n40903 ) ;
  assign n40905 = n40903 | n40904 ;
  assign n40906 = ( x230 & n40902 ) | ( x230 & n40905 ) | ( n40902 & n40905 ) ;
  assign n40907 = ~n40902 & n40906 ;
  assign n40908 = ~x199 & x1091 ;
  assign n40909 = ( ~x200 & n40892 ) | ( ~x200 & n40908 ) | ( n40892 & n40908 ) ;
  assign n40910 = ~x200 & n40909 ;
  assign n40911 = ( ~n15098 & n40897 ) | ( ~n15098 & n40910 ) | ( n40897 & n40910 ) ;
  assign n40912 = ~n15098 & n40911 ;
  assign n40913 = x1091 & ~n40856 ;
  assign n40914 = n40883 | n40913 ;
  assign n40915 = ( n40877 & ~n40878 ) | ( n40877 & n40914 ) | ( ~n40878 & n40914 ) ;
  assign n40916 = ( x230 & n40878 ) | ( x230 & n40915 ) | ( n40878 & n40915 ) ;
  assign n40917 = ( ~n40907 & n40912 ) | ( ~n40907 & n40916 ) | ( n40912 & n40916 ) ;
  assign n40918 = ~n40907 & n40917 ;
  assign n40919 = n40901 ^ x1134 ^ 1'b0 ;
  assign n40920 = ( n40901 & n40918 ) | ( n40901 & n40919 ) | ( n40918 & n40919 ) ;
  assign n40921 = ~x1154 & n36094 ;
  assign n40922 = ( n36143 & n36645 ) | ( n36143 & ~n40921 ) | ( n36645 & ~n40921 ) ;
  assign n40923 = ~n36143 & n40922 ;
  assign n40924 = ~x219 & n40923 ;
  assign n40925 = ~x199 & x1154 ;
  assign n40926 = x200 & ~n40925 ;
  assign n40927 = ( n36209 & n36558 ) | ( n36209 & ~n40926 ) | ( n36558 & ~n40926 ) ;
  assign n40928 = ~n36209 & n40927 ;
  assign n40929 = ( x219 & n36021 ) | ( x219 & n40928 ) | ( n36021 & n40928 ) ;
  assign n40930 = n40928 ^ n36021 ^ 1'b0 ;
  assign n40931 = ( x219 & n40929 ) | ( x219 & n40930 ) | ( n40929 & n40930 ) ;
  assign n40932 = ( x211 & ~n40924 ) | ( x211 & n40931 ) | ( ~n40924 & n40931 ) ;
  assign n40933 = n40924 | n40932 ;
  assign n40934 = x219 & ~n36559 ;
  assign n40935 = x1153 & ~n36216 ;
  assign n40936 = ~x1155 & n40935 ;
  assign n40937 = ( x1154 & n36507 ) | ( x1154 & n40936 ) | ( n36507 & n40936 ) ;
  assign n40938 = n36507 & n40937 ;
  assign n40939 = n40938 ^ x1155 ^ 1'b0 ;
  assign n40940 = ( ~x1155 & n37421 ) | ( ~x1155 & n40939 ) | ( n37421 & n40939 ) ;
  assign n40941 = ( x1155 & n40938 ) | ( x1155 & n40940 ) | ( n40938 & n40940 ) ;
  assign n40942 = x211 & ~n40941 ;
  assign n40943 = ( x211 & n40934 ) | ( x211 & n40942 ) | ( n40934 & n40942 ) ;
  assign n40944 = ( n7318 & n40933 ) | ( n7318 & ~n40943 ) | ( n40933 & ~n40943 ) ;
  assign n40945 = ~n7318 & n40944 ;
  assign n40946 = x219 | n35964 ;
  assign n40947 = ( n35980 & ~n36831 ) | ( n35980 & n40946 ) | ( ~n36831 & n40946 ) ;
  assign n40948 = ~n36831 & n40947 ;
  assign n40949 = n7318 & n40948 ;
  assign n40950 = ( x230 & n40945 ) | ( x230 & ~n40949 ) | ( n40945 & ~n40949 ) ;
  assign n40951 = ~n40945 & n40950 ;
  assign n40952 = n40364 | n40368 ;
  assign n40953 = x267 & ~n40952 ;
  assign n40954 = ~x267 & n38507 ;
  assign n40955 = ~n40056 & n40954 ;
  assign n40956 = ( n38458 & n40953 ) | ( n38458 & ~n40955 ) | ( n40953 & ~n40955 ) ;
  assign n40957 = ~n40953 & n40956 ;
  assign n40958 = x1091 & ~n40948 ;
  assign n40959 = x267 | x1091 ;
  assign n40960 = n38458 | n40959 ;
  assign n40961 = ~n40958 & n40960 ;
  assign n40962 = n7318 & ~n40961 ;
  assign n40963 = ( n7318 & n40957 ) | ( n7318 & n40962 ) | ( n40957 & n40962 ) ;
  assign n40964 = n40075 | n40097 ;
  assign n40965 = n38554 & n40964 ;
  assign n40966 = n38600 & ~n40965 ;
  assign n40967 = x1154 & ~n40679 ;
  assign n40968 = ( x1154 & n40966 ) | ( x1154 & n40967 ) | ( n40966 & n40967 ) ;
  assign n40969 = ~x1154 & n40086 ;
  assign n40970 = x1155 & ~n40969 ;
  assign n40971 = ~n40968 & n40970 ;
  assign n40972 = ( n38571 & n40968 ) | ( n38571 & ~n40971 ) | ( n40968 & ~n40971 ) ;
  assign n40973 = n40094 & n40349 ;
  assign n40974 = x1155 | n40451 ;
  assign n40975 = n40973 | n40974 ;
  assign n40976 = ( ~x211 & n40972 ) | ( ~x211 & n40975 ) | ( n40972 & n40975 ) ;
  assign n40977 = x211 & n40976 ;
  assign n40978 = x1153 & ~n38630 ;
  assign n40979 = x1155 | n40978 ;
  assign n40980 = x1153 | n40646 ;
  assign n40981 = ~n40979 & n40980 ;
  assign n40982 = x1153 & n38591 ;
  assign n40983 = n40453 | n40982 ;
  assign n40984 = x1155 & n40983 ;
  assign n40985 = x1154 & ~n40647 ;
  assign n40986 = ( n40981 & ~n40984 ) | ( n40981 & n40985 ) | ( ~n40984 & n40985 ) ;
  assign n40987 = ~n40981 & n40986 ;
  assign n40988 = n40136 & ~n40979 ;
  assign n40989 = x1154 | n40984 ;
  assign n40990 = n40988 | n40989 ;
  assign n40991 = ( x211 & ~n40987 ) | ( x211 & n40990 ) | ( ~n40987 & n40990 ) ;
  assign n40992 = ~x211 & n40991 ;
  assign n40993 = ( x267 & ~n40977 ) | ( x267 & n40992 ) | ( ~n40977 & n40992 ) ;
  assign n40994 = n40977 | n40993 ;
  assign n40995 = x1154 & ~n40965 ;
  assign n40996 = x1154 | n38525 ;
  assign n40997 = n40143 | n40996 ;
  assign n40998 = ( x1155 & ~n40995 ) | ( x1155 & n40997 ) | ( ~n40995 & n40997 ) ;
  assign n40999 = ~x1155 & n40998 ;
  assign n41000 = x1155 & ~n40153 ;
  assign n41001 = n38553 | n40634 ;
  assign n41002 = ( ~n40141 & n41000 ) | ( ~n40141 & n41001 ) | ( n41000 & n41001 ) ;
  assign n41003 = n40141 & n41002 ;
  assign n41004 = ( x267 & n40999 ) | ( x267 & ~n41003 ) | ( n40999 & ~n41003 ) ;
  assign n41005 = ~n40999 & n41004 ;
  assign n41008 = x1154 & x1155 ;
  assign n41009 = ( n38558 & ~n40342 ) | ( n38558 & n41008 ) | ( ~n40342 & n41008 ) ;
  assign n41010 = ~n38558 & n41009 ;
  assign n41006 = x1154 | n38541 ;
  assign n41007 = n40973 | n41006 ;
  assign n41011 = n41010 ^ n41007 ^ 1'b0 ;
  assign n41012 = ( x211 & ~n41007 ) | ( x211 & n41010 ) | ( ~n41007 & n41010 ) ;
  assign n41013 = ( x211 & ~n41011 ) | ( x211 & n41012 ) | ( ~n41011 & n41012 ) ;
  assign n41014 = n38577 & n40311 ;
  assign n41015 = x1155 | n41014 ;
  assign n41016 = ( ~x267 & n40973 ) | ( ~x267 & n41015 ) | ( n40973 & n41015 ) ;
  assign n41017 = ~x267 & n41016 ;
  assign n41018 = n35963 & ~n40091 ;
  assign n41019 = ( n40324 & ~n40982 ) | ( n40324 & n41018 ) | ( ~n40982 & n41018 ) ;
  assign n41020 = ~n40324 & n41019 ;
  assign n41021 = ( n41013 & n41017 ) | ( n41013 & ~n41020 ) | ( n41017 & ~n41020 ) ;
  assign n41022 = ~n41013 & n41021 ;
  assign n41023 = ( x219 & n41005 ) | ( x219 & n41022 ) | ( n41005 & n41022 ) ;
  assign n41024 = n41022 ^ n41005 ^ 1'b0 ;
  assign n41025 = ( x219 & n41023 ) | ( x219 & n41024 ) | ( n41023 & n41024 ) ;
  assign n41026 = n40597 & n41000 ;
  assign n41027 = ~x1155 & n38600 ;
  assign n41028 = n40983 ^ n38666 ^ n38631 ;
  assign n41029 = n41027 & n41028 ;
  assign n41030 = ( x1154 & n41026 ) | ( x1154 & ~n41029 ) | ( n41026 & ~n41029 ) ;
  assign n41031 = ~n41026 & n41030 ;
  assign n41032 = x1154 | n40097 ;
  assign n41033 = n38651 | n41032 ;
  assign n41034 = ~x1155 & n41033 ;
  assign n41035 = n38545 | n41032 ;
  assign n41036 = n41034 | n41035 ;
  assign n41037 = x211 & ~n41036 ;
  assign n41038 = ( x211 & n41031 ) | ( x211 & n41037 ) | ( n41031 & n41037 ) ;
  assign n41039 = x1154 & ~n41028 ;
  assign n41040 = n41034 & ~n41039 ;
  assign n41041 = n38644 | n40432 ;
  assign n41042 = n41041 ^ x211 ^ 1'b0 ;
  assign n41043 = x1154 & ~n38553 ;
  assign n41044 = x1155 & ~n41043 ;
  assign n41045 = ( n41041 & ~n41042 ) | ( n41041 & n41044 ) | ( ~n41042 & n41044 ) ;
  assign n41046 = ( x211 & n41042 ) | ( x211 & n41045 ) | ( n41042 & n41045 ) ;
  assign n41047 = ( x267 & n41040 ) | ( x267 & n41046 ) | ( n41040 & n41046 ) ;
  assign n41048 = n41046 ^ n41040 ^ 1'b0 ;
  assign n41049 = ( x267 & n41047 ) | ( x267 & n41048 ) | ( n41047 & n41048 ) ;
  assign n41050 = n41049 ^ n41038 ^ 1'b0 ;
  assign n41051 = ( n41038 & n41049 ) | ( n41038 & n41050 ) | ( n41049 & n41050 ) ;
  assign n41052 = ( x219 & ~n41038 ) | ( x219 & n41051 ) | ( ~n41038 & n41051 ) ;
  assign n41053 = ~n41025 & n41052 ;
  assign n41054 = ( n40994 & n41025 ) | ( n40994 & ~n41053 ) | ( n41025 & ~n41053 ) ;
  assign n41055 = ( ~x253 & x254 ) | ( ~x253 & n41054 ) | ( x254 & n41054 ) ;
  assign n41056 = x253 & n41055 ;
  assign n41057 = x1091 & n40923 ;
  assign n41058 = x211 | n41057 ;
  assign n41059 = x1091 & n40721 ;
  assign n41060 = n40188 & n41059 ;
  assign n41061 = x1154 & ~n41060 ;
  assign n41062 = ~x299 & n36506 ;
  assign n41063 = x1091 & ~x1155 ;
  assign n41064 = n41062 & n41063 ;
  assign n41065 = n41061 & ~n41064 ;
  assign n41066 = x1155 & n36559 ;
  assign n41067 = x1154 & ~n41066 ;
  assign n41068 = ( x1155 & n41065 ) | ( x1155 & n41067 ) | ( n41065 & n41067 ) ;
  assign n41069 = x211 & n41068 ;
  assign n41070 = ~n36227 & n40400 ;
  assign n41071 = n37424 & n41070 ;
  assign n41072 = x1154 & ~n41065 ;
  assign n41073 = ( x211 & ~n41071 ) | ( x211 & n41072 ) | ( ~n41071 & n41072 ) ;
  assign n41074 = n41071 | n41073 ;
  assign n41075 = ( x219 & n41069 ) | ( x219 & n41074 ) | ( n41069 & n41074 ) ;
  assign n41076 = ~n41069 & n41075 ;
  assign n41077 = n36507 & n41063 ;
  assign n41078 = ( n35964 & n41060 ) | ( n35964 & ~n41077 ) | ( n41060 & ~n41077 ) ;
  assign n41079 = ~n41060 & n41078 ;
  assign n41080 = x219 | n41079 ;
  assign n41081 = ~n41076 & n41080 ;
  assign n41082 = ( n41058 & n41076 ) | ( n41058 & ~n41081 ) | ( n41076 & ~n41081 ) ;
  assign n41083 = x1155 | n36592 ;
  assign n41084 = ~n36106 & n40175 ;
  assign n41085 = ( n40417 & n41083 ) | ( n40417 & n41084 ) | ( n41083 & n41084 ) ;
  assign n41086 = n41083 & n41085 ;
  assign n41087 = ( x211 & x1154 ) | ( x211 & ~n41086 ) | ( x1154 & ~n41086 ) ;
  assign n41088 = ~x1154 & n41087 ;
  assign n41089 = ( x267 & n41082 ) | ( x267 & ~n41088 ) | ( n41082 & ~n41088 ) ;
  assign n41090 = ~x267 & n41089 ;
  assign n41091 = ~x1155 & n36507 ;
  assign n41092 = ( ~n11550 & n36167 ) | ( ~n11550 & n41091 ) | ( n36167 & n41091 ) ;
  assign n41093 = ~n11550 & n41092 ;
  assign n41094 = ( x1091 & n41067 ) | ( x1091 & n41093 ) | ( n41067 & n41093 ) ;
  assign n41095 = ~n41093 & n41094 ;
  assign n41096 = n40400 & ~n40935 ;
  assign n41097 = n36227 | n38688 ;
  assign n41098 = n41096 & n41097 ;
  assign n41099 = ( x211 & n41095 ) | ( x211 & ~n41098 ) | ( n41095 & ~n41098 ) ;
  assign n41100 = ~n41095 & n41099 ;
  assign n41101 = ~n37425 & n41096 ;
  assign n41102 = x1091 & ~n41062 ;
  assign n41103 = n41061 & n41102 ;
  assign n41104 = ( x219 & n41101 ) | ( x219 & ~n41103 ) | ( n41101 & ~n41103 ) ;
  assign n41105 = ~n41101 & n41104 ;
  assign n41106 = x1155 | n40294 ;
  assign n41107 = n40214 & ~n41106 ;
  assign n41108 = x1155 & ~n40189 ;
  assign n41109 = n38693 & n41108 ;
  assign n41110 = ( x1154 & n41107 ) | ( x1154 & n41109 ) | ( n41107 & n41109 ) ;
  assign n41111 = n41109 ^ n41107 ^ 1'b0 ;
  assign n41112 = ( x1154 & n41110 ) | ( x1154 & n41111 ) | ( n41110 & n41111 ) ;
  assign n41113 = n40389 & n41108 ;
  assign n41114 = x1091 & ~n41083 ;
  assign n41115 = n41113 | n41114 ;
  assign n41116 = n41115 ^ x1154 ^ 1'b0 ;
  assign n41117 = ( x1154 & n41115 ) | ( x1154 & n41116 ) | ( n41115 & n41116 ) ;
  assign n41118 = ( x219 & ~x1154 ) | ( x219 & n41117 ) | ( ~x1154 & n41117 ) ;
  assign n41119 = ( ~n41105 & n41112 ) | ( ~n41105 & n41118 ) | ( n41112 & n41118 ) ;
  assign n41120 = ~n41105 & n41119 ;
  assign n41121 = ( x211 & ~n41100 ) | ( x211 & n41120 ) | ( ~n41100 & n41120 ) ;
  assign n41122 = ~n41100 & n41121 ;
  assign n41123 = ~n41090 & n41122 ;
  assign n41124 = ( x267 & n41090 ) | ( x267 & ~n41123 ) | ( n41090 & ~n41123 ) ;
  assign n41125 = ~n38458 & n41124 ;
  assign n41126 = ( n7318 & ~n41056 ) | ( n7318 & n41125 ) | ( ~n41056 & n41125 ) ;
  assign n41127 = n41056 | n41126 ;
  assign n41128 = ( n38506 & n40963 ) | ( n38506 & n41127 ) | ( n40963 & n41127 ) ;
  assign n41129 = ~n40963 & n41128 ;
  assign n41130 = x1091 ^ x267 ^ 1'b0 ;
  assign n41131 = ( x267 & n40948 ) | ( x267 & n41130 ) | ( n40948 & n41130 ) ;
  assign n41132 = ( n7318 & n38506 ) | ( n7318 & ~n41131 ) | ( n38506 & ~n41131 ) ;
  assign n41133 = n41131 ^ n38506 ^ 1'b0 ;
  assign n41134 = ( n38506 & n41132 ) | ( n38506 & ~n41133 ) | ( n41132 & ~n41133 ) ;
  assign n41135 = n7318 | n41124 ;
  assign n41136 = n41135 ^ n41134 ^ 1'b0 ;
  assign n41137 = ( n41134 & n41135 ) | ( n41134 & n41136 ) | ( n41135 & n41136 ) ;
  assign n41138 = ( x230 & ~n41134 ) | ( x230 & n41137 ) | ( ~n41134 & n41137 ) ;
  assign n41139 = ( ~n40951 & n41129 ) | ( ~n40951 & n41138 ) | ( n41129 & n41138 ) ;
  assign n41140 = ~n40951 & n41139 ;
  assign n41141 = ( n10075 & n10077 ) | ( n10075 & ~n40271 ) | ( n10077 & ~n40271 ) ;
  assign n41142 = x1151 & n41141 ;
  assign n41143 = x1152 | n41142 ;
  assign n41144 = ( x1150 & n40040 ) | ( x1150 & n41143 ) | ( n40040 & n41143 ) ;
  assign n41145 = ~x1150 & n41144 ;
  assign n41146 = n15098 & ~n40209 ;
  assign n41147 = n7318 | n36166 ;
  assign n41148 = ~n41146 & n41147 ;
  assign n41149 = x1151 & ~n41148 ;
  assign n41150 = ( x1152 & ~n41145 ) | ( x1152 & n41149 ) | ( ~n41145 & n41149 ) ;
  assign n41151 = n41150 ^ n41145 ^ 1'b0 ;
  assign n41152 = ( n41145 & ~n41150 ) | ( n41145 & n41151 ) | ( ~n41150 & n41151 ) ;
  assign n41153 = x268 & x1152 ;
  assign n41154 = ~x211 & n15098 ;
  assign n41155 = n7318 | n36106 ;
  assign n41156 = ~n41154 & n41155 ;
  assign n41157 = x1152 & ~n41156 ;
  assign n41159 = x219 & n15098 ;
  assign n41158 = x199 | n15098 ;
  assign n41160 = n41159 ^ n41158 ^ n15098 ;
  assign n41161 = ~n41157 & n41160 ;
  assign n41162 = ~x1151 & n41156 ;
  assign n41163 = ( x1150 & n41161 ) | ( x1150 & ~n41162 ) | ( n41161 & ~n41162 ) ;
  assign n41164 = ~n41161 & n41163 ;
  assign n41165 = ~n41153 & n41164 ;
  assign n41166 = ( x1091 & n41152 ) | ( x1091 & n41165 ) | ( n41152 & n41165 ) ;
  assign n41167 = n41165 ^ n41152 ^ 1'b0 ;
  assign n41168 = ( x1091 & n41166 ) | ( x1091 & n41167 ) | ( n41166 & n41167 ) ;
  assign n41169 = x1152 & n41164 ;
  assign n41170 = x1091 & ~n41169 ;
  assign n41171 = ~n41168 & n41170 ;
  assign n41172 = ( x268 & n41168 ) | ( x268 & ~n41171 ) | ( n41168 & ~n41171 ) ;
  assign n41173 = n41172 ^ n38505 ^ 1'b0 ;
  assign n41174 = ( n38505 & n41172 ) | ( n38505 & n41173 ) | ( n41172 & n41173 ) ;
  assign n41175 = ( x230 & ~n38505 ) | ( x230 & n41174 ) | ( ~n38505 & n41174 ) ;
  assign n41176 = n38647 ^ x219 ^ 1'b0 ;
  assign n41177 = ( n38647 & n40093 ) | ( n38647 & n41176 ) | ( n40093 & n41176 ) ;
  assign n41178 = ( x57 & ~n5193 ) | ( x57 & n41177 ) | ( ~n5193 & n41177 ) ;
  assign n41179 = ~x57 & n41178 ;
  assign n41180 = x219 | n38571 ;
  assign n41181 = ( ~n38540 & n41179 ) | ( ~n38540 & n41180 ) | ( n41179 & n41180 ) ;
  assign n41182 = n38540 & n41181 ;
  assign n41183 = n7318 & ~n40056 ;
  assign n41184 = n41182 ^ n40057 ^ 1'b0 ;
  assign n41185 = ( ~n40057 & n41183 ) | ( ~n40057 & n41184 ) | ( n41183 & n41184 ) ;
  assign n41186 = ( n40057 & n41182 ) | ( n40057 & n41185 ) | ( n41182 & n41185 ) ;
  assign n41187 = ~x1151 & n41186 ;
  assign n41188 = n40071 & n41183 ;
  assign n41189 = n38556 & n40154 ;
  assign n41190 = x219 & n40093 ;
  assign n41191 = n38523 & n41190 ;
  assign n41192 = n41189 | n41191 ;
  assign n41193 = ~n7318 & n41192 ;
  assign n41194 = n41188 | n41193 ;
  assign n41195 = x1151 & n41194 ;
  assign n41196 = ( x1152 & n41187 ) | ( x1152 & ~n41195 ) | ( n41187 & ~n41195 ) ;
  assign n41197 = ~n41187 & n41196 ;
  assign n41198 = n38587 | n40144 ;
  assign n41199 = n41192 & n41198 ;
  assign n41200 = n7318 | n41199 ;
  assign n41201 = x219 & n7318 ;
  assign n41202 = ~n38473 & n41201 ;
  assign n41203 = n40072 | n41202 ;
  assign n41204 = n41200 & ~n41203 ;
  assign n41205 = x1151 & n41204 ;
  assign n41206 = n7318 | n40137 ;
  assign n41207 = n38529 | n41206 ;
  assign n41208 = n40057 & ~n41202 ;
  assign n41209 = n41207 & n41208 ;
  assign n41210 = ~x1151 & n41209 ;
  assign n41211 = ( x1152 & ~n41205 ) | ( x1152 & n41210 ) | ( ~n41205 & n41210 ) ;
  assign n41212 = n41205 | n41211 ;
  assign n41213 = n41212 ^ n41197 ^ 1'b0 ;
  assign n41214 = ( n41197 & n41212 ) | ( n41197 & n41213 ) | ( n41212 & n41213 ) ;
  assign n41215 = ( x268 & ~n41197 ) | ( x268 & n41214 ) | ( ~n41197 & n41214 ) ;
  assign n41216 = n40063 & n41183 ;
  assign n41217 = x219 & ~n38513 ;
  assign n41218 = n40119 | n41217 ;
  assign n41219 = n38515 & n41218 ;
  assign n41220 = n40092 | n41219 ;
  assign n41221 = n7318 | n41220 ;
  assign n41222 = ( ~n7318 & n41216 ) | ( ~n7318 & n41221 ) | ( n41216 & n41221 ) ;
  assign n41223 = ~x1151 & n41222 ;
  assign n41224 = n7318 & ~n40368 ;
  assign n41225 = ~n40047 & n41224 ;
  assign n41226 = n41216 & ~n41225 ;
  assign n41227 = n41188 | n41226 ;
  assign n41228 = n41179 | n41227 ;
  assign n41229 = x1151 & n41228 ;
  assign n41230 = ( x268 & ~n41223 ) | ( x268 & n41229 ) | ( ~n41223 & n41229 ) ;
  assign n41231 = n41223 | n41230 ;
  assign n41232 = x1091 | n38464 ;
  assign n41233 = n7318 | n40079 ;
  assign n41234 = n41232 & ~n41233 ;
  assign n41235 = x219 & n38574 ;
  assign n41236 = n41206 | n41235 ;
  assign n41237 = ~n40364 & n41224 ;
  assign n41238 = ( n41234 & n41236 ) | ( n41234 & ~n41237 ) | ( n41236 & ~n41237 ) ;
  assign n41239 = ~n41234 & n41238 ;
  assign n41240 = x1151 & ~n41239 ;
  assign n41241 = x268 & ~n41240 ;
  assign n41242 = ~n40070 & n41224 ;
  assign n41243 = ~n38473 & n40156 ;
  assign n41244 = ( n41200 & ~n41242 ) | ( n41200 & n41243 ) | ( ~n41242 & n41243 ) ;
  assign n41245 = ~n41242 & n41244 ;
  assign n41246 = x1151 | n41245 ;
  assign n41247 = n41241 & n41246 ;
  assign n41248 = x1152 & ~n41247 ;
  assign n41249 = n41231 & n41248 ;
  assign n41250 = ~n7318 & n38512 ;
  assign n41251 = n41219 & n41250 ;
  assign n41252 = n41226 | n41251 ;
  assign n41253 = x1151 | n41252 ;
  assign n41254 = n40066 & ~n40364 ;
  assign n41255 = n41236 & ~n41254 ;
  assign n41256 = n38468 & ~n41255 ;
  assign n41257 = n41209 | n41256 ;
  assign n41258 = x1151 & ~n41257 ;
  assign n41259 = ( x268 & n41253 ) | ( x268 & ~n41258 ) | ( n41253 & ~n41258 ) ;
  assign n41260 = ~x268 & n41259 ;
  assign n41262 = n40066 & ~n40070 ;
  assign n41263 = n41192 | n41233 ;
  assign n41264 = ~n41262 & n41263 ;
  assign n41265 = x1151 | n41264 ;
  assign n41261 = x1151 | n41255 ;
  assign n41266 = n41265 ^ n41261 ^ n41255 ;
  assign n41267 = x268 & ~n41266 ;
  assign n41268 = ( ~x1152 & n41260 ) | ( ~x1152 & n41267 ) | ( n41260 & n41267 ) ;
  assign n41269 = ~x1152 & n41268 ;
  assign n41270 = ( x1150 & n41249 ) | ( x1150 & n41269 ) | ( n41249 & n41269 ) ;
  assign n41271 = n41269 ^ n41249 ^ 1'b0 ;
  assign n41272 = ( x1150 & n41270 ) | ( x1150 & n41271 ) | ( n41270 & n41271 ) ;
  assign n41273 = x219 & n40141 ;
  assign n41274 = n7318 | n40144 ;
  assign n41275 = ( ~n41225 & n41273 ) | ( ~n41225 & n41274 ) | ( n41273 & n41274 ) ;
  assign n41276 = ~n41225 & n41275 ;
  assign n41277 = ~x1151 & n41276 ;
  assign n41278 = ~n40064 & n41224 ;
  assign n41279 = ( n38654 & n40119 ) | ( n38654 & n41273 ) | ( n40119 & n41273 ) ;
  assign n41280 = ( n7318 & ~n41278 ) | ( n7318 & n41279 ) | ( ~n41278 & n41279 ) ;
  assign n41281 = ~n41278 & n41280 ;
  assign n41282 = x1151 & n41281 ;
  assign n41283 = ( x1152 & n41277 ) | ( x1152 & ~n41282 ) | ( n41277 & ~n41282 ) ;
  assign n41284 = ~n41277 & n41283 ;
  assign n41285 = n38468 | n41255 ;
  assign n41286 = ~x1151 & n41285 ;
  assign n41287 = x1152 | n41286 ;
  assign n41288 = n7318 | n40115 ;
  assign n41289 = n40119 | n41288 ;
  assign n41290 = ~n40067 & n41289 ;
  assign n41291 = x1151 & n41290 ;
  assign n41292 = ( x268 & n41287 ) | ( x268 & n41291 ) | ( n41287 & n41291 ) ;
  assign n41293 = n41291 ^ n41287 ^ 1'b0 ;
  assign n41294 = ( x268 & n41292 ) | ( x268 & n41293 ) | ( n41292 & n41293 ) ;
  assign n41295 = n41294 ^ n41284 ^ 1'b0 ;
  assign n41296 = ( n41284 & n41294 ) | ( n41284 & n41295 ) | ( n41294 & n41295 ) ;
  assign n41297 = ( x1150 & ~n41284 ) | ( x1150 & n41296 ) | ( ~n41284 & n41296 ) ;
  assign n41298 = ~n41272 & n41297 ;
  assign n41299 = ( n41215 & n41272 ) | ( n41215 & ~n41298 ) | ( n41272 & ~n41298 ) ;
  assign n41300 = n41175 ^ n38505 ^ 1'b0 ;
  assign n41301 = ( ~n38505 & n41299 ) | ( ~n38505 & n41300 ) | ( n41299 & n41300 ) ;
  assign n41302 = ( n38505 & n41175 ) | ( n38505 & n41301 ) | ( n41175 & n41301 ) ;
  assign n41303 = x230 & ~n41164 ;
  assign n41304 = ( n41152 & n41302 ) | ( n41152 & ~n41303 ) | ( n41302 & ~n41303 ) ;
  assign n41305 = n41302 ^ n41152 ^ 1'b0 ;
  assign n41306 = ( n41302 & n41304 ) | ( n41302 & ~n41305 ) | ( n41304 & ~n41305 ) ;
  assign n41307 = ~x199 & x1137 ;
  assign n41308 = x200 & ~n41307 ;
  assign n41309 = ~x199 & x1136 ;
  assign n41310 = x199 & x1138 ;
  assign n41311 = x200 | n41310 ;
  assign n41312 = n41309 | n41311 ;
  assign n41313 = ( n15098 & ~n41308 ) | ( n15098 & n41312 ) | ( ~n41308 & n41312 ) ;
  assign n41314 = ~n15098 & n41313 ;
  assign n41315 = ~x211 & x1138 ;
  assign n41316 = x1136 ^ x211 ^ 1'b0 ;
  assign n41317 = ( x1136 & x1137 ) | ( x1136 & n41316 ) | ( x1137 & n41316 ) ;
  assign n41318 = n41315 ^ x219 ^ 1'b0 ;
  assign n41319 = ( n41315 & n41317 ) | ( n41315 & ~n41318 ) | ( n41317 & ~n41318 ) ;
  assign n41320 = n7318 ^ x299 ^ 1'b0 ;
  assign n41321 = ( x299 & n7318 ) | ( x299 & ~n41320 ) | ( n7318 & ~n41320 ) ;
  assign n41322 = ( n41319 & n41320 ) | ( n41319 & n41321 ) | ( n41320 & n41321 ) ;
  assign n41323 = ( x230 & n41314 ) | ( x230 & n41322 ) | ( n41314 & n41322 ) ;
  assign n41324 = n41322 ^ n41314 ^ 1'b0 ;
  assign n41325 = ( x230 & n41323 ) | ( x230 & n41324 ) | ( n41323 & n41324 ) ;
  assign n41326 = ~x817 & n38462 ;
  assign n41327 = x269 & ~n38462 ;
  assign n41328 = ( x1091 & ~n41326 ) | ( x1091 & n41327 ) | ( ~n41326 & n41327 ) ;
  assign n41329 = n41326 | n41328 ;
  assign n41330 = ~x200 & x1091 ;
  assign n41331 = x1138 & n41330 ;
  assign n41332 = x199 & ~n41331 ;
  assign n41333 = ~n15098 & n41332 ;
  assign n41334 = x1138 & n40233 ;
  assign n41335 = n41159 & ~n41334 ;
  assign n41336 = ( n41329 & n41333 ) | ( n41329 & n41335 ) | ( n41333 & n41335 ) ;
  assign n41337 = n41335 ^ n41333 ^ 1'b0 ;
  assign n41338 = ( n41329 & n41336 ) | ( n41329 & n41337 ) | ( n41336 & n41337 ) ;
  assign n41339 = x1091 & n41317 ;
  assign n41340 = n37869 & ~n41339 ;
  assign n41341 = ~x200 & n40889 ;
  assign n41342 = x1137 & n38701 ;
  assign n41343 = n41341 | n41342 ;
  assign n41344 = ( n41158 & ~n41340 ) | ( n41158 & n41343 ) | ( ~n41340 & n41343 ) ;
  assign n41345 = ~n41340 & n41344 ;
  assign n41346 = ~x817 & n38479 ;
  assign n41347 = x1091 | n41346 ;
  assign n41348 = n38479 & ~n41347 ;
  assign n41349 = ( x269 & n41347 ) | ( x269 & ~n41348 ) | ( n41347 & ~n41348 ) ;
  assign n41350 = ( n41338 & ~n41345 ) | ( n41338 & n41349 ) | ( ~n41345 & n41349 ) ;
  assign n41351 = n41345 ^ n41338 ^ 1'b0 ;
  assign n41352 = ( n41338 & n41350 ) | ( n41338 & ~n41351 ) | ( n41350 & ~n41351 ) ;
  assign n41353 = ( x230 & ~n41325 ) | ( x230 & n41352 ) | ( ~n41325 & n41352 ) ;
  assign n41354 = ~n41325 & n41353 ;
  assign n41355 = ~x805 & n38479 ;
  assign n41356 = x1091 | n41355 ;
  assign n41357 = n38479 & ~n41356 ;
  assign n41358 = ( x270 & n41356 ) | ( x270 & ~n41357 ) | ( n41356 & ~n41357 ) ;
  assign n41359 = ~x805 & n38462 ;
  assign n41360 = x1091 | n41359 ;
  assign n41361 = n38462 & ~n41360 ;
  assign n41362 = ( x270 & n41360 ) | ( x270 & ~n41361 ) | ( n41360 & ~n41361 ) ;
  assign n41363 = n41362 ^ x230 ^ 1'b0 ;
  assign n41364 = ~x200 & n40782 ;
  assign n41365 = ( x199 & n15098 ) | ( x199 & ~n41364 ) | ( n15098 & ~n41364 ) ;
  assign n41366 = ~n15098 & n41365 ;
  assign n41367 = n40233 & n40766 ;
  assign n41368 = ~n41366 & n41367 ;
  assign n41369 = ( n41159 & n41366 ) | ( n41159 & ~n41368 ) | ( n41366 & ~n41368 ) ;
  assign n41370 = ( n41362 & ~n41363 ) | ( n41362 & n41369 ) | ( ~n41363 & n41369 ) ;
  assign n41371 = ( x230 & n41363 ) | ( x230 & n41370 ) | ( n41363 & n41370 ) ;
  assign n41372 = x1139 ^ x211 ^ 1'b0 ;
  assign n41373 = ( x1139 & x1140 ) | ( x1139 & n41372 ) | ( x1140 & n41372 ) ;
  assign n41374 = x1091 & n41373 ;
  assign n41375 = n37869 & ~n41374 ;
  assign n41378 = x1139 & n41330 ;
  assign n41376 = x1091 & x1140 ;
  assign n41377 = ~x200 & n41376 ;
  assign n41379 = n41378 ^ n41377 ^ n41376 ;
  assign n41380 = n41158 | n41379 ;
  assign n41381 = ~n41375 & n41380 ;
  assign n41382 = ~n41371 & n41381 ;
  assign n41383 = ( n41358 & n41371 ) | ( n41358 & ~n41382 ) | ( n41371 & ~n41382 ) ;
  assign n41384 = n40766 ^ x219 ^ 1'b0 ;
  assign n41385 = ( n40766 & n41373 ) | ( n40766 & ~n41384 ) | ( n41373 & ~n41384 ) ;
  assign n41386 = ( x230 & n38767 ) | ( x230 & n41385 ) | ( n38767 & n41385 ) ;
  assign n41387 = ~x199 & x1140 ;
  assign n41388 = x200 & ~n41387 ;
  assign n41389 = ~x199 & x1139 ;
  assign n41390 = x199 & x1141 ;
  assign n41391 = x200 | n41390 ;
  assign n41392 = ( ~n41388 & n41389 ) | ( ~n41388 & n41391 ) | ( n41389 & n41391 ) ;
  assign n41393 = ~n41388 & n41392 ;
  assign n41394 = ( x299 & n7318 ) | ( x299 & ~n41393 ) | ( n7318 & ~n41393 ) ;
  assign n41395 = n41393 | n41394 ;
  assign n41396 = n41383 & ~n41395 ;
  assign n41397 = ( n41383 & ~n41386 ) | ( n41383 & n41396 ) | ( ~n41386 & n41396 ) ;
  assign n41398 = x1147 & n40036 ;
  assign n41399 = ( ~x219 & n37647 ) | ( ~x219 & n37667 ) | ( n37647 & n37667 ) ;
  assign n41400 = n41398 | n41399 ;
  assign n41401 = ( n37163 & n37908 ) | ( n37163 & ~n37917 ) | ( n37908 & ~n37917 ) ;
  assign n41402 = ( ~n7318 & n41400 ) | ( ~n7318 & n41401 ) | ( n41400 & n41401 ) ;
  assign n41403 = ~n7318 & n41402 ;
  assign n41404 = n37075 | n39111 ;
  assign n41405 = ~x211 & x1147 ;
  assign n41406 = x219 & ~n41405 ;
  assign n41407 = n7318 & ~n41406 ;
  assign n41408 = n41404 & n41407 ;
  assign n41409 = ( x230 & n41403 ) | ( x230 & ~n41408 ) | ( n41403 & ~n41408 ) ;
  assign n41410 = ~n41403 & n41409 ;
  assign n41411 = n38465 ^ x271 ^ 1'b0 ;
  assign n41412 = ( n38465 & ~n41232 ) | ( n38465 & n41411 ) | ( ~n41232 & n41411 ) ;
  assign n41413 = x219 & ~n41412 ;
  assign n41414 = x1091 & x1146 ;
  assign n41415 = x1091 | n38481 ;
  assign n41416 = n41415 ^ n41412 ^ n41232 ;
  assign n41417 = n41414 | n41416 ;
  assign n41418 = ~x211 & n41414 ;
  assign n41419 = n41417 & ~n41418 ;
  assign n41420 = x1091 & n37075 ;
  assign n41421 = x219 | n41420 ;
  assign n41422 = ( ~n41413 & n41419 ) | ( ~n41413 & n41421 ) | ( n41419 & n41421 ) ;
  assign n41423 = ~n41413 & n41422 ;
  assign n41424 = n40048 & n41405 ;
  assign n41425 = ( n15098 & n41423 ) | ( n15098 & ~n41424 ) | ( n41423 & ~n41424 ) ;
  assign n41426 = ~n41423 & n41425 ;
  assign n41427 = n41412 ^ x199 ^ 1'b0 ;
  assign n41428 = ( n41412 & n41417 ) | ( n41412 & ~n41427 ) | ( n41417 & ~n41427 ) ;
  assign n41429 = x200 & ~n41428 ;
  assign n41430 = x1091 & x1145 ;
  assign n41431 = x199 | n41430 ;
  assign n41432 = n41416 | n41431 ;
  assign n41433 = ( ~x199 & n41412 ) | ( ~x199 & n41427 ) | ( n41412 & n41427 ) ;
  assign n41434 = ( ~n41427 & n41432 ) | ( ~n41427 & n41433 ) | ( n41432 & n41433 ) ;
  assign n41435 = x1147 & n38717 ;
  assign n41436 = x200 | n41435 ;
  assign n41437 = ( ~n41429 & n41434 ) | ( ~n41429 & n41436 ) | ( n41434 & n41436 ) ;
  assign n41438 = ~n41429 & n41437 ;
  assign n41439 = ( n15098 & ~n41426 ) | ( n15098 & n41438 ) | ( ~n41426 & n41438 ) ;
  assign n41440 = ~n41426 & n41439 ;
  assign n41441 = ( x230 & ~n41410 ) | ( x230 & n41440 ) | ( ~n41410 & n41440 ) ;
  assign n41442 = ~n41410 & n41441 ;
  assign n41443 = x1149 & ~x1150 ;
  assign n41444 = n7318 | n36112 ;
  assign n41445 = ( n37869 & ~n41154 ) | ( n37869 & n41444 ) | ( ~n41154 & n41444 ) ;
  assign n41446 = ~n37869 & n41445 ;
  assign n41447 = ( x1149 & n41443 ) | ( x1149 & n41446 ) | ( n41443 & n41446 ) ;
  assign n41448 = n41160 & n41447 ;
  assign n41449 = n7318 & ~n9343 ;
  assign n41450 = n11553 & ~n41449 ;
  assign n41451 = ~x1150 & n41450 ;
  assign n41452 = ( ~x1149 & n41156 ) | ( ~x1149 & n41451 ) | ( n41156 & n41451 ) ;
  assign n41453 = ~x1149 & n41452 ;
  assign n41454 = x1148 & ~n41453 ;
  assign n41455 = ~n41448 & n41454 ;
  assign n41456 = x1150 & n40039 ;
  assign n41457 = x1149 | n41456 ;
  assign n41458 = ~x1148 & n41457 ;
  assign n41459 = ~x1150 & n41141 ;
  assign n41460 = x1149 & ~n41148 ;
  assign n41461 = n41447 | n41460 ;
  assign n41462 = ~n41459 & n41461 ;
  assign n41463 = n41458 & ~n41462 ;
  assign n41464 = ( x230 & n41455 ) | ( x230 & ~n41463 ) | ( n41455 & ~n41463 ) ;
  assign n41465 = ~n41455 & n41464 ;
  assign n41466 = n41458 ^ x283 ^ 1'b0 ;
  assign n41467 = x1150 & n41148 ;
  assign n41468 = x1149 & ~n41459 ;
  assign n41469 = x1091 & ~n41468 ;
  assign n41470 = ( x1091 & n41467 ) | ( x1091 & n41469 ) | ( n41467 & n41469 ) ;
  assign n41471 = ( n41458 & ~n41466 ) | ( n41458 & n41470 ) | ( ~n41466 & n41470 ) ;
  assign n41472 = ( x283 & n41466 ) | ( x283 & n41471 ) | ( n41466 & n41471 ) ;
  assign n41473 = n41472 ^ x1091 ^ 1'b0 ;
  assign n41474 = ( ~x1091 & n41455 ) | ( ~x1091 & n41473 ) | ( n41455 & n41473 ) ;
  assign n41475 = ( x1091 & n41472 ) | ( x1091 & n41474 ) | ( n41472 & n41474 ) ;
  assign n41476 = x1150 & n41228 ;
  assign n41477 = ~x1150 & n41257 ;
  assign n41478 = x1149 & ~n41477 ;
  assign n41479 = ~n41476 & n41478 ;
  assign n41480 = x1150 & n41222 ;
  assign n41481 = ~x1150 & n41252 ;
  assign n41482 = x1149 | n41481 ;
  assign n41483 = n41480 | n41482 ;
  assign n41484 = x1148 & ~n41483 ;
  assign n41485 = ( x1148 & n41479 ) | ( x1148 & n41484 ) | ( n41479 & n41484 ) ;
  assign n41486 = x1150 | n41209 ;
  assign n41487 = ~x1149 & n41486 ;
  assign n41488 = x1150 & ~n41186 ;
  assign n41489 = n41487 & ~n41488 ;
  assign n41490 = x1150 & ~n41194 ;
  assign n41491 = x1149 & ~n41490 ;
  assign n41492 = x1150 | n41204 ;
  assign n41493 = n41491 & n41492 ;
  assign n41494 = ( x1148 & ~n41489 ) | ( x1148 & n41493 ) | ( ~n41489 & n41493 ) ;
  assign n41495 = n41489 | n41494 ;
  assign n41496 = x283 & ~n41495 ;
  assign n41497 = ( x283 & n41485 ) | ( x283 & n41496 ) | ( n41485 & n41496 ) ;
  assign n41498 = ( x272 & n41475 ) | ( x272 & ~n41497 ) | ( n41475 & ~n41497 ) ;
  assign n41499 = ~x272 & n41498 ;
  assign n41500 = n41156 | n41443 ;
  assign n41501 = n41160 & n41500 ;
  assign n41502 = ( x1091 & n41453 ) | ( x1091 & n41501 ) | ( n41453 & n41501 ) ;
  assign n41503 = n41501 ^ n41453 ^ 1'b0 ;
  assign n41504 = ( x1091 & n41502 ) | ( x1091 & n41503 ) | ( n41502 & n41503 ) ;
  assign n41505 = ( x283 & x1148 ) | ( x283 & ~n41504 ) | ( x1148 & ~n41504 ) ;
  assign n41506 = n41505 ^ x1148 ^ 1'b0 ;
  assign n41507 = ( x283 & n41505 ) | ( x283 & ~n41506 ) | ( n41505 & ~n41506 ) ;
  assign n41508 = n15098 & n40396 ;
  assign n41509 = ~n7318 & n38729 ;
  assign n41510 = n41508 | n41509 ;
  assign n41511 = x1150 | n41510 ;
  assign n41512 = x1091 & ~n41148 ;
  assign n41513 = x1150 & ~n41512 ;
  assign n41514 = x1149 & ~n41513 ;
  assign n41515 = n41511 & n41514 ;
  assign n41516 = x1091 & ~n41457 ;
  assign n41517 = ( x1148 & ~n41515 ) | ( x1148 & n41516 ) | ( ~n41515 & n41516 ) ;
  assign n41518 = n41515 | n41517 ;
  assign n41519 = x272 & ~n41518 ;
  assign n41520 = ( x272 & n41507 ) | ( x272 & n41519 ) | ( n41507 & n41519 ) ;
  assign n41521 = x1150 & n41276 ;
  assign n41522 = ~x1150 & n41285 ;
  assign n41523 = ( x1149 & ~n41521 ) | ( x1149 & n41522 ) | ( ~n41521 & n41522 ) ;
  assign n41524 = n41521 | n41523 ;
  assign n41525 = x1150 & n41281 ;
  assign n41526 = ~x1150 & n41290 ;
  assign n41527 = x1149 & ~n41526 ;
  assign n41528 = ~n41525 & n41527 ;
  assign n41529 = ( x1148 & n41524 ) | ( x1148 & ~n41528 ) | ( n41524 & ~n41528 ) ;
  assign n41530 = n41529 ^ n41524 ^ 1'b0 ;
  assign n41531 = ( x1148 & n41529 ) | ( x1148 & ~n41530 ) | ( n41529 & ~n41530 ) ;
  assign n41536 = ~x1150 & n41255 ;
  assign n41537 = x1150 & n41239 ;
  assign n41538 = ( x1149 & n41536 ) | ( x1149 & ~n41537 ) | ( n41536 & ~n41537 ) ;
  assign n41539 = ~n41536 & n41538 ;
  assign n41532 = x1150 & n41245 ;
  assign n41533 = ~x1150 & n41264 ;
  assign n41534 = ( x1149 & ~n41532 ) | ( x1149 & n41533 ) | ( ~n41532 & n41533 ) ;
  assign n41535 = n41532 | n41534 ;
  assign n41540 = n41539 ^ n41535 ^ 1'b0 ;
  assign n41541 = ( x1148 & ~n41535 ) | ( x1148 & n41539 ) | ( ~n41535 & n41539 ) ;
  assign n41542 = ( x1148 & ~n41540 ) | ( x1148 & n41541 ) | ( ~n41540 & n41541 ) ;
  assign n41543 = x283 & ~n41542 ;
  assign n41544 = n41531 & n41543 ;
  assign n41545 = ( x230 & n41520 ) | ( x230 & ~n41544 ) | ( n41520 & ~n41544 ) ;
  assign n41546 = n41545 ^ n41520 ^ 1'b0 ;
  assign n41547 = ( x230 & n41545 ) | ( x230 & ~n41546 ) | ( n41545 & ~n41546 ) ;
  assign n41548 = ( ~n41465 & n41499 ) | ( ~n41465 & n41547 ) | ( n41499 & n41547 ) ;
  assign n41549 = ~n41465 & n41548 ;
  assign n41550 = x1146 & ~n38964 ;
  assign n41551 = ~n41450 & n41550 ;
  assign n41552 = x1148 | n41551 ;
  assign n41553 = n37869 & n38417 ;
  assign n41554 = x1146 | n9353 ;
  assign n41555 = ~n41158 & n41554 ;
  assign n41556 = ( x1147 & n41553 ) | ( x1147 & n41555 ) | ( n41553 & n41555 ) ;
  assign n41557 = n41555 ^ n41553 ^ 1'b0 ;
  assign n41558 = ( x1147 & n41556 ) | ( x1147 & n41557 ) | ( n41556 & n41557 ) ;
  assign n41559 = ( x230 & n41552 ) | ( x230 & n41558 ) | ( n41552 & n41558 ) ;
  assign n41560 = n41558 ^ n41552 ^ 1'b0 ;
  assign n41561 = ( x230 & n41559 ) | ( x230 & n41560 ) | ( n41559 & n41560 ) ;
  assign n41562 = n37775 & n40048 ;
  assign n41563 = x273 | n38483 ;
  assign n41564 = ~n38490 & n41563 ;
  assign n41565 = ~x200 & n41414 ;
  assign n41566 = x199 | n41565 ;
  assign n41567 = n41564 | n41566 ;
  assign n41568 = x273 | n38466 ;
  assign n41569 = ~n38467 & n41568 ;
  assign n41570 = x199 & ~n41569 ;
  assign n41571 = ( x299 & n41567 ) | ( x299 & ~n41570 ) | ( n41567 & ~n41570 ) ;
  assign n41572 = ~x299 & n41571 ;
  assign n41573 = n38718 & ~n41429 ;
  assign n41574 = n41572 | n41573 ;
  assign n41575 = x1091 & n38496 ;
  assign n41576 = x219 & ~n41569 ;
  assign n41577 = x219 | n41418 ;
  assign n41578 = ( n41564 & ~n41576 ) | ( n41564 & n41577 ) | ( ~n41576 & n41577 ) ;
  assign n41579 = ~n41576 & n41578 ;
  assign n41580 = x299 & n41579 ;
  assign n41581 = ( x299 & n41575 ) | ( x299 & n41580 ) | ( n41575 & n41580 ) ;
  assign n41582 = ( ~n7318 & n41574 ) | ( ~n7318 & n41581 ) | ( n41574 & n41581 ) ;
  assign n41583 = ~n7318 & n41582 ;
  assign n41584 = ( x1148 & n41562 ) | ( x1148 & ~n41583 ) | ( n41562 & ~n41583 ) ;
  assign n41585 = ~n41562 & n41584 ;
  assign n41586 = n41572 | n41580 ;
  assign n41587 = ~n38032 & n41586 ;
  assign n41588 = ( x1148 & ~n41585 ) | ( x1148 & n41587 ) | ( ~n41585 & n41587 ) ;
  assign n41589 = ~n41585 & n41588 ;
  assign n41590 = n41589 ^ n7318 ^ 1'b0 ;
  assign n41591 = ( ~n7318 & n41579 ) | ( ~n7318 & n41590 ) | ( n41579 & n41590 ) ;
  assign n41592 = ( n7318 & n41589 ) | ( n7318 & n41591 ) | ( n41589 & n41591 ) ;
  assign n41593 = n10076 | n38579 ;
  assign n41594 = x1091 & n41593 ;
  assign n41595 = ( ~n7318 & n41586 ) | ( ~n7318 & n41594 ) | ( n41586 & n41594 ) ;
  assign n41596 = ~n7318 & n41595 ;
  assign n41597 = x1091 & n40067 ;
  assign n41598 = ( x1147 & n41596 ) | ( x1147 & n41597 ) | ( n41596 & n41597 ) ;
  assign n41599 = n41597 ^ n41596 ^ 1'b0 ;
  assign n41600 = ( x1147 & n41598 ) | ( x1147 & n41599 ) | ( n41598 & n41599 ) ;
  assign n41601 = ( ~x230 & n41592 ) | ( ~x230 & n41600 ) | ( n41592 & n41600 ) ;
  assign n41602 = ~x230 & n41601 ;
  assign n41603 = x1147 & n37869 ;
  assign n41604 = n41154 | n41603 ;
  assign n41605 = x1146 | n9343 ;
  assign n41606 = n41604 & n41605 ;
  assign n41607 = ~x199 & x1147 ;
  assign n41608 = x200 & ~n41607 ;
  assign n41609 = ( n15098 & n41554 ) | ( n15098 & ~n41608 ) | ( n41554 & ~n41608 ) ;
  assign n41610 = ~n15098 & n41609 ;
  assign n41611 = ( x1148 & n41606 ) | ( x1148 & ~n41610 ) | ( n41606 & ~n41610 ) ;
  assign n41612 = ~n41606 & n41611 ;
  assign n41613 = ~n41602 & n41612 ;
  assign n41614 = ( n41561 & n41602 ) | ( n41561 & ~n41613 ) | ( n41602 & ~n41613 ) ;
  assign n41615 = x219 | n36046 ;
  assign n41616 = n37076 | n41615 ;
  assign n41617 = n35995 | n37911 ;
  assign n41618 = ~n38371 & n41617 ;
  assign n41619 = n36026 | n37647 ;
  assign n41620 = n41618 ^ n41616 ^ 1'b0 ;
  assign n41621 = ( ~n41616 & n41619 ) | ( ~n41616 & n41620 ) | ( n41619 & n41620 ) ;
  assign n41622 = ( n41616 & n41618 ) | ( n41616 & n41621 ) | ( n41618 & n41621 ) ;
  assign n41623 = n41622 ^ n7318 ^ 1'b0 ;
  assign n41624 = ( x230 & n7318 ) | ( x230 & ~n41622 ) | ( n7318 & ~n41622 ) ;
  assign n41625 = ( x230 & ~n41623 ) | ( x230 & n41624 ) | ( ~n41623 & n41624 ) ;
  assign n41626 = ~x659 & n38462 ;
  assign n41627 = x274 & ~n38462 ;
  assign n41628 = ( x1091 & ~n41626 ) | ( x1091 & n41627 ) | ( ~n41626 & n41627 ) ;
  assign n41629 = n41626 | n41628 ;
  assign n41630 = x219 & ~n41420 ;
  assign n41631 = n41629 & n41630 ;
  assign n41632 = ~x659 & n38479 ;
  assign n41633 = x1091 | n41632 ;
  assign n41634 = n38479 & ~n41633 ;
  assign n41635 = ( x274 & n41633 ) | ( x274 & ~n41634 ) | ( n41633 & ~n41634 ) ;
  assign n41636 = ~n40804 & n41635 ;
  assign n41637 = x211 | n41636 ;
  assign n41638 = ~n40845 & n41635 ;
  assign n41639 = x211 & ~n41638 ;
  assign n41640 = ( x219 & n41637 ) | ( x219 & ~n41639 ) | ( n41637 & ~n41639 ) ;
  assign n41641 = ~x219 & n41640 ;
  assign n41642 = ( n15098 & n41631 ) | ( n15098 & ~n41641 ) | ( n41631 & ~n41641 ) ;
  assign n41643 = ~n41631 & n41642 ;
  assign n41644 = ~x200 & n41430 ;
  assign n41645 = ( x199 & n41629 ) | ( x199 & n41644 ) | ( n41629 & n41644 ) ;
  assign n41646 = ~n41644 & n41645 ;
  assign n41647 = x200 | n41636 ;
  assign n41648 = x200 & ~n41638 ;
  assign n41649 = ( x199 & n41647 ) | ( x199 & ~n41648 ) | ( n41647 & ~n41648 ) ;
  assign n41650 = ~x199 & n41649 ;
  assign n41651 = ( n15098 & ~n41646 ) | ( n15098 & n41650 ) | ( ~n41646 & n41650 ) ;
  assign n41652 = n41646 | n41651 ;
  assign n41653 = ( x230 & ~n41643 ) | ( x230 & n41652 ) | ( ~n41643 & n41652 ) ;
  assign n41654 = ~x230 & n41653 ;
  assign n41655 = n37643 & n41616 ;
  assign n41656 = ~n41654 & n41655 ;
  assign n41657 = ( n41625 & n41654 ) | ( n41625 & ~n41656 ) | ( n41654 & ~n41656 ) ;
  assign n41658 = x1149 & n41160 ;
  assign n41659 = x1151 & ~n41156 ;
  assign n41660 = n41658 & ~n41659 ;
  assign n41661 = n41156 & n41443 ;
  assign n41662 = n38354 & n40039 ;
  assign n41663 = x1151 | n41141 ;
  assign n41664 = x1150 & ~n41149 ;
  assign n41665 = n41663 & n41664 ;
  assign n41666 = ( x1149 & ~n41662 ) | ( x1149 & n41665 ) | ( ~n41662 & n41665 ) ;
  assign n41667 = n41662 | n41666 ;
  assign n41668 = ( n41660 & ~n41661 ) | ( n41660 & n41667 ) | ( ~n41661 & n41667 ) ;
  assign n41669 = ~n41660 & n41668 ;
  assign n41670 = n41525 ^ n41521 ^ n41276 ;
  assign n41671 = x1151 & n41670 ;
  assign n41672 = n41526 ^ n41522 ^ n41290 ;
  assign n41673 = ~x1151 & n41672 ;
  assign n41674 = ( x275 & n41671 ) | ( x275 & ~n41673 ) | ( n41671 & ~n41673 ) ;
  assign n41675 = ~n41671 & n41674 ;
  assign n41676 = x1151 & ~n41490 ;
  assign n41677 = x1150 | n41186 ;
  assign n41678 = n41676 & n41677 ;
  assign n41679 = ~x1151 & n41486 ;
  assign n41680 = x1150 & ~n41204 ;
  assign n41681 = n41679 & ~n41680 ;
  assign n41682 = ( ~x275 & n41678 ) | ( ~x275 & n41681 ) | ( n41678 & n41681 ) ;
  assign n41683 = ~x275 & n41682 ;
  assign n41684 = ( x1149 & ~n41675 ) | ( x1149 & n41683 ) | ( ~n41675 & n41683 ) ;
  assign n41685 = n41675 | n41684 ;
  assign n41686 = x1151 & ~n41476 ;
  assign n41687 = ~x1150 & n41222 ;
  assign n41688 = n41686 & ~n41687 ;
  assign n41689 = x1150 & n41257 ;
  assign n41690 = ( x1151 & n41481 ) | ( x1151 & ~n41689 ) | ( n41481 & ~n41689 ) ;
  assign n41691 = n41689 | n41690 ;
  assign n41692 = ( x275 & ~n41688 ) | ( x275 & n41691 ) | ( ~n41688 & n41691 ) ;
  assign n41693 = ~x275 & n41692 ;
  assign n41694 = x1151 & ~n41245 ;
  assign n41695 = ( x1150 & n41265 ) | ( x1150 & ~n41694 ) | ( n41265 & ~n41694 ) ;
  assign n41696 = ~x1150 & n41695 ;
  assign n41697 = x1150 & ~n41240 ;
  assign n41698 = n41261 & n41697 ;
  assign n41699 = ( x275 & n41696 ) | ( x275 & ~n41698 ) | ( n41696 & ~n41698 ) ;
  assign n41700 = ~n41696 & n41699 ;
  assign n41701 = ( x1149 & n41693 ) | ( x1149 & ~n41700 ) | ( n41693 & ~n41700 ) ;
  assign n41702 = ~n41693 & n41701 ;
  assign n41703 = n38504 & ~n41702 ;
  assign n41704 = n41685 & n41703 ;
  assign n41705 = ~x1151 & n39082 ;
  assign n41706 = n41510 & n41705 ;
  assign n41707 = ~x1149 & n41149 ;
  assign n41708 = n41660 | n41707 ;
  assign n41709 = x1150 & n41708 ;
  assign n41710 = ~x1149 & x1151 ;
  assign n41711 = n40039 & n41710 ;
  assign n41712 = x1149 & ~n41156 ;
  assign n41713 = ~x1151 & n41450 ;
  assign n41714 = n41712 & ~n41713 ;
  assign n41715 = ( x1150 & ~n41711 ) | ( x1150 & n41714 ) | ( ~n41711 & n41714 ) ;
  assign n41716 = n41711 | n41715 ;
  assign n41717 = x1091 & ~n41716 ;
  assign n41718 = ( x1091 & n41709 ) | ( x1091 & n41717 ) | ( n41709 & n41717 ) ;
  assign n41719 = ( x275 & n41706 ) | ( x275 & n41718 ) | ( n41706 & n41718 ) ;
  assign n41720 = n41718 ^ n41706 ^ 1'b0 ;
  assign n41721 = ( x275 & n41719 ) | ( x275 & n41720 ) | ( n41719 & n41720 ) ;
  assign n41722 = x1091 & n41669 ;
  assign n41723 = x275 | n41722 ;
  assign n41724 = ~n38504 & n41723 ;
  assign n41725 = ( n41704 & ~n41721 ) | ( n41704 & n41724 ) | ( ~n41721 & n41724 ) ;
  assign n41726 = n41721 ^ n41704 ^ 1'b0 ;
  assign n41727 = ( n41704 & n41725 ) | ( n41704 & ~n41726 ) | ( n41725 & ~n41726 ) ;
  assign n41728 = n41669 ^ x230 ^ 1'b0 ;
  assign n41729 = ( n41669 & n41727 ) | ( n41669 & ~n41728 ) | ( n41727 & ~n41728 ) ;
  assign n41730 = n35993 | n37919 ;
  assign n41731 = ~n37908 & n41730 ;
  assign n41732 = ( x230 & n15098 ) | ( x230 & n41731 ) | ( n15098 & n41731 ) ;
  assign n41733 = n41731 ^ n15098 ^ 1'b0 ;
  assign n41734 = ( x230 & n41732 ) | ( x230 & n41733 ) | ( n41732 & n41733 ) ;
  assign n41735 = x276 | n38463 ;
  assign n41736 = ~n41232 & n41735 ;
  assign n41737 = x199 & ~n41565 ;
  assign n41738 = ~n15098 & n41737 ;
  assign n41739 = n41159 & ~n41418 ;
  assign n41740 = ( ~n41736 & n41738 ) | ( ~n41736 & n41739 ) | ( n41738 & n41739 ) ;
  assign n41741 = ~n41736 & n41740 ;
  assign n41742 = x1145 & n38701 ;
  assign n41743 = ( n40846 & n41158 ) | ( n40846 & ~n41742 ) | ( n41158 & ~n41742 ) ;
  assign n41744 = n41742 | n41743 ;
  assign n41745 = n36054 | n37633 ;
  assign n41746 = x1091 & n41745 ;
  assign n41747 = n41746 ^ n41744 ^ 1'b0 ;
  assign n41748 = ( ~n37869 & n41746 ) | ( ~n37869 & n41747 ) | ( n41746 & n41747 ) ;
  assign n41749 = ( n41744 & ~n41747 ) | ( n41744 & n41748 ) | ( ~n41747 & n41748 ) ;
  assign n41750 = x276 | n38480 ;
  assign n41751 = ( ~n41415 & n41749 ) | ( ~n41415 & n41750 ) | ( n41749 & n41750 ) ;
  assign n41752 = n41749 ^ n41415 ^ 1'b0 ;
  assign n41753 = ( n41749 & n41751 ) | ( n41749 & ~n41752 ) | ( n41751 & ~n41752 ) ;
  assign n41754 = ( x230 & ~n41741 ) | ( x230 & n41753 ) | ( ~n41741 & n41753 ) ;
  assign n41755 = ~x230 & n41754 ;
  assign n41756 = ~x219 & n41745 ;
  assign n41757 = x1146 & n38496 ;
  assign n41758 = ( n15098 & n41756 ) | ( n15098 & ~n41757 ) | ( n41756 & ~n41757 ) ;
  assign n41759 = ~n41756 & n41758 ;
  assign n41760 = ~n41755 & n41759 ;
  assign n41761 = ( n41734 & n41755 ) | ( n41734 & ~n41760 ) | ( n41755 & ~n41760 ) ;
  assign n41762 = n35992 | n41387 ;
  assign n41763 = x200 & ~n40772 ;
  assign n41764 = ( n15098 & n41762 ) | ( n15098 & ~n41763 ) | ( n41762 & ~n41763 ) ;
  assign n41765 = n41764 ^ n41762 ^ 1'b0 ;
  assign n41766 = ( n15098 & n41764 ) | ( n15098 & ~n41765 ) | ( n41764 & ~n41765 ) ;
  assign n41767 = x219 & ~n40813 ;
  assign n41768 = ~x211 & x1140 ;
  assign n41769 = x211 & x1141 ;
  assign n41770 = x219 | n41769 ;
  assign n41771 = ( ~n41767 & n41768 ) | ( ~n41767 & n41770 ) | ( n41768 & n41770 ) ;
  assign n41772 = ~n41767 & n41771 ;
  assign n41773 = ( x299 & n7318 ) | ( x299 & ~n41772 ) | ( n7318 & ~n41772 ) ;
  assign n41774 = ~n41772 & n41773 ;
  assign n41775 = x230 & ~n41774 ;
  assign n41776 = n41766 & n41775 ;
  assign n41777 = ~x820 & n38479 ;
  assign n41778 = x1091 | n41777 ;
  assign n41779 = n38479 & ~n41778 ;
  assign n41780 = ( x277 & n41778 ) | ( x277 & ~n41779 ) | ( n41778 & ~n41779 ) ;
  assign n41781 = ~n41376 & n41780 ;
  assign n41782 = x211 | n41781 ;
  assign n41783 = ~n40782 & n41780 ;
  assign n41784 = x211 & ~n41783 ;
  assign n41785 = ( x219 & n41782 ) | ( x219 & ~n41784 ) | ( n41782 & ~n41784 ) ;
  assign n41786 = ~x219 & n41785 ;
  assign n41787 = ~x820 & n38462 ;
  assign n41788 = x1091 | n41787 ;
  assign n41789 = n38462 & ~n41788 ;
  assign n41790 = ( x277 & n41788 ) | ( x277 & ~n41789 ) | ( n41788 & ~n41789 ) ;
  assign n41791 = n40794 | n41767 ;
  assign n41792 = n41790 & n41791 ;
  assign n41793 = ( n15098 & n41786 ) | ( n15098 & ~n41792 ) | ( n41786 & ~n41792 ) ;
  assign n41794 = ~n41786 & n41793 ;
  assign n41795 = x200 | n41781 ;
  assign n41796 = x200 & ~n41783 ;
  assign n41797 = ( x199 & n41795 ) | ( x199 & ~n41796 ) | ( n41795 & ~n41796 ) ;
  assign n41798 = ~x199 & n41797 ;
  assign n41799 = n41790 ^ n15098 ^ 1'b0 ;
  assign n41800 = ~x200 & n40785 ;
  assign n41801 = x199 & ~n41800 ;
  assign n41802 = ( n41790 & ~n41799 ) | ( n41790 & n41801 ) | ( ~n41799 & n41801 ) ;
  assign n41803 = ( n15098 & n41799 ) | ( n15098 & n41802 ) | ( n41799 & n41802 ) ;
  assign n41804 = ( ~n41794 & n41798 ) | ( ~n41794 & n41803 ) | ( n41798 & n41803 ) ;
  assign n41805 = ~n41794 & n41804 ;
  assign n41806 = ( x230 & ~n41776 ) | ( x230 & n41805 ) | ( ~n41776 & n41805 ) ;
  assign n41807 = ~n41776 & n41806 ;
  assign n41808 = ~x199 & x1133 ;
  assign n41809 = x200 & ~n41808 ;
  assign n41810 = x299 | n41809 ;
  assign n41811 = ~x199 & x1132 ;
  assign n41812 = x200 | n41811 ;
  assign n41813 = ~n41810 & n41812 ;
  assign n41814 = x1132 ^ x211 ^ 1'b0 ;
  assign n41815 = ( x1132 & x1133 ) | ( x1132 & n41814 ) | ( x1133 & n41814 ) ;
  assign n41816 = n36026 & n41815 ;
  assign n41817 = ( ~n7318 & n41813 ) | ( ~n7318 & n41816 ) | ( n41813 & n41816 ) ;
  assign n41818 = ~n7318 & n41817 ;
  assign n41819 = n37211 & n41815 ;
  assign n41820 = ( x230 & n41818 ) | ( x230 & ~n41819 ) | ( n41818 & ~n41819 ) ;
  assign n41821 = ~n41818 & n41820 ;
  assign n41822 = ~x976 & n38462 ;
  assign n41823 = x278 | n38462 ;
  assign n41824 = ( x1091 & ~n41822 ) | ( x1091 & n41823 ) | ( ~n41822 & n41823 ) ;
  assign n41825 = ~x1091 & n41824 ;
  assign n41826 = x199 & ~n41825 ;
  assign n41827 = x1091 & ~x1132 ;
  assign n41828 = x976 & n38479 ;
  assign n41829 = x1091 | n41828 ;
  assign n41830 = n38479 & ~n41829 ;
  assign n41831 = ( x278 & n41829 ) | ( x278 & ~n41830 ) | ( n41829 & ~n41830 ) ;
  assign n41832 = ~n41827 & n41831 ;
  assign n41833 = x199 | n41832 ;
  assign n41834 = n41833 ^ n41826 ^ 1'b0 ;
  assign n41835 = ( n41826 & n41833 ) | ( n41826 & n41834 ) | ( n41833 & n41834 ) ;
  assign n41836 = ( x200 & ~n41826 ) | ( x200 & n41835 ) | ( ~n41826 & n41835 ) ;
  assign n41837 = n41825 ^ x199 ^ 1'b0 ;
  assign n41838 = x1091 & ~x1133 ;
  assign n41839 = n41831 & ~n41838 ;
  assign n41840 = ( n41825 & ~n41837 ) | ( n41825 & n41839 ) | ( ~n41837 & n41839 ) ;
  assign n41841 = ( x200 & x299 ) | ( x200 & ~n41840 ) | ( x299 & ~n41840 ) ;
  assign n41842 = n41840 ^ x299 ^ 1'b0 ;
  assign n41843 = ( x299 & n41841 ) | ( x299 & ~n41842 ) | ( n41841 & ~n41842 ) ;
  assign n41844 = n41836 & ~n41843 ;
  assign n41845 = x1091 & ~n41815 ;
  assign n41846 = n41831 & ~n41845 ;
  assign n41847 = n41825 ^ x219 ^ 1'b0 ;
  assign n41848 = ( n41825 & n41846 ) | ( n41825 & ~n41847 ) | ( n41846 & ~n41847 ) ;
  assign n41849 = x299 & n41848 ;
  assign n41850 = ( ~n7318 & n41844 ) | ( ~n7318 & n41849 ) | ( n41844 & n41849 ) ;
  assign n41851 = ~n7318 & n41850 ;
  assign n41852 = n7318 & n41848 ;
  assign n41853 = x230 | n41852 ;
  assign n41854 = ( ~n41821 & n41851 ) | ( ~n41821 & n41853 ) | ( n41851 & n41853 ) ;
  assign n41855 = ~n41821 & n41854 ;
  assign n41860 = ( n37776 & n40038 ) | ( n37776 & n41815 ) | ( n40038 & n41815 ) ;
  assign n41856 = n40276 | n41816 ;
  assign n41857 = ( n9354 & ~n41810 ) | ( n9354 & n41813 ) | ( ~n41810 & n41813 ) ;
  assign n41858 = ( ~n7318 & n41856 ) | ( ~n7318 & n41857 ) | ( n41856 & n41857 ) ;
  assign n41859 = ~n7318 & n41858 ;
  assign n41861 = ( x230 & ~n41859 ) | ( x230 & n41860 ) | ( ~n41859 & n41860 ) ;
  assign n41862 = ~n41860 & n41861 ;
  assign n41863 = n11550 & n40233 ;
  assign n41864 = n41849 | n41863 ;
  assign n41865 = ( n38717 & ~n41843 ) | ( n38717 & n41844 ) | ( ~n41843 & n41844 ) ;
  assign n41866 = ( ~n7318 & n41864 ) | ( ~n7318 & n41865 ) | ( n41864 & n41865 ) ;
  assign n41867 = ~n7318 & n41866 ;
  assign n41868 = n41562 | n41853 ;
  assign n41869 = ( ~n41862 & n41867 ) | ( ~n41862 & n41868 ) | ( n41867 & n41868 ) ;
  assign n41870 = ~n41862 & n41869 ;
  assign n41871 = n41855 ^ x1134 ^ 1'b0 ;
  assign n41872 = ( n41855 & n41870 ) | ( n41855 & n41871 ) | ( n41870 & n41871 ) ;
  assign n41873 = x1135 & n38496 ;
  assign n41874 = ~x211 & x1133 ;
  assign n41875 = x211 | x1133 ;
  assign n41876 = ~x219 & n41875 ;
  assign n41877 = n41873 | n41876 ;
  assign n41878 = ( n41873 & n41874 ) | ( n41873 & n41877 ) | ( n41874 & n41877 ) ;
  assign n41879 = n7318 & n41878 ;
  assign n41880 = x299 & n41878 ;
  assign n41881 = x1133 ^ x199 ^ 1'b0 ;
  assign n41882 = ( x1133 & x1135 ) | ( x1133 & n41881 ) | ( x1135 & n41881 ) ;
  assign n41883 = ( x200 & ~x299 ) | ( x200 & n41882 ) | ( ~x299 & n41882 ) ;
  assign n41884 = ~x200 & n41883 ;
  assign n41885 = ( ~n7318 & n41880 ) | ( ~n7318 & n41884 ) | ( n41880 & n41884 ) ;
  assign n41886 = ~n7318 & n41885 ;
  assign n41887 = ( x230 & n41879 ) | ( x230 & ~n41886 ) | ( n41879 & ~n41886 ) ;
  assign n41888 = ~n41879 & n41887 ;
  assign n41889 = x958 & n38479 ;
  assign n41890 = x1091 | n41889 ;
  assign n41891 = n38479 & ~n41890 ;
  assign n41892 = ( x279 & n41890 ) | ( x279 & ~n41891 ) | ( n41890 & ~n41891 ) ;
  assign n41893 = ~x1133 & n41330 ;
  assign n41894 = x199 | n41893 ;
  assign n41895 = n41892 & ~n41894 ;
  assign n41896 = x279 | n38462 ;
  assign n41897 = ~x958 & n38462 ;
  assign n41898 = ( x1091 & n41896 ) | ( x1091 & ~n41897 ) | ( n41896 & ~n41897 ) ;
  assign n41899 = ~x1091 & n41898 ;
  assign n41900 = x1135 & n41330 ;
  assign n41901 = n41899 | n41900 ;
  assign n41902 = x199 & n41901 ;
  assign n41903 = ( ~n15098 & n41895 ) | ( ~n15098 & n41902 ) | ( n41895 & n41902 ) ;
  assign n41904 = ~n15098 & n41903 ;
  assign n41905 = ~n38701 & n41904 ;
  assign n41906 = x1091 & ~n41874 ;
  assign n41907 = ( x219 & n41892 ) | ( x219 & ~n41906 ) | ( n41892 & ~n41906 ) ;
  assign n41908 = n41907 ^ n41892 ^ 1'b0 ;
  assign n41909 = ( x219 & n41907 ) | ( x219 & ~n41908 ) | ( n41907 & ~n41908 ) ;
  assign n41910 = n41909 ^ x230 ^ 1'b0 ;
  assign n41911 = ( x219 & ~x1135 ) | ( x219 & n40794 ) | ( ~x1135 & n40794 ) ;
  assign n41912 = n41911 ^ n41899 ^ 1'b0 ;
  assign n41913 = ( n15098 & n41899 ) | ( n15098 & ~n41911 ) | ( n41899 & ~n41911 ) ;
  assign n41914 = ( n15098 & ~n41912 ) | ( n15098 & n41913 ) | ( ~n41912 & n41913 ) ;
  assign n41915 = ( n41909 & ~n41910 ) | ( n41909 & n41914 ) | ( ~n41910 & n41914 ) ;
  assign n41916 = ( x230 & n41910 ) | ( x230 & n41915 ) | ( n41910 & n41915 ) ;
  assign n41917 = ( ~n41888 & n41905 ) | ( ~n41888 & n41916 ) | ( n41905 & n41916 ) ;
  assign n41918 = ~n41888 & n41917 ;
  assign n41919 = n15098 & ~n41877 ;
  assign n41920 = ~x200 & x1135 ;
  assign n41921 = x199 & ~n41920 ;
  assign n41922 = x1133 | n9353 ;
  assign n41923 = n41922 ^ n41921 ^ 1'b0 ;
  assign n41924 = ( n41921 & n41922 ) | ( n41921 & n41923 ) | ( n41922 & n41923 ) ;
  assign n41925 = ( n15098 & ~n41921 ) | ( n15098 & n41924 ) | ( ~n41921 & n41924 ) ;
  assign n41926 = x230 & ~n41925 ;
  assign n41927 = ( x230 & n41919 ) | ( x230 & n41926 ) | ( n41919 & n41926 ) ;
  assign n41928 = x1091 & n41875 ;
  assign n41929 = n37869 & n41928 ;
  assign n41930 = n41904 | n41929 ;
  assign n41931 = ( n41916 & ~n41927 ) | ( n41916 & n41930 ) | ( ~n41927 & n41930 ) ;
  assign n41932 = ~n41927 & n41931 ;
  assign n41933 = n41918 ^ x1134 ^ 1'b0 ;
  assign n41934 = ( n41918 & n41932 ) | ( n41918 & n41933 ) | ( n41932 & n41933 ) ;
  assign n41935 = x200 & ~n41309 ;
  assign n41936 = x199 & x1137 ;
  assign n41937 = x200 | n40862 ;
  assign n41938 = ( ~n41935 & n41936 ) | ( ~n41935 & n41937 ) | ( n41936 & n41937 ) ;
  assign n41939 = ~n41935 & n41938 ;
  assign n41940 = n41939 ^ n15098 ^ 1'b0 ;
  assign n41941 = ( x230 & n15098 ) | ( x230 & ~n41939 ) | ( n15098 & ~n41939 ) ;
  assign n41942 = ( x230 & ~n41940 ) | ( x230 & n41941 ) | ( ~n41940 & n41941 ) ;
  assign n41943 = ( x1135 & x1136 ) | ( x1135 & ~n41316 ) | ( x1136 & ~n41316 ) ;
  assign n41944 = x1091 & ~n41943 ;
  assign n41945 = x914 & n38479 ;
  assign n41946 = x280 | n38479 ;
  assign n41947 = ( x1091 & ~n41945 ) | ( x1091 & n41946 ) | ( ~n41945 & n41946 ) ;
  assign n41948 = ~x1091 & n41947 ;
  assign n41949 = ( ~x219 & n41944 ) | ( ~x219 & n41948 ) | ( n41944 & n41948 ) ;
  assign n41950 = ~x219 & n41949 ;
  assign n41951 = ~x914 & n38462 ;
  assign n41952 = x1091 | n41951 ;
  assign n41953 = n38462 & ~n41952 ;
  assign n41954 = ( x280 & n41952 ) | ( x280 & ~n41953 ) | ( n41952 & ~n41953 ) ;
  assign n41955 = n41954 ^ n41950 ^ 1'b0 ;
  assign n41956 = ~x211 & x1137 ;
  assign n41957 = x219 & ~n41956 ;
  assign n41958 = n40794 | n41957 ;
  assign n41959 = ( n41954 & ~n41955 ) | ( n41954 & n41958 ) | ( ~n41955 & n41958 ) ;
  assign n41960 = ( n41950 & n41955 ) | ( n41950 & n41959 ) | ( n41955 & n41959 ) ;
  assign n41961 = ( n41320 & n41321 ) | ( n41320 & n41960 ) | ( n41321 & n41960 ) ;
  assign n41962 = x200 & x1136 ;
  assign n41963 = x1091 & ~n41920 ;
  assign n41964 = ~n41962 & n41963 ;
  assign n41965 = ( x199 & n41948 ) | ( x199 & ~n41964 ) | ( n41948 & ~n41964 ) ;
  assign n41966 = n41964 | n41965 ;
  assign n41967 = x1137 & n41330 ;
  assign n41968 = ( x199 & ~n41954 ) | ( x199 & n41967 ) | ( ~n41954 & n41967 ) ;
  assign n41969 = ( n15098 & n41966 ) | ( n15098 & ~n41968 ) | ( n41966 & ~n41968 ) ;
  assign n41970 = ~n15098 & n41969 ;
  assign n41971 = ( ~x230 & n41961 ) | ( ~x230 & n41970 ) | ( n41961 & n41970 ) ;
  assign n41972 = ~x230 & n41971 ;
  assign n41973 = n41943 ^ x219 ^ 1'b0 ;
  assign n41974 = ( n41943 & n41956 ) | ( n41943 & n41973 ) | ( n41956 & n41973 ) ;
  assign n41975 = ( n41320 & n41321 ) | ( n41320 & n41974 ) | ( n41321 & n41974 ) ;
  assign n41976 = ~n41972 & n41975 ;
  assign n41977 = ( n41942 & n41972 ) | ( n41942 & ~n41976 ) | ( n41972 & ~n41976 ) ;
  assign n41978 = ~x199 & x1138 ;
  assign n41979 = x200 & ~n41978 ;
  assign n41980 = x199 & x1139 ;
  assign n41981 = x200 | n41307 ;
  assign n41982 = n41980 | n41981 ;
  assign n41983 = ( n15098 & ~n41979 ) | ( n15098 & n41982 ) | ( ~n41979 & n41982 ) ;
  assign n41984 = ~n15098 & n41983 ;
  assign n41985 = ~x211 & x1139 ;
  assign n41986 = n41985 ^ x219 ^ 1'b0 ;
  assign n41987 = n41956 ^ n41315 ^ x1138 ;
  assign n41988 = ( n41985 & ~n41986 ) | ( n41985 & n41987 ) | ( ~n41986 & n41987 ) ;
  assign n41989 = ( n41320 & n41321 ) | ( n41320 & n41988 ) | ( n41321 & n41988 ) ;
  assign n41990 = ( x230 & n41984 ) | ( x230 & n41989 ) | ( n41984 & n41989 ) ;
  assign n41991 = n41989 ^ n41984 ^ 1'b0 ;
  assign n41992 = ( x230 & n41990 ) | ( x230 & n41991 ) | ( n41990 & n41991 ) ;
  assign n41993 = ~x830 & n38479 ;
  assign n41994 = x1091 | n41993 ;
  assign n41995 = n38479 & ~n41994 ;
  assign n41996 = ( x281 & n41994 ) | ( x281 & ~n41995 ) | ( n41994 & ~n41995 ) ;
  assign n41997 = ~x830 & n38462 ;
  assign n41998 = x281 & ~n38462 ;
  assign n41999 = ( x1091 & ~n41997 ) | ( x1091 & n41998 ) | ( ~n41997 & n41998 ) ;
  assign n42000 = n41997 | n41999 ;
  assign n42001 = x199 & ~n41378 ;
  assign n42002 = ~n15098 & n42001 ;
  assign n42003 = x1139 & n40233 ;
  assign n42004 = n41159 & ~n42003 ;
  assign n42005 = ( n42000 & n42002 ) | ( n42000 & n42004 ) | ( n42002 & n42004 ) ;
  assign n42006 = n42004 ^ n42002 ^ 1'b0 ;
  assign n42007 = ( n42000 & n42005 ) | ( n42000 & n42006 ) | ( n42005 & n42006 ) ;
  assign n42008 = x1091 & n41987 ;
  assign n42009 = n37869 & ~n42008 ;
  assign n42010 = x1138 & n38701 ;
  assign n42011 = n41967 | n42010 ;
  assign n42012 = n41158 | n42011 ;
  assign n42013 = ~n42009 & n42012 ;
  assign n42014 = ~n42007 & n42013 ;
  assign n42015 = ( n41996 & n42007 ) | ( n41996 & ~n42014 ) | ( n42007 & ~n42014 ) ;
  assign n42016 = ( x230 & ~n41992 ) | ( x230 & n42015 ) | ( ~n41992 & n42015 ) ;
  assign n42017 = ~n41992 & n42016 ;
  assign n42018 = x200 & ~n41389 ;
  assign n42019 = x199 & x1140 ;
  assign n42020 = x200 | n41978 ;
  assign n42021 = n42019 | n42020 ;
  assign n42022 = ( n15098 & ~n42018 ) | ( n15098 & n42021 ) | ( ~n42018 & n42021 ) ;
  assign n42023 = ~n15098 & n42022 ;
  assign n42024 = ( x1138 & x1139 ) | ( x1138 & ~n41372 ) | ( x1139 & ~n41372 ) ;
  assign n42025 = n41768 ^ x219 ^ 1'b0 ;
  assign n42026 = ( n41768 & n42024 ) | ( n41768 & ~n42025 ) | ( n42024 & ~n42025 ) ;
  assign n42027 = ( n41320 & n41321 ) | ( n41320 & n42026 ) | ( n41321 & n42026 ) ;
  assign n42028 = ( x230 & n42023 ) | ( x230 & n42027 ) | ( n42023 & n42027 ) ;
  assign n42029 = n42027 ^ n42023 ^ 1'b0 ;
  assign n42030 = ( x230 & n42028 ) | ( x230 & n42029 ) | ( n42028 & n42029 ) ;
  assign n42031 = ~x836 & n38479 ;
  assign n42032 = x1091 | n42031 ;
  assign n42033 = n38479 & ~n42032 ;
  assign n42034 = ( x282 & n42032 ) | ( x282 & ~n42033 ) | ( n42032 & ~n42033 ) ;
  assign n42035 = ~x836 & n38462 ;
  assign n42036 = x282 & ~n38462 ;
  assign n42037 = ( x1091 & ~n42035 ) | ( x1091 & n42036 ) | ( ~n42035 & n42036 ) ;
  assign n42038 = n42035 | n42037 ;
  assign n42039 = ( x199 & n15098 ) | ( x199 & ~n41377 ) | ( n15098 & ~n41377 ) ;
  assign n42040 = ~n15098 & n42039 ;
  assign n42041 = x1140 & n40233 ;
  assign n42042 = n41159 & ~n42041 ;
  assign n42043 = ( n42038 & n42040 ) | ( n42038 & n42042 ) | ( n42040 & n42042 ) ;
  assign n42044 = n42042 ^ n42040 ^ 1'b0 ;
  assign n42045 = ( n42038 & n42043 ) | ( n42038 & n42044 ) | ( n42043 & n42044 ) ;
  assign n42046 = x1091 & n42024 ;
  assign n42047 = n37869 & ~n42046 ;
  assign n42048 = x1139 & n38701 ;
  assign n42049 = n41331 | n42048 ;
  assign n42050 = n41158 | n42049 ;
  assign n42051 = ~n42047 & n42050 ;
  assign n42052 = ~n42045 & n42051 ;
  assign n42053 = ( n42034 & n42045 ) | ( n42034 & ~n42052 ) | ( n42045 & ~n42052 ) ;
  assign n42054 = ( x230 & ~n42030 ) | ( x230 & n42053 ) | ( ~n42030 & n42053 ) ;
  assign n42055 = ~n42030 & n42054 ;
  assign n42056 = x1147 & ~n41450 ;
  assign n42057 = x1149 & n40039 ;
  assign n42058 = ( ~x1148 & n42056 ) | ( ~x1148 & n42057 ) | ( n42056 & n42057 ) ;
  assign n42059 = ~x1148 & n42058 ;
  assign n42060 = n41460 & ~n42056 ;
  assign n42061 = x1149 | n41141 ;
  assign n42062 = x1147 & ~n41160 ;
  assign n42063 = n42061 | n42062 ;
  assign n42064 = ( x1148 & n42060 ) | ( x1148 & n42063 ) | ( n42060 & n42063 ) ;
  assign n42065 = ~n42060 & n42064 ;
  assign n42066 = ( x230 & n42059 ) | ( x230 & ~n42065 ) | ( n42059 & ~n42065 ) ;
  assign n42067 = ~n42059 & n42066 ;
  assign n42068 = x1147 | n41209 ;
  assign n42069 = x1147 & ~n41252 ;
  assign n42070 = ( x1149 & n42068 ) | ( x1149 & ~n42069 ) | ( n42068 & ~n42069 ) ;
  assign n42071 = ~x1149 & n42070 ;
  assign n42072 = x1147 & ~n41222 ;
  assign n42073 = x1147 | n41186 ;
  assign n42074 = ( x1149 & n42072 ) | ( x1149 & n42073 ) | ( n42072 & n42073 ) ;
  assign n42075 = ~n42072 & n42074 ;
  assign n42076 = ( x1148 & ~n42071 ) | ( x1148 & n42075 ) | ( ~n42071 & n42075 ) ;
  assign n42077 = n42071 | n42076 ;
  assign n42078 = x1147 & ~n41257 ;
  assign n42079 = x1149 | n42078 ;
  assign n42080 = ( x1147 & n41204 ) | ( x1147 & ~n42079 ) | ( n41204 & ~n42079 ) ;
  assign n42081 = ~n42079 & n42080 ;
  assign n42082 = x1147 & ~n41228 ;
  assign n42083 = x1147 | n41194 ;
  assign n42084 = ( x1149 & n42082 ) | ( x1149 & n42083 ) | ( n42082 & n42083 ) ;
  assign n42085 = ~n42082 & n42084 ;
  assign n42086 = ( x1148 & n42081 ) | ( x1148 & ~n42085 ) | ( n42081 & ~n42085 ) ;
  assign n42087 = ~n42081 & n42086 ;
  assign n42088 = ( x283 & n42077 ) | ( x283 & ~n42087 ) | ( n42077 & ~n42087 ) ;
  assign n42089 = ~x283 & n42088 ;
  assign n42090 = x1147 & n41255 ;
  assign n42091 = x1148 & ~n42090 ;
  assign n42092 = ~x1147 & n41290 ;
  assign n42093 = ( x1149 & n42091 ) | ( x1149 & ~n42092 ) | ( n42091 & ~n42092 ) ;
  assign n42094 = n42093 ^ n42091 ^ 1'b0 ;
  assign n42095 = ( x1149 & n42093 ) | ( x1149 & ~n42094 ) | ( n42093 & ~n42094 ) ;
  assign n42096 = x1147 & n41264 ;
  assign n42097 = ~x1147 & n41285 ;
  assign n42098 = ( x1148 & ~n42096 ) | ( x1148 & n42097 ) | ( ~n42096 & n42097 ) ;
  assign n42099 = n42096 | n42098 ;
  assign n42100 = x283 & ~n42099 ;
  assign n42101 = ( x283 & n42095 ) | ( x283 & n42100 ) | ( n42095 & n42100 ) ;
  assign n42102 = ~x1147 & n41281 ;
  assign n42103 = x1147 & n41239 ;
  assign n42104 = ( x1148 & n42102 ) | ( x1148 & ~n42103 ) | ( n42102 & ~n42103 ) ;
  assign n42105 = ~n42102 & n42104 ;
  assign n42106 = x1147 & n41245 ;
  assign n42107 = ~x1147 & n41276 ;
  assign n42108 = ( x1148 & ~n42106 ) | ( x1148 & n42107 ) | ( ~n42106 & n42107 ) ;
  assign n42109 = n42106 | n42108 ;
  assign n42110 = ( x1149 & n42105 ) | ( x1149 & n42109 ) | ( n42105 & n42109 ) ;
  assign n42111 = ~n42105 & n42110 ;
  assign n42112 = ( x230 & n42101 ) | ( x230 & ~n42111 ) | ( n42101 & ~n42111 ) ;
  assign n42113 = n42112 ^ n42101 ^ 1'b0 ;
  assign n42114 = ( x230 & n42112 ) | ( x230 & ~n42113 ) | ( n42112 & ~n42113 ) ;
  assign n42115 = ( ~n42067 & n42089 ) | ( ~n42067 & n42114 ) | ( n42089 & n42114 ) ;
  assign n42116 = ~n42067 & n42115 ;
  assign n42117 = x1143 & n40529 ;
  assign n42118 = n37871 & n42117 ;
  assign n42119 = ( x284 & n40529 ) | ( x284 & ~n42118 ) | ( n40529 & ~n42118 ) ;
  assign n42120 = ~n42118 & n42119 ;
  assign n42121 = ~n2070 & n8992 ;
  assign n42122 = ~n11179 & n42121 ;
  assign n42123 = x286 & n42122 ;
  assign n42124 = x288 & x289 ;
  assign n42125 = n42123 & n42124 ;
  assign n42126 = x285 & n42125 ;
  assign n42127 = n7318 | n42126 ;
  assign n42128 = ~n7318 & n42121 ;
  assign n42129 = ( x285 & n42125 ) | ( x285 & n42128 ) | ( n42125 & n42128 ) ;
  assign n42130 = ~n42127 & n42129 ;
  assign n42131 = ~n7318 & n42125 ;
  assign n42132 = ~x286 & n11179 ;
  assign n42133 = ~x288 & n42132 ;
  assign n42134 = ~x289 & n42133 ;
  assign n42135 = ( x285 & n42131 ) | ( x285 & ~n42134 ) | ( n42131 & ~n42134 ) ;
  assign n42136 = ~n42131 & n42135 ;
  assign n42137 = ( ~x793 & n42130 ) | ( ~x793 & n42136 ) | ( n42130 & n42136 ) ;
  assign n42138 = ~x793 & n42137 ;
  assign n42139 = ~x288 & n6611 ;
  assign n42140 = n11179 & n42139 ;
  assign n42141 = ~x286 & n42140 ;
  assign n42142 = ( ~x286 & n7318 ) | ( ~x286 & n42140 ) | ( n7318 & n42140 ) ;
  assign n42143 = ( x793 & ~n42141 ) | ( x793 & n42142 ) | ( ~n42141 & n42142 ) ;
  assign n42144 = x288 & ~n42123 ;
  assign n42145 = x286 | n42122 ;
  assign n42146 = n42144 & n42145 ;
  assign n42147 = ~n42121 & n42132 ;
  assign n42148 = n11179 & ~n42121 ;
  assign n42149 = x286 & ~n42148 ;
  assign n42150 = n42147 | n42149 ;
  assign n42151 = ( x288 & n6611 ) | ( x288 & n42150 ) | ( n6611 & n42150 ) ;
  assign n42152 = ~x288 & n42151 ;
  assign n42153 = ( x57 & n5193 ) | ( x57 & ~n42152 ) | ( n5193 & ~n42152 ) ;
  assign n42154 = n42152 | n42153 ;
  assign n42155 = ( ~n42143 & n42146 ) | ( ~n42143 & n42154 ) | ( n42146 & n42154 ) ;
  assign n42156 = ~n42143 & n42155 ;
  assign n42157 = ~x287 & x457 ;
  assign n42158 = x332 | n42157 ;
  assign n42159 = n11179 ^ x288 ^ 1'b0 ;
  assign n42160 = ( x288 & n42139 ) | ( x288 & n42159 ) | ( n42139 & n42159 ) ;
  assign n42161 = n42128 & n42160 ;
  assign n42162 = x793 | n42161 ;
  assign n42163 = ( n42128 & n42160 ) | ( n42128 & ~n42162 ) | ( n42160 & ~n42162 ) ;
  assign n42164 = ~n42162 & n42163 ;
  assign n42165 = x285 & ~x289 ;
  assign n42166 = n42133 & n42165 ;
  assign n42167 = ( ~x289 & n7318 ) | ( ~x289 & n42141 ) | ( n7318 & n42141 ) ;
  assign n42168 = ( x793 & ~n42166 ) | ( x793 & n42167 ) | ( ~n42166 & n42167 ) ;
  assign n42169 = ~x289 & n42144 ;
  assign n42170 = n42147 & n42165 ;
  assign n42171 = x289 & ~n42147 ;
  assign n42172 = ( x288 & ~n42170 ) | ( x288 & n42171 ) | ( ~n42170 & n42171 ) ;
  assign n42173 = n42170 | n42172 ;
  assign n42174 = ( n42125 & ~n42169 ) | ( n42125 & n42173 ) | ( ~n42169 & n42173 ) ;
  assign n42175 = ~n42125 & n42174 ;
  assign n42176 = ( n7318 & ~n42168 ) | ( n7318 & n42175 ) | ( ~n42168 & n42175 ) ;
  assign n42177 = ~n42168 & n42176 ;
  assign n42178 = x1048 ^ x476 ^ 1'b0 ;
  assign n42179 = ( x290 & x1048 ) | ( x290 & n42178 ) | ( x1048 & n42178 ) ;
  assign n42180 = x1049 ^ x476 ^ 1'b0 ;
  assign n42181 = ( x291 & x1049 ) | ( x291 & n42180 ) | ( x1049 & n42180 ) ;
  assign n42182 = x1084 ^ x476 ^ 1'b0 ;
  assign n42183 = ( x292 & x1084 ) | ( x292 & n42182 ) | ( x1084 & n42182 ) ;
  assign n42184 = x1059 ^ x476 ^ 1'b0 ;
  assign n42185 = ( x293 & x1059 ) | ( x293 & n42184 ) | ( x1059 & n42184 ) ;
  assign n42186 = x1072 ^ x476 ^ 1'b0 ;
  assign n42187 = ( x294 & x1072 ) | ( x294 & n42186 ) | ( x1072 & n42186 ) ;
  assign n42188 = x1053 ^ x476 ^ 1'b0 ;
  assign n42189 = ( x295 & x1053 ) | ( x295 & n42188 ) | ( x1053 & n42188 ) ;
  assign n42190 = x1037 ^ x476 ^ 1'b0 ;
  assign n42191 = ( x296 & x1037 ) | ( x296 & n42190 ) | ( x1037 & n42190 ) ;
  assign n42192 = x1044 ^ x476 ^ 1'b0 ;
  assign n42193 = ( x297 & x1044 ) | ( x297 & n42192 ) | ( x1044 & n42192 ) ;
  assign n42194 = x1044 ^ x478 ^ 1'b0 ;
  assign n42195 = ( x298 & x1044 ) | ( x298 & n42194 ) | ( x1044 & n42194 ) ;
  assign n42196 = x54 | n11639 ;
  assign n42197 = n11912 & ~n42196 ;
  assign n42198 = n1292 & ~n42197 ;
  assign n42199 = ( x54 & n42197 ) | ( x54 & ~n42198 ) | ( n42197 & ~n42198 ) ;
  assign n42200 = ( n2054 & ~n7448 ) | ( n2054 & n42199 ) | ( ~n7448 & n42199 ) ;
  assign n42201 = ~n2054 & n42200 ;
  assign n42202 = n9903 ^ x39 ^ 1'b0 ;
  assign n42203 = ( n9903 & n42201 ) | ( n9903 & ~n42202 ) | ( n42201 & ~n42202 ) ;
  assign n42204 = x57 & ~x59 ;
  assign n42205 = ~n8663 & n42204 ;
  assign n42206 = ~x312 & n42205 ;
  assign n42207 = x300 & ~n42206 ;
  assign n42208 = ~x300 & n42206 ;
  assign n42209 = x55 | n42208 ;
  assign n42210 = n42207 | n42209 ;
  assign n42211 = x301 | n42209 ;
  assign n42212 = ~x55 & x301 ;
  assign n42213 = n42208 & n42212 ;
  assign n42214 = n42211 & ~n42213 ;
  assign n42215 = ~x215 & n2125 ;
  assign n42216 = ~x273 & n42215 ;
  assign n42217 = x833 & n6810 ;
  assign n42218 = ~x937 & n42217 ;
  assign n42219 = n42216 | n42218 ;
  assign n42220 = ( n41320 & n41321 ) | ( n41320 & n42219 ) | ( n41321 & n42219 ) ;
  assign n42221 = x273 & n2161 ;
  assign n42222 = n4870 | n7318 ;
  assign n42223 = x937 & n2170 ;
  assign n42224 = ( ~n42221 & n42222 ) | ( ~n42221 & n42223 ) | ( n42222 & n42223 ) ;
  assign n42225 = n42221 | n42224 ;
  assign n42226 = ~n42220 & n42225 ;
  assign n42227 = ( n1359 & n42220 ) | ( n1359 & ~n42226 ) | ( n42220 & ~n42226 ) ;
  assign n42228 = ~n2264 & n15098 ;
  assign n42229 = n42225 & ~n42228 ;
  assign n42230 = ~n42227 & n42229 ;
  assign n42231 = ( x237 & n42227 ) | ( x237 & ~n42230 ) | ( n42227 & ~n42230 ) ;
  assign n42232 = ~n4865 & n15098 ;
  assign n42233 = n42222 & ~n42232 ;
  assign n42234 = ( ~x1148 & n42231 ) | ( ~x1148 & n42233 ) | ( n42231 & n42233 ) ;
  assign n42235 = n42231 ^ x1148 ^ 1'b0 ;
  assign n42236 = ( n42231 & n42234 ) | ( n42231 & ~n42235 ) | ( n42234 & ~n42235 ) ;
  assign n42237 = x1049 ^ x478 ^ 1'b0 ;
  assign n42238 = ( x303 & x1049 ) | ( x303 & n42237 ) | ( x1049 & n42237 ) ;
  assign n42239 = x1048 ^ x478 ^ 1'b0 ;
  assign n42240 = ( x304 & x1048 ) | ( x304 & n42239 ) | ( x1048 & n42239 ) ;
  assign n42241 = x1084 ^ x478 ^ 1'b0 ;
  assign n42242 = ( x305 & x1084 ) | ( x305 & n42241 ) | ( x1084 & n42241 ) ;
  assign n42243 = x1059 ^ x478 ^ 1'b0 ;
  assign n42244 = ( x306 & x1059 ) | ( x306 & n42243 ) | ( x1059 & n42243 ) ;
  assign n42245 = x1053 ^ x478 ^ 1'b0 ;
  assign n42246 = ( x307 & x1053 ) | ( x307 & n42245 ) | ( x1053 & n42245 ) ;
  assign n42247 = x1037 ^ x478 ^ 1'b0 ;
  assign n42248 = ( x308 & x1037 ) | ( x308 & n42247 ) | ( x1037 & n42247 ) ;
  assign n42249 = x1072 ^ x478 ^ 1'b0 ;
  assign n42250 = ( x309 & x1072 ) | ( x309 & n42249 ) | ( x1072 & n42249 ) ;
  assign n42251 = ~x271 & n2161 ;
  assign n42252 = x222 & ~x934 ;
  assign n42253 = n42251 | n42252 ;
  assign n42254 = n42222 | n42253 ;
  assign n42255 = n2263 & n42232 ;
  assign n42256 = x271 & n2125 ;
  assign n42257 = x934 & n2022 ;
  assign n42258 = n42256 | n42257 ;
  assign n42259 = n42255 & n42258 ;
  assign n42260 = ( n42228 & n42254 ) | ( n42228 & ~n42259 ) | ( n42254 & ~n42259 ) ;
  assign n42261 = ~n42228 & n42260 ;
  assign n42262 = n1359 & ~n42222 ;
  assign n42263 = n42255 | n42262 ;
  assign n42264 = ~x1147 & n42263 ;
  assign n42265 = ~n42261 & n42264 ;
  assign n42266 = n42232 & ~n42258 ;
  assign n42267 = n1360 | n15098 ;
  assign n42268 = x1147 & n42267 ;
  assign n42269 = ~n42222 & n42253 ;
  assign n42270 = ( n42266 & n42268 ) | ( n42266 & ~n42269 ) | ( n42268 & ~n42269 ) ;
  assign n42271 = ~n42266 & n42270 ;
  assign n42272 = ( x233 & n42265 ) | ( x233 & n42271 ) | ( n42265 & n42271 ) ;
  assign n42273 = n42271 ^ n42265 ^ 1'b0 ;
  assign n42274 = ( x233 & n42272 ) | ( x233 & n42273 ) | ( n42272 & n42273 ) ;
  assign n42275 = x1147 & n42233 ;
  assign n42276 = n42261 & ~n42275 ;
  assign n42277 = ( x233 & ~n42274 ) | ( x233 & n42276 ) | ( ~n42274 & n42276 ) ;
  assign n42278 = ~n42274 & n42277 ;
  assign n42279 = x55 | x311 ;
  assign n42280 = n42213 ^ x311 ^ 1'b0 ;
  assign n42281 = ( ~x311 & n42279 ) | ( ~x311 & n42280 ) | ( n42279 & n42280 ) ;
  assign n42282 = n42205 ^ x312 ^ 1'b0 ;
  assign n42283 = ~x55 & n42282 ;
  assign n42284 = n8966 | n11950 ;
  assign n42285 = n5023 & ~n11954 ;
  assign n42286 = ( n8761 & n42284 ) | ( n8761 & ~n42285 ) | ( n42284 & ~n42285 ) ;
  assign n42287 = ~n8761 & n42286 ;
  assign n42288 = x954 ^ x313 ^ 1'b0 ;
  assign n42289 = ( ~x313 & n42287 ) | ( ~x313 & n42288 ) | ( n42287 & n42288 ) ;
  assign n42290 = ~x39 & n13104 ;
  assign n42291 = ( n1205 & n2036 ) | ( n1205 & n13787 ) | ( n2036 & n13787 ) ;
  assign n42292 = ( ~n13897 & n42290 ) | ( ~n13897 & n42291 ) | ( n42290 & n42291 ) ;
  assign n42293 = ~n13897 & n42292 ;
  assign n42294 = ( n2096 & n8758 ) | ( n2096 & ~n42293 ) | ( n8758 & ~n42293 ) ;
  assign n42295 = n42293 | n42294 ;
  assign n42296 = n42295 ^ n13270 ^ 1'b0 ;
  assign n42297 = n5459 | n7448 ;
  assign n42298 = ( n13270 & n42296 ) | ( n13270 & ~n42297 ) | ( n42296 & ~n42297 ) ;
  assign n42299 = ( n42295 & ~n42296 ) | ( n42295 & n42298 ) | ( ~n42296 & n42298 ) ;
  assign n42300 = ( n13255 & n13256 ) | ( n13255 & ~n42299 ) | ( n13256 & ~n42299 ) ;
  assign n42301 = n42299 | n42300 ;
  assign n42302 = ~x340 & n42128 ;
  assign n42303 = n42302 ^ x1080 ^ 1'b0 ;
  assign n42304 = ( x315 & x1080 ) | ( x315 & ~n42303 ) | ( x1080 & ~n42303 ) ;
  assign n42305 = n42302 ^ x1047 ^ 1'b0 ;
  assign n42306 = ( x316 & x1047 ) | ( x316 & ~n42305 ) | ( x1047 & ~n42305 ) ;
  assign n42307 = ~x330 & n42128 ;
  assign n42308 = n42307 ^ x1078 ^ 1'b0 ;
  assign n42309 = ( x317 & x1078 ) | ( x317 & ~n42308 ) | ( x1078 & ~n42308 ) ;
  assign n42310 = ~x341 & n42128 ;
  assign n42311 = n42310 ^ x1074 ^ 1'b0 ;
  assign n42312 = ( x318 & x1074 ) | ( x318 & ~n42311 ) | ( x1074 & ~n42311 ) ;
  assign n42313 = n42310 ^ x1072 ^ 1'b0 ;
  assign n42314 = ( x319 & x1072 ) | ( x319 & ~n42313 ) | ( x1072 & ~n42313 ) ;
  assign n42315 = n42302 ^ x1048 ^ 1'b0 ;
  assign n42316 = ( x320 & x1048 ) | ( x320 & ~n42315 ) | ( x1048 & ~n42315 ) ;
  assign n42317 = n42302 ^ x1058 ^ 1'b0 ;
  assign n42318 = ( x321 & x1058 ) | ( x321 & ~n42317 ) | ( x1058 & ~n42317 ) ;
  assign n42319 = n42302 ^ x1051 ^ 1'b0 ;
  assign n42320 = ( x322 & x1051 ) | ( x322 & ~n42319 ) | ( x1051 & ~n42319 ) ;
  assign n42321 = n42302 ^ x1065 ^ 1'b0 ;
  assign n42322 = ( x323 & x1065 ) | ( x323 & ~n42321 ) | ( x1065 & ~n42321 ) ;
  assign n42323 = n42310 ^ x1086 ^ 1'b0 ;
  assign n42324 = ( x324 & x1086 ) | ( x324 & ~n42323 ) | ( x1086 & ~n42323 ) ;
  assign n42325 = n42310 ^ x1063 ^ 1'b0 ;
  assign n42326 = ( x325 & x1063 ) | ( x325 & ~n42325 ) | ( x1063 & ~n42325 ) ;
  assign n42327 = n42310 ^ x1057 ^ 1'b0 ;
  assign n42328 = ( x326 & x1057 ) | ( x326 & ~n42327 ) | ( x1057 & ~n42327 ) ;
  assign n42329 = n42302 ^ x1040 ^ 1'b0 ;
  assign n42330 = ( x327 & x1040 ) | ( x327 & ~n42329 ) | ( x1040 & ~n42329 ) ;
  assign n42331 = n42310 ^ x1058 ^ 1'b0 ;
  assign n42332 = ( x328 & x1058 ) | ( x328 & ~n42331 ) | ( x1058 & ~n42331 ) ;
  assign n42333 = n42310 ^ x1043 ^ 1'b0 ;
  assign n42334 = ( x329 & x1043 ) | ( x329 & ~n42333 ) | ( x1043 & ~n42333 ) ;
  assign n42335 = x1092 & ~n8670 ;
  assign n42336 = n42121 ^ x340 ^ 1'b0 ;
  assign n42337 = ( x330 & x340 ) | ( x330 & ~n42336 ) | ( x340 & ~n42336 ) ;
  assign n42338 = ( n7318 & n42335 ) | ( n7318 & ~n42337 ) | ( n42335 & ~n42337 ) ;
  assign n42339 = ~n7318 & n42338 ;
  assign n42340 = n7318 & n42335 ;
  assign n42341 = ( ~x330 & n42339 ) | ( ~x330 & n42340 ) | ( n42339 & n42340 ) ;
  assign n42342 = n42339 ^ x330 ^ 1'b0 ;
  assign n42343 = ( n42339 & n42341 ) | ( n42339 & ~n42342 ) | ( n42341 & ~n42342 ) ;
  assign n42344 = n42121 ^ x341 ^ 1'b0 ;
  assign n42345 = ( x331 & x341 ) | ( x331 & ~n42344 ) | ( x341 & ~n42344 ) ;
  assign n42346 = ( n7318 & n42335 ) | ( n7318 & ~n42345 ) | ( n42335 & ~n42345 ) ;
  assign n42347 = ~n7318 & n42346 ;
  assign n42348 = ( ~x331 & n42340 ) | ( ~x331 & n42347 ) | ( n42340 & n42347 ) ;
  assign n42349 = n42347 ^ x331 ^ 1'b0 ;
  assign n42350 = ( n42347 & n42348 ) | ( n42347 & ~n42349 ) | ( n42348 & ~n42349 ) ;
  assign n42351 = x39 & n8962 ;
  assign n42352 = n9608 & ~n11657 ;
  assign n42353 = x332 & ~n8108 ;
  assign n42354 = n9608 | n11592 ;
  assign n42355 = ~n6387 & n42354 ;
  assign n42356 = x70 | n42355 ;
  assign n42357 = n42353 & n42356 ;
  assign n42358 = ( ~x39 & n42352 ) | ( ~x39 & n42357 ) | ( n42352 & n42357 ) ;
  assign n42359 = ~x39 & n42358 ;
  assign n42360 = ( x38 & ~n42351 ) | ( x38 & n42359 ) | ( ~n42351 & n42359 ) ;
  assign n42361 = n42351 | n42360 ;
  assign n42362 = ( n5053 & ~n8793 ) | ( n5053 & n42361 ) | ( ~n8793 & n42361 ) ;
  assign n42363 = ~n5053 & n42362 ;
  assign n42364 = n42310 ^ x1040 ^ 1'b0 ;
  assign n42365 = ( x333 & x1040 ) | ( x333 & ~n42364 ) | ( x1040 & ~n42364 ) ;
  assign n42366 = n42310 ^ x1065 ^ 1'b0 ;
  assign n42367 = ( x334 & x1065 ) | ( x334 & ~n42366 ) | ( x1065 & ~n42366 ) ;
  assign n42368 = n42310 ^ x1069 ^ 1'b0 ;
  assign n42369 = ( x335 & x1069 ) | ( x335 & ~n42368 ) | ( x1069 & ~n42368 ) ;
  assign n42370 = n42307 ^ x1070 ^ 1'b0 ;
  assign n42371 = ( x336 & x1070 ) | ( x336 & ~n42370 ) | ( x1070 & ~n42370 ) ;
  assign n42372 = n42307 ^ x1044 ^ 1'b0 ;
  assign n42373 = ( x337 & x1044 ) | ( x337 & ~n42372 ) | ( x1044 & ~n42372 ) ;
  assign n42374 = n42307 ^ x1072 ^ 1'b0 ;
  assign n42375 = ( x338 & x1072 ) | ( x338 & ~n42374 ) | ( x1072 & ~n42374 ) ;
  assign n42376 = n42307 ^ x1086 ^ 1'b0 ;
  assign n42377 = ( x339 & x1086 ) | ( x339 & ~n42376 ) | ( x1086 & ~n42376 ) ;
  assign n42378 = ~x331 & n42121 ;
  assign n42379 = ~n7318 & n42335 ;
  assign n42380 = x340 | n42121 ;
  assign n42381 = n42379 & n42380 ;
  assign n42382 = ~n42378 & n42381 ;
  assign n42383 = n42382 ^ x340 ^ 1'b0 ;
  assign n42384 = ( ~x340 & n42340 ) | ( ~x340 & n42383 ) | ( n42340 & n42383 ) ;
  assign n42385 = ( x340 & n42382 ) | ( x340 & n42384 ) | ( n42382 & n42384 ) ;
  assign n42386 = n42310 ^ n42307 ^ x341 ;
  assign n42387 = ( x1092 & n8670 ) | ( x1092 & ~n42386 ) | ( n8670 & ~n42386 ) ;
  assign n42388 = ~n8670 & n42387 ;
  assign n42389 = n42302 ^ x1049 ^ 1'b0 ;
  assign n42390 = ( x342 & x1049 ) | ( x342 & ~n42389 ) | ( x1049 & ~n42389 ) ;
  assign n42391 = n42302 ^ x1062 ^ 1'b0 ;
  assign n42392 = ( x343 & x1062 ) | ( x343 & ~n42391 ) | ( x1062 & ~n42391 ) ;
  assign n42393 = n42302 ^ x1069 ^ 1'b0 ;
  assign n42394 = ( x344 & x1069 ) | ( x344 & ~n42393 ) | ( x1069 & ~n42393 ) ;
  assign n42395 = n42302 ^ x1039 ^ 1'b0 ;
  assign n42396 = ( x345 & x1039 ) | ( x345 & ~n42395 ) | ( x1039 & ~n42395 ) ;
  assign n42397 = n42302 ^ x1067 ^ 1'b0 ;
  assign n42398 = ( x346 & x1067 ) | ( x346 & ~n42397 ) | ( x1067 & ~n42397 ) ;
  assign n42399 = n42302 ^ x1055 ^ 1'b0 ;
  assign n42400 = ( x347 & x1055 ) | ( x347 & ~n42399 ) | ( x1055 & ~n42399 ) ;
  assign n42401 = n42302 ^ x1087 ^ 1'b0 ;
  assign n42402 = ( x348 & x1087 ) | ( x348 & ~n42401 ) | ( x1087 & ~n42401 ) ;
  assign n42403 = n42302 ^ x1043 ^ 1'b0 ;
  assign n42404 = ( x349 & x1043 ) | ( x349 & ~n42403 ) | ( x1043 & ~n42403 ) ;
  assign n42405 = n42302 ^ x1035 ^ 1'b0 ;
  assign n42406 = ( x350 & x1035 ) | ( x350 & ~n42405 ) | ( x1035 & ~n42405 ) ;
  assign n42407 = n42302 ^ x1079 ^ 1'b0 ;
  assign n42408 = ( x351 & x1079 ) | ( x351 & ~n42407 ) | ( x1079 & ~n42407 ) ;
  assign n42409 = n42302 ^ x1078 ^ 1'b0 ;
  assign n42410 = ( x352 & x1078 ) | ( x352 & ~n42409 ) | ( x1078 & ~n42409 ) ;
  assign n42411 = n42302 ^ x1063 ^ 1'b0 ;
  assign n42412 = ( x353 & x1063 ) | ( x353 & ~n42411 ) | ( x1063 & ~n42411 ) ;
  assign n42413 = n42302 ^ x1045 ^ 1'b0 ;
  assign n42414 = ( x354 & x1045 ) | ( x354 & ~n42413 ) | ( x1045 & ~n42413 ) ;
  assign n42415 = n42302 ^ x1084 ^ 1'b0 ;
  assign n42416 = ( x355 & x1084 ) | ( x355 & ~n42415 ) | ( x1084 & ~n42415 ) ;
  assign n42417 = n42302 ^ x1081 ^ 1'b0 ;
  assign n42418 = ( x356 & x1081 ) | ( x356 & ~n42417 ) | ( x1081 & ~n42417 ) ;
  assign n42419 = n42302 ^ x1076 ^ 1'b0 ;
  assign n42420 = ( x357 & x1076 ) | ( x357 & ~n42419 ) | ( x1076 & ~n42419 ) ;
  assign n42421 = n42302 ^ x1071 ^ 1'b0 ;
  assign n42422 = ( x358 & x1071 ) | ( x358 & ~n42421 ) | ( x1071 & ~n42421 ) ;
  assign n42423 = n42302 ^ x1068 ^ 1'b0 ;
  assign n42424 = ( x359 & x1068 ) | ( x359 & ~n42423 ) | ( x1068 & ~n42423 ) ;
  assign n42425 = n42302 ^ x1042 ^ 1'b0 ;
  assign n42426 = ( x360 & x1042 ) | ( x360 & ~n42425 ) | ( x1042 & ~n42425 ) ;
  assign n42427 = n42302 ^ x1059 ^ 1'b0 ;
  assign n42428 = ( x361 & x1059 ) | ( x361 & ~n42427 ) | ( x1059 & ~n42427 ) ;
  assign n42429 = n42302 ^ x1070 ^ 1'b0 ;
  assign n42430 = ( x362 & x1070 ) | ( x362 & ~n42429 ) | ( x1070 & ~n42429 ) ;
  assign n42431 = n42307 ^ x1049 ^ 1'b0 ;
  assign n42432 = ( x363 & x1049 ) | ( x363 & ~n42431 ) | ( x1049 & ~n42431 ) ;
  assign n42433 = n42307 ^ x1062 ^ 1'b0 ;
  assign n42434 = ( x364 & x1062 ) | ( x364 & ~n42433 ) | ( x1062 & ~n42433 ) ;
  assign n42435 = n42307 ^ x1065 ^ 1'b0 ;
  assign n42436 = ( x365 & x1065 ) | ( x365 & ~n42435 ) | ( x1065 & ~n42435 ) ;
  assign n42437 = n42307 ^ x1069 ^ 1'b0 ;
  assign n42438 = ( x366 & x1069 ) | ( x366 & ~n42437 ) | ( x1069 & ~n42437 ) ;
  assign n42439 = n42307 ^ x1039 ^ 1'b0 ;
  assign n42440 = ( x367 & x1039 ) | ( x367 & ~n42439 ) | ( x1039 & ~n42439 ) ;
  assign n42441 = n42307 ^ x1067 ^ 1'b0 ;
  assign n42442 = ( x368 & x1067 ) | ( x368 & ~n42441 ) | ( x1067 & ~n42441 ) ;
  assign n42443 = n42307 ^ x1080 ^ 1'b0 ;
  assign n42444 = ( x369 & x1080 ) | ( x369 & ~n42443 ) | ( x1080 & ~n42443 ) ;
  assign n42445 = n42307 ^ x1055 ^ 1'b0 ;
  assign n42446 = ( x370 & x1055 ) | ( x370 & ~n42445 ) | ( x1055 & ~n42445 ) ;
  assign n42447 = n42307 ^ x1051 ^ 1'b0 ;
  assign n42448 = ( x371 & x1051 ) | ( x371 & ~n42447 ) | ( x1051 & ~n42447 ) ;
  assign n42449 = n42307 ^ x1048 ^ 1'b0 ;
  assign n42450 = ( x372 & x1048 ) | ( x372 & ~n42449 ) | ( x1048 & ~n42449 ) ;
  assign n42451 = n42307 ^ x1087 ^ 1'b0 ;
  assign n42452 = ( x373 & x1087 ) | ( x373 & ~n42451 ) | ( x1087 & ~n42451 ) ;
  assign n42453 = n42307 ^ x1035 ^ 1'b0 ;
  assign n42454 = ( x374 & x1035 ) | ( x374 & ~n42453 ) | ( x1035 & ~n42453 ) ;
  assign n42455 = n42307 ^ x1047 ^ 1'b0 ;
  assign n42456 = ( x375 & x1047 ) | ( x375 & ~n42455 ) | ( x1047 & ~n42455 ) ;
  assign n42457 = n42307 ^ x1079 ^ 1'b0 ;
  assign n42458 = ( x376 & x1079 ) | ( x376 & ~n42457 ) | ( x1079 & ~n42457 ) ;
  assign n42459 = n42307 ^ x1074 ^ 1'b0 ;
  assign n42460 = ( x377 & x1074 ) | ( x377 & ~n42459 ) | ( x1074 & ~n42459 ) ;
  assign n42461 = n42307 ^ x1063 ^ 1'b0 ;
  assign n42462 = ( x378 & x1063 ) | ( x378 & ~n42461 ) | ( x1063 & ~n42461 ) ;
  assign n42463 = n42307 ^ x1045 ^ 1'b0 ;
  assign n42464 = ( x379 & x1045 ) | ( x379 & ~n42463 ) | ( x1045 & ~n42463 ) ;
  assign n42465 = n42307 ^ x1084 ^ 1'b0 ;
  assign n42466 = ( x380 & x1084 ) | ( x380 & ~n42465 ) | ( x1084 & ~n42465 ) ;
  assign n42467 = n42307 ^ x1081 ^ 1'b0 ;
  assign n42468 = ( x381 & x1081 ) | ( x381 & ~n42467 ) | ( x1081 & ~n42467 ) ;
  assign n42469 = n42307 ^ x1076 ^ 1'b0 ;
  assign n42470 = ( x382 & x1076 ) | ( x382 & ~n42469 ) | ( x1076 & ~n42469 ) ;
  assign n42471 = n42307 ^ x1071 ^ 1'b0 ;
  assign n42472 = ( x383 & x1071 ) | ( x383 & ~n42471 ) | ( x1071 & ~n42471 ) ;
  assign n42473 = n42307 ^ x1068 ^ 1'b0 ;
  assign n42474 = ( x384 & x1068 ) | ( x384 & ~n42473 ) | ( x1068 & ~n42473 ) ;
  assign n42475 = n42307 ^ x1042 ^ 1'b0 ;
  assign n42476 = ( x385 & x1042 ) | ( x385 & ~n42475 ) | ( x1042 & ~n42475 ) ;
  assign n42477 = n42307 ^ x1059 ^ 1'b0 ;
  assign n42478 = ( x386 & x1059 ) | ( x386 & ~n42477 ) | ( x1059 & ~n42477 ) ;
  assign n42479 = n42307 ^ x1053 ^ 1'b0 ;
  assign n42480 = ( x387 & x1053 ) | ( x387 & ~n42479 ) | ( x1053 & ~n42479 ) ;
  assign n42481 = n42307 ^ x1037 ^ 1'b0 ;
  assign n42482 = ( x388 & x1037 ) | ( x388 & ~n42481 ) | ( x1037 & ~n42481 ) ;
  assign n42483 = n42307 ^ x1036 ^ 1'b0 ;
  assign n42484 = ( x389 & x1036 ) | ( x389 & ~n42483 ) | ( x1036 & ~n42483 ) ;
  assign n42485 = n42310 ^ x1049 ^ 1'b0 ;
  assign n42486 = ( x390 & x1049 ) | ( x390 & ~n42485 ) | ( x1049 & ~n42485 ) ;
  assign n42487 = n42310 ^ x1062 ^ 1'b0 ;
  assign n42488 = ( x391 & x1062 ) | ( x391 & ~n42487 ) | ( x1062 & ~n42487 ) ;
  assign n42489 = n42310 ^ x1039 ^ 1'b0 ;
  assign n42490 = ( x392 & x1039 ) | ( x392 & ~n42489 ) | ( x1039 & ~n42489 ) ;
  assign n42491 = n42310 ^ x1067 ^ 1'b0 ;
  assign n42492 = ( x393 & x1067 ) | ( x393 & ~n42491 ) | ( x1067 & ~n42491 ) ;
  assign n42493 = n42310 ^ x1080 ^ 1'b0 ;
  assign n42494 = ( x394 & x1080 ) | ( x394 & ~n42493 ) | ( x1080 & ~n42493 ) ;
  assign n42495 = n42310 ^ x1055 ^ 1'b0 ;
  assign n42496 = ( x395 & x1055 ) | ( x395 & ~n42495 ) | ( x1055 & ~n42495 ) ;
  assign n42497 = n42310 ^ x1051 ^ 1'b0 ;
  assign n42498 = ( x396 & x1051 ) | ( x396 & ~n42497 ) | ( x1051 & ~n42497 ) ;
  assign n42499 = n42310 ^ x1048 ^ 1'b0 ;
  assign n42500 = ( x397 & x1048 ) | ( x397 & ~n42499 ) | ( x1048 & ~n42499 ) ;
  assign n42501 = n42310 ^ x1087 ^ 1'b0 ;
  assign n42502 = ( x398 & x1087 ) | ( x398 & ~n42501 ) | ( x1087 & ~n42501 ) ;
  assign n42503 = n42310 ^ x1047 ^ 1'b0 ;
  assign n42504 = ( x399 & x1047 ) | ( x399 & ~n42503 ) | ( x1047 & ~n42503 ) ;
  assign n42505 = n42310 ^ x1035 ^ 1'b0 ;
  assign n42506 = ( x400 & x1035 ) | ( x400 & ~n42505 ) | ( x1035 & ~n42505 ) ;
  assign n42507 = n42310 ^ x1079 ^ 1'b0 ;
  assign n42508 = ( x401 & x1079 ) | ( x401 & ~n42507 ) | ( x1079 & ~n42507 ) ;
  assign n42509 = n42310 ^ x1078 ^ 1'b0 ;
  assign n42510 = ( x402 & x1078 ) | ( x402 & ~n42509 ) | ( x1078 & ~n42509 ) ;
  assign n42511 = n42310 ^ x1045 ^ 1'b0 ;
  assign n42512 = ( x403 & x1045 ) | ( x403 & ~n42511 ) | ( x1045 & ~n42511 ) ;
  assign n42513 = n42310 ^ x1084 ^ 1'b0 ;
  assign n42514 = ( x404 & x1084 ) | ( x404 & ~n42513 ) | ( x1084 & ~n42513 ) ;
  assign n42515 = n42310 ^ x1081 ^ 1'b0 ;
  assign n42516 = ( x405 & x1081 ) | ( x405 & ~n42515 ) | ( x1081 & ~n42515 ) ;
  assign n42517 = n42310 ^ x1076 ^ 1'b0 ;
  assign n42518 = ( x406 & x1076 ) | ( x406 & ~n42517 ) | ( x1076 & ~n42517 ) ;
  assign n42519 = n42310 ^ x1071 ^ 1'b0 ;
  assign n42520 = ( x407 & x1071 ) | ( x407 & ~n42519 ) | ( x1071 & ~n42519 ) ;
  assign n42521 = n42310 ^ x1068 ^ 1'b0 ;
  assign n42522 = ( x408 & x1068 ) | ( x408 & ~n42521 ) | ( x1068 & ~n42521 ) ;
  assign n42523 = n42310 ^ x1042 ^ 1'b0 ;
  assign n42524 = ( x409 & x1042 ) | ( x409 & ~n42523 ) | ( x1042 & ~n42523 ) ;
  assign n42525 = n42310 ^ x1059 ^ 1'b0 ;
  assign n42526 = ( x410 & x1059 ) | ( x410 & ~n42525 ) | ( x1059 & ~n42525 ) ;
  assign n42527 = n42310 ^ x1053 ^ 1'b0 ;
  assign n42528 = ( x411 & x1053 ) | ( x411 & ~n42527 ) | ( x1053 & ~n42527 ) ;
  assign n42529 = n42310 ^ x1037 ^ 1'b0 ;
  assign n42530 = ( x412 & x1037 ) | ( x412 & ~n42529 ) | ( x1037 & ~n42529 ) ;
  assign n42531 = n42310 ^ x1036 ^ 1'b0 ;
  assign n42532 = ( x413 & x1036 ) | ( x413 & ~n42531 ) | ( x1036 & ~n42531 ) ;
  assign n42533 = ~n7318 & n42378 ;
  assign n42534 = n42533 ^ x1049 ^ 1'b0 ;
  assign n42535 = ( x414 & x1049 ) | ( x414 & ~n42534 ) | ( x1049 & ~n42534 ) ;
  assign n42536 = n42533 ^ x1062 ^ 1'b0 ;
  assign n42537 = ( x415 & x1062 ) | ( x415 & ~n42536 ) | ( x1062 & ~n42536 ) ;
  assign n42538 = n42533 ^ x1069 ^ 1'b0 ;
  assign n42539 = ( x416 & x1069 ) | ( x416 & ~n42538 ) | ( x1069 & ~n42538 ) ;
  assign n42540 = n42533 ^ x1039 ^ 1'b0 ;
  assign n42541 = ( x417 & x1039 ) | ( x417 & ~n42540 ) | ( x1039 & ~n42540 ) ;
  assign n42542 = n42533 ^ x1067 ^ 1'b0 ;
  assign n42543 = ( x418 & x1067 ) | ( x418 & ~n42542 ) | ( x1067 & ~n42542 ) ;
  assign n42544 = n42533 ^ x1080 ^ 1'b0 ;
  assign n42545 = ( x419 & x1080 ) | ( x419 & ~n42544 ) | ( x1080 & ~n42544 ) ;
  assign n42546 = n42533 ^ x1055 ^ 1'b0 ;
  assign n42547 = ( x420 & x1055 ) | ( x420 & ~n42546 ) | ( x1055 & ~n42546 ) ;
  assign n42548 = n42533 ^ x1051 ^ 1'b0 ;
  assign n42549 = ( x421 & x1051 ) | ( x421 & ~n42548 ) | ( x1051 & ~n42548 ) ;
  assign n42550 = n42533 ^ x1048 ^ 1'b0 ;
  assign n42551 = ( x422 & x1048 ) | ( x422 & ~n42550 ) | ( x1048 & ~n42550 ) ;
  assign n42552 = n42533 ^ x1087 ^ 1'b0 ;
  assign n42553 = ( x423 & x1087 ) | ( x423 & ~n42552 ) | ( x1087 & ~n42552 ) ;
  assign n42554 = n42533 ^ x1047 ^ 1'b0 ;
  assign n42555 = ( x424 & x1047 ) | ( x424 & ~n42554 ) | ( x1047 & ~n42554 ) ;
  assign n42556 = n42533 ^ x1035 ^ 1'b0 ;
  assign n42557 = ( x425 & x1035 ) | ( x425 & ~n42556 ) | ( x1035 & ~n42556 ) ;
  assign n42558 = n42533 ^ x1079 ^ 1'b0 ;
  assign n42559 = ( x426 & x1079 ) | ( x426 & ~n42558 ) | ( x1079 & ~n42558 ) ;
  assign n42560 = n42533 ^ x1078 ^ 1'b0 ;
  assign n42561 = ( x427 & x1078 ) | ( x427 & ~n42560 ) | ( x1078 & ~n42560 ) ;
  assign n42562 = n42533 ^ x1045 ^ 1'b0 ;
  assign n42563 = ( x428 & x1045 ) | ( x428 & ~n42562 ) | ( x1045 & ~n42562 ) ;
  assign n42564 = n42533 ^ x1084 ^ 1'b0 ;
  assign n42565 = ( x429 & x1084 ) | ( x429 & ~n42564 ) | ( x1084 & ~n42564 ) ;
  assign n42566 = n42533 ^ x1076 ^ 1'b0 ;
  assign n42567 = ( x430 & x1076 ) | ( x430 & ~n42566 ) | ( x1076 & ~n42566 ) ;
  assign n42568 = n42533 ^ x1071 ^ 1'b0 ;
  assign n42569 = ( x431 & x1071 ) | ( x431 & ~n42568 ) | ( x1071 & ~n42568 ) ;
  assign n42570 = n42533 ^ x1068 ^ 1'b0 ;
  assign n42571 = ( x432 & x1068 ) | ( x432 & ~n42570 ) | ( x1068 & ~n42570 ) ;
  assign n42572 = n42533 ^ x1042 ^ 1'b0 ;
  assign n42573 = ( x433 & x1042 ) | ( x433 & ~n42572 ) | ( x1042 & ~n42572 ) ;
  assign n42574 = n42533 ^ x1059 ^ 1'b0 ;
  assign n42575 = ( x434 & x1059 ) | ( x434 & ~n42574 ) | ( x1059 & ~n42574 ) ;
  assign n42576 = n42533 ^ x1053 ^ 1'b0 ;
  assign n42577 = ( x435 & x1053 ) | ( x435 & ~n42576 ) | ( x1053 & ~n42576 ) ;
  assign n42578 = n42533 ^ x1037 ^ 1'b0 ;
  assign n42579 = ( x436 & x1037 ) | ( x436 & ~n42578 ) | ( x1037 & ~n42578 ) ;
  assign n42580 = n42533 ^ x1070 ^ 1'b0 ;
  assign n42581 = ( x437 & x1070 ) | ( x437 & ~n42580 ) | ( x1070 & ~n42580 ) ;
  assign n42582 = n42533 ^ x1036 ^ 1'b0 ;
  assign n42583 = ( x438 & x1036 ) | ( x438 & ~n42582 ) | ( x1036 & ~n42582 ) ;
  assign n42584 = n42307 ^ x1057 ^ 1'b0 ;
  assign n42585 = ( x439 & x1057 ) | ( x439 & ~n42584 ) | ( x1057 & ~n42584 ) ;
  assign n42586 = n42307 ^ x1043 ^ 1'b0 ;
  assign n42587 = ( x440 & x1043 ) | ( x440 & ~n42586 ) | ( x1043 & ~n42586 ) ;
  assign n42588 = n42302 ^ x1044 ^ 1'b0 ;
  assign n42589 = ( x441 & x1044 ) | ( x441 & ~n42588 ) | ( x1044 & ~n42588 ) ;
  assign n42590 = n42307 ^ x1058 ^ 1'b0 ;
  assign n42591 = ( x442 & x1058 ) | ( x442 & ~n42590 ) | ( x1058 & ~n42590 ) ;
  assign n42592 = n42533 ^ x1044 ^ 1'b0 ;
  assign n42593 = ( x443 & x1044 ) | ( x443 & ~n42592 ) | ( x1044 & ~n42592 ) ;
  assign n42594 = n42533 ^ x1072 ^ 1'b0 ;
  assign n42595 = ( x444 & x1072 ) | ( x444 & ~n42594 ) | ( x1072 & ~n42594 ) ;
  assign n42596 = n42533 ^ x1081 ^ 1'b0 ;
  assign n42597 = ( x445 & x1081 ) | ( x445 & ~n42596 ) | ( x1081 & ~n42596 ) ;
  assign n42598 = n42533 ^ x1086 ^ 1'b0 ;
  assign n42599 = ( x446 & x1086 ) | ( x446 & ~n42598 ) | ( x1086 & ~n42598 ) ;
  assign n42600 = n42307 ^ x1040 ^ 1'b0 ;
  assign n42601 = ( x447 & x1040 ) | ( x447 & ~n42600 ) | ( x1040 & ~n42600 ) ;
  assign n42602 = n42533 ^ x1074 ^ 1'b0 ;
  assign n42603 = ( x448 & x1074 ) | ( x448 & ~n42602 ) | ( x1074 & ~n42602 ) ;
  assign n42604 = n42533 ^ x1057 ^ 1'b0 ;
  assign n42605 = ( x449 & x1057 ) | ( x449 & ~n42604 ) | ( x1057 & ~n42604 ) ;
  assign n42606 = n42302 ^ x1036 ^ 1'b0 ;
  assign n42607 = ( x450 & x1036 ) | ( x450 & ~n42606 ) | ( x1036 & ~n42606 ) ;
  assign n42608 = n42533 ^ x1063 ^ 1'b0 ;
  assign n42609 = ( x451 & x1063 ) | ( x451 & ~n42608 ) | ( x1063 & ~n42608 ) ;
  assign n42610 = n42302 ^ x1053 ^ 1'b0 ;
  assign n42611 = ( x452 & x1053 ) | ( x452 & ~n42610 ) | ( x1053 & ~n42610 ) ;
  assign n42612 = n42533 ^ x1040 ^ 1'b0 ;
  assign n42613 = ( x453 & x1040 ) | ( x453 & ~n42612 ) | ( x1040 & ~n42612 ) ;
  assign n42614 = n42533 ^ x1043 ^ 1'b0 ;
  assign n42615 = ( x454 & x1043 ) | ( x454 & ~n42614 ) | ( x1043 & ~n42614 ) ;
  assign n42616 = n42302 ^ x1037 ^ 1'b0 ;
  assign n42617 = ( x455 & x1037 ) | ( x455 & ~n42616 ) | ( x1037 & ~n42616 ) ;
  assign n42618 = n42310 ^ x1044 ^ 1'b0 ;
  assign n42619 = ( x456 & x1044 ) | ( x456 & ~n42618 ) | ( x1044 & ~n42618 ) ;
  assign n42620 = x594 & x600 ;
  assign n42621 = x990 & n42620 ;
  assign n42622 = x600 & ~x810 ;
  assign n42623 = x804 & ~n42622 ;
  assign n42624 = ~x815 & n42623 ;
  assign n42625 = n42621 & n42624 ;
  assign n42630 = ~x599 & x810 ;
  assign n42631 = x596 & ~n42630 ;
  assign n42632 = x804 & ~n42631 ;
  assign n42633 = ( x595 & x815 ) | ( x595 & n42632 ) | ( x815 & n42632 ) ;
  assign n42634 = ~n42632 & n42633 ;
  assign n42627 = x804 | x810 ;
  assign n42635 = ( x595 & n42627 ) | ( x595 & ~n42634 ) | ( n42627 & ~n42634 ) ;
  assign n42636 = ~n42634 & n42635 ;
  assign n42637 = x597 & n42620 ;
  assign n42638 = ( x601 & n42636 ) | ( x601 & n42637 ) | ( n42636 & n42637 ) ;
  assign n42639 = ~n42636 & n42638 ;
  assign n42626 = x815 | n42623 ;
  assign n42628 = ~x601 & n42627 ;
  assign n42629 = n42626 | n42628 ;
  assign n42640 = n42639 ^ n42629 ^ 1'b0 ;
  assign n42641 = ( x605 & ~n42629 ) | ( x605 & n42639 ) | ( ~n42629 & n42639 ) ;
  assign n42642 = ( x605 & ~n42640 ) | ( x605 & n42641 ) | ( ~n42640 & n42641 ) ;
  assign n42643 = ( x821 & n42625 ) | ( x821 & n42642 ) | ( n42625 & n42642 ) ;
  assign n42644 = n42642 ^ n42625 ^ 1'b0 ;
  assign n42645 = ( x821 & n42643 ) | ( x821 & n42644 ) | ( n42643 & n42644 ) ;
  assign n42646 = n42302 ^ x1072 ^ 1'b0 ;
  assign n42647 = ( x458 & x1072 ) | ( x458 & ~n42646 ) | ( x1072 & ~n42646 ) ;
  assign n42648 = n42533 ^ x1058 ^ 1'b0 ;
  assign n42649 = ( x459 & x1058 ) | ( x459 & ~n42648 ) | ( x1058 & ~n42648 ) ;
  assign n42650 = n42302 ^ x1086 ^ 1'b0 ;
  assign n42651 = ( x460 & x1086 ) | ( x460 & ~n42650 ) | ( x1086 & ~n42650 ) ;
  assign n42652 = n42302 ^ x1057 ^ 1'b0 ;
  assign n42653 = ( x461 & x1057 ) | ( x461 & ~n42652 ) | ( x1057 & ~n42652 ) ;
  assign n42654 = n42302 ^ x1074 ^ 1'b0 ;
  assign n42655 = ( x462 & x1074 ) | ( x462 & ~n42654 ) | ( x1074 & ~n42654 ) ;
  assign n42656 = n42310 ^ x1070 ^ 1'b0 ;
  assign n42657 = ( x463 & x1070 ) | ( x463 & ~n42656 ) | ( x1070 & ~n42656 ) ;
  assign n42658 = n42533 ^ x1065 ^ 1'b0 ;
  assign n42659 = ( x464 & x1065 ) | ( x464 & ~n42658 ) | ( x1065 & ~n42658 ) ;
  assign n42660 = x926 & n42217 ;
  assign n42661 = ~x243 & n42215 ;
  assign n42662 = n7318 & ~n42661 ;
  assign n42663 = x1157 & n4865 ;
  assign n42664 = ( n42660 & n42662 ) | ( n42660 & ~n42663 ) | ( n42662 & ~n42663 ) ;
  assign n42665 = ~n42660 & n42664 ;
  assign n42666 = n2291 & ~n10054 ;
  assign n42667 = ~x243 & x1157 ;
  assign n42668 = x926 & n42667 ;
  assign n42669 = ~n42666 & n42668 ;
  assign n42670 = n10031 | n10034 ;
  assign n42671 = ~x243 & n42670 ;
  assign n42672 = x299 | n2170 ;
  assign n42673 = ~n10053 & n42672 ;
  assign n42674 = n42667 | n42673 ;
  assign n42675 = n42671 | n42674 ;
  assign n42676 = n4870 & ~n4872 ;
  assign n42677 = x926 & ~n42676 ;
  assign n42678 = x1157 & n42676 ;
  assign n42679 = ( n42671 & ~n42677 ) | ( n42671 & n42678 ) | ( ~n42677 & n42678 ) ;
  assign n42680 = n42677 | n42679 ;
  assign n42681 = ( n42669 & n42675 ) | ( n42669 & n42680 ) | ( n42675 & n42680 ) ;
  assign n42682 = ~n42669 & n42681 ;
  assign n42683 = ( n7318 & ~n42665 ) | ( n7318 & n42682 ) | ( ~n42665 & n42682 ) ;
  assign n42684 = ~n42665 & n42683 ;
  assign n42685 = n15098 ^ n2264 ^ 1'b0 ;
  assign n42686 = ( n1360 & n2264 ) | ( n1360 & ~n42685 ) | ( n2264 & ~n42685 ) ;
  assign n42687 = x943 & x1151 ;
  assign n42688 = ~n42686 & n42687 ;
  assign n42689 = n7318 ^ n2022 ^ 1'b0 ;
  assign n42690 = ( n2022 & n42673 ) | ( n2022 & ~n42689 ) | ( n42673 & ~n42689 ) ;
  assign n42691 = x275 | n42690 ;
  assign n42692 = n42215 ^ n7318 ^ 1'b0 ;
  assign n42693 = ( n42215 & n42670 ) | ( n42215 & ~n42692 ) | ( n42670 & ~n42692 ) ;
  assign n42694 = x943 | n42693 ;
  assign n42695 = n42233 | n42694 ;
  assign n42696 = ( n42688 & n42691 ) | ( n42688 & n42695 ) | ( n42691 & n42695 ) ;
  assign n42697 = ~n42688 & n42696 ;
  assign n42698 = x943 & ~n42263 ;
  assign n42699 = n42694 & ~n42698 ;
  assign n42700 = n42699 ^ x1151 ^ 1'b0 ;
  assign n42701 = ( x1151 & n42699 ) | ( x1151 & ~n42700 ) | ( n42699 & ~n42700 ) ;
  assign n42702 = ( n42697 & n42700 ) | ( n42697 & n42701 ) | ( n42700 & n42701 ) ;
  assign n42703 = n7472 | n8757 ;
  assign n42704 = n15261 | n42703 ;
  assign n42705 = x102 | n11879 ;
  assign n42706 = ( n15258 & ~n42704 ) | ( n15258 & n42705 ) | ( ~n42704 & n42705 ) ;
  assign n42707 = ~n15258 & n42706 ;
  assign n42708 = x40 & ~x287 ;
  assign n42709 = n39972 & n42708 ;
  assign n42710 = n42709 ^ n42707 ^ 1'b0 ;
  assign n42711 = n42707 ^ n5022 ^ 1'b0 ;
  assign n42712 = ( n42707 & n42710 ) | ( n42707 & ~n42711 ) | ( n42710 & ~n42711 ) ;
  assign n42713 = ~n6490 & n42712 ;
  assign n42714 = n6490 & n42710 ;
  assign n42715 = ( x1091 & n42713 ) | ( x1091 & ~n42714 ) | ( n42713 & ~n42714 ) ;
  assign n42716 = ~n42713 & n42715 ;
  assign n42717 = n42707 ^ n6425 ^ 1'b0 ;
  assign n42718 = ( n42707 & n42710 ) | ( n42707 & ~n42717 ) | ( n42710 & ~n42717 ) ;
  assign n42719 = x1093 & n42718 ;
  assign n42720 = ~x1093 & n42712 ;
  assign n42721 = x1091 | n42720 ;
  assign n42722 = ( ~n42716 & n42719 ) | ( ~n42716 & n42721 ) | ( n42719 & n42721 ) ;
  assign n42723 = ~n42716 & n42722 ;
  assign n42724 = ( n1207 & n42297 ) | ( n1207 & ~n42723 ) | ( n42297 & ~n42723 ) ;
  assign n42725 = n42723 | n42724 ;
  assign n42726 = ~n35897 & n42709 ;
  assign n42727 = n42726 ^ n42725 ^ 1'b0 ;
  assign n42728 = ( ~n8760 & n42726 ) | ( ~n8760 & n42727 ) | ( n42726 & n42727 ) ;
  assign n42729 = ( n42725 & ~n42727 ) | ( n42725 & n42728 ) | ( ~n42727 & n42728 ) ;
  assign n42730 = x38 & ~x39 ;
  assign n42731 = ( n7455 & ~n8793 ) | ( n7455 & n42730 ) | ( ~n8793 & n42730 ) ;
  assign n42732 = ~n7455 & n42731 ;
  assign n42733 = ~n9977 & n42732 ;
  assign n42734 = ( x468 & n9977 ) | ( x468 & ~n42733 ) | ( n9977 & ~n42733 ) ;
  assign n42735 = x942 & n42217 ;
  assign n42736 = ~x263 & n42215 ;
  assign n42737 = n7318 & ~n42736 ;
  assign n42738 = x1156 & n4865 ;
  assign n42739 = ( n42735 & n42737 ) | ( n42735 & ~n42738 ) | ( n42737 & ~n42738 ) ;
  assign n42740 = ~n42735 & n42739 ;
  assign n42741 = ~x263 & x1156 ;
  assign n42742 = x942 & n42741 ;
  assign n42743 = ~n42666 & n42742 ;
  assign n42744 = ~x263 & n42670 ;
  assign n42745 = n42673 | n42741 ;
  assign n42746 = n42744 | n42745 ;
  assign n42747 = x942 & ~n42676 ;
  assign n42748 = x1156 & n42676 ;
  assign n42749 = ( n42744 & ~n42747 ) | ( n42744 & n42748 ) | ( ~n42747 & n42748 ) ;
  assign n42750 = n42747 | n42749 ;
  assign n42751 = ( n42743 & n42746 ) | ( n42743 & n42750 ) | ( n42746 & n42750 ) ;
  assign n42752 = ~n42743 & n42751 ;
  assign n42753 = ( n7318 & ~n42740 ) | ( n7318 & n42752 ) | ( ~n42740 & n42752 ) ;
  assign n42754 = ~n42740 & n42753 ;
  assign n42755 = x925 & n42217 ;
  assign n42756 = x267 & n42215 ;
  assign n42757 = n7318 & ~n42756 ;
  assign n42758 = x1155 & n4865 ;
  assign n42759 = ( n42755 & n42757 ) | ( n42755 & ~n42758 ) | ( n42757 & ~n42758 ) ;
  assign n42760 = ~n42755 & n42759 ;
  assign n42761 = x267 & x1155 ;
  assign n42762 = x925 & n42761 ;
  assign n42763 = ~n42666 & n42762 ;
  assign n42764 = x267 & n42670 ;
  assign n42765 = n42673 | n42761 ;
  assign n42766 = n42764 | n42765 ;
  assign n42767 = x925 & ~n42676 ;
  assign n42768 = x1155 & n42676 ;
  assign n42769 = ( n42764 & ~n42767 ) | ( n42764 & n42768 ) | ( ~n42767 & n42768 ) ;
  assign n42770 = n42767 | n42769 ;
  assign n42771 = ( n42763 & n42766 ) | ( n42763 & n42770 ) | ( n42766 & n42770 ) ;
  assign n42772 = ~n42763 & n42771 ;
  assign n42773 = ( n7318 & ~n42760 ) | ( n7318 & n42772 ) | ( ~n42760 & n42772 ) ;
  assign n42774 = ~n42760 & n42773 ;
  assign n42775 = x941 & n42217 ;
  assign n42776 = x253 & n42215 ;
  assign n42777 = n7318 & ~n42776 ;
  assign n42778 = x1153 & n4865 ;
  assign n42779 = ( n42775 & n42777 ) | ( n42775 & ~n42778 ) | ( n42777 & ~n42778 ) ;
  assign n42780 = ~n42775 & n42779 ;
  assign n42781 = x253 & x1153 ;
  assign n42782 = x941 & n42781 ;
  assign n42783 = ~n42666 & n42782 ;
  assign n42784 = x253 & n42670 ;
  assign n42785 = n42673 | n42781 ;
  assign n42786 = n42784 | n42785 ;
  assign n42787 = x941 & ~n42676 ;
  assign n42788 = x1153 & n42676 ;
  assign n42789 = ( n42784 & ~n42787 ) | ( n42784 & n42788 ) | ( ~n42787 & n42788 ) ;
  assign n42790 = n42787 | n42789 ;
  assign n42791 = ( n42783 & n42786 ) | ( n42783 & n42790 ) | ( n42786 & n42790 ) ;
  assign n42792 = ~n42783 & n42791 ;
  assign n42793 = ( n7318 & ~n42780 ) | ( n7318 & n42792 ) | ( ~n42780 & n42792 ) ;
  assign n42794 = ~n42780 & n42793 ;
  assign n42795 = x923 & n42217 ;
  assign n42796 = x254 & n42215 ;
  assign n42797 = n7318 & ~n42796 ;
  assign n42798 = x1154 & n4865 ;
  assign n42799 = ( n42795 & n42797 ) | ( n42795 & ~n42798 ) | ( n42797 & ~n42798 ) ;
  assign n42800 = ~n42795 & n42799 ;
  assign n42801 = x254 & x1154 ;
  assign n42802 = x923 & n42801 ;
  assign n42803 = ~n42666 & n42802 ;
  assign n42804 = x254 & n42670 ;
  assign n42805 = n42673 | n42801 ;
  assign n42806 = n42804 | n42805 ;
  assign n42807 = x923 & ~n42676 ;
  assign n42808 = x1154 & n42676 ;
  assign n42809 = ( n42804 & ~n42807 ) | ( n42804 & n42808 ) | ( ~n42807 & n42808 ) ;
  assign n42810 = n42807 | n42809 ;
  assign n42811 = ( n42803 & n42806 ) | ( n42803 & n42810 ) | ( n42806 & n42810 ) ;
  assign n42812 = ~n42803 & n42811 ;
  assign n42813 = ( n7318 & ~n42800 ) | ( n7318 & n42812 ) | ( ~n42800 & n42812 ) ;
  assign n42814 = ~n42800 & n42813 ;
  assign n42815 = x922 & x1152 ;
  assign n42816 = ~n42686 & n42815 ;
  assign n42817 = x922 | n42693 ;
  assign n42818 = n42233 | n42817 ;
  assign n42819 = x268 | n42690 ;
  assign n42820 = ( n42816 & n42818 ) | ( n42816 & n42819 ) | ( n42818 & n42819 ) ;
  assign n42821 = ~n42816 & n42820 ;
  assign n42822 = x922 & ~n42263 ;
  assign n42823 = n42817 & ~n42822 ;
  assign n42824 = n42823 ^ x1152 ^ 1'b0 ;
  assign n42825 = ( x1152 & n42823 ) | ( x1152 & ~n42824 ) | ( n42823 & ~n42824 ) ;
  assign n42826 = ( n42821 & n42824 ) | ( n42821 & n42825 ) | ( n42824 & n42825 ) ;
  assign n42827 = x931 & x1150 ;
  assign n42828 = ~n42686 & n42827 ;
  assign n42829 = x272 | n42690 ;
  assign n42830 = x931 | n42693 ;
  assign n42831 = n42233 | n42830 ;
  assign n42832 = ( n42828 & n42829 ) | ( n42828 & n42831 ) | ( n42829 & n42831 ) ;
  assign n42833 = ~n42828 & n42832 ;
  assign n42834 = x931 & ~n42263 ;
  assign n42835 = n42830 & ~n42834 ;
  assign n42836 = n42835 ^ x1150 ^ 1'b0 ;
  assign n42837 = ( x1150 & n42835 ) | ( x1150 & ~n42836 ) | ( n42835 & ~n42836 ) ;
  assign n42838 = ( n42833 & n42836 ) | ( n42833 & n42837 ) | ( n42836 & n42837 ) ;
  assign n42839 = x936 & x1149 ;
  assign n42840 = ~n42686 & n42839 ;
  assign n42841 = x936 | n42693 ;
  assign n42842 = n42233 | n42841 ;
  assign n42843 = x283 | n42690 ;
  assign n42844 = ( n42840 & n42842 ) | ( n42840 & n42843 ) | ( n42842 & n42843 ) ;
  assign n42845 = ~n42840 & n42844 ;
  assign n42846 = x936 & ~n42263 ;
  assign n42847 = n42841 & ~n42846 ;
  assign n42848 = n42847 ^ x1149 ^ 1'b0 ;
  assign n42849 = ( x1149 & n42847 ) | ( x1149 & ~n42848 ) | ( n42847 & ~n42848 ) ;
  assign n42850 = ( n42845 & n42848 ) | ( n42845 & n42849 ) | ( n42848 & n42849 ) ;
  assign n42851 = n2070 | n8757 ;
  assign n42852 = ~n8746 & n10077 ;
  assign n42853 = ~n8742 & n42852 ;
  assign n42854 = ( n10077 & n11536 ) | ( n10077 & ~n42853 ) | ( n11536 & ~n42853 ) ;
  assign n42855 = ~n42853 & n42854 ;
  assign n42856 = ( n11540 & n42851 ) | ( n11540 & ~n42855 ) | ( n42851 & ~n42855 ) ;
  assign n42857 = ~n42851 & n42856 ;
  assign n42858 = x71 & n10077 ;
  assign n42859 = ( ~n7318 & n42857 ) | ( ~n7318 & n42858 ) | ( n42857 & n42858 ) ;
  assign n42860 = ~n7318 & n42859 ;
  assign n42861 = n7318 & n10075 ;
  assign n42862 = n42860 ^ x71 ^ 1'b0 ;
  assign n42863 = ( ~x71 & n42861 ) | ( ~x71 & n42862 ) | ( n42861 & n42862 ) ;
  assign n42864 = ( x71 & n42860 ) | ( x71 & n42863 ) | ( n42860 & n42863 ) ;
  assign n42865 = x71 & ~n41450 ;
  assign n42866 = n32360 ^ x248 ^ 1'b0 ;
  assign n42867 = ( x248 & x481 ) | ( x248 & ~n42866 ) | ( x481 & ~n42866 ) ;
  assign n42868 = n32372 ^ x249 ^ 1'b0 ;
  assign n42869 = ( x249 & x482 ) | ( x249 & ~n42868 ) | ( x482 & ~n42868 ) ;
  assign n42870 = n32491 ^ x242 ^ 1'b0 ;
  assign n42871 = ( x242 & x483 ) | ( x242 & ~n42870 ) | ( x483 & ~n42870 ) ;
  assign n42872 = n32491 ^ x249 ^ 1'b0 ;
  assign n42873 = ( x249 & x484 ) | ( x249 & ~n42872 ) | ( x484 & ~n42872 ) ;
  assign n42874 = n33661 ^ x234 ^ 1'b0 ;
  assign n42875 = ( x234 & x485 ) | ( x234 & ~n42874 ) | ( x485 & ~n42874 ) ;
  assign n42876 = n33661 ^ x244 ^ 1'b0 ;
  assign n42877 = ( x244 & x486 ) | ( x244 & ~n42876 ) | ( x486 & ~n42876 ) ;
  assign n42878 = n32360 ^ x246 ^ 1'b0 ;
  assign n42879 = ( x246 & x487 ) | ( x246 & ~n42878 ) | ( x487 & ~n42878 ) ;
  assign n42880 = n32360 ^ x239 ^ 1'b0 ;
  assign n42881 = ( ~x239 & x488 ) | ( ~x239 & n42880 ) | ( x488 & n42880 ) ;
  assign n42882 = n33661 ^ x242 ^ 1'b0 ;
  assign n42883 = ( x242 & x489 ) | ( x242 & ~n42882 ) | ( x489 & ~n42882 ) ;
  assign n42884 = n32491 ^ x241 ^ 1'b0 ;
  assign n42885 = ( x241 & x490 ) | ( x241 & ~n42884 ) | ( x490 & ~n42884 ) ;
  assign n42886 = n32491 ^ x238 ^ 1'b0 ;
  assign n42887 = ( x238 & x491 ) | ( x238 & ~n42886 ) | ( x491 & ~n42886 ) ;
  assign n42888 = n32491 ^ x240 ^ 1'b0 ;
  assign n42889 = ( x240 & x492 ) | ( x240 & ~n42888 ) | ( x492 & ~n42888 ) ;
  assign n42890 = n32491 ^ x244 ^ 1'b0 ;
  assign n42891 = ( x244 & x493 ) | ( x244 & ~n42890 ) | ( x493 & ~n42890 ) ;
  assign n42892 = n32491 ^ x239 ^ 1'b0 ;
  assign n42893 = ( ~x239 & x494 ) | ( ~x239 & n42892 ) | ( x494 & n42892 ) ;
  assign n42894 = n32491 ^ x235 ^ 1'b0 ;
  assign n42895 = ( x235 & x495 ) | ( x235 & ~n42894 ) | ( x495 & ~n42894 ) ;
  assign n42896 = n32485 ^ x249 ^ 1'b0 ;
  assign n42897 = ( x249 & x496 ) | ( x249 & ~n42896 ) | ( x496 & ~n42896 ) ;
  assign n42898 = n32485 ^ x239 ^ 1'b0 ;
  assign n42899 = ( ~x239 & x497 ) | ( ~x239 & n42898 ) | ( x497 & n42898 ) ;
  assign n42900 = n32372 ^ x238 ^ 1'b0 ;
  assign n42901 = ( x238 & x498 ) | ( x238 & ~n42900 ) | ( x498 & ~n42900 ) ;
  assign n42902 = n32485 ^ x246 ^ 1'b0 ;
  assign n42903 = ( x246 & x499 ) | ( x246 & ~n42902 ) | ( x499 & ~n42902 ) ;
  assign n42904 = n32485 ^ x241 ^ 1'b0 ;
  assign n42905 = ( x241 & x500 ) | ( x241 & ~n42904 ) | ( x500 & ~n42904 ) ;
  assign n42906 = n32485 ^ x248 ^ 1'b0 ;
  assign n42907 = ( x248 & x501 ) | ( x248 & ~n42906 ) | ( x501 & ~n42906 ) ;
  assign n42908 = n32485 ^ x247 ^ 1'b0 ;
  assign n42909 = ( x247 & x502 ) | ( x247 & ~n42908 ) | ( x502 & ~n42908 ) ;
  assign n42910 = n32485 ^ x245 ^ 1'b0 ;
  assign n42911 = ( x245 & x503 ) | ( x245 & ~n42910 ) | ( x503 & ~n42910 ) ;
  assign n42912 = n32480 ^ x242 ^ 1'b0 ;
  assign n42913 = ( x242 & x504 ) | ( x242 & ~n42912 ) | ( x504 & ~n42912 ) ;
  assign n42914 = x234 & n32479 ;
  assign n42915 = ~x505 & n32363 ;
  assign n42916 = n42914 & n42915 ;
  assign n42917 = n15098 ^ n5292 ^ 1'b0 ;
  assign n42918 = ( n5201 & n5292 ) | ( n5201 & ~n42917 ) | ( n5292 & ~n42917 ) ;
  assign n42919 = ~x234 & n42918 ;
  assign n42920 = n32485 & n42919 ;
  assign n42921 = ~n42916 & n42920 ;
  assign n42922 = ( x505 & n42916 ) | ( x505 & ~n42921 ) | ( n42916 & ~n42921 ) ;
  assign n42923 = n32480 ^ x241 ^ 1'b0 ;
  assign n42924 = ( x241 & x506 ) | ( x241 & ~n42923 ) | ( x506 & ~n42923 ) ;
  assign n42925 = n32480 ^ x238 ^ 1'b0 ;
  assign n42926 = ( x238 & x507 ) | ( x238 & ~n42925 ) | ( x507 & ~n42925 ) ;
  assign n42927 = n32480 ^ x247 ^ 1'b0 ;
  assign n42928 = ( x247 & x508 ) | ( x247 & ~n42927 ) | ( x508 & ~n42927 ) ;
  assign n42929 = n32480 ^ x245 ^ 1'b0 ;
  assign n42930 = ( x245 & x509 ) | ( x245 & ~n42929 ) | ( x509 & ~n42929 ) ;
  assign n42931 = n32360 ^ x242 ^ 1'b0 ;
  assign n42932 = ( x242 & x510 ) | ( x242 & ~n42931 ) | ( x510 & ~n42931 ) ;
  assign n42933 = ~n5497 & n15098 ;
  assign n42934 = n5530 | n7318 ;
  assign n42935 = ~n42933 & n42934 ;
  assign n42936 = ~x234 & n42935 ;
  assign n42937 = n42936 ^ n32360 ^ 1'b0 ;
  assign n42938 = ( x511 & ~n42936 ) | ( x511 & n42937 ) | ( ~n42936 & n42937 ) ;
  assign n42939 = n32360 ^ x235 ^ 1'b0 ;
  assign n42940 = ( x235 & x512 ) | ( x235 & ~n42939 ) | ( x512 & ~n42939 ) ;
  assign n42941 = n32360 ^ x244 ^ 1'b0 ;
  assign n42942 = ( x244 & x513 ) | ( x244 & ~n42941 ) | ( x513 & ~n42941 ) ;
  assign n42943 = n32360 ^ x245 ^ 1'b0 ;
  assign n42944 = ( x245 & x514 ) | ( x245 & ~n42943 ) | ( x514 & ~n42943 ) ;
  assign n42945 = n32360 ^ x240 ^ 1'b0 ;
  assign n42946 = ( x240 & x515 ) | ( x240 & ~n42945 ) | ( x515 & ~n42945 ) ;
  assign n42947 = n32360 ^ x247 ^ 1'b0 ;
  assign n42948 = ( x247 & x516 ) | ( x247 & ~n42947 ) | ( x516 & ~n42947 ) ;
  assign n42949 = n32360 ^ x238 ^ 1'b0 ;
  assign n42950 = ( x238 & x517 ) | ( x238 & ~n42949 ) | ( x517 & ~n42949 ) ;
  assign n42951 = x234 & n32359 ;
  assign n42952 = ~x518 & n32363 ;
  assign n42953 = n42951 & n42952 ;
  assign n42954 = n32366 & n42936 ;
  assign n42955 = ~n42953 & n42954 ;
  assign n42956 = ( x518 & n42953 ) | ( x518 & ~n42955 ) | ( n42953 & ~n42955 ) ;
  assign n42957 = n32366 ^ x239 ^ 1'b0 ;
  assign n42958 = ( ~x239 & x519 ) | ( ~x239 & n42957 ) | ( x519 & n42957 ) ;
  assign n42959 = n32366 ^ x246 ^ 1'b0 ;
  assign n42960 = ( x246 & x520 ) | ( x246 & ~n42959 ) | ( x520 & ~n42959 ) ;
  assign n42961 = n32366 ^ x248 ^ 1'b0 ;
  assign n42962 = ( x248 & x521 ) | ( x248 & ~n42961 ) | ( x521 & ~n42961 ) ;
  assign n42963 = n32366 ^ x238 ^ 1'b0 ;
  assign n42964 = ( x238 & x522 ) | ( x238 & ~n42963 ) | ( x522 & ~n42963 ) ;
  assign n42965 = ~x523 & n32488 ;
  assign n42966 = n42951 & n42965 ;
  assign n42967 = n33689 & n42936 ;
  assign n42968 = ~n42966 & n42967 ;
  assign n42969 = ( x523 & n42966 ) | ( x523 & ~n42968 ) | ( n42966 & ~n42968 ) ;
  assign n42970 = n33689 ^ x239 ^ 1'b0 ;
  assign n42971 = ( ~x239 & x524 ) | ( ~x239 & n42970 ) | ( x524 & n42970 ) ;
  assign n42972 = n33689 ^ x245 ^ 1'b0 ;
  assign n42973 = ( x245 & x525 ) | ( x245 & ~n42972 ) | ( x525 & ~n42972 ) ;
  assign n42974 = n33689 ^ x246 ^ 1'b0 ;
  assign n42975 = ( x246 & x526 ) | ( x246 & ~n42974 ) | ( x526 & ~n42974 ) ;
  assign n42976 = n33689 ^ x247 ^ 1'b0 ;
  assign n42977 = ( x247 & x527 ) | ( x247 & ~n42976 ) | ( x527 & ~n42976 ) ;
  assign n42978 = n33689 ^ x249 ^ 1'b0 ;
  assign n42979 = ( x249 & x528 ) | ( x249 & ~n42978 ) | ( x528 & ~n42978 ) ;
  assign n42980 = n33689 ^ x238 ^ 1'b0 ;
  assign n42981 = ( x238 & x529 ) | ( x238 & ~n42980 ) | ( x529 & ~n42980 ) ;
  assign n42982 = n33689 ^ x240 ^ 1'b0 ;
  assign n42983 = ( x240 & x530 ) | ( x240 & ~n42982 ) | ( x530 & ~n42982 ) ;
  assign n42984 = n32372 ^ x235 ^ 1'b0 ;
  assign n42985 = ( x235 & x531 ) | ( x235 & ~n42984 ) | ( x531 & ~n42984 ) ;
  assign n42986 = n32372 ^ x247 ^ 1'b0 ;
  assign n42987 = ( x247 & x532 ) | ( x247 & ~n42986 ) | ( x532 & ~n42986 ) ;
  assign n42988 = n32480 ^ x235 ^ 1'b0 ;
  assign n42989 = ( x235 & x533 ) | ( x235 & ~n42988 ) | ( x533 & ~n42988 ) ;
  assign n42990 = n32480 ^ x239 ^ 1'b0 ;
  assign n42991 = ( ~x239 & x534 ) | ( ~x239 & n42990 ) | ( x534 & n42990 ) ;
  assign n42992 = n32480 ^ x240 ^ 1'b0 ;
  assign n42993 = ( x240 & x535 ) | ( x240 & ~n42992 ) | ( x535 & ~n42992 ) ;
  assign n42994 = n32480 ^ x246 ^ 1'b0 ;
  assign n42995 = ( x246 & x536 ) | ( x246 & ~n42994 ) | ( x536 & ~n42994 ) ;
  assign n42996 = n32480 ^ x248 ^ 1'b0 ;
  assign n42997 = ( x248 & x537 ) | ( x248 & ~n42996 ) | ( x537 & ~n42996 ) ;
  assign n42998 = n32480 ^ x249 ^ 1'b0 ;
  assign n42999 = ( x249 & x538 ) | ( x249 & ~n42998 ) | ( x538 & ~n42998 ) ;
  assign n43000 = n32485 ^ x242 ^ 1'b0 ;
  assign n43001 = ( x242 & x539 ) | ( x242 & ~n43000 ) | ( x539 & ~n43000 ) ;
  assign n43002 = n32485 ^ x235 ^ 1'b0 ;
  assign n43003 = ( x235 & x540 ) | ( x235 & ~n43002 ) | ( x540 & ~n43002 ) ;
  assign n43004 = n32485 ^ x244 ^ 1'b0 ;
  assign n43005 = ( x244 & x541 ) | ( x244 & ~n43004 ) | ( x541 & ~n43004 ) ;
  assign n43006 = n32485 ^ x240 ^ 1'b0 ;
  assign n43007 = ( x240 & x542 ) | ( x240 & ~n43006 ) | ( x542 & ~n43006 ) ;
  assign n43008 = n32485 ^ x238 ^ 1'b0 ;
  assign n43009 = ( x238 & x543 ) | ( x238 & ~n43008 ) | ( x543 & ~n43008 ) ;
  assign n43010 = ~x544 & n32488 ;
  assign n43011 = n42914 & n43010 ;
  assign n43012 = n32491 & n42919 ;
  assign n43013 = ~n43011 & n43012 ;
  assign n43014 = ( x544 & n43011 ) | ( x544 & ~n43013 ) | ( n43011 & ~n43013 ) ;
  assign n43015 = n32491 ^ x245 ^ 1'b0 ;
  assign n43016 = ( x245 & x545 ) | ( x245 & ~n43015 ) | ( x545 & ~n43015 ) ;
  assign n43017 = n32491 ^ x246 ^ 1'b0 ;
  assign n43018 = ( x246 & x546 ) | ( x246 & ~n43017 ) | ( x546 & ~n43017 ) ;
  assign n43019 = n32491 ^ x247 ^ 1'b0 ;
  assign n43020 = ( x247 & x547 ) | ( x247 & ~n43019 ) | ( x547 & ~n43019 ) ;
  assign n43021 = n32491 ^ x248 ^ 1'b0 ;
  assign n43022 = ( x248 & x548 ) | ( x248 & ~n43021 ) | ( x548 & ~n43021 ) ;
  assign n43023 = n33661 ^ x235 ^ 1'b0 ;
  assign n43024 = ( x235 & x549 ) | ( x235 & ~n43023 ) | ( x549 & ~n43023 ) ;
  assign n43025 = n33661 ^ x239 ^ 1'b0 ;
  assign n43026 = ( ~x239 & x550 ) | ( ~x239 & n43025 ) | ( x550 & n43025 ) ;
  assign n43027 = n33661 ^ x240 ^ 1'b0 ;
  assign n43028 = ( x240 & x551 ) | ( x240 & ~n43027 ) | ( x551 & ~n43027 ) ;
  assign n43029 = n33661 ^ x247 ^ 1'b0 ;
  assign n43030 = ( x247 & x552 ) | ( x247 & ~n43029 ) | ( x552 & ~n43029 ) ;
  assign n43031 = n33661 ^ x241 ^ 1'b0 ;
  assign n43032 = ( x241 & x553 ) | ( x241 & ~n43031 ) | ( x553 & ~n43031 ) ;
  assign n43033 = n33661 ^ x248 ^ 1'b0 ;
  assign n43034 = ( x248 & x554 ) | ( x248 & ~n43033 ) | ( x554 & ~n43033 ) ;
  assign n43035 = n33661 ^ x249 ^ 1'b0 ;
  assign n43036 = ( x249 & x555 ) | ( x249 & ~n43035 ) | ( x555 & ~n43035 ) ;
  assign n43037 = n32372 ^ x242 ^ 1'b0 ;
  assign n43038 = ( x242 & x556 ) | ( x242 & ~n43037 ) | ( x556 & ~n43037 ) ;
  assign n43039 = ~x557 & n32351 ;
  assign n43040 = n42914 & n43039 ;
  assign n43041 = n32480 & n42919 ;
  assign n43042 = ~n43040 & n43041 ;
  assign n43043 = ( x557 & n43040 ) | ( x557 & ~n43042 ) | ( n43040 & ~n43042 ) ;
  assign n43044 = n32480 ^ x244 ^ 1'b0 ;
  assign n43045 = ( x244 & x558 ) | ( x244 & ~n43044 ) | ( x558 & ~n43044 ) ;
  assign n43046 = n32360 ^ x241 ^ 1'b0 ;
  assign n43047 = ( x241 & x559 ) | ( x241 & ~n43046 ) | ( x559 & ~n43046 ) ;
  assign n43048 = n32372 ^ x240 ^ 1'b0 ;
  assign n43049 = ( x240 & x560 ) | ( x240 & ~n43048 ) | ( x560 & ~n43048 ) ;
  assign n43050 = n32366 ^ x247 ^ 1'b0 ;
  assign n43051 = ( x247 & x561 ) | ( x247 & ~n43050 ) | ( x561 & ~n43050 ) ;
  assign n43052 = n32372 ^ x241 ^ 1'b0 ;
  assign n43053 = ( x241 & x562 ) | ( x241 & ~n43052 ) | ( x562 & ~n43052 ) ;
  assign n43054 = n33661 ^ x246 ^ 1'b0 ;
  assign n43055 = ( x246 & x563 ) | ( x246 & ~n43054 ) | ( x563 & ~n43054 ) ;
  assign n43056 = n32372 ^ x246 ^ 1'b0 ;
  assign n43057 = ( x246 & x564 ) | ( x246 & ~n43056 ) | ( x564 & ~n43056 ) ;
  assign n43058 = n32372 ^ x248 ^ 1'b0 ;
  assign n43059 = ( x248 & x565 ) | ( x248 & ~n43058 ) | ( x565 & ~n43058 ) ;
  assign n43060 = n32372 ^ x244 ^ 1'b0 ;
  assign n43061 = ( x244 & x566 ) | ( x244 & ~n43060 ) | ( x566 & ~n43060 ) ;
  assign n43062 = ~x567 & x1092 ;
  assign n43063 = ~x1093 & n43062 ;
  assign n43064 = x1157 | n43063 ;
  assign n43065 = x680 & n16124 ;
  assign n43066 = n17083 | n43065 ;
  assign n43067 = ( ~n17083 & n43063 ) | ( ~n17083 & n43066 ) | ( n43063 & n43066 ) ;
  assign n43068 = ~n17088 & n43067 ;
  assign n43069 = ~n17093 & n43068 ;
  assign n43070 = ~x647 & n43069 ;
  assign n43071 = n43064 | n43070 ;
  assign n43072 = n16339 & n43063 ;
  assign n43073 = x603 & ~n15659 ;
  assign n43074 = n15547 & ~n18309 ;
  assign n43075 = ( n18315 & n43073 ) | ( n18315 & n43074 ) | ( n43073 & n43074 ) ;
  assign n43076 = ~n18315 & n43075 ;
  assign n43077 = x789 | n43063 ;
  assign n43078 = n43076 | n43077 ;
  assign n43079 = x619 & n43076 ;
  assign n43080 = n43063 | n43079 ;
  assign n43081 = x1159 & n43080 ;
  assign n43082 = ~x619 & n43076 ;
  assign n43083 = ( ~x1159 & n43063 ) | ( ~x1159 & n43082 ) | ( n43063 & n43082 ) ;
  assign n43084 = ~x1159 & n43083 ;
  assign n43085 = ( x789 & n43081 ) | ( x789 & ~n43084 ) | ( n43081 & ~n43084 ) ;
  assign n43086 = ~n43081 & n43085 ;
  assign n43087 = n43078 & ~n43086 ;
  assign n43088 = n43063 ^ n16518 ^ 1'b0 ;
  assign n43089 = ( n43063 & n43087 ) | ( n43063 & ~n43088 ) | ( n43087 & ~n43088 ) ;
  assign n43090 = ~n16339 & n43089 ;
  assign n43091 = n43072 | n43090 ;
  assign n43092 = ~x647 & n43091 ;
  assign n43093 = x628 & n43068 ;
  assign n43094 = n43063 | n43093 ;
  assign n43095 = ( x1156 & ~n17240 ) | ( x1156 & n43094 ) | ( ~n17240 & n43094 ) ;
  assign n43096 = ( x629 & n17240 ) | ( x629 & n43095 ) | ( n17240 & n43095 ) ;
  assign n43097 = n43096 ^ n16557 ^ 1'b0 ;
  assign n43098 = ( ~n16557 & n43089 ) | ( ~n16557 & n43097 ) | ( n43089 & n43097 ) ;
  assign n43099 = ( n16557 & n43096 ) | ( n16557 & n43098 ) | ( n43096 & n43098 ) ;
  assign n43100 = n16556 & n43089 ;
  assign n43101 = ~x628 & n43068 ;
  assign n43102 = ( ~x1156 & n43063 ) | ( ~x1156 & n43101 ) | ( n43063 & n43101 ) ;
  assign n43103 = ~x1156 & n43102 ;
  assign n43104 = ( x629 & n43100 ) | ( x629 & ~n43103 ) | ( n43100 & ~n43103 ) ;
  assign n43105 = ~n43100 & n43104 ;
  assign n43106 = x792 & ~n43105 ;
  assign n43107 = n43099 & n43106 ;
  assign n43108 = ~n17087 & n43067 ;
  assign n43109 = n16278 & n43086 ;
  assign n43110 = n43108 & ~n43109 ;
  assign n43111 = ( ~n16519 & n43087 ) | ( ~n16519 & n43110 ) | ( n43087 & n43110 ) ;
  assign n43112 = ~n16519 & n43111 ;
  assign n43113 = n43112 ^ x788 ^ 1'b0 ;
  assign n43114 = ~n16279 & n43108 ;
  assign n43115 = ~x641 & n43114 ;
  assign n43116 = n43063 | n43115 ;
  assign n43117 = n16454 & n43116 ;
  assign n43118 = x641 & n43114 ;
  assign n43119 = n43063 | n43118 ;
  assign n43120 = n43117 ^ n16453 ^ 1'b0 ;
  assign n43121 = ( ~n16453 & n43119 ) | ( ~n16453 & n43120 ) | ( n43119 & n43120 ) ;
  assign n43122 = ( n16453 & n43117 ) | ( n16453 & n43121 ) | ( n43117 & n43121 ) ;
  assign n43123 = n43122 ^ n32751 ^ 1'b0 ;
  assign n43124 = ( ~n32751 & n43087 ) | ( ~n32751 & n43123 ) | ( n43087 & n43123 ) ;
  assign n43125 = ( n32751 & n43122 ) | ( n32751 & n43124 ) | ( n43122 & n43124 ) ;
  assign n43126 = ( x788 & ~n43113 ) | ( x788 & n43125 ) | ( ~n43113 & n43125 ) ;
  assign n43127 = ( n43112 & n43113 ) | ( n43112 & n43126 ) | ( n43113 & n43126 ) ;
  assign n43128 = ( ~n18482 & n43107 ) | ( ~n18482 & n43127 ) | ( n43107 & n43127 ) ;
  assign n43129 = n43107 ^ n18482 ^ 1'b0 ;
  assign n43130 = ( n43107 & n43128 ) | ( n43107 & ~n43129 ) | ( n43128 & ~n43129 ) ;
  assign n43131 = x647 & n43130 ;
  assign n43132 = ( x1157 & n43092 ) | ( x1157 & ~n43131 ) | ( n43092 & ~n43131 ) ;
  assign n43133 = ~n43092 & n43132 ;
  assign n43134 = x630 & ~n43133 ;
  assign n43135 = n43071 & n43134 ;
  assign n43136 = ~x647 & n43130 ;
  assign n43137 = x647 & n43091 ;
  assign n43138 = ( x1157 & ~n43136 ) | ( x1157 & n43137 ) | ( ~n43136 & n43137 ) ;
  assign n43139 = n43136 | n43138 ;
  assign n43140 = x1157 & ~n43063 ;
  assign n43141 = x647 & n43069 ;
  assign n43142 = n43140 & ~n43141 ;
  assign n43143 = ( x630 & n43139 ) | ( x630 & ~n43142 ) | ( n43139 & ~n43142 ) ;
  assign n43144 = ~x630 & n43143 ;
  assign n43145 = ( x787 & n43135 ) | ( x787 & ~n43144 ) | ( n43135 & ~n43144 ) ;
  assign n43146 = ~n43135 & n43145 ;
  assign n43147 = ( x787 & n43130 ) | ( x787 & ~n43146 ) | ( n43130 & ~n43146 ) ;
  assign n43148 = ~n43146 & n43147 ;
  assign n43149 = x644 & ~n43148 ;
  assign n43150 = ~n17273 & n43069 ;
  assign n43151 = n43063 | n43150 ;
  assign n43152 = x644 | n43151 ;
  assign n43153 = ( x715 & n43149 ) | ( x715 & n43152 ) | ( n43149 & n43152 ) ;
  assign n43154 = ~n43149 & n43153 ;
  assign n43155 = ~n16376 & n43090 ;
  assign n43156 = x644 & n43155 ;
  assign n43157 = ( ~x715 & n43063 ) | ( ~x715 & n43156 ) | ( n43063 & n43156 ) ;
  assign n43158 = ~x715 & n43157 ;
  assign n43159 = ( x1160 & n43154 ) | ( x1160 & ~n43158 ) | ( n43154 & ~n43158 ) ;
  assign n43160 = ~n43154 & n43159 ;
  assign n43161 = ~x644 & n43148 ;
  assign n43162 = x644 & n43151 ;
  assign n43163 = ( x715 & ~n43161 ) | ( x715 & n43162 ) | ( ~n43161 & n43162 ) ;
  assign n43164 = n43161 | n43163 ;
  assign n43165 = ~x644 & n43155 ;
  assign n43166 = x715 & ~n43063 ;
  assign n43167 = ~n43165 & n43166 ;
  assign n43168 = ( x1160 & n43164 ) | ( x1160 & ~n43167 ) | ( n43164 & ~n43167 ) ;
  assign n43169 = n43168 ^ n43164 ^ 1'b0 ;
  assign n43170 = ( x1160 & n43168 ) | ( x1160 & ~n43169 ) | ( n43168 & ~n43169 ) ;
  assign n43171 = ( x790 & n43160 ) | ( x790 & n43170 ) | ( n43160 & n43170 ) ;
  assign n43172 = ~n43160 & n43171 ;
  assign n43173 = ( ~x790 & n43148 ) | ( ~x790 & n43172 ) | ( n43148 & n43172 ) ;
  assign n43174 = n43172 ^ x790 ^ 1'b0 ;
  assign n43175 = ( n43172 & n43173 ) | ( n43172 & ~n43174 ) | ( n43173 & ~n43174 ) ;
  assign n43176 = n43062 ^ x230 ^ 1'b0 ;
  assign n43177 = ( n43062 & n43175 ) | ( n43062 & n43176 ) | ( n43175 & n43176 ) ;
  assign n43178 = n32372 ^ x245 ^ 1'b0 ;
  assign n43179 = ( x245 & x568 ) | ( x245 & ~n43178 ) | ( x568 & ~n43178 ) ;
  assign n43180 = n32372 ^ x239 ^ 1'b0 ;
  assign n43181 = ( ~x239 & x569 ) | ( ~x239 & n43180 ) | ( x569 & n43180 ) ;
  assign n43182 = x570 | n32369 ;
  assign n43183 = n42951 & ~n43182 ;
  assign n43184 = n32372 & n42936 ;
  assign n43185 = ~n43183 & n43184 ;
  assign n43186 = ( x570 & n43183 ) | ( x570 & ~n43185 ) | ( n43183 & ~n43185 ) ;
  assign n43187 = n33689 ^ x241 ^ 1'b0 ;
  assign n43188 = ( x241 & x571 ) | ( x241 & ~n43187 ) | ( x571 & ~n43187 ) ;
  assign n43189 = n33689 ^ x244 ^ 1'b0 ;
  assign n43190 = ( x244 & x572 ) | ( x244 & ~n43189 ) | ( x572 & ~n43189 ) ;
  assign n43191 = n33689 ^ x242 ^ 1'b0 ;
  assign n43192 = ( x242 & x573 ) | ( x242 & ~n43191 ) | ( x573 & ~n43191 ) ;
  assign n43193 = n32366 ^ x241 ^ 1'b0 ;
  assign n43194 = ( x241 & x574 ) | ( x241 & ~n43193 ) | ( x574 & ~n43193 ) ;
  assign n43195 = n33689 ^ x235 ^ 1'b0 ;
  assign n43196 = ( x235 & x575 ) | ( x235 & ~n43195 ) | ( x575 & ~n43195 ) ;
  assign n43197 = n33689 ^ x248 ^ 1'b0 ;
  assign n43198 = ( x248 & x576 ) | ( x248 & ~n43197 ) | ( x576 & ~n43197 ) ;
  assign n43199 = n33661 ^ x238 ^ 1'b0 ;
  assign n43200 = ( x238 & x577 ) | ( x238 & ~n43199 ) | ( x577 & ~n43199 ) ;
  assign n43201 = n32366 ^ x249 ^ 1'b0 ;
  assign n43202 = ( x249 & x578 ) | ( x249 & ~n43201 ) | ( x578 & ~n43201 ) ;
  assign n43203 = n32360 ^ x249 ^ 1'b0 ;
  assign n43204 = ( x249 & x579 ) | ( x249 & ~n43203 ) | ( x579 & ~n43203 ) ;
  assign n43205 = n33661 ^ x245 ^ 1'b0 ;
  assign n43206 = ( x245 & x580 ) | ( x245 & ~n43205 ) | ( x580 & ~n43205 ) ;
  assign n43207 = n32366 ^ x235 ^ 1'b0 ;
  assign n43208 = ( x235 & x581 ) | ( x235 & ~n43207 ) | ( x581 & ~n43207 ) ;
  assign n43209 = n32366 ^ x240 ^ 1'b0 ;
  assign n43210 = ( x240 & x582 ) | ( x240 & ~n43209 ) | ( x582 & ~n43209 ) ;
  assign n43211 = n32366 ^ x245 ^ 1'b0 ;
  assign n43212 = ( x245 & x584 ) | ( x245 & ~n43211 ) | ( x584 & ~n43211 ) ;
  assign n43213 = n32366 ^ x244 ^ 1'b0 ;
  assign n43214 = ( x244 & x585 ) | ( x244 & ~n43213 ) | ( x585 & ~n43213 ) ;
  assign n43215 = n32366 ^ x242 ^ 1'b0 ;
  assign n43216 = ( x242 & x586 ) | ( x242 & ~n43215 ) | ( x586 & ~n43215 ) ;
  assign n43217 = x230 & n15524 ;
  assign n43218 = ( n18309 & ~n33075 ) | ( n18309 & n43217 ) | ( ~n33075 & n43217 ) ;
  assign n43219 = ~n18309 & n43218 ;
  assign n43220 = ( n18321 & ~n28311 ) | ( n18321 & n43219 ) | ( ~n28311 & n43219 ) ;
  assign n43221 = ~n18321 & n43220 ;
  assign n43222 = ( ~x230 & x587 ) | ( ~x230 & n43221 ) | ( x587 & n43221 ) ;
  assign n43223 = n43221 ^ x230 ^ 1'b0 ;
  assign n43224 = ( n43221 & n43222 ) | ( n43221 & ~n43223 ) | ( n43222 & ~n43223 ) ;
  assign n43225 = ~x123 & n10860 ;
  assign n43226 = ~x591 & n43225 ;
  assign n43227 = x588 | n43225 ;
  assign n43228 = ( n42335 & n43226 ) | ( n42335 & n43227 ) | ( n43226 & n43227 ) ;
  assign n43229 = ~n43226 & n43228 ;
  assign n43230 = ~x201 & n42935 ;
  assign n43231 = ~x204 & n42918 ;
  assign n43232 = ( x233 & n43230 ) | ( x233 & ~n43231 ) | ( n43230 & ~n43231 ) ;
  assign n43233 = ~n43230 & n43232 ;
  assign n43234 = ~x202 & n42935 ;
  assign n43235 = ~x205 & n42918 ;
  assign n43236 = x233 | n43235 ;
  assign n43237 = ( ~n43233 & n43234 ) | ( ~n43233 & n43236 ) | ( n43234 & n43236 ) ;
  assign n43238 = ~n43233 & n43237 ;
  assign n43239 = ~x220 & n42935 ;
  assign n43240 = ~x206 & n42918 ;
  assign n43241 = ( x233 & n43239 ) | ( x233 & ~n43240 ) | ( n43239 & ~n43240 ) ;
  assign n43242 = ~n43239 & n43241 ;
  assign n43243 = ~x203 & n42935 ;
  assign n43244 = ~x218 & n42918 ;
  assign n43245 = x233 | n43244 ;
  assign n43246 = ( ~n43242 & n43243 ) | ( ~n43242 & n43245 ) | ( n43243 & n43245 ) ;
  assign n43247 = ~n43242 & n43246 ;
  assign n43248 = n43238 ^ x237 ^ 1'b0 ;
  assign n43249 = ( n43238 & n43247 ) | ( n43238 & ~n43248 ) | ( n43247 & ~n43248 ) ;
  assign n43250 = x588 & n43225 ;
  assign n43251 = x590 & ~n43225 ;
  assign n43252 = ( n42335 & n43250 ) | ( n42335 & ~n43251 ) | ( n43250 & ~n43251 ) ;
  assign n43253 = ~n43250 & n43252 ;
  assign n43254 = ~x592 & n43225 ;
  assign n43255 = x591 | n43225 ;
  assign n43256 = ( n42335 & n43254 ) | ( n42335 & n43255 ) | ( n43254 & n43255 ) ;
  assign n43257 = ~n43254 & n43256 ;
  assign n43258 = ~x590 & n43225 ;
  assign n43259 = x592 | n43225 ;
  assign n43260 = ( n42335 & n43258 ) | ( n42335 & n43259 ) | ( n43258 & n43259 ) ;
  assign n43261 = ~n43258 & n43260 ;
  assign n43262 = x542 ^ x240 ^ 1'b0 ;
  assign n43263 = x496 ^ x249 ^ 1'b0 ;
  assign n43264 = x499 ^ x246 ^ 1'b0 ;
  assign n43265 = x501 ^ x248 ^ 1'b0 ;
  assign n43266 = ( ~n43263 & n43264 ) | ( ~n43263 & n43265 ) | ( n43264 & n43265 ) ;
  assign n43267 = n43263 | n43266 ;
  assign n43268 = x234 & n42918 ;
  assign n43269 = ~n43267 & n43268 ;
  assign n43270 = ( x505 & n43267 ) | ( x505 & ~n43269 ) | ( n43267 & ~n43269 ) ;
  assign n43271 = ( x505 & n42919 ) | ( x505 & ~n43270 ) | ( n42919 & ~n43270 ) ;
  assign n43272 = ~n43270 & n43271 ;
  assign n43273 = x241 | x500 ;
  assign n43274 = x241 & x500 ;
  assign n43275 = n43273 & ~n43274 ;
  assign n43276 = n43272 & ~n43275 ;
  assign n43277 = ~n43262 & n43276 ;
  assign n43278 = x497 & n43277 ;
  assign n43279 = x239 | n43278 ;
  assign n43280 = ~x497 & n43277 ;
  assign n43281 = x239 & ~n43280 ;
  assign n43282 = n43279 & ~n43281 ;
  assign n43283 = x539 & n43282 ;
  assign n43284 = x242 & ~n43283 ;
  assign n43285 = ~x539 & n43282 ;
  assign n43286 = x242 | n43285 ;
  assign n43287 = ~n43284 & n43286 ;
  assign n43288 = x540 & n43287 ;
  assign n43289 = x235 & ~n43288 ;
  assign n43290 = ~x540 & n43287 ;
  assign n43291 = x235 | n43290 ;
  assign n43292 = ~n43289 & n43291 ;
  assign n43293 = x541 ^ x244 ^ 1'b0 ;
  assign n43294 = n43292 & ~n43293 ;
  assign n43295 = x503 ^ x245 ^ 1'b0 ;
  assign n43296 = n43294 & ~n43295 ;
  assign n43297 = ~x502 & n43296 ;
  assign n43298 = x247 | n43297 ;
  assign n43299 = x502 & n43296 ;
  assign n43300 = x247 & ~n43299 ;
  assign n43301 = n43298 & ~n43300 ;
  assign n43302 = x238 & n43301 ;
  assign n43303 = x520 ^ x246 ^ 1'b0 ;
  assign n43304 = x578 ^ x249 ^ 1'b0 ;
  assign n43305 = x521 ^ x248 ^ 1'b0 ;
  assign n43306 = n43304 | n43305 ;
  assign n43307 = x574 ^ x241 ^ 1'b0 ;
  assign n43308 = ( ~n43303 & n43306 ) | ( ~n43303 & n43307 ) | ( n43306 & n43307 ) ;
  assign n43309 = n43303 | n43308 ;
  assign n43310 = x234 & n42935 ;
  assign n43311 = ~n43309 & n43310 ;
  assign n43312 = ( x518 & n43309 ) | ( x518 & ~n43311 ) | ( n43309 & ~n43311 ) ;
  assign n43313 = ( x518 & n42936 ) | ( x518 & ~n43312 ) | ( n42936 & ~n43312 ) ;
  assign n43314 = ~n43312 & n43313 ;
  assign n43315 = x582 & n43314 ;
  assign n43316 = x240 & ~n43315 ;
  assign n43317 = ~x582 & n43314 ;
  assign n43318 = x240 | n43317 ;
  assign n43319 = ~n43316 & n43318 ;
  assign n43320 = x519 ^ x239 ^ 1'b0 ;
  assign n43321 = n43319 & n43320 ;
  assign n43322 = x586 ^ x242 ^ 1'b0 ;
  assign n43323 = n43321 & ~n43322 ;
  assign n43324 = x581 ^ x235 ^ 1'b0 ;
  assign n43325 = n43323 & ~n43324 ;
  assign n43326 = x585 & n43325 ;
  assign n43327 = x244 & ~n43326 ;
  assign n43328 = ~x585 & n43325 ;
  assign n43329 = x244 | n43328 ;
  assign n43330 = ~n43327 & n43329 ;
  assign n43331 = x584 & n43330 ;
  assign n43332 = x245 & ~n43331 ;
  assign n43333 = ~x584 & n43330 ;
  assign n43334 = x245 | n43333 ;
  assign n43335 = ~n43332 & n43334 ;
  assign n43336 = x247 | x561 ;
  assign n43337 = x247 & x561 ;
  assign n43338 = n43336 & ~n43337 ;
  assign n43339 = n43335 & ~n43338 ;
  assign n43340 = ~x238 & n43339 ;
  assign n43341 = ( x522 & ~n43302 ) | ( x522 & n43340 ) | ( ~n43302 & n43340 ) ;
  assign n43342 = n43302 | n43341 ;
  assign n43343 = x584 & n43294 ;
  assign n43344 = x245 | n43343 ;
  assign n43345 = x585 & n43292 ;
  assign n43346 = x244 | n43345 ;
  assign n43347 = x540 & n43323 ;
  assign n43348 = x235 | n43347 ;
  assign n43349 = x539 & n43321 ;
  assign n43350 = x242 | n43349 ;
  assign n43351 = x582 & n43276 ;
  assign n43352 = x240 | n43351 ;
  assign n43353 = ~x500 & n43276 ;
  assign n43354 = n43272 & n43274 ;
  assign n43355 = ( n43314 & ~n43353 ) | ( n43314 & n43354 ) | ( ~n43353 & n43354 ) ;
  assign n43356 = n43353 | n43355 ;
  assign n43357 = ~x582 & n43356 ;
  assign n43358 = ( ~n43316 & n43352 ) | ( ~n43316 & n43357 ) | ( n43352 & n43357 ) ;
  assign n43359 = ~n43316 & n43358 ;
  assign n43360 = n43359 ^ x542 ^ 1'b0 ;
  assign n43361 = ( n43276 & n43318 ) | ( n43276 & n43319 ) | ( n43318 & n43319 ) ;
  assign n43362 = ( n43359 & n43360 ) | ( n43359 & n43361 ) | ( n43360 & n43361 ) ;
  assign n43363 = ~x497 & n43362 ;
  assign n43364 = x497 & n43319 ;
  assign n43365 = x239 & ~n43364 ;
  assign n43366 = n43279 & ~n43365 ;
  assign n43367 = ( n43279 & n43363 ) | ( n43279 & n43366 ) | ( n43363 & n43366 ) ;
  assign n43368 = ~x497 & n43319 ;
  assign n43369 = x239 | n43368 ;
  assign n43370 = x497 & n43362 ;
  assign n43371 = ( ~n43281 & n43369 ) | ( ~n43281 & n43370 ) | ( n43369 & n43370 ) ;
  assign n43372 = ~n43281 & n43371 ;
  assign n43373 = n43367 ^ x519 ^ 1'b0 ;
  assign n43374 = ( n43367 & n43372 ) | ( n43367 & n43373 ) | ( n43372 & n43373 ) ;
  assign n43375 = ~x539 & n43374 ;
  assign n43376 = ( ~n43284 & n43350 ) | ( ~n43284 & n43375 ) | ( n43350 & n43375 ) ;
  assign n43377 = ~n43284 & n43376 ;
  assign n43378 = x539 & n43374 ;
  assign n43379 = ~x539 & n43321 ;
  assign n43380 = x242 & ~n43379 ;
  assign n43381 = n43286 & ~n43380 ;
  assign n43382 = ( n43286 & n43378 ) | ( n43286 & n43381 ) | ( n43378 & n43381 ) ;
  assign n43383 = n43377 ^ x586 ^ 1'b0 ;
  assign n43384 = ( n43377 & n43382 ) | ( n43377 & n43383 ) | ( n43382 & n43383 ) ;
  assign n43385 = ~x540 & n43384 ;
  assign n43386 = ( ~n43289 & n43348 ) | ( ~n43289 & n43385 ) | ( n43348 & n43385 ) ;
  assign n43387 = ~n43289 & n43386 ;
  assign n43388 = x540 & n43384 ;
  assign n43389 = ~x540 & n43323 ;
  assign n43390 = x235 & ~n43389 ;
  assign n43391 = n43291 & ~n43390 ;
  assign n43392 = ( n43291 & n43388 ) | ( n43291 & n43391 ) | ( n43388 & n43391 ) ;
  assign n43393 = n43387 ^ x581 ^ 1'b0 ;
  assign n43394 = ( n43387 & n43392 ) | ( n43387 & n43393 ) | ( n43392 & n43393 ) ;
  assign n43395 = ~x585 & n43394 ;
  assign n43396 = ( ~n43327 & n43346 ) | ( ~n43327 & n43395 ) | ( n43346 & n43395 ) ;
  assign n43397 = ~n43327 & n43396 ;
  assign n43398 = x585 & n43394 ;
  assign n43399 = ~x585 & n43292 ;
  assign n43400 = x244 & ~n43399 ;
  assign n43401 = n43329 & ~n43400 ;
  assign n43402 = ( n43329 & n43398 ) | ( n43329 & n43401 ) | ( n43398 & n43401 ) ;
  assign n43403 = n43397 ^ x541 ^ 1'b0 ;
  assign n43404 = ( n43397 & n43402 ) | ( n43397 & n43403 ) | ( n43402 & n43403 ) ;
  assign n43405 = ~x584 & n43404 ;
  assign n43406 = ( ~n43332 & n43344 ) | ( ~n43332 & n43405 ) | ( n43344 & n43405 ) ;
  assign n43407 = ~n43332 & n43406 ;
  assign n43408 = ~x584 & n43294 ;
  assign n43409 = x584 & n43404 ;
  assign n43410 = ( x245 & n43408 ) | ( x245 & ~n43409 ) | ( n43408 & ~n43409 ) ;
  assign n43411 = ~n43408 & n43410 ;
  assign n43412 = ( x245 & n43333 ) | ( x245 & ~n43411 ) | ( n43333 & ~n43411 ) ;
  assign n43413 = ~n43411 & n43412 ;
  assign n43414 = n43407 ^ x503 ^ 1'b0 ;
  assign n43415 = ( n43407 & n43413 ) | ( n43407 & n43414 ) | ( n43413 & n43414 ) ;
  assign n43416 = x502 & ~n43415 ;
  assign n43417 = x502 | n43335 ;
  assign n43418 = ( x561 & n43416 ) | ( x561 & n43417 ) | ( n43416 & n43417 ) ;
  assign n43419 = ~n43416 & n43418 ;
  assign n43420 = ( n43300 & n43337 ) | ( n43300 & ~n43419 ) | ( n43337 & ~n43419 ) ;
  assign n43421 = ~n43419 & n43420 ;
  assign n43422 = n43298 & n43336 ;
  assign n43423 = x502 & ~n43335 ;
  assign n43424 = x561 | n43423 ;
  assign n43425 = ( n43415 & n43416 ) | ( n43415 & ~n43424 ) | ( n43416 & ~n43424 ) ;
  assign n43426 = ( ~n43421 & n43422 ) | ( ~n43421 & n43425 ) | ( n43422 & n43425 ) ;
  assign n43427 = ~n43421 & n43426 ;
  assign n43428 = x238 & n43427 ;
  assign n43429 = x522 & ~n43428 ;
  assign n43430 = x543 & ~n43429 ;
  assign n43431 = n43342 & n43430 ;
  assign n43432 = x238 & n43339 ;
  assign n43433 = x522 & ~n43432 ;
  assign n43434 = ~x238 & n43301 ;
  assign n43435 = ( x543 & n43433 ) | ( x543 & ~n43434 ) | ( n43433 & ~n43434 ) ;
  assign n43436 = n43435 ^ n43433 ^ 1'b0 ;
  assign n43437 = ( x543 & n43435 ) | ( x543 & ~n43436 ) | ( n43435 & ~n43436 ) ;
  assign n43438 = ~x238 & n43427 ;
  assign n43439 = ( x522 & ~n43437 ) | ( x522 & n43438 ) | ( ~n43437 & n43438 ) ;
  assign n43440 = ~n43437 & n43439 ;
  assign n43441 = ( ~x233 & n43431 ) | ( ~x233 & n43440 ) | ( n43431 & n43440 ) ;
  assign n43442 = ~x233 & n43441 ;
  assign n43443 = x536 ^ x246 ^ 1'b0 ;
  assign n43444 = x557 | n42919 ;
  assign n43445 = x557 & ~n43268 ;
  assign n43446 = ( n43443 & n43444 ) | ( n43443 & ~n43445 ) | ( n43444 & ~n43445 ) ;
  assign n43447 = ~n43443 & n43446 ;
  assign n43448 = ~x538 & n43447 ;
  assign n43449 = x538 & n43447 ;
  assign n43450 = n43448 ^ x249 ^ 1'b0 ;
  assign n43451 = ( n43448 & n43449 ) | ( n43448 & n43450 ) | ( n43449 & n43450 ) ;
  assign n43452 = ~x537 & n43451 ;
  assign n43453 = x248 | n43452 ;
  assign n43454 = x537 & n43451 ;
  assign n43455 = x248 & ~n43454 ;
  assign n43456 = n43453 & ~n43455 ;
  assign n43457 = x506 ^ x241 ^ 1'b0 ;
  assign n43458 = n43456 & ~n43457 ;
  assign n43459 = x535 ^ x240 ^ 1'b0 ;
  assign n43460 = n43458 & ~n43459 ;
  assign n43461 = x534 & n43460 ;
  assign n43462 = x239 | n43461 ;
  assign n43463 = ~x534 & n43460 ;
  assign n43464 = x239 & ~n43463 ;
  assign n43465 = n43462 & ~n43464 ;
  assign n43466 = x504 & n43465 ;
  assign n43467 = x242 & ~n43466 ;
  assign n43468 = ~x504 & n43465 ;
  assign n43469 = x242 | n43468 ;
  assign n43470 = ~n43467 & n43469 ;
  assign n43471 = x533 & n43470 ;
  assign n43472 = x235 & ~n43471 ;
  assign n43473 = ~x533 & n43470 ;
  assign n43474 = x235 | n43473 ;
  assign n43475 = ~n43472 & n43474 ;
  assign n43476 = x558 & n43475 ;
  assign n43477 = x244 & ~n43476 ;
  assign n43478 = ~x558 & n43475 ;
  assign n43479 = x244 | n43478 ;
  assign n43480 = ~n43477 & n43479 ;
  assign n43481 = x509 & n43480 ;
  assign n43482 = x245 & ~n43481 ;
  assign n43483 = ~x509 & n43480 ;
  assign n43484 = x245 | n43483 ;
  assign n43485 = ~n43482 & n43484 ;
  assign n43486 = x508 & n43485 ;
  assign n43487 = x247 & ~n43486 ;
  assign n43488 = ~x508 & n43485 ;
  assign n43489 = x247 | n43488 ;
  assign n43490 = ~n43487 & n43489 ;
  assign n43491 = x238 & n43490 ;
  assign n43492 = x481 ^ x248 ^ 1'b0 ;
  assign n43493 = x487 ^ x246 ^ 1'b0 ;
  assign n43494 = x511 | n42936 ;
  assign n43495 = x511 & ~n43310 ;
  assign n43496 = ( n43493 & n43494 ) | ( n43493 & ~n43495 ) | ( n43494 & ~n43495 ) ;
  assign n43497 = ~n43493 & n43496 ;
  assign n43498 = x579 ^ x249 ^ 1'b0 ;
  assign n43499 = n43497 & ~n43498 ;
  assign n43500 = ~n43492 & n43499 ;
  assign n43501 = x559 & n43500 ;
  assign n43502 = x241 & ~n43501 ;
  assign n43503 = ~x559 & n43500 ;
  assign n43504 = x241 | n43503 ;
  assign n43505 = ~n43502 & n43504 ;
  assign n43506 = x515 & n43505 ;
  assign n43507 = x240 & ~n43506 ;
  assign n43508 = ~x515 & n43505 ;
  assign n43509 = x240 | n43508 ;
  assign n43510 = ~n43507 & n43509 ;
  assign n43511 = x488 ^ x239 ^ 1'b0 ;
  assign n43512 = n43510 & n43511 ;
  assign n43513 = x510 ^ x242 ^ 1'b0 ;
  assign n43514 = n43512 & ~n43513 ;
  assign n43515 = x512 ^ x235 ^ 1'b0 ;
  assign n43516 = n43514 & ~n43515 ;
  assign n43517 = x513 ^ x244 ^ 1'b0 ;
  assign n43518 = n43516 & ~n43517 ;
  assign n43519 = x514 ^ x245 ^ 1'b0 ;
  assign n43520 = n43518 & ~n43519 ;
  assign n43521 = x516 ^ x247 ^ 1'b0 ;
  assign n43522 = n43520 & ~n43521 ;
  assign n43523 = ~x238 & n43522 ;
  assign n43524 = ( x517 & ~n43491 ) | ( x517 & n43523 ) | ( ~n43491 & n43523 ) ;
  assign n43525 = n43491 | n43524 ;
  assign n43526 = ~x508 & n43520 ;
  assign n43527 = x509 & n43518 ;
  assign n43528 = x245 | n43527 ;
  assign n43529 = x558 & n43516 ;
  assign n43530 = x244 | n43529 ;
  assign n43531 = x533 & n43514 ;
  assign n43532 = x235 | n43531 ;
  assign n43533 = x504 & n43512 ;
  assign n43534 = x242 | n43533 ;
  assign n43535 = x515 & n43458 ;
  assign n43536 = x240 | n43535 ;
  assign n43537 = x559 & n43456 ;
  assign n43538 = x241 | n43537 ;
  assign n43539 = x537 & n43499 ;
  assign n43540 = x248 | n43539 ;
  assign n43541 = x249 | n43448 ;
  assign n43542 = n43497 & n43541 ;
  assign n43543 = n43499 ^ x579 ^ 1'b0 ;
  assign n43544 = ( n43499 & n43542 ) | ( n43499 & n43543 ) | ( n43542 & n43543 ) ;
  assign n43545 = x249 & ~n43449 ;
  assign n43546 = ~n43544 & n43545 ;
  assign n43547 = ( n43541 & n43544 ) | ( n43541 & ~n43546 ) | ( n43544 & ~n43546 ) ;
  assign n43548 = ~x537 & n43547 ;
  assign n43549 = ( ~n43455 & n43540 ) | ( ~n43455 & n43548 ) | ( n43540 & n43548 ) ;
  assign n43550 = ~n43455 & n43549 ;
  assign n43551 = x537 & n43547 ;
  assign n43552 = ~x537 & n43499 ;
  assign n43553 = x248 & ~n43552 ;
  assign n43554 = n43453 & ~n43553 ;
  assign n43555 = ( n43453 & n43551 ) | ( n43453 & n43554 ) | ( n43551 & n43554 ) ;
  assign n43556 = n43550 ^ x481 ^ 1'b0 ;
  assign n43557 = ( n43550 & n43555 ) | ( n43550 & n43556 ) | ( n43555 & n43556 ) ;
  assign n43558 = ~x559 & n43557 ;
  assign n43559 = ( ~n43502 & n43538 ) | ( ~n43502 & n43558 ) | ( n43538 & n43558 ) ;
  assign n43560 = ~n43502 & n43559 ;
  assign n43561 = x559 & n43557 ;
  assign n43562 = ~x559 & n43456 ;
  assign n43563 = x241 & ~n43562 ;
  assign n43564 = n43504 & ~n43563 ;
  assign n43565 = ( n43504 & n43561 ) | ( n43504 & n43564 ) | ( n43561 & n43564 ) ;
  assign n43566 = n43560 ^ x506 ^ 1'b0 ;
  assign n43567 = ( n43560 & n43565 ) | ( n43560 & n43566 ) | ( n43565 & n43566 ) ;
  assign n43568 = ~x515 & n43567 ;
  assign n43569 = ( ~n43507 & n43536 ) | ( ~n43507 & n43568 ) | ( n43536 & n43568 ) ;
  assign n43570 = ~n43507 & n43569 ;
  assign n43571 = ~x515 & n43458 ;
  assign n43572 = x515 & n43567 ;
  assign n43573 = ( x240 & n43571 ) | ( x240 & ~n43572 ) | ( n43571 & ~n43572 ) ;
  assign n43574 = ~n43571 & n43573 ;
  assign n43575 = ( x240 & n43508 ) | ( x240 & ~n43574 ) | ( n43508 & ~n43574 ) ;
  assign n43576 = ~n43574 & n43575 ;
  assign n43577 = n43570 ^ x535 ^ 1'b0 ;
  assign n43578 = ( n43570 & n43576 ) | ( n43570 & n43577 ) | ( n43576 & n43577 ) ;
  assign n43579 = ~x534 & n43578 ;
  assign n43580 = x534 & n43510 ;
  assign n43581 = x239 & ~n43580 ;
  assign n43582 = n43462 & ~n43581 ;
  assign n43583 = ( n43462 & n43579 ) | ( n43462 & n43582 ) | ( n43579 & n43582 ) ;
  assign n43584 = ~x534 & n43510 ;
  assign n43585 = x239 | n43584 ;
  assign n43586 = x534 & n43578 ;
  assign n43587 = ( ~n43464 & n43585 ) | ( ~n43464 & n43586 ) | ( n43585 & n43586 ) ;
  assign n43588 = ~n43464 & n43587 ;
  assign n43589 = n43583 ^ x488 ^ 1'b0 ;
  assign n43590 = ( n43583 & n43588 ) | ( n43583 & n43589 ) | ( n43588 & n43589 ) ;
  assign n43591 = ~x504 & n43590 ;
  assign n43592 = ( ~n43467 & n43534 ) | ( ~n43467 & n43591 ) | ( n43534 & n43591 ) ;
  assign n43593 = ~n43467 & n43592 ;
  assign n43594 = x504 & n43590 ;
  assign n43595 = ~x504 & n43512 ;
  assign n43596 = x242 & ~n43595 ;
  assign n43597 = n43469 & ~n43596 ;
  assign n43598 = ( n43469 & n43594 ) | ( n43469 & n43597 ) | ( n43594 & n43597 ) ;
  assign n43599 = n43593 ^ x510 ^ 1'b0 ;
  assign n43600 = ( n43593 & n43598 ) | ( n43593 & n43599 ) | ( n43598 & n43599 ) ;
  assign n43601 = ~x533 & n43600 ;
  assign n43602 = ( ~n43472 & n43532 ) | ( ~n43472 & n43601 ) | ( n43532 & n43601 ) ;
  assign n43603 = ~n43472 & n43602 ;
  assign n43604 = x533 & n43600 ;
  assign n43605 = ~x533 & n43514 ;
  assign n43606 = x235 & ~n43605 ;
  assign n43607 = n43474 & ~n43606 ;
  assign n43608 = ( n43474 & n43604 ) | ( n43474 & n43607 ) | ( n43604 & n43607 ) ;
  assign n43609 = n43603 ^ x512 ^ 1'b0 ;
  assign n43610 = ( n43603 & n43608 ) | ( n43603 & n43609 ) | ( n43608 & n43609 ) ;
  assign n43611 = ~x558 & n43610 ;
  assign n43612 = ( ~n43477 & n43530 ) | ( ~n43477 & n43611 ) | ( n43530 & n43611 ) ;
  assign n43613 = ~n43477 & n43612 ;
  assign n43614 = x558 & n43610 ;
  assign n43615 = ~x558 & n43516 ;
  assign n43616 = x244 & ~n43615 ;
  assign n43617 = n43479 & ~n43616 ;
  assign n43618 = ( n43479 & n43614 ) | ( n43479 & n43617 ) | ( n43614 & n43617 ) ;
  assign n43619 = n43613 ^ x513 ^ 1'b0 ;
  assign n43620 = ( n43613 & n43618 ) | ( n43613 & n43619 ) | ( n43618 & n43619 ) ;
  assign n43621 = ~x509 & n43620 ;
  assign n43622 = ( ~n43482 & n43528 ) | ( ~n43482 & n43621 ) | ( n43528 & n43621 ) ;
  assign n43623 = ~n43482 & n43622 ;
  assign n43624 = x509 & n43620 ;
  assign n43625 = ~x509 & n43518 ;
  assign n43626 = x245 & ~n43625 ;
  assign n43627 = n43484 & ~n43626 ;
  assign n43628 = ( n43484 & n43624 ) | ( n43484 & n43627 ) | ( n43624 & n43627 ) ;
  assign n43629 = n43623 ^ x514 ^ 1'b0 ;
  assign n43630 = ( n43623 & n43628 ) | ( n43623 & n43629 ) | ( n43628 & n43629 ) ;
  assign n43631 = x508 & n43630 ;
  assign n43632 = ( x247 & n43526 ) | ( x247 & ~n43631 ) | ( n43526 & ~n43631 ) ;
  assign n43633 = ~n43526 & n43632 ;
  assign n43634 = x516 & ~n43489 ;
  assign n43635 = ( x516 & n43633 ) | ( x516 & n43634 ) | ( n43633 & n43634 ) ;
  assign n43636 = x508 & n43520 ;
  assign n43637 = x247 | n43636 ;
  assign n43638 = ~x508 & n43630 ;
  assign n43639 = ( ~n43487 & n43637 ) | ( ~n43487 & n43638 ) | ( n43637 & n43638 ) ;
  assign n43640 = ~n43487 & n43639 ;
  assign n43641 = ( x516 & ~n43635 ) | ( x516 & n43640 ) | ( ~n43635 & n43640 ) ;
  assign n43642 = ~n43635 & n43641 ;
  assign n43643 = x238 & n43642 ;
  assign n43644 = x517 & ~n43643 ;
  assign n43645 = x507 & ~n43644 ;
  assign n43646 = n43525 & n43645 ;
  assign n43647 = x238 & n43522 ;
  assign n43648 = x517 & ~n43647 ;
  assign n43649 = ~x238 & n43490 ;
  assign n43650 = ( x507 & n43648 ) | ( x507 & ~n43649 ) | ( n43648 & ~n43649 ) ;
  assign n43651 = n43650 ^ n43648 ^ 1'b0 ;
  assign n43652 = ( x507 & n43650 ) | ( x507 & ~n43651 ) | ( n43650 & ~n43651 ) ;
  assign n43653 = ~x238 & n43642 ;
  assign n43654 = ( x517 & ~n43652 ) | ( x517 & n43653 ) | ( ~n43652 & n43653 ) ;
  assign n43655 = ~n43652 & n43654 ;
  assign n43656 = ( x233 & n43646 ) | ( x233 & n43655 ) | ( n43646 & n43655 ) ;
  assign n43657 = n43655 ^ n43646 ^ 1'b0 ;
  assign n43658 = ( x233 & n43656 ) | ( x233 & n43657 ) | ( n43656 & n43657 ) ;
  assign n43659 = ( x237 & n43442 ) | ( x237 & ~n43658 ) | ( n43442 & ~n43658 ) ;
  assign n43660 = ~n43442 & n43659 ;
  assign n43661 = x237 ^ x233 ^ 1'b0 ;
  assign n43662 = ~x246 & x564 ;
  assign n43663 = n43662 ^ x249 ^ 1'b0 ;
  assign n43664 = ( x249 & x482 ) | ( x249 & n43663 ) | ( x482 & n43663 ) ;
  assign n43665 = n43664 ^ n43662 ^ x482 ;
  assign n43666 = n43665 ^ x241 ^ 1'b0 ;
  assign n43667 = ( x241 & x562 ) | ( x241 & n43666 ) | ( x562 & n43666 ) ;
  assign n43668 = n43667 ^ n43665 ^ x562 ;
  assign n43669 = n43310 & ~n43668 ;
  assign n43670 = ( x570 & n43668 ) | ( x570 & ~n43669 ) | ( n43668 & ~n43669 ) ;
  assign n43671 = ( x570 & n42936 ) | ( x570 & ~n43670 ) | ( n42936 & ~n43670 ) ;
  assign n43672 = ~n43670 & n43671 ;
  assign n43673 = x565 ^ x248 ^ 1'b0 ;
  assign n43674 = x246 & ~x564 ;
  assign n43675 = x560 & ~n43674 ;
  assign n43676 = ~n43673 & n43675 ;
  assign n43677 = x240 & ~n43676 ;
  assign n43678 = ( x240 & ~n43672 ) | ( x240 & n43677 ) | ( ~n43672 & n43677 ) ;
  assign n43679 = x560 ^ x240 ^ 1'b0 ;
  assign n43680 = n43673 | n43674 ;
  assign n43681 = ( n43672 & n43679 ) | ( n43672 & ~n43680 ) | ( n43679 & ~n43680 ) ;
  assign n43682 = ~n43679 & n43681 ;
  assign n43683 = ( x240 & ~n43678 ) | ( x240 & n43682 ) | ( ~n43678 & n43682 ) ;
  assign n43684 = ~n43678 & n43683 ;
  assign n43685 = x569 ^ x239 ^ 1'b0 ;
  assign n43686 = n43684 & n43685 ;
  assign n43687 = x242 | x556 ;
  assign n43688 = x242 & x556 ;
  assign n43689 = n43687 & ~n43688 ;
  assign n43690 = n43686 & ~n43689 ;
  assign n43691 = x531 ^ x235 ^ 1'b0 ;
  assign n43692 = n43690 & ~n43691 ;
  assign n43693 = x566 ^ x244 ^ 1'b0 ;
  assign n43694 = n43692 & ~n43693 ;
  assign n43695 = x568 & n43694 ;
  assign n43696 = x245 & ~n43695 ;
  assign n43697 = ~x568 & n43694 ;
  assign n43698 = x245 | n43697 ;
  assign n43699 = ~n43696 & n43698 ;
  assign n43700 = ~x552 & n43699 ;
  assign n43701 = x553 ^ x241 ^ 1'b0 ;
  assign n43702 = x551 ^ x240 ^ 1'b0 ;
  assign n43703 = x555 ^ x249 ^ 1'b0 ;
  assign n43704 = ( ~n43701 & n43702 ) | ( ~n43701 & n43703 ) | ( n43702 & n43703 ) ;
  assign n43705 = n43701 | n43704 ;
  assign n43706 = x554 ^ x248 ^ 1'b0 ;
  assign n43707 = x563 ^ x246 ^ 1'b0 ;
  assign n43708 = ( ~n43705 & n43706 ) | ( ~n43705 & n43707 ) | ( n43706 & n43707 ) ;
  assign n43709 = n43705 | n43708 ;
  assign n43710 = n43268 & ~n43709 ;
  assign n43711 = ( x485 & n43709 ) | ( x485 & ~n43710 ) | ( n43709 & ~n43710 ) ;
  assign n43712 = ( x485 & n42919 ) | ( x485 & ~n43711 ) | ( n42919 & ~n43711 ) ;
  assign n43713 = ~n43711 & n43712 ;
  assign n43714 = x550 & n43713 ;
  assign n43715 = ~x550 & n43713 ;
  assign n43716 = n43714 ^ x239 ^ 1'b0 ;
  assign n43717 = ( n43714 & n43715 ) | ( n43714 & n43716 ) | ( n43715 & n43716 ) ;
  assign n43718 = ~x489 & n43717 ;
  assign n43719 = x242 | n43718 ;
  assign n43720 = x489 & n43717 ;
  assign n43721 = x242 & ~n43720 ;
  assign n43722 = n43719 & ~n43721 ;
  assign n43723 = x549 & n43722 ;
  assign n43724 = x235 & ~n43723 ;
  assign n43725 = ~x549 & n43722 ;
  assign n43726 = x235 | n43725 ;
  assign n43727 = ~n43724 & n43726 ;
  assign n43728 = x486 & n43727 ;
  assign n43729 = x244 & ~n43728 ;
  assign n43730 = ~x486 & n43727 ;
  assign n43731 = x244 | n43730 ;
  assign n43732 = ~n43729 & n43731 ;
  assign n43733 = x568 & n43732 ;
  assign n43734 = x245 | n43733 ;
  assign n43735 = x486 & n43692 ;
  assign n43736 = x244 | n43735 ;
  assign n43737 = x549 & n43690 ;
  assign n43738 = x235 | n43737 ;
  assign n43739 = x489 | n43686 ;
  assign n43740 = x239 & ~n43715 ;
  assign n43741 = x569 & ~n43740 ;
  assign n43742 = n43684 & n43741 ;
  assign n43743 = x239 & ~x569 ;
  assign n43744 = n43682 & n43743 ;
  assign n43745 = ( n43717 & ~n43742 ) | ( n43717 & n43744 ) | ( ~n43742 & n43744 ) ;
  assign n43746 = n43742 | n43745 ;
  assign n43747 = x489 & ~n43746 ;
  assign n43748 = x556 & ~n43747 ;
  assign n43749 = n43739 & n43748 ;
  assign n43750 = n43721 & ~n43749 ;
  assign n43751 = x489 | n43746 ;
  assign n43752 = x489 & ~n43686 ;
  assign n43753 = ( x556 & n43751 ) | ( x556 & ~n43752 ) | ( n43751 & ~n43752 ) ;
  assign n43754 = ~x556 & n43753 ;
  assign n43755 = n43687 & n43719 ;
  assign n43756 = ( ~n43750 & n43754 ) | ( ~n43750 & n43755 ) | ( n43754 & n43755 ) ;
  assign n43757 = ~n43750 & n43756 ;
  assign n43758 = ~x549 & n43757 ;
  assign n43759 = ( ~n43724 & n43738 ) | ( ~n43724 & n43758 ) | ( n43738 & n43758 ) ;
  assign n43760 = ~n43724 & n43759 ;
  assign n43761 = x549 & n43757 ;
  assign n43762 = ~x549 & n43690 ;
  assign n43763 = x235 & ~n43762 ;
  assign n43764 = n43726 & ~n43763 ;
  assign n43765 = ( n43726 & n43761 ) | ( n43726 & n43764 ) | ( n43761 & n43764 ) ;
  assign n43766 = n43760 ^ x531 ^ 1'b0 ;
  assign n43767 = ( n43760 & n43765 ) | ( n43760 & n43766 ) | ( n43765 & n43766 ) ;
  assign n43768 = ~x486 & n43767 ;
  assign n43769 = ( ~n43729 & n43736 ) | ( ~n43729 & n43768 ) | ( n43736 & n43768 ) ;
  assign n43770 = ~n43729 & n43769 ;
  assign n43771 = x486 & n43767 ;
  assign n43772 = ~x486 & n43692 ;
  assign n43773 = x244 & ~n43772 ;
  assign n43774 = n43731 & ~n43773 ;
  assign n43775 = ( n43731 & n43771 ) | ( n43731 & n43774 ) | ( n43771 & n43774 ) ;
  assign n43776 = n43770 ^ x566 ^ 1'b0 ;
  assign n43777 = ( n43770 & n43775 ) | ( n43770 & n43776 ) | ( n43775 & n43776 ) ;
  assign n43778 = ~x568 & n43777 ;
  assign n43779 = ( ~n43696 & n43734 ) | ( ~n43696 & n43778 ) | ( n43734 & n43778 ) ;
  assign n43780 = ~n43696 & n43779 ;
  assign n43781 = ~x568 & n43732 ;
  assign n43782 = x568 & n43777 ;
  assign n43783 = ( x245 & n43781 ) | ( x245 & ~n43782 ) | ( n43781 & ~n43782 ) ;
  assign n43784 = ~n43781 & n43783 ;
  assign n43785 = ( x245 & n43697 ) | ( x245 & ~n43784 ) | ( n43697 & ~n43784 ) ;
  assign n43786 = ~n43784 & n43785 ;
  assign n43787 = n43780 ^ x580 ^ 1'b0 ;
  assign n43788 = ( n43780 & n43786 ) | ( n43780 & n43787 ) | ( n43786 & n43787 ) ;
  assign n43789 = x552 & n43788 ;
  assign n43790 = ( x247 & n43700 ) | ( x247 & ~n43789 ) | ( n43700 & ~n43789 ) ;
  assign n43791 = ~n43700 & n43790 ;
  assign n43792 = x580 ^ x245 ^ 1'b0 ;
  assign n43793 = n43732 & ~n43792 ;
  assign n43794 = ~x552 & n43793 ;
  assign n43795 = x247 | n43794 ;
  assign n43796 = x532 & ~n43795 ;
  assign n43797 = ( x532 & n43791 ) | ( x532 & n43796 ) | ( n43791 & n43796 ) ;
  assign n43798 = x552 & n43793 ;
  assign n43799 = x247 & ~n43798 ;
  assign n43800 = x552 & n43699 ;
  assign n43801 = x247 | n43800 ;
  assign n43802 = ~x552 & n43788 ;
  assign n43803 = ( ~n43799 & n43801 ) | ( ~n43799 & n43802 ) | ( n43801 & n43802 ) ;
  assign n43804 = ~n43799 & n43803 ;
  assign n43805 = ( x532 & ~n43797 ) | ( x532 & n43804 ) | ( ~n43797 & n43804 ) ;
  assign n43806 = ~n43797 & n43805 ;
  assign n43807 = ~x238 & n43806 ;
  assign n43808 = x577 | n43807 ;
  assign n43809 = n43795 & ~n43799 ;
  assign n43810 = ~x238 & n43809 ;
  assign n43811 = x532 ^ x247 ^ 1'b0 ;
  assign n43812 = n43699 & ~n43811 ;
  assign n43813 = x238 & n43812 ;
  assign n43814 = ( x577 & ~n43810 ) | ( x577 & n43813 ) | ( ~n43810 & n43813 ) ;
  assign n43815 = n43810 | n43814 ;
  assign n43816 = x238 & n43806 ;
  assign n43817 = x577 & ~n43816 ;
  assign n43818 = x498 & ~n43817 ;
  assign n43819 = n43815 & n43818 ;
  assign n43820 = ~x238 & n43812 ;
  assign n43821 = x577 & ~n43820 ;
  assign n43822 = x238 & n43809 ;
  assign n43823 = ( x498 & n43821 ) | ( x498 & ~n43822 ) | ( n43821 & ~n43822 ) ;
  assign n43824 = n43823 ^ n43821 ^ 1'b0 ;
  assign n43825 = ( x498 & n43823 ) | ( x498 & ~n43824 ) | ( n43823 & ~n43824 ) ;
  assign n43826 = ~n43819 & n43825 ;
  assign n43827 = ( n43808 & n43819 ) | ( n43808 & ~n43826 ) | ( n43819 & ~n43826 ) ;
  assign n43828 = ( x233 & ~n43661 ) | ( x233 & n43827 ) | ( ~n43661 & n43827 ) ;
  assign n43829 = ( ~x233 & x237 ) | ( ~x233 & n43828 ) | ( x237 & n43828 ) ;
  assign n43830 = x490 ^ x241 ^ 1'b0 ;
  assign n43831 = x484 ^ x249 ^ 1'b0 ;
  assign n43832 = x546 ^ x246 ^ 1'b0 ;
  assign n43833 = x548 ^ x248 ^ 1'b0 ;
  assign n43834 = ( ~n43831 & n43832 ) | ( ~n43831 & n43833 ) | ( n43832 & n43833 ) ;
  assign n43835 = n43831 | n43834 ;
  assign n43836 = ( x544 & n42919 ) | ( x544 & ~n43835 ) | ( n42919 & ~n43835 ) ;
  assign n43837 = ~n43835 & n43836 ;
  assign n43838 = n43837 ^ n43268 ^ 1'b0 ;
  assign n43839 = ( ~x544 & n43268 ) | ( ~x544 & n43838 ) | ( n43268 & n43838 ) ;
  assign n43840 = ( n43837 & ~n43838 ) | ( n43837 & n43839 ) | ( ~n43838 & n43839 ) ;
  assign n43841 = ~n43830 & n43840 ;
  assign n43842 = x240 | x492 ;
  assign n43843 = x240 & x492 ;
  assign n43844 = n43842 & ~n43843 ;
  assign n43845 = n43841 & ~n43844 ;
  assign n43846 = x494 & n43845 ;
  assign n43847 = x239 | n43846 ;
  assign n43848 = ~x494 & n43845 ;
  assign n43849 = x239 & ~n43848 ;
  assign n43850 = n43847 & ~n43849 ;
  assign n43851 = x483 & n43850 ;
  assign n43852 = x242 & ~n43851 ;
  assign n43853 = ~x483 & n43850 ;
  assign n43854 = x242 | n43853 ;
  assign n43855 = ~n43852 & n43854 ;
  assign n43856 = x495 & n43855 ;
  assign n43857 = x235 & ~n43856 ;
  assign n43858 = ~x495 & n43855 ;
  assign n43859 = x235 | n43858 ;
  assign n43860 = ~n43857 & n43859 ;
  assign n43861 = x493 ^ x244 ^ 1'b0 ;
  assign n43862 = n43860 & ~n43861 ;
  assign n43863 = x545 & n43862 ;
  assign n43864 = x245 & ~n43863 ;
  assign n43865 = ~x545 & n43862 ;
  assign n43866 = x245 | n43865 ;
  assign n43867 = ~n43864 & n43866 ;
  assign n43868 = x547 & n43867 ;
  assign n43869 = x247 & ~n43868 ;
  assign n43870 = ~x547 & n43867 ;
  assign n43871 = x247 | n43870 ;
  assign n43872 = ~n43869 & n43871 ;
  assign n43873 = x238 & n43872 ;
  assign n43874 = x528 ^ x249 ^ 1'b0 ;
  assign n43875 = x526 ^ x246 ^ 1'b0 ;
  assign n43876 = x576 ^ x248 ^ 1'b0 ;
  assign n43877 = ( ~n43874 & n43875 ) | ( ~n43874 & n43876 ) | ( n43875 & n43876 ) ;
  assign n43878 = n43874 | n43877 ;
  assign n43879 = n43310 & ~n43878 ;
  assign n43880 = ( x523 & n43878 ) | ( x523 & ~n43879 ) | ( n43878 & ~n43879 ) ;
  assign n43881 = ( x523 & n42936 ) | ( x523 & ~n43880 ) | ( n42936 & ~n43880 ) ;
  assign n43882 = ~n43880 & n43881 ;
  assign n43883 = x571 & n43882 ;
  assign n43884 = x241 & ~n43883 ;
  assign n43885 = ~x571 & n43882 ;
  assign n43886 = x241 | n43885 ;
  assign n43887 = ~n43884 & n43886 ;
  assign n43888 = ~x530 & n43887 ;
  assign n43889 = x240 | n43888 ;
  assign n43890 = x530 & n43887 ;
  assign n43891 = x240 & ~n43890 ;
  assign n43892 = n43889 & ~n43891 ;
  assign n43893 = x524 ^ x239 ^ 1'b0 ;
  assign n43894 = n43892 & n43893 ;
  assign n43895 = x573 ^ x242 ^ 1'b0 ;
  assign n43896 = n43894 & ~n43895 ;
  assign n43897 = x575 ^ x235 ^ 1'b0 ;
  assign n43898 = n43896 & ~n43897 ;
  assign n43899 = x572 & n43898 ;
  assign n43900 = x244 & ~n43899 ;
  assign n43901 = ~x572 & n43898 ;
  assign n43902 = x244 | n43901 ;
  assign n43903 = ~n43900 & n43902 ;
  assign n43904 = x525 ^ x245 ^ 1'b0 ;
  assign n43905 = n43903 & ~n43904 ;
  assign n43906 = x527 ^ x247 ^ 1'b0 ;
  assign n43907 = n43905 & ~n43906 ;
  assign n43908 = ~x238 & n43907 ;
  assign n43909 = ( x529 & ~n43873 ) | ( x529 & n43908 ) | ( ~n43873 & n43908 ) ;
  assign n43910 = n43873 | n43909 ;
  assign n43911 = x547 & n43905 ;
  assign n43912 = x247 | n43911 ;
  assign n43913 = x545 & n43903 ;
  assign n43914 = x245 | n43913 ;
  assign n43915 = x572 & n43860 ;
  assign n43916 = x244 | n43915 ;
  assign n43917 = x495 & n43896 ;
  assign n43918 = x235 | n43917 ;
  assign n43919 = x483 & n43894 ;
  assign n43920 = x242 | n43919 ;
  assign n43921 = ( n43840 & ~n43884 ) | ( n43840 & n43887 ) | ( ~n43884 & n43887 ) ;
  assign n43922 = n43921 ^ x490 ^ 1'b0 ;
  assign n43923 = ( n43840 & n43886 ) | ( n43840 & n43887 ) | ( n43886 & n43887 ) ;
  assign n43924 = ( n43921 & n43922 ) | ( n43921 & n43923 ) | ( n43922 & n43923 ) ;
  assign n43925 = x530 & ~n43924 ;
  assign n43926 = x530 | n43841 ;
  assign n43927 = ( x492 & n43925 ) | ( x492 & n43926 ) | ( n43925 & n43926 ) ;
  assign n43928 = ~n43925 & n43927 ;
  assign n43929 = ( n43843 & n43891 ) | ( n43843 & ~n43928 ) | ( n43891 & ~n43928 ) ;
  assign n43930 = ~n43928 & n43929 ;
  assign n43931 = n43842 & n43889 ;
  assign n43932 = x530 & ~n43841 ;
  assign n43933 = x492 | n43932 ;
  assign n43934 = ( x530 & n43924 ) | ( x530 & ~n43933 ) | ( n43924 & ~n43933 ) ;
  assign n43935 = ~n43933 & n43934 ;
  assign n43936 = ( ~n43930 & n43931 ) | ( ~n43930 & n43935 ) | ( n43931 & n43935 ) ;
  assign n43937 = ~n43930 & n43936 ;
  assign n43938 = ~x494 & n43937 ;
  assign n43939 = x494 & n43892 ;
  assign n43940 = x239 & ~n43939 ;
  assign n43941 = n43847 & ~n43940 ;
  assign n43942 = ( n43847 & n43938 ) | ( n43847 & n43941 ) | ( n43938 & n43941 ) ;
  assign n43943 = ~x494 & n43892 ;
  assign n43944 = x239 | n43943 ;
  assign n43945 = x494 & n43937 ;
  assign n43946 = ( ~n43849 & n43944 ) | ( ~n43849 & n43945 ) | ( n43944 & n43945 ) ;
  assign n43947 = ~n43849 & n43946 ;
  assign n43948 = n43942 ^ x524 ^ 1'b0 ;
  assign n43949 = ( n43942 & n43947 ) | ( n43942 & n43948 ) | ( n43947 & n43948 ) ;
  assign n43950 = ~x483 & n43949 ;
  assign n43951 = ( ~n43852 & n43920 ) | ( ~n43852 & n43950 ) | ( n43920 & n43950 ) ;
  assign n43952 = ~n43852 & n43951 ;
  assign n43953 = x483 & n43949 ;
  assign n43954 = ~x483 & n43894 ;
  assign n43955 = x242 & ~n43954 ;
  assign n43956 = n43854 & ~n43955 ;
  assign n43957 = ( n43854 & n43953 ) | ( n43854 & n43956 ) | ( n43953 & n43956 ) ;
  assign n43958 = n43952 ^ x573 ^ 1'b0 ;
  assign n43959 = ( n43952 & n43957 ) | ( n43952 & n43958 ) | ( n43957 & n43958 ) ;
  assign n43960 = ~x495 & n43959 ;
  assign n43961 = ( ~n43857 & n43918 ) | ( ~n43857 & n43960 ) | ( n43918 & n43960 ) ;
  assign n43962 = ~n43857 & n43961 ;
  assign n43963 = x495 & n43959 ;
  assign n43964 = ~x495 & n43896 ;
  assign n43965 = x235 & ~n43964 ;
  assign n43966 = n43859 & ~n43965 ;
  assign n43967 = ( n43859 & n43963 ) | ( n43859 & n43966 ) | ( n43963 & n43966 ) ;
  assign n43968 = n43962 ^ x575 ^ 1'b0 ;
  assign n43969 = ( n43962 & n43967 ) | ( n43962 & n43968 ) | ( n43967 & n43968 ) ;
  assign n43970 = ~x572 & n43969 ;
  assign n43971 = ( ~n43900 & n43916 ) | ( ~n43900 & n43970 ) | ( n43916 & n43970 ) ;
  assign n43972 = ~n43900 & n43971 ;
  assign n43973 = ~x572 & n43860 ;
  assign n43974 = x572 & n43969 ;
  assign n43975 = ( x244 & n43973 ) | ( x244 & ~n43974 ) | ( n43973 & ~n43974 ) ;
  assign n43976 = ~n43973 & n43975 ;
  assign n43977 = ( x244 & n43901 ) | ( x244 & ~n43976 ) | ( n43901 & ~n43976 ) ;
  assign n43978 = ~n43976 & n43977 ;
  assign n43979 = n43972 ^ x493 ^ 1'b0 ;
  assign n43980 = ( n43972 & n43978 ) | ( n43972 & n43979 ) | ( n43978 & n43979 ) ;
  assign n43981 = ~x545 & n43980 ;
  assign n43982 = ( ~n43864 & n43914 ) | ( ~n43864 & n43981 ) | ( n43914 & n43981 ) ;
  assign n43983 = ~n43864 & n43982 ;
  assign n43984 = x545 & n43980 ;
  assign n43985 = ~x545 & n43903 ;
  assign n43986 = x245 & ~n43985 ;
  assign n43987 = n43866 & ~n43986 ;
  assign n43988 = ( n43866 & n43984 ) | ( n43866 & n43987 ) | ( n43984 & n43987 ) ;
  assign n43989 = n43983 ^ x525 ^ 1'b0 ;
  assign n43990 = ( n43983 & n43988 ) | ( n43983 & n43989 ) | ( n43988 & n43989 ) ;
  assign n43991 = ~x547 & n43990 ;
  assign n43992 = ( ~n43869 & n43912 ) | ( ~n43869 & n43991 ) | ( n43912 & n43991 ) ;
  assign n43993 = ~n43869 & n43992 ;
  assign n43994 = ~x547 & n43905 ;
  assign n43995 = x547 & n43990 ;
  assign n43996 = ( x247 & n43994 ) | ( x247 & ~n43995 ) | ( n43994 & ~n43995 ) ;
  assign n43997 = ~n43994 & n43996 ;
  assign n43998 = ( x247 & n43870 ) | ( x247 & ~n43997 ) | ( n43870 & ~n43997 ) ;
  assign n43999 = ~n43997 & n43998 ;
  assign n44000 = n43993 ^ x527 ^ 1'b0 ;
  assign n44001 = ( n43993 & n43999 ) | ( n43993 & n44000 ) | ( n43999 & n44000 ) ;
  assign n44002 = x238 & n44001 ;
  assign n44003 = x529 & ~n44002 ;
  assign n44004 = x491 & ~n44003 ;
  assign n44005 = n43910 & n44004 ;
  assign n44006 = x238 & n43907 ;
  assign n44007 = x529 & ~n44006 ;
  assign n44008 = ~x238 & n43872 ;
  assign n44009 = ( x491 & n44007 ) | ( x491 & ~n44008 ) | ( n44007 & ~n44008 ) ;
  assign n44010 = n44009 ^ n44007 ^ 1'b0 ;
  assign n44011 = ( x491 & n44009 ) | ( x491 & ~n44010 ) | ( n44009 & ~n44010 ) ;
  assign n44012 = ~x238 & n44001 ;
  assign n44013 = ( x529 & ~n44011 ) | ( x529 & n44012 ) | ( ~n44011 & n44012 ) ;
  assign n44014 = ~n44011 & n44013 ;
  assign n44015 = ( x233 & n44005 ) | ( x233 & n44014 ) | ( n44005 & n44014 ) ;
  assign n44016 = n44014 ^ n44005 ^ 1'b0 ;
  assign n44017 = ( x233 & n44015 ) | ( x233 & n44016 ) | ( n44015 & n44016 ) ;
  assign n44018 = ( ~n43660 & n43829 ) | ( ~n43660 & n44017 ) | ( n43829 & n44017 ) ;
  assign n44019 = ~n43660 & n44018 ;
  assign n44020 = ~x806 & n42621 ;
  assign n44021 = x332 | x806 ;
  assign n44022 = x990 & ~n44021 ;
  assign n44023 = x600 & n44022 ;
  assign n44024 = ~x332 & x594 ;
  assign n44025 = ( ~n44020 & n44023 ) | ( ~n44020 & n44024 ) | ( n44023 & n44024 ) ;
  assign n44026 = ~n44020 & n44025 ;
  assign n44027 = x601 & n42637 ;
  assign n44028 = x605 & ~x806 ;
  assign n44029 = n44027 & n44028 ;
  assign n44030 = n44029 ^ x332 ^ 1'b0 ;
  assign n44031 = ( x595 & ~n44029 ) | ( x595 & n44030 ) | ( ~n44029 & n44030 ) ;
  assign n44032 = n44031 ^ n44030 ^ 1'b0 ;
  assign n44033 = ~x332 & x596 ;
  assign n44034 = x595 & n42637 ;
  assign n44035 = n44022 & n44034 ;
  assign n44036 = n44035 ^ x596 ^ 1'b0 ;
  assign n44037 = ( ~x596 & n44033 ) | ( ~x596 & n44036 ) | ( n44033 & n44036 ) ;
  assign n44038 = n44020 ^ x332 ^ 1'b0 ;
  assign n44039 = ( x597 & ~n44020 ) | ( x597 & n44038 ) | ( ~n44020 & n44038 ) ;
  assign n44040 = n44039 ^ n44038 ^ 1'b0 ;
  assign n44041 = x740 & x780 ;
  assign n44042 = n5081 & n44041 ;
  assign n44043 = x882 | n7318 ;
  assign n44044 = x947 & ~n44043 ;
  assign n44045 = ~n44042 & n44044 ;
  assign n44046 = ( x598 & n44042 ) | ( x598 & ~n44045 ) | ( n44042 & ~n44045 ) ;
  assign n44047 = ~x332 & x599 ;
  assign n44048 = x596 & n44035 ;
  assign n44049 = n44048 ^ x599 ^ 1'b0 ;
  assign n44050 = ( ~x599 & n44047 ) | ( ~x599 & n44049 ) | ( n44047 & n44049 ) ;
  assign n44051 = ~x332 & x600 ;
  assign n44052 = n44022 ^ x600 ^ 1'b0 ;
  assign n44053 = ( ~x600 & n44051 ) | ( ~x600 & n44052 ) | ( n44051 & n44052 ) ;
  assign n44054 = ~x601 & x806 ;
  assign n44055 = x806 | x989 ;
  assign n44056 = ( x332 & ~n44054 ) | ( x332 & n44055 ) | ( ~n44054 & n44055 ) ;
  assign n44057 = ~x332 & n44056 ;
  assign n44058 = x230 & n15777 ;
  assign n44059 = ~n16559 & n44058 ;
  assign n44060 = x790 ^ x715 ^ 1'b0 ;
  assign n44061 = ( x715 & ~x1160 ) | ( x715 & n44060 ) | ( ~x1160 & n44060 ) ;
  assign n44062 = n44061 ^ n44060 ^ 1'b0 ;
  assign n44063 = ( n17083 & n17273 ) | ( n17083 & ~n44062 ) | ( n17273 & ~n44062 ) ;
  assign n44064 = n44062 | n44063 ;
  assign n44065 = ( n17088 & n44059 ) | ( n17088 & ~n44064 ) | ( n44059 & ~n44064 ) ;
  assign n44066 = ~n17088 & n44065 ;
  assign n44067 = ( ~x230 & x602 ) | ( ~x230 & n44066 ) | ( x602 & n44066 ) ;
  assign n44068 = n44066 ^ x230 ^ 1'b0 ;
  assign n44069 = ( n44066 & n44067 ) | ( n44066 & ~n44068 ) | ( n44067 & ~n44068 ) ;
  assign n44070 = ~x980 & x1038 ;
  assign n44071 = x1060 & n44070 ;
  assign n44072 = x952 & ~x1061 ;
  assign n44073 = n44071 & n44072 ;
  assign n44074 = x832 & n44073 ;
  assign n44075 = x603 | n44074 ;
  assign n44076 = x871 | x872 ;
  assign n44077 = x966 & n44076 ;
  assign n44078 = x832 & ~x1100 ;
  assign n44079 = n44073 & n44078 ;
  assign n44080 = x966 | n44079 ;
  assign n44081 = ~n44077 & n44080 ;
  assign n44082 = ( n44075 & n44077 ) | ( n44075 & ~n44081 ) | ( n44077 & ~n44081 ) ;
  assign n44083 = ~x299 & x983 ;
  assign n44084 = x907 & n44083 ;
  assign n44085 = x604 & ~n44084 ;
  assign n44086 = x823 & ~n15383 ;
  assign n44087 = n44086 ^ x779 ^ 1'b0 ;
  assign n44088 = ( ~x779 & n44085 ) | ( ~x779 & n44087 ) | ( n44085 & n44087 ) ;
  assign n44089 = ~x605 & n44021 ;
  assign n44090 = x332 | n44028 ;
  assign n44091 = n44089 | n44090 ;
  assign n44092 = n44074 ^ x1104 ^ 1'b0 ;
  assign n44093 = ( x606 & x1104 ) | ( x606 & ~n44092 ) | ( x1104 & ~n44092 ) ;
  assign n44094 = n44093 ^ x966 ^ 1'b0 ;
  assign n44095 = ( x837 & n44093 ) | ( x837 & n44094 ) | ( n44093 & n44094 ) ;
  assign n44096 = x607 | n44074 ;
  assign n44097 = ~x1107 & n44074 ;
  assign n44098 = ( x966 & n44096 ) | ( x966 & ~n44097 ) | ( n44096 & ~n44097 ) ;
  assign n44099 = ~x966 & n44098 ;
  assign n44100 = x608 | n44074 ;
  assign n44101 = ~x1116 & n44074 ;
  assign n44102 = ( x966 & n44100 ) | ( x966 & ~n44101 ) | ( n44100 & ~n44101 ) ;
  assign n44103 = ~x966 & n44102 ;
  assign n44104 = x609 | n44074 ;
  assign n44105 = ~x1118 & n44074 ;
  assign n44106 = ( x966 & n44104 ) | ( x966 & ~n44105 ) | ( n44104 & ~n44105 ) ;
  assign n44107 = ~x966 & n44106 ;
  assign n44108 = x610 | n44074 ;
  assign n44109 = ~x1113 & n44074 ;
  assign n44110 = ( x966 & n44108 ) | ( x966 & ~n44109 ) | ( n44108 & ~n44109 ) ;
  assign n44111 = ~x966 & n44110 ;
  assign n44112 = x611 | n44074 ;
  assign n44113 = ~x1114 & n44074 ;
  assign n44114 = ( x966 & n44112 ) | ( x966 & ~n44113 ) | ( n44112 & ~n44113 ) ;
  assign n44115 = ~x966 & n44114 ;
  assign n44116 = x612 | n44074 ;
  assign n44117 = ~x1111 & n44074 ;
  assign n44118 = ( x966 & n44116 ) | ( x966 & ~n44117 ) | ( n44116 & ~n44117 ) ;
  assign n44119 = ~x966 & n44118 ;
  assign n44120 = x613 | n44074 ;
  assign n44121 = ~x1115 & n44074 ;
  assign n44122 = ( x966 & n44120 ) | ( x966 & ~n44121 ) | ( n44120 & ~n44121 ) ;
  assign n44123 = ~x966 & n44122 ;
  assign n44124 = ~x1102 & n44074 ;
  assign n44125 = x614 | n44074 ;
  assign n44126 = ( x966 & ~n44124 ) | ( x966 & n44125 ) | ( ~n44124 & n44125 ) ;
  assign n44127 = ~x966 & n44126 ;
  assign n44128 = n44127 ^ x871 ^ 1'b0 ;
  assign n44129 = ( ~x871 & x966 ) | ( ~x871 & n44128 ) | ( x966 & n44128 ) ;
  assign n44130 = ( x871 & n44127 ) | ( x871 & n44129 ) | ( n44127 & n44129 ) ;
  assign n44131 = x779 & x797 ;
  assign n44132 = n5078 & n44131 ;
  assign n44133 = x907 & ~n44043 ;
  assign n44134 = ( x615 & ~n44132 ) | ( x615 & n44133 ) | ( ~n44132 & n44133 ) ;
  assign n44135 = ~n44132 & n44134 ;
  assign n44136 = ~x1101 & n44074 ;
  assign n44137 = x616 | n44074 ;
  assign n44138 = ( x966 & ~n44136 ) | ( x966 & n44137 ) | ( ~n44136 & n44137 ) ;
  assign n44139 = ~x966 & n44138 ;
  assign n44140 = n44139 ^ x872 ^ 1'b0 ;
  assign n44141 = ( ~x872 & x966 ) | ( ~x872 & n44140 ) | ( x966 & n44140 ) ;
  assign n44142 = ( x872 & n44139 ) | ( x872 & n44141 ) | ( n44139 & n44141 ) ;
  assign n44143 = n44074 ^ x1105 ^ 1'b0 ;
  assign n44144 = ( x617 & x1105 ) | ( x617 & ~n44143 ) | ( x1105 & ~n44143 ) ;
  assign n44145 = n44144 ^ x966 ^ 1'b0 ;
  assign n44146 = ( x850 & n44144 ) | ( x850 & n44145 ) | ( n44144 & n44145 ) ;
  assign n44147 = x618 | n44074 ;
  assign n44148 = ~x1117 & n44074 ;
  assign n44149 = ( x966 & n44147 ) | ( x966 & ~n44148 ) | ( n44147 & ~n44148 ) ;
  assign n44150 = ~x966 & n44149 ;
  assign n44151 = x619 | n44074 ;
  assign n44152 = ~x1122 & n44074 ;
  assign n44153 = ( x966 & n44151 ) | ( x966 & ~n44152 ) | ( n44151 & ~n44152 ) ;
  assign n44154 = ~x966 & n44153 ;
  assign n44155 = x620 | n44074 ;
  assign n44156 = ~x1112 & n44074 ;
  assign n44157 = ( x966 & n44155 ) | ( x966 & ~n44156 ) | ( n44155 & ~n44156 ) ;
  assign n44158 = ~x966 & n44157 ;
  assign n44159 = x621 | n44074 ;
  assign n44160 = ~x1108 & n44074 ;
  assign n44161 = ( x966 & n44159 ) | ( x966 & ~n44160 ) | ( n44159 & ~n44160 ) ;
  assign n44162 = ~x966 & n44161 ;
  assign n44163 = x622 | n44074 ;
  assign n44164 = ~x1109 & n44074 ;
  assign n44165 = ( x966 & n44163 ) | ( x966 & ~n44164 ) | ( n44163 & ~n44164 ) ;
  assign n44166 = ~x966 & n44165 ;
  assign n44167 = x623 | n44074 ;
  assign n44168 = ~x1106 & n44074 ;
  assign n44169 = ( x966 & n44167 ) | ( x966 & ~n44168 ) | ( n44167 & ~n44168 ) ;
  assign n44170 = ~x966 & n44169 ;
  assign n44171 = x947 & n44083 ;
  assign n44172 = x624 & ~n44171 ;
  assign n44173 = x831 & ~n15527 ;
  assign n44174 = n44173 ^ x780 ^ 1'b0 ;
  assign n44175 = ( ~x780 & n44172 ) | ( ~x780 & n44174 ) | ( n44172 & n44174 ) ;
  assign n44176 = x832 & ~x973 ;
  assign n44177 = ~x1054 & x1066 ;
  assign n44178 = ( ~x1088 & n44176 ) | ( ~x1088 & n44177 ) | ( n44176 & n44177 ) ;
  assign n44179 = x1088 & n44178 ;
  assign n44180 = ~x953 & n44179 ;
  assign n44181 = x625 | n44180 ;
  assign n44182 = ~x1116 & n44180 ;
  assign n44183 = ( x962 & n44181 ) | ( x962 & ~n44182 ) | ( n44181 & ~n44182 ) ;
  assign n44184 = ~x962 & n44183 ;
  assign n44185 = x626 | n44074 ;
  assign n44186 = ~x1121 & n44074 ;
  assign n44187 = ( x966 & n44185 ) | ( x966 & ~n44186 ) | ( n44185 & ~n44186 ) ;
  assign n44188 = ~x966 & n44187 ;
  assign n44189 = x627 | n44180 ;
  assign n44190 = ~x1117 & n44180 ;
  assign n44191 = ( x962 & n44189 ) | ( x962 & ~n44190 ) | ( n44189 & ~n44190 ) ;
  assign n44192 = ~x962 & n44191 ;
  assign n44193 = x628 | n44180 ;
  assign n44194 = ~x1119 & n44180 ;
  assign n44195 = ( x962 & n44193 ) | ( x962 & ~n44194 ) | ( n44193 & ~n44194 ) ;
  assign n44196 = ~x962 & n44195 ;
  assign n44197 = x629 | n44074 ;
  assign n44198 = ~x1119 & n44074 ;
  assign n44199 = ( x966 & n44197 ) | ( x966 & ~n44198 ) | ( n44197 & ~n44198 ) ;
  assign n44200 = ~x966 & n44199 ;
  assign n44201 = x630 | n44074 ;
  assign n44202 = ~x1120 & n44074 ;
  assign n44203 = ( x966 & n44201 ) | ( x966 & ~n44202 ) | ( n44201 & ~n44202 ) ;
  assign n44204 = ~x966 & n44203 ;
  assign n44205 = ~x1113 & n44180 ;
  assign n44206 = x962 | n44205 ;
  assign n44207 = n44180 & ~n44206 ;
  assign n44208 = ( x631 & n44206 ) | ( x631 & ~n44207 ) | ( n44206 & ~n44207 ) ;
  assign n44209 = ~x1115 & n44180 ;
  assign n44210 = x962 | n44209 ;
  assign n44211 = n44180 & ~n44210 ;
  assign n44212 = ( x632 & n44210 ) | ( x632 & ~n44211 ) | ( n44210 & ~n44211 ) ;
  assign n44213 = x633 | n44074 ;
  assign n44214 = ~x1110 & n44074 ;
  assign n44215 = ( x966 & n44213 ) | ( x966 & ~n44214 ) | ( n44213 & ~n44214 ) ;
  assign n44216 = ~x966 & n44215 ;
  assign n44217 = x634 | n44180 ;
  assign n44218 = ~x1110 & n44180 ;
  assign n44219 = ( x962 & n44217 ) | ( x962 & ~n44218 ) | ( n44217 & ~n44218 ) ;
  assign n44220 = ~x962 & n44219 ;
  assign n44221 = ~x1112 & n44180 ;
  assign n44222 = x962 | n44221 ;
  assign n44223 = n44180 & ~n44222 ;
  assign n44224 = ( x635 & n44222 ) | ( x635 & ~n44223 ) | ( n44222 & ~n44223 ) ;
  assign n44225 = x636 | n44074 ;
  assign n44226 = ~x1127 & n44074 ;
  assign n44227 = ( x966 & n44225 ) | ( x966 & ~n44226 ) | ( n44225 & ~n44226 ) ;
  assign n44228 = ~x966 & n44227 ;
  assign n44229 = x637 | n44180 ;
  assign n44230 = ~x1105 & n44180 ;
  assign n44231 = ( x962 & n44229 ) | ( x962 & ~n44230 ) | ( n44229 & ~n44230 ) ;
  assign n44232 = ~x962 & n44231 ;
  assign n44233 = x638 | n44180 ;
  assign n44234 = ~x1107 & n44180 ;
  assign n44235 = ( x962 & n44233 ) | ( x962 & ~n44234 ) | ( n44233 & ~n44234 ) ;
  assign n44236 = ~x962 & n44235 ;
  assign n44237 = x639 | n44180 ;
  assign n44238 = ~x1109 & n44180 ;
  assign n44239 = ( x962 & n44237 ) | ( x962 & ~n44238 ) | ( n44237 & ~n44238 ) ;
  assign n44240 = ~x962 & n44239 ;
  assign n44241 = x640 | n44074 ;
  assign n44242 = ~x1128 & n44074 ;
  assign n44243 = ( x966 & n44241 ) | ( x966 & ~n44242 ) | ( n44241 & ~n44242 ) ;
  assign n44244 = ~x966 & n44243 ;
  assign n44245 = x641 | n44180 ;
  assign n44246 = ~x1121 & n44180 ;
  assign n44247 = ( x962 & n44245 ) | ( x962 & ~n44246 ) | ( n44245 & ~n44246 ) ;
  assign n44248 = ~x962 & n44247 ;
  assign n44249 = x642 | n44074 ;
  assign n44250 = ~x1103 & n44074 ;
  assign n44251 = ( x966 & n44249 ) | ( x966 & ~n44250 ) | ( n44249 & ~n44250 ) ;
  assign n44252 = ~x966 & n44251 ;
  assign n44253 = x643 | n44180 ;
  assign n44254 = ~x1104 & n44180 ;
  assign n44255 = ( x962 & n44253 ) | ( x962 & ~n44254 ) | ( n44253 & ~n44254 ) ;
  assign n44256 = ~x962 & n44255 ;
  assign n44257 = x644 | n44074 ;
  assign n44258 = ~x1123 & n44074 ;
  assign n44259 = ( x966 & n44257 ) | ( x966 & ~n44258 ) | ( n44257 & ~n44258 ) ;
  assign n44260 = ~x966 & n44259 ;
  assign n44261 = x645 | n44074 ;
  assign n44262 = ~x1125 & n44074 ;
  assign n44263 = ( x966 & n44261 ) | ( x966 & ~n44262 ) | ( n44261 & ~n44262 ) ;
  assign n44264 = ~x966 & n44263 ;
  assign n44265 = ~x1114 & n44180 ;
  assign n44266 = x962 | n44265 ;
  assign n44267 = n44180 & ~n44266 ;
  assign n44268 = ( x646 & n44266 ) | ( x646 & ~n44267 ) | ( n44266 & ~n44267 ) ;
  assign n44269 = x647 | n44180 ;
  assign n44270 = ~x1120 & n44180 ;
  assign n44271 = ( x962 & n44269 ) | ( x962 & ~n44270 ) | ( n44269 & ~n44270 ) ;
  assign n44272 = ~x962 & n44271 ;
  assign n44273 = x648 | n44180 ;
  assign n44274 = ~x1122 & n44180 ;
  assign n44275 = ( x962 & n44273 ) | ( x962 & ~n44274 ) | ( n44273 & ~n44274 ) ;
  assign n44276 = ~x962 & n44275 ;
  assign n44277 = ~x1126 & n44180 ;
  assign n44278 = x962 | n44277 ;
  assign n44279 = n44180 & ~n44278 ;
  assign n44280 = ( x649 & n44278 ) | ( x649 & ~n44279 ) | ( n44278 & ~n44279 ) ;
  assign n44281 = ~x1127 & n44180 ;
  assign n44282 = x962 | n44281 ;
  assign n44283 = n44180 & ~n44282 ;
  assign n44284 = ( x650 & n44282 ) | ( x650 & ~n44283 ) | ( n44282 & ~n44283 ) ;
  assign n44285 = x651 | n44074 ;
  assign n44286 = ~x1130 & n44074 ;
  assign n44287 = ( x966 & n44285 ) | ( x966 & ~n44286 ) | ( n44285 & ~n44286 ) ;
  assign n44288 = ~x966 & n44287 ;
  assign n44289 = x652 | n44074 ;
  assign n44290 = ~x1131 & n44074 ;
  assign n44291 = ( x966 & n44289 ) | ( x966 & ~n44290 ) | ( n44289 & ~n44290 ) ;
  assign n44292 = ~x966 & n44291 ;
  assign n44293 = x653 | n44074 ;
  assign n44294 = ~x1129 & n44074 ;
  assign n44295 = ( x966 & n44293 ) | ( x966 & ~n44294 ) | ( n44293 & ~n44294 ) ;
  assign n44296 = ~x966 & n44295 ;
  assign n44297 = ~x1130 & n44180 ;
  assign n44298 = x962 | n44297 ;
  assign n44299 = n44180 & ~n44298 ;
  assign n44300 = ( x654 & n44298 ) | ( x654 & ~n44299 ) | ( n44298 & ~n44299 ) ;
  assign n44301 = ~x1124 & n44180 ;
  assign n44302 = x962 | n44301 ;
  assign n44303 = n44180 & ~n44302 ;
  assign n44304 = ( x655 & n44302 ) | ( x655 & ~n44303 ) | ( n44302 & ~n44303 ) ;
  assign n44305 = x656 | n44074 ;
  assign n44306 = ~x1126 & n44074 ;
  assign n44307 = ( x966 & n44305 ) | ( x966 & ~n44306 ) | ( n44305 & ~n44306 ) ;
  assign n44308 = ~x966 & n44307 ;
  assign n44309 = ~x1131 & n44180 ;
  assign n44310 = x962 | n44309 ;
  assign n44311 = n44180 & ~n44310 ;
  assign n44312 = ( x657 & n44310 ) | ( x657 & ~n44311 ) | ( n44310 & ~n44311 ) ;
  assign n44313 = x658 | n44074 ;
  assign n44314 = ~x1124 & n44074 ;
  assign n44315 = ( x966 & n44313 ) | ( x966 & ~n44314 ) | ( n44313 & ~n44314 ) ;
  assign n44316 = ~x966 & n44315 ;
  assign n44317 = x266 & x992 ;
  assign n44318 = ~x280 & n44317 ;
  assign n44319 = ~x269 & n44318 ;
  assign n44320 = ~x281 & n44319 ;
  assign n44321 = x270 | x277 ;
  assign n44322 = x282 | n44321 ;
  assign n44323 = n44320 & ~n44322 ;
  assign n44324 = ~x264 & n44323 ;
  assign n44325 = ~x265 & n44324 ;
  assign n44326 = n44325 ^ x274 ^ 1'b0 ;
  assign n44327 = x660 | n44180 ;
  assign n44328 = ~x1118 & n44180 ;
  assign n44329 = ( x962 & n44327 ) | ( x962 & ~n44328 ) | ( n44327 & ~n44328 ) ;
  assign n44330 = ~x962 & n44329 ;
  assign n44331 = x661 | n44180 ;
  assign n44332 = ~x1101 & n44180 ;
  assign n44333 = ( x962 & n44331 ) | ( x962 & ~n44332 ) | ( n44331 & ~n44332 ) ;
  assign n44334 = ~x962 & n44333 ;
  assign n44335 = x662 | n44180 ;
  assign n44336 = ~x1102 & n44180 ;
  assign n44337 = ( x962 & n44335 ) | ( x962 & ~n44336 ) | ( n44335 & ~n44336 ) ;
  assign n44338 = ~x962 & n44337 ;
  assign n44339 = ~x591 & x592 ;
  assign n44340 = x365 & n44339 ;
  assign n44341 = x334 & x591 ;
  assign n44342 = ~x592 & n44341 ;
  assign n44343 = ( ~x590 & n44340 ) | ( ~x590 & n44342 ) | ( n44340 & n44342 ) ;
  assign n44344 = ~x590 & n44343 ;
  assign n44345 = x590 & ~x592 ;
  assign n44346 = x591 | x592 ;
  assign n44347 = ( x592 & n44345 ) | ( x592 & ~n44346 ) | ( n44345 & ~n44346 ) ;
  assign n44348 = x323 & n44347 ;
  assign n44349 = ( x588 & ~n44344 ) | ( x588 & n44348 ) | ( ~n44344 & n44348 ) ;
  assign n44350 = n44344 | n44349 ;
  assign n44351 = x199 & ~x1065 ;
  assign n44352 = x223 | x224 ;
  assign n44353 = x199 | x257 ;
  assign n44354 = ( n44351 & n44352 ) | ( n44351 & n44353 ) | ( n44352 & n44353 ) ;
  assign n44355 = ~n44351 & n44354 ;
  assign n44356 = x592 | n7276 ;
  assign n44357 = x464 & ~n44356 ;
  assign n44358 = x588 & ~n44357 ;
  assign n44359 = n44352 | n44358 ;
  assign n44360 = ~n44355 & n44359 ;
  assign n44361 = ( n44350 & n44355 ) | ( n44350 & ~n44360 ) | ( n44355 & ~n44360 ) ;
  assign n44362 = x1137 | x1138 ;
  assign n44363 = x815 | x1136 ;
  assign n44364 = ~x633 & x1136 ;
  assign n44365 = ( x1135 & n44363 ) | ( x1135 & ~n44364 ) | ( n44363 & ~n44364 ) ;
  assign n44366 = ~x1135 & n44365 ;
  assign n44367 = ~x634 & x1136 ;
  assign n44368 = ~n44366 & n44367 ;
  assign n44369 = x1135 & x1136 ;
  assign n44370 = ( x784 & x1135 ) | ( x784 & n44369 ) | ( x1135 & n44369 ) ;
  assign n44371 = ( n44366 & ~n44368 ) | ( n44366 & n44370 ) | ( ~n44368 & n44370 ) ;
  assign n44372 = ( x1134 & ~n44362 ) | ( x1134 & n44371 ) | ( ~n44362 & n44371 ) ;
  assign n44373 = ~x1134 & n44372 ;
  assign n44374 = x1135 & ~n44362 ;
  assign n44375 = x1136 & ~n44374 ;
  assign n44376 = ~x766 & n44375 ;
  assign n44377 = ~x700 & x1135 ;
  assign n44378 = x1135 & ~x1136 ;
  assign n44379 = x1134 & ~n44362 ;
  assign n44380 = ~n44378 & n44379 ;
  assign n44381 = x855 | x1136 ;
  assign n44382 = ( n44377 & n44380 ) | ( n44377 & n44381 ) | ( n44380 & n44381 ) ;
  assign n44383 = ~n44377 & n44382 ;
  assign n44384 = n44383 ^ n44376 ^ 1'b0 ;
  assign n44385 = ( n44376 & n44383 ) | ( n44376 & n44384 ) | ( n44383 & n44384 ) ;
  assign n44386 = ( n44373 & ~n44376 ) | ( n44373 & n44385 ) | ( ~n44376 & n44385 ) ;
  assign n44387 = n44361 ^ n10841 ^ 1'b0 ;
  assign n44388 = ( n44361 & n44386 ) | ( n44361 & n44387 ) | ( n44386 & n44387 ) ;
  assign n44389 = ~x727 & x1135 ;
  assign n44390 = x772 | x1135 ;
  assign n44391 = ( x1136 & n44389 ) | ( x1136 & n44390 ) | ( n44389 & n44390 ) ;
  assign n44392 = ~n44389 & n44391 ;
  assign n44393 = x1135 | x1136 ;
  assign n44394 = x872 & ~n44393 ;
  assign n44395 = ( x1134 & n44392 ) | ( x1134 & ~n44394 ) | ( n44392 & ~n44394 ) ;
  assign n44396 = ~n44392 & n44395 ;
  assign n44397 = x614 & ~x1135 ;
  assign n44398 = x662 & x1135 ;
  assign n44399 = ( x1136 & n44397 ) | ( x1136 & ~n44398 ) | ( n44397 & ~n44398 ) ;
  assign n44400 = ~n44397 & n44399 ;
  assign n44401 = ( x811 & x1136 ) | ( x811 & ~n44378 ) | ( x1136 & ~n44378 ) ;
  assign n44402 = x785 & x1135 ;
  assign n44403 = n44401 | n44402 ;
  assign n44404 = n44403 ^ n44400 ^ 1'b0 ;
  assign n44405 = ( n44400 & n44403 ) | ( n44400 & n44404 ) | ( n44403 & n44404 ) ;
  assign n44406 = ( x1134 & ~n44400 ) | ( x1134 & n44405 ) | ( ~n44400 & n44405 ) ;
  assign n44407 = n10841 & ~n44362 ;
  assign n44408 = ( n44396 & n44406 ) | ( n44396 & n44407 ) | ( n44406 & n44407 ) ;
  assign n44409 = ~n44396 & n44408 ;
  assign n44410 = x380 & ~x591 ;
  assign n44411 = x592 & ~n44410 ;
  assign n44412 = ~x590 & x592 ;
  assign n44413 = x588 | n44412 ;
  assign n44414 = ~x590 & x591 ;
  assign n44415 = x404 & n44414 ;
  assign n44416 = ( ~n44411 & n44413 ) | ( ~n44411 & n44415 ) | ( n44413 & n44415 ) ;
  assign n44417 = ~n44411 & n44416 ;
  assign n44418 = n44417 ^ x355 ^ 1'b0 ;
  assign n44419 = ( ~x355 & n44347 ) | ( ~x355 & n44418 ) | ( n44347 & n44418 ) ;
  assign n44420 = ( x355 & n44417 ) | ( x355 & n44419 ) | ( n44417 & n44419 ) ;
  assign n44421 = x199 | x292 ;
  assign n44422 = x199 & ~x1084 ;
  assign n44423 = n44352 & ~n44422 ;
  assign n44424 = n44421 & n44423 ;
  assign n44425 = x429 & ~n44356 ;
  assign n44426 = x588 & ~n44425 ;
  assign n44427 = n44352 | n44426 ;
  assign n44428 = ~n44424 & n44427 ;
  assign n44429 = ( n44420 & n44424 ) | ( n44420 & ~n44428 ) | ( n44424 & ~n44428 ) ;
  assign n44430 = ( ~n10841 & n44409 ) | ( ~n10841 & n44429 ) | ( n44409 & n44429 ) ;
  assign n44431 = n44409 ^ n10841 ^ 1'b0 ;
  assign n44432 = ( n44409 & n44430 ) | ( n44409 & ~n44431 ) | ( n44430 & ~n44431 ) ;
  assign n44433 = x665 | n44180 ;
  assign n44434 = ~x1108 & n44180 ;
  assign n44435 = ( x962 & n44433 ) | ( x962 & ~n44434 ) | ( n44433 & ~n44434 ) ;
  assign n44436 = ~x962 & n44435 ;
  assign n44437 = x337 & ~x591 ;
  assign n44438 = x592 & ~n44437 ;
  assign n44439 = x456 & n44414 ;
  assign n44440 = ( n44413 & ~n44438 ) | ( n44413 & n44439 ) | ( ~n44438 & n44439 ) ;
  assign n44441 = ~n44438 & n44440 ;
  assign n44442 = n44441 ^ x441 ^ 1'b0 ;
  assign n44443 = ( ~x441 & n44347 ) | ( ~x441 & n44442 ) | ( n44347 & n44442 ) ;
  assign n44444 = ( x441 & n44441 ) | ( x441 & n44443 ) | ( n44441 & n44443 ) ;
  assign n44445 = x443 & ~n44356 ;
  assign n44446 = x588 & ~n44445 ;
  assign n44447 = ( n44352 & n44444 ) | ( n44352 & ~n44446 ) | ( n44444 & ~n44446 ) ;
  assign n44448 = ~n44352 & n44447 ;
  assign n44449 = x199 | x297 ;
  assign n44450 = x199 & ~x1044 ;
  assign n44451 = n44352 & ~n44450 ;
  assign n44452 = n44449 & n44451 ;
  assign n44453 = ( ~n10841 & n44448 ) | ( ~n10841 & n44452 ) | ( n44448 & n44452 ) ;
  assign n44454 = ~n10841 & n44453 ;
  assign n44455 = x873 | x1136 ;
  assign n44456 = ~x691 & x1135 ;
  assign n44457 = n44455 & ~n44456 ;
  assign n44458 = ~x764 & n44375 ;
  assign n44459 = n44380 & ~n44458 ;
  assign n44460 = n44457 & n44459 ;
  assign n44461 = x1134 | n44362 ;
  assign n44462 = ~x638 & x1135 ;
  assign n44463 = x607 | x1135 ;
  assign n44464 = ( x1136 & n44462 ) | ( x1136 & n44463 ) | ( n44462 & n44463 ) ;
  assign n44465 = ~n44462 & n44464 ;
  assign n44466 = ~x790 & x1135 ;
  assign n44467 = x1136 | n44466 ;
  assign n44468 = x799 & ~x1135 ;
  assign n44469 = ( ~n44465 & n44467 ) | ( ~n44465 & n44468 ) | ( n44467 & n44468 ) ;
  assign n44470 = ~n44465 & n44469 ;
  assign n44471 = ( ~n44460 & n44461 ) | ( ~n44460 & n44470 ) | ( n44461 & n44470 ) ;
  assign n44472 = ~n44460 & n44471 ;
  assign n44473 = ~n44454 & n44472 ;
  assign n44474 = ( n10841 & n44454 ) | ( n10841 & ~n44473 ) | ( n44454 & ~n44473 ) ;
  assign n44475 = x792 & ~x1136 ;
  assign n44476 = x681 & x1136 ;
  assign n44477 = ( x1135 & n44475 ) | ( x1135 & ~n44476 ) | ( n44475 & ~n44476 ) ;
  assign n44478 = ~n44475 & n44477 ;
  assign n44479 = x809 | x1136 ;
  assign n44480 = x642 & x1136 ;
  assign n44481 = ( x1135 & n44479 ) | ( x1135 & ~n44480 ) | ( n44479 & ~n44480 ) ;
  assign n44482 = ~x1135 & n44481 ;
  assign n44483 = ( ~x1134 & n44478 ) | ( ~x1134 & n44482 ) | ( n44478 & n44482 ) ;
  assign n44484 = ~x1134 & n44483 ;
  assign n44485 = ~x699 & x1135 ;
  assign n44486 = x763 | x1135 ;
  assign n44487 = ( x1136 & n44485 ) | ( x1136 & n44486 ) | ( n44485 & n44486 ) ;
  assign n44488 = ~n44485 & n44487 ;
  assign n44489 = x871 & ~n44393 ;
  assign n44490 = ( x1134 & n44488 ) | ( x1134 & ~n44489 ) | ( n44488 & ~n44489 ) ;
  assign n44491 = ~n44488 & n44490 ;
  assign n44492 = ( n44407 & n44484 ) | ( n44407 & ~n44491 ) | ( n44484 & ~n44491 ) ;
  assign n44493 = ~n44484 & n44492 ;
  assign n44494 = x338 & ~x591 ;
  assign n44495 = x592 & ~n44494 ;
  assign n44496 = x319 & n44414 ;
  assign n44497 = ( n44413 & ~n44495 ) | ( n44413 & n44496 ) | ( ~n44495 & n44496 ) ;
  assign n44498 = ~n44495 & n44497 ;
  assign n44499 = n44498 ^ x458 ^ 1'b0 ;
  assign n44500 = ( ~x458 & n44347 ) | ( ~x458 & n44499 ) | ( n44347 & n44499 ) ;
  assign n44501 = ( x458 & n44498 ) | ( x458 & n44500 ) | ( n44498 & n44500 ) ;
  assign n44502 = x199 | x294 ;
  assign n44503 = x199 & ~x1072 ;
  assign n44504 = n44352 & ~n44503 ;
  assign n44505 = n44502 & n44504 ;
  assign n44506 = x444 & ~n44356 ;
  assign n44507 = x588 & ~n44506 ;
  assign n44508 = n44352 | n44507 ;
  assign n44509 = ~n44505 & n44508 ;
  assign n44510 = ( n44501 & n44505 ) | ( n44501 & ~n44509 ) | ( n44505 & ~n44509 ) ;
  assign n44511 = ( ~n10841 & n44493 ) | ( ~n10841 & n44510 ) | ( n44493 & n44510 ) ;
  assign n44512 = n44493 ^ n10841 ^ 1'b0 ;
  assign n44513 = ( n44493 & n44511 ) | ( n44493 & ~n44512 ) | ( n44511 & ~n44512 ) ;
  assign n44514 = ~x680 & x1135 ;
  assign n44515 = x603 | x1135 ;
  assign n44516 = ( x1136 & n44514 ) | ( x1136 & n44515 ) | ( n44514 & n44515 ) ;
  assign n44517 = ~n44514 & n44516 ;
  assign n44518 = x981 | x1135 ;
  assign n44519 = ~x778 & x1135 ;
  assign n44520 = ( x1136 & n44518 ) | ( x1136 & ~n44519 ) | ( n44518 & ~n44519 ) ;
  assign n44521 = ~x1136 & n44520 ;
  assign n44522 = ( ~n44461 & n44517 ) | ( ~n44461 & n44521 ) | ( n44517 & n44521 ) ;
  assign n44523 = ~n44461 & n44522 ;
  assign n44524 = ~x759 & n44375 ;
  assign n44525 = ~x696 & x1135 ;
  assign n44526 = x837 | x1136 ;
  assign n44527 = ( n44380 & n44525 ) | ( n44380 & n44526 ) | ( n44525 & n44526 ) ;
  assign n44528 = ~n44525 & n44527 ;
  assign n44529 = n44528 ^ n44524 ^ 1'b0 ;
  assign n44530 = ( n44524 & n44528 ) | ( n44524 & n44529 ) | ( n44528 & n44529 ) ;
  assign n44531 = ( n44523 & ~n44524 ) | ( n44523 & n44530 ) | ( ~n44524 & n44530 ) ;
  assign n44532 = x363 & ~x591 ;
  assign n44533 = x592 & ~n44532 ;
  assign n44534 = x390 & n44414 ;
  assign n44535 = ( n44413 & ~n44533 ) | ( n44413 & n44534 ) | ( ~n44533 & n44534 ) ;
  assign n44536 = ~n44533 & n44535 ;
  assign n44537 = n44536 ^ x342 ^ 1'b0 ;
  assign n44538 = ( ~x342 & n44347 ) | ( ~x342 & n44537 ) | ( n44347 & n44537 ) ;
  assign n44539 = ( x342 & n44536 ) | ( x342 & n44538 ) | ( n44536 & n44538 ) ;
  assign n44540 = x199 | x291 ;
  assign n44541 = x199 & ~x1049 ;
  assign n44542 = n44352 & ~n44541 ;
  assign n44543 = n44540 & n44542 ;
  assign n44544 = x414 & ~n44356 ;
  assign n44545 = x588 & ~n44544 ;
  assign n44546 = n44352 | n44545 ;
  assign n44547 = ~n44543 & n44546 ;
  assign n44548 = ( n44539 & n44543 ) | ( n44539 & ~n44547 ) | ( n44543 & ~n44547 ) ;
  assign n44549 = n44531 ^ n10841 ^ 1'b0 ;
  assign n44550 = ( n44531 & n44548 ) | ( n44531 & ~n44549 ) | ( n44548 & ~n44549 ) ;
  assign n44551 = ~x1125 & n44180 ;
  assign n44552 = x962 | n44551 ;
  assign n44553 = n44180 & ~n44552 ;
  assign n44554 = ( x669 & n44552 ) | ( x669 & ~n44553 ) | ( n44552 & ~n44553 ) ;
  assign n44555 = x364 & n44339 ;
  assign n44556 = x391 & x591 ;
  assign n44557 = ~x592 & n44556 ;
  assign n44558 = ( ~x590 & n44555 ) | ( ~x590 & n44557 ) | ( n44555 & n44557 ) ;
  assign n44559 = ~x590 & n44558 ;
  assign n44560 = x343 & n44347 ;
  assign n44561 = ( x588 & ~n44559 ) | ( x588 & n44560 ) | ( ~n44559 & n44560 ) ;
  assign n44562 = n44559 | n44561 ;
  assign n44563 = x199 | x258 ;
  assign n44564 = x199 & ~x1062 ;
  assign n44565 = n44352 & ~n44564 ;
  assign n44566 = n44563 & n44565 ;
  assign n44567 = x415 & ~n44356 ;
  assign n44568 = x588 & ~n44567 ;
  assign n44569 = n44352 | n44568 ;
  assign n44570 = ~n44566 & n44569 ;
  assign n44571 = ( n44562 & n44566 ) | ( n44562 & ~n44570 ) | ( n44566 & ~n44570 ) ;
  assign n44572 = x1136 & ~n44362 ;
  assign n44573 = x852 | x1136 ;
  assign n44574 = x723 & x1135 ;
  assign n44575 = n44573 & ~n44574 ;
  assign n44576 = x745 & n44375 ;
  assign n44577 = n44380 & ~n44576 ;
  assign n44578 = n44575 & n44577 ;
  assign n44579 = x695 & x1135 ;
  assign n44580 = x1134 | n44579 ;
  assign n44581 = ( x612 & x1135 ) | ( x612 & ~n44580 ) | ( x1135 & ~n44580 ) ;
  assign n44582 = ~n44580 & n44581 ;
  assign n44583 = n44578 ^ n44572 ^ 1'b0 ;
  assign n44584 = ( ~n44572 & n44582 ) | ( ~n44572 & n44583 ) | ( n44582 & n44583 ) ;
  assign n44585 = ( n44572 & n44578 ) | ( n44572 & n44584 ) | ( n44578 & n44584 ) ;
  assign n44586 = n44571 ^ n10841 ^ 1'b0 ;
  assign n44587 = ( n44571 & n44585 ) | ( n44571 & n44586 ) | ( n44585 & n44586 ) ;
  assign n44588 = x447 & n44339 ;
  assign n44589 = x333 & x591 ;
  assign n44590 = ~x592 & n44589 ;
  assign n44591 = ( ~x590 & n44588 ) | ( ~x590 & n44590 ) | ( n44588 & n44590 ) ;
  assign n44592 = ~x590 & n44591 ;
  assign n44593 = x327 & n44347 ;
  assign n44594 = ( x588 & ~n44592 ) | ( x588 & n44593 ) | ( ~n44592 & n44593 ) ;
  assign n44595 = n44592 | n44594 ;
  assign n44596 = x199 | x261 ;
  assign n44597 = x199 & ~x1040 ;
  assign n44598 = n44352 & ~n44597 ;
  assign n44599 = n44596 & n44598 ;
  assign n44600 = x453 & ~n44356 ;
  assign n44601 = x588 & ~n44600 ;
  assign n44602 = n44352 | n44601 ;
  assign n44603 = ~n44599 & n44602 ;
  assign n44604 = ( n44595 & n44599 ) | ( n44595 & ~n44603 ) | ( n44599 & ~n44603 ) ;
  assign n44605 = x865 | x1136 ;
  assign n44606 = x724 & x1135 ;
  assign n44607 = n44605 & ~n44606 ;
  assign n44608 = x741 & n44375 ;
  assign n44609 = n44380 & ~n44608 ;
  assign n44610 = n44607 & n44609 ;
  assign n44611 = x646 & x1135 ;
  assign n44612 = x1134 | n44611 ;
  assign n44613 = ( x611 & x1135 ) | ( x611 & ~n44612 ) | ( x1135 & ~n44612 ) ;
  assign n44614 = ~n44612 & n44613 ;
  assign n44615 = n44610 ^ n44572 ^ 1'b0 ;
  assign n44616 = ( ~n44572 & n44614 ) | ( ~n44572 & n44615 ) | ( n44614 & n44615 ) ;
  assign n44617 = ( n44572 & n44610 ) | ( n44572 & n44616 ) | ( n44610 & n44616 ) ;
  assign n44618 = n44604 ^ n10841 ^ 1'b0 ;
  assign n44619 = ( n44604 & n44617 ) | ( n44604 & n44618 ) | ( n44617 & n44618 ) ;
  assign n44620 = ~x661 & x1135 ;
  assign n44621 = x616 | x1135 ;
  assign n44622 = ( x1136 & n44620 ) | ( x1136 & n44621 ) | ( n44620 & n44621 ) ;
  assign n44623 = ~n44620 & n44622 ;
  assign n44624 = x808 | x1135 ;
  assign n44625 = ~x781 & x1135 ;
  assign n44626 = ( x1136 & n44624 ) | ( x1136 & ~n44625 ) | ( n44624 & ~n44625 ) ;
  assign n44627 = ~x1136 & n44626 ;
  assign n44628 = ( ~n44461 & n44623 ) | ( ~n44461 & n44627 ) | ( n44623 & n44627 ) ;
  assign n44629 = ~n44461 & n44628 ;
  assign n44630 = ~x758 & n44375 ;
  assign n44631 = ~x736 & x1135 ;
  assign n44632 = x850 | x1136 ;
  assign n44633 = ( n44380 & n44631 ) | ( n44380 & n44632 ) | ( n44631 & n44632 ) ;
  assign n44634 = ~n44631 & n44633 ;
  assign n44635 = n44634 ^ n44630 ^ 1'b0 ;
  assign n44636 = ( n44630 & n44634 ) | ( n44630 & n44635 ) | ( n44634 & n44635 ) ;
  assign n44637 = ( n44629 & ~n44630 ) | ( n44629 & n44636 ) | ( ~n44630 & n44636 ) ;
  assign n44638 = x372 & ~x591 ;
  assign n44639 = x592 & ~n44638 ;
  assign n44640 = x397 & n44414 ;
  assign n44641 = ( n44413 & ~n44639 ) | ( n44413 & n44640 ) | ( ~n44639 & n44640 ) ;
  assign n44642 = ~n44639 & n44641 ;
  assign n44643 = n44642 ^ x320 ^ 1'b0 ;
  assign n44644 = ( ~x320 & n44347 ) | ( ~x320 & n44643 ) | ( n44347 & n44643 ) ;
  assign n44645 = ( x320 & n44642 ) | ( x320 & n44644 ) | ( n44642 & n44644 ) ;
  assign n44646 = x199 | x290 ;
  assign n44647 = x199 & ~x1048 ;
  assign n44648 = n44352 & ~n44647 ;
  assign n44649 = n44646 & n44648 ;
  assign n44650 = x422 & ~n44356 ;
  assign n44651 = x588 & ~n44650 ;
  assign n44652 = n44352 | n44651 ;
  assign n44653 = ~n44649 & n44652 ;
  assign n44654 = ( n44645 & n44649 ) | ( n44645 & ~n44653 ) | ( n44649 & ~n44653 ) ;
  assign n44655 = n44637 ^ n10841 ^ 1'b0 ;
  assign n44656 = ( n44637 & n44654 ) | ( n44637 & ~n44655 ) | ( n44654 & ~n44655 ) ;
  assign n44657 = x387 & ~x591 ;
  assign n44658 = x592 & ~n44657 ;
  assign n44659 = x411 & n44414 ;
  assign n44660 = ( n44413 & ~n44658 ) | ( n44413 & n44659 ) | ( ~n44658 & n44659 ) ;
  assign n44661 = ~n44658 & n44660 ;
  assign n44662 = n44661 ^ x452 ^ 1'b0 ;
  assign n44663 = ( ~x452 & n44347 ) | ( ~x452 & n44662 ) | ( n44347 & n44662 ) ;
  assign n44664 = ( x452 & n44661 ) | ( x452 & n44663 ) | ( n44661 & n44663 ) ;
  assign n44665 = x435 & ~n44356 ;
  assign n44666 = x588 & ~n44665 ;
  assign n44667 = ( n44352 & n44664 ) | ( n44352 & ~n44666 ) | ( n44664 & ~n44666 ) ;
  assign n44668 = ~n44352 & n44667 ;
  assign n44669 = x199 | x295 ;
  assign n44670 = x199 & ~x1053 ;
  assign n44671 = n44352 & ~n44670 ;
  assign n44672 = n44669 & n44671 ;
  assign n44673 = ( ~n10841 & n44668 ) | ( ~n10841 & n44672 ) | ( n44668 & n44672 ) ;
  assign n44674 = ~n10841 & n44673 ;
  assign n44675 = x866 | x1136 ;
  assign n44676 = ~x706 & x1135 ;
  assign n44677 = n44675 & ~n44676 ;
  assign n44678 = ~x749 & n44375 ;
  assign n44679 = n44380 & ~n44678 ;
  assign n44680 = n44677 & n44679 ;
  assign n44681 = ~x637 & x1135 ;
  assign n44682 = x617 | x1135 ;
  assign n44683 = ( x1136 & n44681 ) | ( x1136 & n44682 ) | ( n44681 & n44682 ) ;
  assign n44684 = ~n44681 & n44683 ;
  assign n44685 = ~x788 & x1135 ;
  assign n44686 = x1136 | n44685 ;
  assign n44687 = x814 & ~x1135 ;
  assign n44688 = ( ~n44684 & n44686 ) | ( ~n44684 & n44687 ) | ( n44686 & n44687 ) ;
  assign n44689 = ~n44684 & n44688 ;
  assign n44690 = ( n44461 & ~n44680 ) | ( n44461 & n44689 ) | ( ~n44680 & n44689 ) ;
  assign n44691 = ~n44680 & n44690 ;
  assign n44692 = ~n44674 & n44691 ;
  assign n44693 = ( n10841 & n44674 ) | ( n10841 & ~n44692 ) | ( n44674 & ~n44692 ) ;
  assign n44694 = ~x735 & x1135 ;
  assign n44695 = x743 | x1135 ;
  assign n44696 = ( x1136 & n44694 ) | ( x1136 & n44695 ) | ( n44694 & n44695 ) ;
  assign n44697 = ~n44694 & n44696 ;
  assign n44698 = x859 & ~n44393 ;
  assign n44699 = ( x1134 & n44697 ) | ( x1134 & ~n44698 ) | ( n44697 & ~n44698 ) ;
  assign n44700 = ~n44697 & n44699 ;
  assign n44701 = x622 & ~x1135 ;
  assign n44702 = x639 & x1135 ;
  assign n44703 = ( x1136 & n44701 ) | ( x1136 & ~n44702 ) | ( n44701 & ~n44702 ) ;
  assign n44704 = ~n44701 & n44703 ;
  assign n44705 = x783 & x1135 ;
  assign n44706 = ( x804 & x1136 ) | ( x804 & ~n44378 ) | ( x1136 & ~n44378 ) ;
  assign n44707 = n44705 | n44706 ;
  assign n44708 = n44707 ^ n44704 ^ 1'b0 ;
  assign n44709 = ( n44704 & n44707 ) | ( n44704 & n44708 ) | ( n44707 & n44708 ) ;
  assign n44710 = ( x1134 & ~n44704 ) | ( x1134 & n44709 ) | ( ~n44704 & n44709 ) ;
  assign n44711 = ( n44407 & n44700 ) | ( n44407 & n44710 ) | ( n44700 & n44710 ) ;
  assign n44712 = ~n44700 & n44711 ;
  assign n44713 = x463 & x591 ;
  assign n44714 = ~x592 & n44713 ;
  assign n44715 = x336 & n44339 ;
  assign n44716 = ( ~x590 & n44714 ) | ( ~x590 & n44715 ) | ( n44714 & n44715 ) ;
  assign n44717 = ~x590 & n44716 ;
  assign n44718 = x362 & n44347 ;
  assign n44719 = ( x588 & ~n44717 ) | ( x588 & n44718 ) | ( ~n44717 & n44718 ) ;
  assign n44720 = n44717 | n44719 ;
  assign n44721 = x199 | x256 ;
  assign n44722 = x199 & ~x1070 ;
  assign n44723 = n44352 & ~n44722 ;
  assign n44724 = n44721 & n44723 ;
  assign n44725 = x437 & ~n44356 ;
  assign n44726 = x588 & ~n44725 ;
  assign n44727 = n44352 | n44726 ;
  assign n44728 = ~n44724 & n44727 ;
  assign n44729 = ( n44720 & n44724 ) | ( n44720 & ~n44728 ) | ( n44724 & ~n44728 ) ;
  assign n44730 = ( ~n10841 & n44712 ) | ( ~n10841 & n44729 ) | ( n44712 & n44729 ) ;
  assign n44731 = n44712 ^ n10841 ^ 1'b0 ;
  assign n44732 = ( n44712 & n44730 ) | ( n44712 & ~n44731 ) | ( n44730 & ~n44731 ) ;
  assign n44733 = x388 & ~x591 ;
  assign n44734 = x592 & ~n44733 ;
  assign n44735 = x412 & n44414 ;
  assign n44736 = ( n44413 & ~n44734 ) | ( n44413 & n44735 ) | ( ~n44734 & n44735 ) ;
  assign n44737 = ~n44734 & n44736 ;
  assign n44738 = n44737 ^ x455 ^ 1'b0 ;
  assign n44739 = ( ~x455 & n44347 ) | ( ~x455 & n44738 ) | ( n44347 & n44738 ) ;
  assign n44740 = ( x455 & n44737 ) | ( x455 & n44739 ) | ( n44737 & n44739 ) ;
  assign n44741 = x436 & ~n44356 ;
  assign n44742 = x588 & ~n44741 ;
  assign n44743 = ( n44352 & n44740 ) | ( n44352 & ~n44742 ) | ( n44740 & ~n44742 ) ;
  assign n44744 = ~n44352 & n44743 ;
  assign n44745 = x199 | x296 ;
  assign n44746 = x199 & ~x1037 ;
  assign n44747 = n44352 & ~n44746 ;
  assign n44748 = n44745 & n44747 ;
  assign n44749 = ( ~n10841 & n44744 ) | ( ~n10841 & n44748 ) | ( n44744 & n44748 ) ;
  assign n44750 = ~n10841 & n44749 ;
  assign n44751 = ~x623 & n44375 ;
  assign n44752 = ~x710 & x1135 ;
  assign n44753 = x1136 & ~n44752 ;
  assign n44754 = x789 & n44378 ;
  assign n44755 = x803 | x1135 ;
  assign n44756 = ( n44753 & ~n44754 ) | ( n44753 & n44755 ) | ( ~n44754 & n44755 ) ;
  assign n44757 = ~n44753 & n44756 ;
  assign n44758 = ( n44461 & ~n44751 ) | ( n44461 & n44757 ) | ( ~n44751 & n44757 ) ;
  assign n44759 = n44751 | n44758 ;
  assign n44760 = ~x730 & x1135 ;
  assign n44761 = x748 | x1135 ;
  assign n44762 = ( x1136 & n44760 ) | ( x1136 & n44761 ) | ( n44760 & n44761 ) ;
  assign n44763 = ~n44760 & n44762 ;
  assign n44764 = n44393 & ~n44763 ;
  assign n44765 = ( x876 & n44763 ) | ( x876 & ~n44764 ) | ( n44763 & ~n44764 ) ;
  assign n44766 = ( n44379 & ~n44759 ) | ( n44379 & n44765 ) | ( ~n44759 & n44765 ) ;
  assign n44767 = n44766 ^ n44759 ^ 1'b0 ;
  assign n44768 = ( n44759 & ~n44766 ) | ( n44759 & n44767 ) | ( ~n44766 & n44767 ) ;
  assign n44769 = ~n44750 & n44768 ;
  assign n44770 = ( n10841 & n44750 ) | ( n10841 & ~n44769 ) | ( n44750 & ~n44769 ) ;
  assign n44771 = x386 & ~x591 ;
  assign n44772 = x592 & ~n44771 ;
  assign n44773 = x410 & n44414 ;
  assign n44774 = ( n44413 & ~n44772 ) | ( n44413 & n44773 ) | ( ~n44772 & n44773 ) ;
  assign n44775 = ~n44772 & n44774 ;
  assign n44776 = n44775 ^ x361 ^ 1'b0 ;
  assign n44777 = ( ~x361 & n44347 ) | ( ~x361 & n44776 ) | ( n44347 & n44776 ) ;
  assign n44778 = ( x361 & n44775 ) | ( x361 & n44777 ) | ( n44775 & n44777 ) ;
  assign n44779 = x434 & ~n44356 ;
  assign n44780 = x588 & ~n44779 ;
  assign n44781 = ( n44352 & n44778 ) | ( n44352 & ~n44780 ) | ( n44778 & ~n44780 ) ;
  assign n44782 = ~n44352 & n44781 ;
  assign n44783 = x199 | x293 ;
  assign n44784 = x199 & ~x1059 ;
  assign n44785 = n44352 & ~n44784 ;
  assign n44786 = n44783 & n44785 ;
  assign n44787 = ( ~n10841 & n44782 ) | ( ~n10841 & n44786 ) | ( n44782 & n44786 ) ;
  assign n44788 = ~n10841 & n44787 ;
  assign n44789 = x881 | x1136 ;
  assign n44790 = ~x729 & x1135 ;
  assign n44791 = n44789 & ~n44790 ;
  assign n44792 = ~x746 & n44375 ;
  assign n44793 = n44380 & ~n44792 ;
  assign n44794 = n44791 & n44793 ;
  assign n44795 = ~x643 & x1135 ;
  assign n44796 = x606 | x1135 ;
  assign n44797 = ( x1136 & n44795 ) | ( x1136 & n44796 ) | ( n44795 & n44796 ) ;
  assign n44798 = ~n44795 & n44797 ;
  assign n44799 = ~x787 & x1135 ;
  assign n44800 = x1136 | n44799 ;
  assign n44801 = x812 & ~x1135 ;
  assign n44802 = ( ~n44798 & n44800 ) | ( ~n44798 & n44801 ) | ( n44800 & n44801 ) ;
  assign n44803 = ~n44798 & n44802 ;
  assign n44804 = ( n44461 & ~n44794 ) | ( n44461 & n44803 ) | ( ~n44794 & n44803 ) ;
  assign n44805 = ~n44794 & n44804 ;
  assign n44806 = ~n44788 & n44805 ;
  assign n44807 = ( n10841 & n44788 ) | ( n10841 & ~n44806 ) | ( n44788 & ~n44806 ) ;
  assign n44808 = x366 & n44339 ;
  assign n44809 = x335 & x591 ;
  assign n44810 = ~x592 & n44809 ;
  assign n44811 = ( ~x590 & n44808 ) | ( ~x590 & n44810 ) | ( n44808 & n44810 ) ;
  assign n44812 = ~x590 & n44811 ;
  assign n44813 = x344 & n44347 ;
  assign n44814 = ( x588 & ~n44812 ) | ( x588 & n44813 ) | ( ~n44812 & n44813 ) ;
  assign n44815 = n44812 | n44814 ;
  assign n44816 = x199 | x259 ;
  assign n44817 = x199 & ~x1069 ;
  assign n44818 = n44352 & ~n44817 ;
  assign n44819 = n44816 & n44818 ;
  assign n44820 = x416 & ~n44356 ;
  assign n44821 = x588 & ~n44820 ;
  assign n44822 = n44352 | n44821 ;
  assign n44823 = ~n44819 & n44822 ;
  assign n44824 = ( n44815 & n44819 ) | ( n44815 & ~n44823 ) | ( n44819 & ~n44823 ) ;
  assign n44825 = x870 | x1136 ;
  assign n44826 = x704 & x1135 ;
  assign n44827 = n44825 & ~n44826 ;
  assign n44828 = x742 & n44375 ;
  assign n44829 = n44380 & ~n44828 ;
  assign n44830 = n44827 & n44829 ;
  assign n44831 = x635 & x1135 ;
  assign n44832 = x1134 | n44831 ;
  assign n44833 = ( x620 & x1135 ) | ( x620 & ~n44832 ) | ( x1135 & ~n44832 ) ;
  assign n44834 = ~n44832 & n44833 ;
  assign n44835 = n44830 ^ n44572 ^ 1'b0 ;
  assign n44836 = ( ~n44572 & n44834 ) | ( ~n44572 & n44835 ) | ( n44834 & n44835 ) ;
  assign n44837 = ( n44572 & n44830 ) | ( n44572 & n44836 ) | ( n44830 & n44836 ) ;
  assign n44838 = n44824 ^ n10841 ^ 1'b0 ;
  assign n44839 = ( n44824 & n44837 ) | ( n44824 & n44838 ) | ( n44837 & n44838 ) ;
  assign n44840 = x368 & n44339 ;
  assign n44841 = x393 & x591 ;
  assign n44842 = ~x592 & n44841 ;
  assign n44843 = ( ~x590 & n44840 ) | ( ~x590 & n44842 ) | ( n44840 & n44842 ) ;
  assign n44844 = ~x590 & n44843 ;
  assign n44845 = x346 & n44347 ;
  assign n44846 = ( x588 & ~n44844 ) | ( x588 & n44845 ) | ( ~n44844 & n44845 ) ;
  assign n44847 = n44844 | n44846 ;
  assign n44848 = x199 | x260 ;
  assign n44849 = x199 & ~x1067 ;
  assign n44850 = n44352 & ~n44849 ;
  assign n44851 = n44848 & n44850 ;
  assign n44852 = x418 & ~n44356 ;
  assign n44853 = x588 & ~n44852 ;
  assign n44854 = n44352 | n44853 ;
  assign n44855 = ~n44851 & n44854 ;
  assign n44856 = ( n44847 & n44851 ) | ( n44847 & ~n44855 ) | ( n44851 & ~n44855 ) ;
  assign n44857 = x856 | x1136 ;
  assign n44858 = x688 & x1135 ;
  assign n44859 = n44857 & ~n44858 ;
  assign n44860 = x760 & n44375 ;
  assign n44861 = n44380 & ~n44860 ;
  assign n44862 = n44859 & n44861 ;
  assign n44863 = x632 & x1135 ;
  assign n44864 = x1134 | n44863 ;
  assign n44865 = ( x613 & x1135 ) | ( x613 & ~n44864 ) | ( x1135 & ~n44864 ) ;
  assign n44866 = ~n44864 & n44865 ;
  assign n44867 = n44862 ^ n44572 ^ 1'b0 ;
  assign n44868 = ( ~n44572 & n44866 ) | ( ~n44572 & n44867 ) | ( n44866 & n44867 ) ;
  assign n44869 = ( n44572 & n44862 ) | ( n44572 & n44868 ) | ( n44862 & n44868 ) ;
  assign n44870 = n44856 ^ n10841 ^ 1'b0 ;
  assign n44871 = ( n44856 & n44869 ) | ( n44856 & n44870 ) | ( n44869 & n44870 ) ;
  assign n44872 = x389 & n44339 ;
  assign n44873 = x413 & x591 ;
  assign n44874 = ~x592 & n44873 ;
  assign n44875 = ( ~x590 & n44872 ) | ( ~x590 & n44874 ) | ( n44872 & n44874 ) ;
  assign n44876 = ~x590 & n44875 ;
  assign n44877 = x450 & n44347 ;
  assign n44878 = ( x588 & ~n44876 ) | ( x588 & n44877 ) | ( ~n44876 & n44877 ) ;
  assign n44879 = n44876 | n44878 ;
  assign n44880 = x199 | x255 ;
  assign n44881 = x199 & ~x1036 ;
  assign n44882 = n44352 & ~n44881 ;
  assign n44883 = n44880 & n44882 ;
  assign n44884 = x438 & ~n44356 ;
  assign n44885 = x588 & ~n44884 ;
  assign n44886 = n44352 | n44885 ;
  assign n44887 = ~n44883 & n44886 ;
  assign n44888 = ( n44879 & n44883 ) | ( n44879 & ~n44887 ) | ( n44883 & ~n44887 ) ;
  assign n44889 = ~x665 & x1136 ;
  assign n44890 = x791 | x1136 ;
  assign n44891 = ( x1135 & n44889 ) | ( x1135 & n44890 ) | ( n44889 & n44890 ) ;
  assign n44892 = ~n44889 & n44891 ;
  assign n44893 = x810 | x1136 ;
  assign n44894 = ~x621 & x1136 ;
  assign n44895 = ( x1135 & n44893 ) | ( x1135 & ~n44894 ) | ( n44893 & ~n44894 ) ;
  assign n44896 = ~x1135 & n44895 ;
  assign n44897 = ( ~n44461 & n44892 ) | ( ~n44461 & n44896 ) | ( n44892 & n44896 ) ;
  assign n44898 = ~n44461 & n44897 ;
  assign n44899 = ~x739 & n44375 ;
  assign n44900 = ~x690 & x1135 ;
  assign n44901 = x874 | x1136 ;
  assign n44902 = ( n44380 & n44900 ) | ( n44380 & n44901 ) | ( n44900 & n44901 ) ;
  assign n44903 = ~n44900 & n44902 ;
  assign n44904 = n44903 ^ n44899 ^ 1'b0 ;
  assign n44905 = ( n44899 & n44903 ) | ( n44899 & n44904 ) | ( n44903 & n44904 ) ;
  assign n44906 = ( n44898 & ~n44899 ) | ( n44898 & n44905 ) | ( ~n44899 & n44905 ) ;
  assign n44907 = n44888 ^ n10841 ^ 1'b0 ;
  assign n44908 = ( n44888 & n44906 ) | ( n44888 & n44907 ) | ( n44906 & n44907 ) ;
  assign n44909 = x680 | n44180 ;
  assign n44910 = ~x1100 & n44180 ;
  assign n44911 = ( x962 & n44909 ) | ( x962 & ~n44910 ) | ( n44909 & ~n44910 ) ;
  assign n44912 = ~x962 & n44911 ;
  assign n44913 = x681 | n44180 ;
  assign n44914 = ~x1103 & n44180 ;
  assign n44915 = ( x962 & n44913 ) | ( x962 & ~n44914 ) | ( n44913 & ~n44914 ) ;
  assign n44916 = ~x962 & n44915 ;
  assign n44917 = x392 & x591 ;
  assign n44918 = ~x592 & n44917 ;
  assign n44919 = x367 & n44339 ;
  assign n44920 = ( ~x590 & n44918 ) | ( ~x590 & n44919 ) | ( n44918 & n44919 ) ;
  assign n44921 = ~x590 & n44920 ;
  assign n44922 = x345 & n44347 ;
  assign n44923 = ( x588 & ~n44921 ) | ( x588 & n44922 ) | ( ~n44921 & n44922 ) ;
  assign n44924 = n44921 | n44923 ;
  assign n44925 = x199 | x251 ;
  assign n44926 = x199 & ~x1039 ;
  assign n44927 = n44352 & ~n44926 ;
  assign n44928 = n44925 & n44927 ;
  assign n44929 = x417 & ~n44356 ;
  assign n44930 = x588 & ~n44929 ;
  assign n44931 = n44352 | n44930 ;
  assign n44932 = ~n44928 & n44931 ;
  assign n44933 = ( n44924 & n44928 ) | ( n44924 & ~n44932 ) | ( n44928 & ~n44932 ) ;
  assign n44934 = x848 | x1136 ;
  assign n44935 = x686 & x1135 ;
  assign n44936 = n44934 & ~n44935 ;
  assign n44937 = x757 & n44375 ;
  assign n44938 = n44380 & ~n44937 ;
  assign n44939 = n44936 & n44938 ;
  assign n44940 = x631 & x1135 ;
  assign n44941 = x1134 | n44940 ;
  assign n44942 = ( x610 & x1135 ) | ( x610 & ~n44941 ) | ( x1135 & ~n44941 ) ;
  assign n44943 = ~n44941 & n44942 ;
  assign n44944 = n44939 ^ n44572 ^ 1'b0 ;
  assign n44945 = ( ~n44572 & n44943 ) | ( ~n44572 & n44944 ) | ( n44943 & n44944 ) ;
  assign n44946 = ( n44572 & n44939 ) | ( n44572 & n44945 ) | ( n44939 & n44945 ) ;
  assign n44947 = n44933 ^ n10841 ^ 1'b0 ;
  assign n44948 = ( n44933 & n44946 ) | ( n44933 & n44947 ) | ( n44946 & n44947 ) ;
  assign n44949 = x953 & n44179 ;
  assign n44950 = ~x1130 & n44949 ;
  assign n44951 = x962 | n44950 ;
  assign n44952 = n44949 & ~n44951 ;
  assign n44953 = ( x684 & n44951 ) | ( x684 & ~n44952 ) | ( n44951 & ~n44952 ) ;
  assign n44954 = x199 & ~x1076 ;
  assign n44955 = ( n40509 & n44352 ) | ( n40509 & n44954 ) | ( n44352 & n44954 ) ;
  assign n44956 = ~n44954 & n44955 ;
  assign n44957 = x588 & ~x590 ;
  assign n44958 = x406 & ~x592 ;
  assign n44959 = n44414 & n44958 ;
  assign n44960 = x357 & n44345 ;
  assign n44961 = x382 & n44412 ;
  assign n44962 = ( ~x591 & n44960 ) | ( ~x591 & n44961 ) | ( n44960 & n44961 ) ;
  assign n44963 = ~x591 & n44962 ;
  assign n44964 = ( ~x588 & n44959 ) | ( ~x588 & n44963 ) | ( n44959 & n44963 ) ;
  assign n44965 = ~x588 & n44964 ;
  assign n44966 = x430 & ~n44346 ;
  assign n44967 = n44965 ^ n44957 ^ 1'b0 ;
  assign n44968 = ( ~n44957 & n44966 ) | ( ~n44957 & n44967 ) | ( n44966 & n44967 ) ;
  assign n44969 = ( n44957 & n44965 ) | ( n44957 & n44968 ) | ( n44965 & n44968 ) ;
  assign n44970 = ( ~n44352 & n44956 ) | ( ~n44352 & n44969 ) | ( n44956 & n44969 ) ;
  assign n44971 = n44956 ^ n44352 ^ 1'b0 ;
  assign n44972 = ( n44956 & n44970 ) | ( n44956 & ~n44971 ) | ( n44970 & ~n44971 ) ;
  assign n44973 = x1136 & n44362 ;
  assign n44974 = x657 & x1135 ;
  assign n44975 = x652 | x1135 ;
  assign n44976 = ( x1136 & n44974 ) | ( x1136 & n44975 ) | ( n44974 & n44975 ) ;
  assign n44977 = ~n44974 & n44976 ;
  assign n44978 = x813 & ~n44362 ;
  assign n44979 = n44393 | n44978 ;
  assign n44980 = ( ~n44393 & n44977 ) | ( ~n44393 & n44979 ) | ( n44977 & n44979 ) ;
  assign n44981 = ( x1134 & ~n44973 ) | ( x1134 & n44980 ) | ( ~n44973 & n44980 ) ;
  assign n44982 = ~x1134 & n44981 ;
  assign n44983 = x728 & x1135 ;
  assign n44984 = x744 & ~x1135 ;
  assign n44985 = ( x1136 & n44983 ) | ( x1136 & ~n44984 ) | ( n44983 & ~n44984 ) ;
  assign n44986 = ~n44983 & n44985 ;
  assign n44987 = n44393 & ~n44986 ;
  assign n44988 = ( x860 & n44986 ) | ( x860 & ~n44987 ) | ( n44986 & ~n44987 ) ;
  assign n44989 = n44982 ^ n44379 ^ 1'b0 ;
  assign n44990 = ( ~n44379 & n44988 ) | ( ~n44379 & n44989 ) | ( n44988 & n44989 ) ;
  assign n44991 = ( n44379 & n44982 ) | ( n44379 & n44990 ) | ( n44982 & n44990 ) ;
  assign n44992 = n44972 ^ n10841 ^ 1'b0 ;
  assign n44993 = ( n44972 & n44991 ) | ( n44972 & n44992 ) | ( n44991 & n44992 ) ;
  assign n44994 = ~x1113 & n44949 ;
  assign n44995 = x962 | n44994 ;
  assign n44996 = n44949 & ~n44995 ;
  assign n44997 = ( x686 & n44995 ) | ( x686 & ~n44996 ) | ( n44995 & ~n44996 ) ;
  assign n44998 = x687 | n44949 ;
  assign n44999 = ~x1127 & n44949 ;
  assign n45000 = ( x962 & n44998 ) | ( x962 & ~n44999 ) | ( n44998 & ~n44999 ) ;
  assign n45001 = ~x962 & n45000 ;
  assign n45002 = ~x1115 & n44949 ;
  assign n45003 = x962 | n45002 ;
  assign n45004 = n44949 & ~n45003 ;
  assign n45005 = ( x688 & n45003 ) | ( x688 & ~n45004 ) | ( n45003 & ~n45004 ) ;
  assign n45006 = x199 & ~x1079 ;
  assign n45007 = x199 | n40487 ;
  assign n45008 = ( n44352 & n45006 ) | ( n44352 & n45007 ) | ( n45006 & n45007 ) ;
  assign n45009 = ~n45006 & n45008 ;
  assign n45010 = x401 & ~x592 ;
  assign n45011 = n44414 & n45010 ;
  assign n45012 = x351 & n44345 ;
  assign n45013 = x376 & n44412 ;
  assign n45014 = ( ~x591 & n45012 ) | ( ~x591 & n45013 ) | ( n45012 & n45013 ) ;
  assign n45015 = ~x591 & n45014 ;
  assign n45016 = ( ~x588 & n45011 ) | ( ~x588 & n45015 ) | ( n45011 & n45015 ) ;
  assign n45017 = ~x588 & n45016 ;
  assign n45018 = x426 & ~n44346 ;
  assign n45019 = n45017 ^ n44957 ^ 1'b0 ;
  assign n45020 = ( ~n44957 & n45018 ) | ( ~n44957 & n45019 ) | ( n45018 & n45019 ) ;
  assign n45021 = ( n44957 & n45017 ) | ( n44957 & n45020 ) | ( n45017 & n45020 ) ;
  assign n45022 = ( ~n44352 & n45009 ) | ( ~n44352 & n45021 ) | ( n45009 & n45021 ) ;
  assign n45023 = n45009 ^ n44352 ^ 1'b0 ;
  assign n45024 = ( n45009 & n45022 ) | ( n45009 & ~n45023 ) | ( n45022 & ~n45023 ) ;
  assign n45025 = x843 | x1136 ;
  assign n45026 = ~x703 & x1135 ;
  assign n45027 = n45025 & ~n45026 ;
  assign n45028 = x752 & n44375 ;
  assign n45029 = n44380 & ~n45028 ;
  assign n45030 = n45027 & n45029 ;
  assign n45031 = x655 & x1135 ;
  assign n45032 = x658 | x1135 ;
  assign n45033 = ( x1136 & n45031 ) | ( x1136 & n45032 ) | ( n45031 & n45032 ) ;
  assign n45034 = ~n45031 & n45033 ;
  assign n45035 = n44393 & ~n45034 ;
  assign n45036 = ( x798 & n45034 ) | ( x798 & ~n45035 ) | ( n45034 & ~n45035 ) ;
  assign n45037 = ( ~n44461 & n45030 ) | ( ~n44461 & n45036 ) | ( n45030 & n45036 ) ;
  assign n45038 = n45030 ^ n44461 ^ 1'b0 ;
  assign n45039 = ( n45030 & n45037 ) | ( n45030 & ~n45038 ) | ( n45037 & ~n45038 ) ;
  assign n45040 = n45024 ^ n10841 ^ 1'b0 ;
  assign n45041 = ( n45024 & n45039 ) | ( n45024 & n45040 ) | ( n45039 & n45040 ) ;
  assign n45042 = x690 | n44949 ;
  assign n45043 = ~x1108 & n44949 ;
  assign n45044 = ( x962 & n45042 ) | ( x962 & ~n45043 ) | ( n45042 & ~n45043 ) ;
  assign n45045 = ~x962 & n45044 ;
  assign n45046 = x691 | n44949 ;
  assign n45047 = ~x1107 & n44949 ;
  assign n45048 = ( x962 & n45046 ) | ( x962 & ~n45047 ) | ( n45046 & ~n45047 ) ;
  assign n45049 = ~x962 & n45048 ;
  assign n45050 = x801 & ~n44393 ;
  assign n45051 = x649 & x1135 ;
  assign n45052 = x656 | x1135 ;
  assign n45053 = ( x1136 & n45051 ) | ( x1136 & n45052 ) | ( n45051 & n45052 ) ;
  assign n45054 = ~n45051 & n45053 ;
  assign n45055 = ( x1134 & ~n45050 ) | ( x1134 & n45054 ) | ( ~n45050 & n45054 ) ;
  assign n45056 = n45050 | n45055 ;
  assign n45057 = ~x726 & x1135 ;
  assign n45058 = x770 & ~x1135 ;
  assign n45059 = ( x1136 & n45057 ) | ( x1136 & ~n45058 ) | ( n45057 & ~n45058 ) ;
  assign n45060 = ~n45057 & n45059 ;
  assign n45061 = x844 & ~n44393 ;
  assign n45062 = ( x1134 & n45060 ) | ( x1134 & ~n45061 ) | ( n45060 & ~n45061 ) ;
  assign n45063 = ~n45060 & n45062 ;
  assign n45064 = n44407 & ~n45063 ;
  assign n45065 = n45056 & n45064 ;
  assign n45066 = x199 & ~x1078 ;
  assign n45067 = x199 | n40495 ;
  assign n45068 = ( n44352 & n45066 ) | ( n44352 & n45067 ) | ( n45066 & n45067 ) ;
  assign n45069 = ~n45066 & n45068 ;
  assign n45070 = x402 & ~x592 ;
  assign n45071 = n44414 & n45070 ;
  assign n45072 = x352 & n44345 ;
  assign n45073 = x317 & n44412 ;
  assign n45074 = ( ~x591 & n45072 ) | ( ~x591 & n45073 ) | ( n45072 & n45073 ) ;
  assign n45075 = ~x591 & n45074 ;
  assign n45076 = ( ~x588 & n45071 ) | ( ~x588 & n45075 ) | ( n45071 & n45075 ) ;
  assign n45077 = ~x588 & n45076 ;
  assign n45078 = x427 & ~n44346 ;
  assign n45079 = n45077 ^ n44957 ^ 1'b0 ;
  assign n45080 = ( ~n44957 & n45078 ) | ( ~n44957 & n45079 ) | ( n45078 & n45079 ) ;
  assign n45081 = ( n44957 & n45077 ) | ( n44957 & n45080 ) | ( n45077 & n45080 ) ;
  assign n45082 = ( ~n44352 & n45069 ) | ( ~n44352 & n45081 ) | ( n45069 & n45081 ) ;
  assign n45083 = n45069 ^ n44352 ^ 1'b0 ;
  assign n45084 = ( n45069 & n45082 ) | ( n45069 & ~n45083 ) | ( n45082 & ~n45083 ) ;
  assign n45085 = ( ~n10841 & n45065 ) | ( ~n10841 & n45084 ) | ( n45065 & n45084 ) ;
  assign n45086 = n45065 ^ n10841 ^ 1'b0 ;
  assign n45087 = ( n45065 & n45085 ) | ( n45065 & ~n45086 ) | ( n45085 & ~n45086 ) ;
  assign n45088 = ~x1129 & n44180 ;
  assign n45089 = x962 | n45088 ;
  assign n45090 = n44180 & ~n45089 ;
  assign n45091 = ( x693 & n45089 ) | ( x693 & ~n45090 ) | ( n45089 & ~n45090 ) ;
  assign n45092 = ~x1128 & n44949 ;
  assign n45093 = x962 | n45092 ;
  assign n45094 = n44949 & ~n45093 ;
  assign n45095 = ( x694 & n45093 ) | ( x694 & ~n45094 ) | ( n45093 & ~n45094 ) ;
  assign n45096 = ~x1111 & n44180 ;
  assign n45097 = x962 | n45096 ;
  assign n45098 = n44180 & ~n45097 ;
  assign n45099 = ( x695 & n45097 ) | ( x695 & ~n45098 ) | ( n45097 & ~n45098 ) ;
  assign n45100 = x696 | n44949 ;
  assign n45101 = ~x1100 & n44949 ;
  assign n45102 = ( x962 & n45100 ) | ( x962 & ~n45101 ) | ( n45100 & ~n45101 ) ;
  assign n45103 = ~x962 & n45102 ;
  assign n45104 = ~x1129 & n44949 ;
  assign n45105 = x962 | n45104 ;
  assign n45106 = n44949 & ~n45105 ;
  assign n45107 = ( x697 & n45105 ) | ( x697 & ~n45106 ) | ( n45105 & ~n45106 ) ;
  assign n45108 = ~x1116 & n44949 ;
  assign n45109 = x962 | n45108 ;
  assign n45110 = n44949 & ~n45109 ;
  assign n45111 = ( x698 & n45109 ) | ( x698 & ~n45110 ) | ( n45109 & ~n45110 ) ;
  assign n45112 = x699 | n44949 ;
  assign n45113 = ~x1103 & n44949 ;
  assign n45114 = ( x962 & n45112 ) | ( x962 & ~n45113 ) | ( n45112 & ~n45113 ) ;
  assign n45115 = ~x962 & n45114 ;
  assign n45116 = x700 | n44949 ;
  assign n45117 = ~x1110 & n44949 ;
  assign n45118 = ( x962 & n45116 ) | ( x962 & ~n45117 ) | ( n45116 & ~n45117 ) ;
  assign n45119 = ~x962 & n45118 ;
  assign n45120 = ~x1123 & n44949 ;
  assign n45121 = x962 | n45120 ;
  assign n45122 = n44949 & ~n45121 ;
  assign n45123 = ( x701 & n45121 ) | ( x701 & ~n45122 ) | ( n45121 & ~n45122 ) ;
  assign n45124 = ~x1117 & n44949 ;
  assign n45125 = x962 | n45124 ;
  assign n45126 = n44949 & ~n45125 ;
  assign n45127 = ( x702 & n45125 ) | ( x702 & ~n45126 ) | ( n45125 & ~n45126 ) ;
  assign n45128 = x703 | n44949 ;
  assign n45129 = ~x1124 & n44949 ;
  assign n45130 = ( x962 & n45128 ) | ( x962 & ~n45129 ) | ( n45128 & ~n45129 ) ;
  assign n45131 = ~x962 & n45130 ;
  assign n45132 = ~x1112 & n44949 ;
  assign n45133 = x962 | n45132 ;
  assign n45134 = n44949 & ~n45133 ;
  assign n45135 = ( x704 & n45133 ) | ( x704 & ~n45134 ) | ( n45133 & ~n45134 ) ;
  assign n45136 = x705 | n44949 ;
  assign n45137 = ~x1125 & n44949 ;
  assign n45138 = ( x962 & n45136 ) | ( x962 & ~n45137 ) | ( n45136 & ~n45137 ) ;
  assign n45139 = ~x962 & n45138 ;
  assign n45140 = x706 | n44949 ;
  assign n45141 = ~x1105 & n44949 ;
  assign n45142 = ( x962 & n45140 ) | ( x962 & ~n45141 ) | ( n45140 & ~n45141 ) ;
  assign n45143 = ~x962 & n45142 ;
  assign n45144 = x395 & x591 ;
  assign n45145 = ~x592 & n45144 ;
  assign n45146 = x370 & n44339 ;
  assign n45147 = ( ~x590 & n45145 ) | ( ~x590 & n45146 ) | ( n45145 & n45146 ) ;
  assign n45148 = ~x590 & n45147 ;
  assign n45149 = n45148 ^ x347 ^ 1'b0 ;
  assign n45150 = ( ~x347 & n44347 ) | ( ~x347 & n45149 ) | ( n44347 & n45149 ) ;
  assign n45151 = ( x347 & n45148 ) | ( x347 & n45150 ) | ( n45148 & n45150 ) ;
  assign n45152 = x199 & ~x1055 ;
  assign n45153 = n44352 & ~n45152 ;
  assign n45154 = ( x304 & x1048 ) | ( x304 & ~n40490 ) | ( x1048 & ~n40490 ) ;
  assign n45155 = x199 | n45154 ;
  assign n45156 = n45153 & n45155 ;
  assign n45157 = n44352 | n44356 ;
  assign n45158 = x420 & x588 ;
  assign n45159 = n45158 ^ n45157 ^ 1'b0 ;
  assign n45160 = ( n45157 & n45158 ) | ( n45157 & n45159 ) | ( n45158 & n45159 ) ;
  assign n45161 = ( n45156 & ~n45157 ) | ( n45156 & n45160 ) | ( ~n45157 & n45160 ) ;
  assign n45162 = x588 | n44352 ;
  assign n45163 = ~n45161 & n45162 ;
  assign n45164 = ( n45151 & n45161 ) | ( n45151 & ~n45163 ) | ( n45161 & ~n45163 ) ;
  assign n45165 = x847 | x1136 ;
  assign n45166 = x702 & x1135 ;
  assign n45167 = n45165 & ~n45166 ;
  assign n45168 = x753 & n44375 ;
  assign n45169 = n44380 & ~n45168 ;
  assign n45170 = n45167 & n45169 ;
  assign n45171 = ~x627 & x1135 ;
  assign n45172 = x1134 | n45171 ;
  assign n45173 = ( x618 & x1135 ) | ( x618 & ~n45172 ) | ( x1135 & ~n45172 ) ;
  assign n45174 = ~n45172 & n45173 ;
  assign n45175 = n45170 ^ n44572 ^ 1'b0 ;
  assign n45176 = ( ~n44572 & n45174 ) | ( ~n44572 & n45175 ) | ( n45174 & n45175 ) ;
  assign n45177 = ( n44572 & n45170 ) | ( n44572 & n45176 ) | ( n45170 & n45176 ) ;
  assign n45178 = n45164 ^ n10841 ^ 1'b0 ;
  assign n45179 = ( n45164 & n45177 ) | ( n45164 & n45178 ) | ( n45177 & n45178 ) ;
  assign n45180 = n44362 | n44378 ;
  assign n45181 = x709 & x1135 ;
  assign n45182 = x1134 & ~n45181 ;
  assign n45183 = x857 | x1136 ;
  assign n45184 = ( n45180 & n45182 ) | ( n45180 & n45183 ) | ( n45182 & n45183 ) ;
  assign n45185 = ~n45180 & n45184 ;
  assign n45186 = ( x754 & n44375 ) | ( x754 & ~n45185 ) | ( n44375 & ~n45185 ) ;
  assign n45187 = n45186 ^ n45185 ^ 1'b0 ;
  assign n45188 = ( n45185 & ~n45186 ) | ( n45185 & n45187 ) | ( ~n45186 & n45187 ) ;
  assign n45189 = x609 | x1135 ;
  assign n45190 = ~x660 & x1135 ;
  assign n45191 = ( x1134 & n45189 ) | ( x1134 & ~n45190 ) | ( n45189 & ~n45190 ) ;
  assign n45192 = ~x1134 & n45191 ;
  assign n45193 = n44572 & n45192 ;
  assign n45194 = ( n10841 & n45188 ) | ( n10841 & ~n45193 ) | ( n45188 & ~n45193 ) ;
  assign n45195 = ~n45188 & n45194 ;
  assign n45196 = x321 & ~n44352 ;
  assign n45197 = n44347 & n45196 ;
  assign n45198 = x592 | n44352 ;
  assign n45199 = x328 & x591 ;
  assign n45200 = ~n45198 & n45199 ;
  assign n45201 = n44339 & ~n44352 ;
  assign n45202 = x442 & n45201 ;
  assign n45203 = ( ~x590 & n45200 ) | ( ~x590 & n45202 ) | ( n45200 & n45202 ) ;
  assign n45204 = ~x590 & n45203 ;
  assign n45205 = ( ~x588 & n45197 ) | ( ~x588 & n45204 ) | ( n45197 & n45204 ) ;
  assign n45206 = ~x588 & n45205 ;
  assign n45207 = n44346 | n44352 ;
  assign n45208 = x459 & n44957 ;
  assign n45209 = ~n45207 & n45208 ;
  assign n45210 = x199 & ~x1058 ;
  assign n45211 = n44352 & ~n45210 ;
  assign n45212 = x305 ^ x200 ^ 1'b0 ;
  assign n45213 = ( x305 & x1084 ) | ( x305 & n45212 ) | ( x1084 & n45212 ) ;
  assign n45214 = x199 | n45213 ;
  assign n45215 = n45211 & n45214 ;
  assign n45216 = ( n10841 & ~n45209 ) | ( n10841 & n45215 ) | ( ~n45209 & n45215 ) ;
  assign n45217 = n45209 | n45216 ;
  assign n45218 = ( ~n45195 & n45206 ) | ( ~n45195 & n45217 ) | ( n45206 & n45217 ) ;
  assign n45219 = ~n45195 & n45218 ;
  assign n45220 = ~x1118 & n44949 ;
  assign n45221 = x962 | n45220 ;
  assign n45222 = n44949 & ~n45221 ;
  assign n45223 = ( x709 & n45221 ) | ( x709 & ~n45222 ) | ( n45221 & ~n45222 ) ;
  assign n45224 = x710 | n44180 ;
  assign n45225 = ~x1106 & n44180 ;
  assign n45226 = ( x962 & n45224 ) | ( x962 & ~n45225 ) | ( n45224 & ~n45225 ) ;
  assign n45227 = ~x962 & n45226 ;
  assign n45228 = x398 & x591 ;
  assign n45229 = ~x592 & n45228 ;
  assign n45230 = x373 & n44339 ;
  assign n45231 = ( ~x590 & n45229 ) | ( ~x590 & n45230 ) | ( n45229 & n45230 ) ;
  assign n45232 = ~x590 & n45231 ;
  assign n45233 = x348 & n44347 ;
  assign n45234 = ( ~n45162 & n45232 ) | ( ~n45162 & n45233 ) | ( n45232 & n45233 ) ;
  assign n45235 = ~n45162 & n45234 ;
  assign n45236 = x199 & ~x1087 ;
  assign n45237 = n44352 & ~n45236 ;
  assign n45238 = ( x306 & x1059 ) | ( x306 & ~n40502 ) | ( x1059 & ~n40502 ) ;
  assign n45239 = x199 | n45238 ;
  assign n45240 = n45237 & n45239 ;
  assign n45241 = x423 & x588 ;
  assign n45242 = ~n45157 & n45241 ;
  assign n45243 = ( ~n45235 & n45240 ) | ( ~n45235 & n45242 ) | ( n45240 & n45242 ) ;
  assign n45244 = n45235 | n45243 ;
  assign n45245 = x858 | x1136 ;
  assign n45246 = x725 & x1135 ;
  assign n45247 = n45245 & ~n45246 ;
  assign n45248 = x755 & n44375 ;
  assign n45249 = n44380 & ~n45248 ;
  assign n45250 = n45247 & n45249 ;
  assign n45251 = ~x647 & x1135 ;
  assign n45252 = x1134 | n45251 ;
  assign n45253 = ( x630 & x1135 ) | ( x630 & ~n45252 ) | ( x1135 & ~n45252 ) ;
  assign n45254 = ~n45252 & n45253 ;
  assign n45255 = n45250 ^ n44572 ^ 1'b0 ;
  assign n45256 = ( ~n44572 & n45254 ) | ( ~n44572 & n45255 ) | ( n45254 & n45255 ) ;
  assign n45257 = ( n44572 & n45250 ) | ( n44572 & n45256 ) | ( n45250 & n45256 ) ;
  assign n45258 = n45244 ^ n10841 ^ 1'b0 ;
  assign n45259 = ( n45244 & n45257 ) | ( n45244 & n45258 ) | ( n45257 & n45258 ) ;
  assign n45260 = x400 & x591 ;
  assign n45261 = ~x592 & n45260 ;
  assign n45262 = x374 & n44339 ;
  assign n45263 = ( ~x590 & n45261 ) | ( ~x590 & n45262 ) | ( n45261 & n45262 ) ;
  assign n45264 = ~x590 & n45263 ;
  assign n45265 = x350 & n44347 ;
  assign n45266 = ( ~x588 & n45264 ) | ( ~x588 & n45265 ) | ( n45264 & n45265 ) ;
  assign n45267 = ~x588 & n45266 ;
  assign n45268 = x425 & ~n44346 ;
  assign n45269 = n44957 & n45268 ;
  assign n45270 = ( n44352 & ~n45267 ) | ( n44352 & n45269 ) | ( ~n45267 & n45269 ) ;
  assign n45271 = n45267 | n45270 ;
  assign n45272 = ~x715 & x1135 ;
  assign n45273 = x1134 | n45272 ;
  assign n45274 = ( x644 & x1135 ) | ( x644 & ~n45273 ) | ( x1135 & ~n45273 ) ;
  assign n45275 = ~n45273 & n45274 ;
  assign n45276 = n44572 & n45275 ;
  assign n45277 = x751 & n44375 ;
  assign n45278 = x701 & x1135 ;
  assign n45279 = x1134 & ~n45278 ;
  assign n45280 = x842 | x1136 ;
  assign n45281 = n45279 & n45280 ;
  assign n45282 = ( n45180 & ~n45277 ) | ( n45180 & n45281 ) | ( ~n45277 & n45281 ) ;
  assign n45283 = ~n45180 & n45282 ;
  assign n45284 = ( n10841 & n45276 ) | ( n10841 & n45283 ) | ( n45276 & n45283 ) ;
  assign n45285 = n45283 ^ n45276 ^ 1'b0 ;
  assign n45286 = ( n10841 & n45284 ) | ( n10841 & n45285 ) | ( n45284 & n45285 ) ;
  assign n45287 = x1044 & n10073 ;
  assign n45288 = x298 & ~n9353 ;
  assign n45289 = x199 & x1035 ;
  assign n45290 = n44352 & ~n45289 ;
  assign n45291 = ( n45287 & ~n45288 ) | ( n45287 & n45290 ) | ( ~n45288 & n45290 ) ;
  assign n45292 = ~n45287 & n45291 ;
  assign n45293 = ( x1163 & n7441 ) | ( x1163 & ~n45292 ) | ( n7441 & ~n45292 ) ;
  assign n45294 = n45292 | n45293 ;
  assign n45295 = ~n45286 & n45294 ;
  assign n45296 = ( n45271 & n45286 ) | ( n45271 & ~n45295 ) | ( n45286 & ~n45295 ) ;
  assign n45297 = x396 & x591 ;
  assign n45298 = ~x592 & n45297 ;
  assign n45299 = x371 & n44339 ;
  assign n45300 = ( ~x590 & n45298 ) | ( ~x590 & n45299 ) | ( n45298 & n45299 ) ;
  assign n45301 = ~x590 & n45300 ;
  assign n45302 = x322 & n44347 ;
  assign n45303 = ( ~n45162 & n45301 ) | ( ~n45162 & n45302 ) | ( n45301 & n45302 ) ;
  assign n45304 = ~n45162 & n45303 ;
  assign n45305 = x199 & ~x1051 ;
  assign n45306 = n44352 & ~n45305 ;
  assign n45307 = x309 ^ x200 ^ 1'b0 ;
  assign n45308 = ( x309 & x1072 ) | ( x309 & n45307 ) | ( x1072 & n45307 ) ;
  assign n45309 = x199 | n45308 ;
  assign n45310 = n45306 & n45309 ;
  assign n45311 = x421 & x588 ;
  assign n45312 = ~n45157 & n45311 ;
  assign n45313 = ( ~n45304 & n45310 ) | ( ~n45304 & n45312 ) | ( n45310 & n45312 ) ;
  assign n45314 = n45304 | n45313 ;
  assign n45315 = x854 | x1136 ;
  assign n45316 = x734 & x1135 ;
  assign n45317 = n45315 & ~n45316 ;
  assign n45318 = x756 & n44375 ;
  assign n45319 = n44380 & ~n45318 ;
  assign n45320 = n45317 & n45319 ;
  assign n45321 = ~x628 & x1135 ;
  assign n45322 = x1134 | n45321 ;
  assign n45323 = ( x629 & x1135 ) | ( x629 & ~n45322 ) | ( x1135 & ~n45322 ) ;
  assign n45324 = ~n45322 & n45323 ;
  assign n45325 = n45320 ^ n44572 ^ 1'b0 ;
  assign n45326 = ( ~n44572 & n45324 ) | ( ~n44572 & n45325 ) | ( n45324 & n45325 ) ;
  assign n45327 = ( n44572 & n45320 ) | ( n44572 & n45326 ) | ( n45320 & n45326 ) ;
  assign n45328 = n45314 ^ n10841 ^ 1'b0 ;
  assign n45329 = ( n45314 & n45327 ) | ( n45314 & n45328 ) | ( n45327 & n45328 ) ;
  assign n45330 = x199 & ~x1057 ;
  assign n45331 = ( n39964 & n44352 ) | ( n39964 & n45330 ) | ( n44352 & n45330 ) ;
  assign n45332 = ~n45330 & n45331 ;
  assign n45333 = x326 & ~x592 ;
  assign n45334 = n44414 & n45333 ;
  assign n45335 = x461 & n44345 ;
  assign n45336 = x439 & n44412 ;
  assign n45337 = ( ~x591 & n45335 ) | ( ~x591 & n45336 ) | ( n45335 & n45336 ) ;
  assign n45338 = ~x591 & n45337 ;
  assign n45339 = ( ~x588 & n45334 ) | ( ~x588 & n45338 ) | ( n45334 & n45338 ) ;
  assign n45340 = ~x588 & n45339 ;
  assign n45341 = x449 & ~n44346 ;
  assign n45342 = n45340 ^ n44957 ^ 1'b0 ;
  assign n45343 = ( ~n44957 & n45341 ) | ( ~n44957 & n45342 ) | ( n45341 & n45342 ) ;
  assign n45344 = ( n44957 & n45340 ) | ( n44957 & n45343 ) | ( n45340 & n45343 ) ;
  assign n45345 = ( ~n44352 & n45332 ) | ( ~n44352 & n45344 ) | ( n45332 & n45344 ) ;
  assign n45346 = n45332 ^ n44352 ^ 1'b0 ;
  assign n45347 = ( n45332 & n45345 ) | ( n45332 & ~n45346 ) | ( n45345 & ~n45346 ) ;
  assign n45348 = x693 & x1135 ;
  assign n45349 = x653 | x1135 ;
  assign n45350 = ( x1136 & n45348 ) | ( x1136 & n45349 ) | ( n45348 & n45349 ) ;
  assign n45351 = ~n45348 & n45350 ;
  assign n45352 = x816 & ~n44362 ;
  assign n45353 = n44393 | n45352 ;
  assign n45354 = ( ~n44393 & n45351 ) | ( ~n44393 & n45353 ) | ( n45351 & n45353 ) ;
  assign n45355 = ( x1134 & ~n44973 ) | ( x1134 & n45354 ) | ( ~n44973 & n45354 ) ;
  assign n45356 = ~x1134 & n45355 ;
  assign n45357 = x697 & x1135 ;
  assign n45358 = x762 & ~x1135 ;
  assign n45359 = ( x1136 & n45357 ) | ( x1136 & ~n45358 ) | ( n45357 & ~n45358 ) ;
  assign n45360 = ~n45357 & n45359 ;
  assign n45361 = n44393 & ~n45360 ;
  assign n45362 = ( x867 & n45360 ) | ( x867 & ~n45361 ) | ( n45360 & ~n45361 ) ;
  assign n45363 = n45356 ^ n44379 ^ 1'b0 ;
  assign n45364 = ( ~n44379 & n45362 ) | ( ~n44379 & n45363 ) | ( n45362 & n45363 ) ;
  assign n45365 = ( n44379 & n45356 ) | ( n44379 & n45364 ) | ( n45356 & n45364 ) ;
  assign n45366 = n45347 ^ n10841 ^ 1'b0 ;
  assign n45367 = ( n45347 & n45365 ) | ( n45347 & n45366 ) | ( n45365 & n45366 ) ;
  assign n45368 = x715 | n44180 ;
  assign n45369 = ~x1123 & n44180 ;
  assign n45370 = ( x962 & n45368 ) | ( x962 & ~n45369 ) | ( n45368 & ~n45369 ) ;
  assign n45371 = ~x962 & n45370 ;
  assign n45372 = x738 & x1135 ;
  assign n45373 = x1134 & ~n45372 ;
  assign n45374 = x845 | x1136 ;
  assign n45375 = ( n45180 & n45373 ) | ( n45180 & n45374 ) | ( n45373 & n45374 ) ;
  assign n45376 = ~n45180 & n45375 ;
  assign n45377 = ( x761 & n44375 ) | ( x761 & ~n45376 ) | ( n44375 & ~n45376 ) ;
  assign n45378 = n45377 ^ n45376 ^ 1'b0 ;
  assign n45379 = ( n45376 & ~n45377 ) | ( n45376 & n45378 ) | ( ~n45377 & n45378 ) ;
  assign n45380 = x626 | x1135 ;
  assign n45381 = ~x641 & x1135 ;
  assign n45382 = ( x1134 & n45380 ) | ( x1134 & ~n45381 ) | ( n45380 & ~n45381 ) ;
  assign n45383 = ~x1134 & n45382 ;
  assign n45384 = n44572 & n45383 ;
  assign n45385 = ( n10841 & n45379 ) | ( n10841 & ~n45384 ) | ( n45379 & ~n45384 ) ;
  assign n45386 = ~n45379 & n45385 ;
  assign n45387 = x349 & ~n44352 ;
  assign n45388 = n44347 & n45387 ;
  assign n45389 = x329 & x591 ;
  assign n45390 = ~n45198 & n45389 ;
  assign n45391 = x440 & n45201 ;
  assign n45392 = ( ~x590 & n45390 ) | ( ~x590 & n45391 ) | ( n45390 & n45391 ) ;
  assign n45393 = ~x590 & n45392 ;
  assign n45394 = ( ~x588 & n45388 ) | ( ~x588 & n45393 ) | ( n45388 & n45393 ) ;
  assign n45395 = ~x588 & n45394 ;
  assign n45396 = x454 & n44957 ;
  assign n45397 = ~n45207 & n45396 ;
  assign n45398 = x199 & ~x1043 ;
  assign n45399 = n44352 & ~n45398 ;
  assign n45400 = x307 ^ x200 ^ 1'b0 ;
  assign n45401 = ( x307 & x1053 ) | ( x307 & n45400 ) | ( x1053 & n45400 ) ;
  assign n45402 = x199 | n45401 ;
  assign n45403 = n45399 & n45402 ;
  assign n45404 = ( n10841 & ~n45397 ) | ( n10841 & n45403 ) | ( ~n45397 & n45403 ) ;
  assign n45405 = n45397 | n45404 ;
  assign n45406 = ( ~n45386 & n45395 ) | ( ~n45386 & n45405 ) | ( n45395 & n45405 ) ;
  assign n45407 = ~n45386 & n45406 ;
  assign n45408 = x318 & x591 ;
  assign n45409 = ~x592 & n45408 ;
  assign n45410 = ~x591 & n6637 ;
  assign n45411 = ( ~x590 & n45409 ) | ( ~x590 & n45410 ) | ( n45409 & n45410 ) ;
  assign n45412 = ~x590 & n45411 ;
  assign n45413 = x462 & n44347 ;
  assign n45414 = ( ~n45162 & n45412 ) | ( ~n45162 & n45413 ) | ( n45412 & n45413 ) ;
  assign n45415 = ~n45162 & n45414 ;
  assign n45416 = x448 & x588 ;
  assign n45417 = ~n45157 & n45416 ;
  assign n45418 = x199 & ~x1074 ;
  assign n45419 = x199 | n40491 ;
  assign n45420 = ( n44352 & n45418 ) | ( n44352 & n45419 ) | ( n45418 & n45419 ) ;
  assign n45421 = ~n45418 & n45420 ;
  assign n45422 = ( ~n45415 & n45417 ) | ( ~n45415 & n45421 ) | ( n45417 & n45421 ) ;
  assign n45423 = n45415 | n45422 ;
  assign n45424 = x669 & x1135 ;
  assign n45425 = x645 | x1135 ;
  assign n45426 = ( x1136 & n45424 ) | ( x1136 & n45425 ) | ( n45424 & n45425 ) ;
  assign n45427 = ~n45424 & n45426 ;
  assign n45428 = x800 & ~n44393 ;
  assign n45429 = ( ~n44461 & n45427 ) | ( ~n44461 & n45428 ) | ( n45427 & n45428 ) ;
  assign n45430 = ~n44461 & n45429 ;
  assign n45431 = x768 & n44375 ;
  assign n45432 = ~x705 & x1135 ;
  assign n45433 = x1134 & ~n45432 ;
  assign n45434 = x839 | x1136 ;
  assign n45435 = ( n45180 & n45433 ) | ( n45180 & n45434 ) | ( n45433 & n45434 ) ;
  assign n45436 = ~n45180 & n45435 ;
  assign n45437 = ( n45430 & ~n45431 ) | ( n45430 & n45436 ) | ( ~n45431 & n45436 ) ;
  assign n45438 = n45431 ^ n45430 ^ 1'b0 ;
  assign n45439 = ( n45430 & n45437 ) | ( n45430 & ~n45438 ) | ( n45437 & ~n45438 ) ;
  assign n45440 = n45423 ^ n10841 ^ 1'b0 ;
  assign n45441 = ( n45423 & n45439 ) | ( n45423 & n45440 ) | ( n45439 & n45440 ) ;
  assign n45442 = x698 & x1135 ;
  assign n45443 = x1134 & ~n45442 ;
  assign n45444 = x853 | x1136 ;
  assign n45445 = ( n45180 & n45443 ) | ( n45180 & n45444 ) | ( n45443 & n45444 ) ;
  assign n45446 = ~n45180 & n45445 ;
  assign n45447 = ( x767 & n44375 ) | ( x767 & ~n45446 ) | ( n44375 & ~n45446 ) ;
  assign n45448 = n45447 ^ n45446 ^ 1'b0 ;
  assign n45449 = ( n45446 & ~n45447 ) | ( n45446 & n45448 ) | ( ~n45447 & n45448 ) ;
  assign n45450 = x608 | x1135 ;
  assign n45451 = ~x625 & x1135 ;
  assign n45452 = ( x1134 & n45450 ) | ( x1134 & ~n45451 ) | ( n45450 & ~n45451 ) ;
  assign n45453 = ~x1134 & n45452 ;
  assign n45454 = n44572 & n45453 ;
  assign n45455 = ( n10841 & n45449 ) | ( n10841 & ~n45454 ) | ( n45449 & ~n45454 ) ;
  assign n45456 = ~n45449 & n45455 ;
  assign n45457 = x315 & ~n44352 ;
  assign n45458 = n44347 & n45457 ;
  assign n45459 = x394 & x591 ;
  assign n45460 = ~n45198 & n45459 ;
  assign n45461 = x369 & n45201 ;
  assign n45462 = ( ~x590 & n45460 ) | ( ~x590 & n45461 ) | ( n45460 & n45461 ) ;
  assign n45463 = ~x590 & n45462 ;
  assign n45464 = ( ~x588 & n45458 ) | ( ~x588 & n45463 ) | ( n45458 & n45463 ) ;
  assign n45465 = ~x588 & n45464 ;
  assign n45466 = x419 & n44957 ;
  assign n45467 = ~n45207 & n45466 ;
  assign n45468 = x199 & ~x1080 ;
  assign n45469 = n44352 & ~n45468 ;
  assign n45470 = x303 ^ x200 ^ 1'b0 ;
  assign n45471 = ( x303 & x1049 ) | ( x303 & n45470 ) | ( x1049 & n45470 ) ;
  assign n45472 = x199 | n45471 ;
  assign n45473 = n45469 & n45472 ;
  assign n45474 = ( n10841 & ~n45467 ) | ( n10841 & n45473 ) | ( ~n45467 & n45473 ) ;
  assign n45475 = n45467 | n45474 ;
  assign n45476 = ( ~n45456 & n45465 ) | ( ~n45456 & n45475 ) | ( n45465 & n45475 ) ;
  assign n45477 = ~n45456 & n45476 ;
  assign n45478 = x378 & n44339 ;
  assign n45479 = x325 & x591 ;
  assign n45480 = ~x592 & n45479 ;
  assign n45481 = ( ~x590 & n45478 ) | ( ~x590 & n45480 ) | ( n45478 & n45480 ) ;
  assign n45482 = ~x590 & n45481 ;
  assign n45483 = x353 & n44347 ;
  assign n45484 = ( ~n45162 & n45482 ) | ( ~n45162 & n45483 ) | ( n45482 & n45483 ) ;
  assign n45485 = ~n45162 & n45484 ;
  assign n45486 = x451 & x588 ;
  assign n45487 = ~n45157 & n45486 ;
  assign n45488 = x199 & ~x1063 ;
  assign n45489 = x199 | n40499 ;
  assign n45490 = ( n44352 & n45488 ) | ( n44352 & n45489 ) | ( n45488 & n45489 ) ;
  assign n45491 = ~n45488 & n45490 ;
  assign n45492 = ( ~n45485 & n45487 ) | ( ~n45485 & n45491 ) | ( n45487 & n45491 ) ;
  assign n45493 = n45485 | n45492 ;
  assign n45494 = x650 & x1135 ;
  assign n45495 = x636 | x1135 ;
  assign n45496 = ( x1136 & n45494 ) | ( x1136 & n45495 ) | ( n45494 & n45495 ) ;
  assign n45497 = ~n45494 & n45496 ;
  assign n45498 = x807 & ~n44393 ;
  assign n45499 = ( ~n44461 & n45497 ) | ( ~n44461 & n45498 ) | ( n45497 & n45498 ) ;
  assign n45500 = ~n44461 & n45499 ;
  assign n45501 = x774 & n44375 ;
  assign n45502 = ~x687 & x1135 ;
  assign n45503 = x1134 & ~n45502 ;
  assign n45504 = x868 | x1136 ;
  assign n45505 = ( n45180 & n45503 ) | ( n45180 & n45504 ) | ( n45503 & n45504 ) ;
  assign n45506 = ~n45180 & n45505 ;
  assign n45507 = ( n45500 & ~n45501 ) | ( n45500 & n45506 ) | ( ~n45501 & n45506 ) ;
  assign n45508 = n45501 ^ n45500 ^ 1'b0 ;
  assign n45509 = ( n45500 & n45507 ) | ( n45500 & ~n45508 ) | ( n45507 & ~n45508 ) ;
  assign n45510 = n45493 ^ n10841 ^ 1'b0 ;
  assign n45511 = ( n45493 & n45509 ) | ( n45493 & n45510 ) | ( n45509 & n45510 ) ;
  assign n45512 = x199 & ~x1081 ;
  assign n45513 = ( n40515 & n44352 ) | ( n40515 & n45512 ) | ( n44352 & n45512 ) ;
  assign n45514 = ~n45512 & n45513 ;
  assign n45515 = x405 & ~x592 ;
  assign n45516 = n44414 & n45515 ;
  assign n45517 = x356 & n44345 ;
  assign n45518 = x381 & n44412 ;
  assign n45519 = ( ~x591 & n45517 ) | ( ~x591 & n45518 ) | ( n45517 & n45518 ) ;
  assign n45520 = ~x591 & n45519 ;
  assign n45521 = ( ~x588 & n45516 ) | ( ~x588 & n45520 ) | ( n45516 & n45520 ) ;
  assign n45522 = ~x588 & n45521 ;
  assign n45523 = x445 & ~n44346 ;
  assign n45524 = n45522 ^ n44957 ^ 1'b0 ;
  assign n45525 = ( ~n44957 & n45523 ) | ( ~n44957 & n45524 ) | ( n45523 & n45524 ) ;
  assign n45526 = ( n44957 & n45522 ) | ( n44957 & n45525 ) | ( n45522 & n45525 ) ;
  assign n45527 = ( ~n44352 & n45514 ) | ( ~n44352 & n45526 ) | ( n45514 & n45526 ) ;
  assign n45528 = n45514 ^ n44352 ^ 1'b0 ;
  assign n45529 = ( n45514 & n45527 ) | ( n45514 & ~n45528 ) | ( n45527 & ~n45528 ) ;
  assign n45530 = x654 & x1135 ;
  assign n45531 = x651 | x1135 ;
  assign n45532 = ( x1136 & n45530 ) | ( x1136 & n45531 ) | ( n45530 & n45531 ) ;
  assign n45533 = ~n45530 & n45532 ;
  assign n45534 = x794 & ~n44362 ;
  assign n45535 = n44393 | n45534 ;
  assign n45536 = ( ~n44393 & n45533 ) | ( ~n44393 & n45535 ) | ( n45533 & n45535 ) ;
  assign n45537 = ( x1134 & ~n44973 ) | ( x1134 & n45536 ) | ( ~n44973 & n45536 ) ;
  assign n45538 = ~x1134 & n45537 ;
  assign n45539 = x684 & x1135 ;
  assign n45540 = x750 & ~x1135 ;
  assign n45541 = ( x1136 & n45539 ) | ( x1136 & ~n45540 ) | ( n45539 & ~n45540 ) ;
  assign n45542 = ~n45539 & n45541 ;
  assign n45543 = n44393 & ~n45542 ;
  assign n45544 = ( x880 & n45542 ) | ( x880 & ~n45543 ) | ( n45542 & ~n45543 ) ;
  assign n45545 = n45538 ^ n44379 ^ 1'b0 ;
  assign n45546 = ( ~n44379 & n45544 ) | ( ~n44379 & n45545 ) | ( n45544 & n45545 ) ;
  assign n45547 = ( n44379 & n45538 ) | ( n44379 & n45546 ) | ( n45538 & n45546 ) ;
  assign n45548 = n45529 ^ n10841 ^ 1'b0 ;
  assign n45549 = ( n45529 & n45547 ) | ( n45529 & n45548 ) | ( n45547 & n45548 ) ;
  assign n45550 = x773 | x801 ;
  assign n45551 = x773 & x801 ;
  assign n45552 = n45550 & ~n45551 ;
  assign n45553 = x800 ^ x771 ^ 1'b0 ;
  assign n45554 = x794 ^ x769 ^ 1'b0 ;
  assign n45555 = x798 ^ x765 ^ 1'b0 ;
  assign n45556 = x807 & ~n45555 ;
  assign n45557 = x747 & n45556 ;
  assign n45558 = x747 | x807 ;
  assign n45559 = n45555 | n45558 ;
  assign n45560 = ~n45557 & n45559 ;
  assign n45561 = n45554 | n45560 ;
  assign n45562 = n45553 | n45561 ;
  assign n45563 = n45552 | n45562 ;
  assign n45564 = x721 & x813 ;
  assign n45565 = ~n45563 & n45564 ;
  assign n45566 = ~n45553 & n45556 ;
  assign n45567 = x721 | x813 ;
  assign n45568 = x794 & x801 ;
  assign n45569 = ~n45567 & n45568 ;
  assign n45570 = n45566 & n45569 ;
  assign n45571 = ( x816 & n45565 ) | ( x816 & n45570 ) | ( n45565 & n45570 ) ;
  assign n45572 = n45570 ^ n45565 ^ 1'b0 ;
  assign n45573 = ( x816 & n45571 ) | ( x816 & n45572 ) | ( n45571 & n45572 ) ;
  assign n45574 = x747 & x773 ;
  assign n45575 = x769 & n45574 ;
  assign n45576 = x775 ^ x721 ^ 1'b0 ;
  assign n45577 = ( x721 & ~n45575 ) | ( x721 & n45576 ) | ( ~n45575 & n45576 ) ;
  assign n45578 = n45577 ^ n45576 ^ 1'b0 ;
  assign n45579 = x795 & ~n45578 ;
  assign n45580 = ( x795 & n45573 ) | ( x795 & n45579 ) | ( n45573 & n45579 ) ;
  assign n45581 = ~x945 & x988 ;
  assign n45582 = x731 & n45581 ;
  assign n45583 = x721 & ~x775 ;
  assign n45584 = n45578 | n45583 ;
  assign n45585 = ( n45580 & n45582 ) | ( n45580 & n45584 ) | ( n45582 & n45584 ) ;
  assign n45586 = ~n45580 & n45585 ;
  assign n45587 = x775 | x816 ;
  assign n45588 = x775 & x816 ;
  assign n45589 = n45587 & ~n45588 ;
  assign n45590 = n45565 & ~n45589 ;
  assign n45591 = n45583 & ~n45590 ;
  assign n45592 = x721 & ~n45582 ;
  assign n45593 = x731 | x795 ;
  assign n45594 = x731 & x795 ;
  assign n45595 = n45593 & ~n45594 ;
  assign n45596 = n45590 & ~n45595 ;
  assign n45597 = n45592 & ~n45596 ;
  assign n45598 = ( ~n45586 & n45591 ) | ( ~n45586 & n45597 ) | ( n45591 & n45597 ) ;
  assign n45599 = n45586 | n45598 ;
  assign n45600 = x199 & ~x1045 ;
  assign n45601 = x199 | n40503 ;
  assign n45602 = ( n44352 & n45600 ) | ( n44352 & n45601 ) | ( n45600 & n45601 ) ;
  assign n45603 = ~n45600 & n45602 ;
  assign n45604 = x428 & x588 ;
  assign n45605 = ( ~n45157 & n45603 ) | ( ~n45157 & n45604 ) | ( n45603 & n45604 ) ;
  assign n45606 = n45603 ^ n45157 ^ 1'b0 ;
  assign n45607 = ( n45603 & n45605 ) | ( n45603 & ~n45606 ) | ( n45605 & ~n45606 ) ;
  assign n45608 = x403 & x591 ;
  assign n45609 = ~x592 & n45608 ;
  assign n45610 = x379 & n44339 ;
  assign n45611 = ( ~x590 & n45609 ) | ( ~x590 & n45610 ) | ( n45609 & n45610 ) ;
  assign n45612 = ~x590 & n45611 ;
  assign n45613 = x354 & n44347 ;
  assign n45614 = ( ~n45162 & n45612 ) | ( ~n45162 & n45613 ) | ( n45612 & n45613 ) ;
  assign n45615 = ~n45162 & n45614 ;
  assign n45616 = ( ~n10841 & n45607 ) | ( ~n10841 & n45615 ) | ( n45607 & n45615 ) ;
  assign n45617 = ~n10841 & n45616 ;
  assign n45618 = x694 & x1134 ;
  assign n45619 = n44369 & ~n45618 ;
  assign n45620 = x640 | x1134 ;
  assign n45621 = x776 & x1134 ;
  assign n45622 = x1136 & ~n45621 ;
  assign n45623 = n45620 & n45622 ;
  assign n45624 = ~x851 & x1134 ;
  assign n45625 = x795 | x1134 ;
  assign n45626 = ( x1136 & ~n45624 ) | ( x1136 & n45625 ) | ( ~n45624 & n45625 ) ;
  assign n45627 = ~x1136 & n45626 ;
  assign n45628 = ( ~x1135 & n45623 ) | ( ~x1135 & n45627 ) | ( n45623 & n45627 ) ;
  assign n45629 = ~x1135 & n45628 ;
  assign n45630 = x732 & ~x1134 ;
  assign n45631 = ~n45629 & n45630 ;
  assign n45632 = ( n45619 & n45629 ) | ( n45619 & ~n45631 ) | ( n45629 & ~n45631 ) ;
  assign n45633 = n45617 ^ n44407 ^ 1'b0 ;
  assign n45634 = ( ~n44407 & n45632 ) | ( ~n44407 & n45633 ) | ( n45632 & n45633 ) ;
  assign n45635 = ( n44407 & n45617 ) | ( n44407 & n45634 ) | ( n45617 & n45634 ) ;
  assign n45636 = ~x1111 & n44949 ;
  assign n45637 = x962 | n45636 ;
  assign n45638 = n44949 & ~n45637 ;
  assign n45639 = ( x723 & n45637 ) | ( x723 & ~n45638 ) | ( n45637 & ~n45638 ) ;
  assign n45640 = ~x1114 & n44949 ;
  assign n45641 = x962 | n45640 ;
  assign n45642 = n44949 & ~n45641 ;
  assign n45643 = ( x724 & n45641 ) | ( x724 & ~n45642 ) | ( n45641 & ~n45642 ) ;
  assign n45644 = ~x1120 & n44949 ;
  assign n45645 = x962 | n45644 ;
  assign n45646 = n44949 & ~n45645 ;
  assign n45647 = ( x725 & n45645 ) | ( x725 & ~n45646 ) | ( n45645 & ~n45646 ) ;
  assign n45648 = x726 | n44949 ;
  assign n45649 = ~x1126 & n44949 ;
  assign n45650 = ( x962 & n45648 ) | ( x962 & ~n45649 ) | ( n45648 & ~n45649 ) ;
  assign n45651 = ~x962 & n45650 ;
  assign n45652 = x727 | n44949 ;
  assign n45653 = ~x1102 & n44949 ;
  assign n45654 = ( x962 & n45652 ) | ( x962 & ~n45653 ) | ( n45652 & ~n45653 ) ;
  assign n45655 = ~x962 & n45654 ;
  assign n45656 = ~x1131 & n44949 ;
  assign n45657 = x962 | n45656 ;
  assign n45658 = n44949 & ~n45657 ;
  assign n45659 = ( x728 & n45657 ) | ( x728 & ~n45658 ) | ( n45657 & ~n45658 ) ;
  assign n45660 = x729 | n44949 ;
  assign n45661 = ~x1104 & n44949 ;
  assign n45662 = ( x962 & n45660 ) | ( x962 & ~n45661 ) | ( n45660 & ~n45661 ) ;
  assign n45663 = ~x962 & n45662 ;
  assign n45664 = x730 | n44949 ;
  assign n45665 = ~x1106 & n44949 ;
  assign n45666 = ( x962 & n45664 ) | ( x962 & ~n45665 ) | ( n45664 & ~n45665 ) ;
  assign n45667 = ~x962 & n45666 ;
  assign n45668 = ~n45564 & n45567 ;
  assign n45669 = n45589 | n45668 ;
  assign n45670 = ~x795 & x801 ;
  assign n45671 = ( n45554 & ~n45669 ) | ( n45554 & n45670 ) | ( ~n45669 & n45670 ) ;
  assign n45672 = ~n45554 & n45671 ;
  assign n45673 = n45574 & ~n45672 ;
  assign n45674 = ( ~n45566 & n45574 ) | ( ~n45566 & n45673 ) | ( n45574 & n45673 ) ;
  assign n45675 = ( x731 & n45581 ) | ( x731 & n45674 ) | ( n45581 & n45674 ) ;
  assign n45676 = n45581 & n45675 ;
  assign n45677 = n45563 | n45668 ;
  assign n45678 = x795 & ~n45589 ;
  assign n45679 = ~n45677 & n45678 ;
  assign n45680 = ~n45676 & n45679 ;
  assign n45681 = ( x731 & n45676 ) | ( x731 & ~n45680 ) | ( n45676 & ~n45680 ) ;
  assign n45682 = n45574 | n45679 ;
  assign n45683 = ( n45582 & ~n45681 ) | ( n45582 & n45682 ) | ( ~n45681 & n45682 ) ;
  assign n45684 = n45683 ^ n45681 ^ 1'b0 ;
  assign n45685 = ( n45681 & ~n45683 ) | ( n45681 & n45684 ) | ( ~n45683 & n45684 ) ;
  assign n45686 = ~x1128 & n44180 ;
  assign n45687 = x962 | n45686 ;
  assign n45688 = n44180 & ~n45687 ;
  assign n45689 = ( x732 & n45687 ) | ( x732 & ~n45688 ) | ( n45687 & ~n45688 ) ;
  assign n45690 = x737 & x1135 ;
  assign n45691 = x1134 & ~n45690 ;
  assign n45692 = x838 | x1136 ;
  assign n45693 = ( n45180 & n45691 ) | ( n45180 & n45692 ) | ( n45691 & n45692 ) ;
  assign n45694 = ~n45180 & n45693 ;
  assign n45695 = ( x777 & n44375 ) | ( x777 & ~n45694 ) | ( n44375 & ~n45694 ) ;
  assign n45696 = n45695 ^ n45694 ^ 1'b0 ;
  assign n45697 = ( n45694 & ~n45695 ) | ( n45694 & n45696 ) | ( ~n45695 & n45696 ) ;
  assign n45698 = x619 | x1135 ;
  assign n45699 = ~x648 & x1135 ;
  assign n45700 = ( x1134 & n45698 ) | ( x1134 & ~n45699 ) | ( n45698 & ~n45699 ) ;
  assign n45701 = ~x1134 & n45700 ;
  assign n45702 = n44572 & n45701 ;
  assign n45703 = ( n10841 & n45697 ) | ( n10841 & ~n45702 ) | ( n45697 & ~n45702 ) ;
  assign n45704 = ~n45697 & n45703 ;
  assign n45705 = x316 & ~n44352 ;
  assign n45706 = n44347 & n45705 ;
  assign n45707 = x399 & x591 ;
  assign n45708 = ~n45198 & n45707 ;
  assign n45709 = x375 & n45201 ;
  assign n45710 = ( ~x590 & n45708 ) | ( ~x590 & n45709 ) | ( n45708 & n45709 ) ;
  assign n45711 = ~x590 & n45710 ;
  assign n45712 = ( ~x588 & n45706 ) | ( ~x588 & n45711 ) | ( n45706 & n45711 ) ;
  assign n45713 = ~x588 & n45712 ;
  assign n45714 = x424 & n44957 ;
  assign n45715 = ~n45207 & n45714 ;
  assign n45716 = x199 & ~x1047 ;
  assign n45717 = n44352 & ~n45716 ;
  assign n45718 = x308 ^ x200 ^ 1'b0 ;
  assign n45719 = ( x308 & x1037 ) | ( x308 & n45718 ) | ( x1037 & n45718 ) ;
  assign n45720 = x199 | n45719 ;
  assign n45721 = n45717 & n45720 ;
  assign n45722 = ( n10841 & ~n45715 ) | ( n10841 & n45721 ) | ( ~n45715 & n45721 ) ;
  assign n45723 = n45715 | n45722 ;
  assign n45724 = ( ~n45704 & n45713 ) | ( ~n45704 & n45723 ) | ( n45713 & n45723 ) ;
  assign n45725 = ~n45704 & n45724 ;
  assign n45726 = ~x1119 & n44949 ;
  assign n45727 = x962 | n45726 ;
  assign n45728 = n44949 & ~n45727 ;
  assign n45729 = ( x734 & n45727 ) | ( x734 & ~n45728 ) | ( n45727 & ~n45728 ) ;
  assign n45730 = x735 | n44949 ;
  assign n45731 = ~x1109 & n44949 ;
  assign n45732 = ( x962 & n45730 ) | ( x962 & ~n45731 ) | ( n45730 & ~n45731 ) ;
  assign n45733 = ~x962 & n45732 ;
  assign n45734 = x736 | n44949 ;
  assign n45735 = ~x1101 & n44949 ;
  assign n45736 = ( x962 & n45734 ) | ( x962 & ~n45735 ) | ( n45734 & ~n45735 ) ;
  assign n45737 = ~x962 & n45736 ;
  assign n45738 = ~x1122 & n44949 ;
  assign n45739 = x962 | n45738 ;
  assign n45740 = n44949 & ~n45739 ;
  assign n45741 = ( x737 & n45739 ) | ( x737 & ~n45740 ) | ( n45739 & ~n45740 ) ;
  assign n45742 = ~x1121 & n44949 ;
  assign n45743 = x962 | n45742 ;
  assign n45744 = n44949 & ~n45743 ;
  assign n45745 = ( x738 & n45743 ) | ( x738 & ~n45744 ) | ( n45743 & ~n45744 ) ;
  assign n45746 = x952 | x1061 ;
  assign n45747 = n44071 & ~n45746 ;
  assign n45748 = x832 & n45747 ;
  assign n45749 = x1108 & n45748 ;
  assign n45750 = x966 | n45749 ;
  assign n45751 = n45748 & ~n45750 ;
  assign n45752 = ( x739 & n45750 ) | ( x739 & ~n45751 ) | ( n45750 & ~n45751 ) ;
  assign n45753 = x741 | n45748 ;
  assign n45754 = x1114 & n45748 ;
  assign n45755 = ( x966 & n45753 ) | ( x966 & ~n45754 ) | ( n45753 & ~n45754 ) ;
  assign n45756 = ~x966 & n45755 ;
  assign n45757 = x742 | n45748 ;
  assign n45758 = x1112 & n45748 ;
  assign n45759 = ( x966 & n45757 ) | ( x966 & ~n45758 ) | ( n45757 & ~n45758 ) ;
  assign n45760 = ~x966 & n45759 ;
  assign n45761 = x1109 & n45748 ;
  assign n45762 = x966 | n45761 ;
  assign n45763 = n45748 & ~n45762 ;
  assign n45764 = ( x743 & n45762 ) | ( x743 & ~n45763 ) | ( n45762 & ~n45763 ) ;
  assign n45765 = x1131 & n45748 ;
  assign n45766 = x744 | n45748 ;
  assign n45767 = ( x966 & ~n45765 ) | ( x966 & n45766 ) | ( ~n45765 & n45766 ) ;
  assign n45768 = ~x966 & n45767 ;
  assign n45769 = x745 | n45748 ;
  assign n45770 = x1111 & n45748 ;
  assign n45771 = ( x966 & n45769 ) | ( x966 & ~n45770 ) | ( n45769 & ~n45770 ) ;
  assign n45772 = ~x966 & n45771 ;
  assign n45773 = x1104 & n45748 ;
  assign n45774 = x966 | n45773 ;
  assign n45775 = n45748 & ~n45774 ;
  assign n45776 = ( x746 & n45774 ) | ( x746 & ~n45775 ) | ( n45774 & ~n45775 ) ;
  assign n45777 = x773 & n45581 ;
  assign n45778 = n45777 ^ x747 ^ 1'b0 ;
  assign n45779 = n45595 | n45669 ;
  assign n45780 = n45553 | n45554 ;
  assign n45781 = n45779 | n45780 ;
  assign n45782 = n45781 ^ n45778 ^ 1'b0 ;
  assign n45783 = n45552 | n45777 ;
  assign n45784 = n45556 & ~n45783 ;
  assign n45785 = n45559 & ~n45784 ;
  assign n45786 = ( x801 & n45784 ) | ( x801 & ~n45785 ) | ( n45784 & ~n45785 ) ;
  assign n45787 = ( n45781 & n45782 ) | ( n45781 & ~n45786 ) | ( n45782 & ~n45786 ) ;
  assign n45788 = ( n45778 & ~n45782 ) | ( n45778 & n45787 ) | ( ~n45782 & n45787 ) ;
  assign n45789 = x1106 & n45748 ;
  assign n45790 = x966 | n45789 ;
  assign n45791 = n45748 & ~n45790 ;
  assign n45792 = ( x748 & n45790 ) | ( x748 & ~n45791 ) | ( n45790 & ~n45791 ) ;
  assign n45793 = x1105 & n45748 ;
  assign n45794 = x966 | n45793 ;
  assign n45795 = n45748 & ~n45794 ;
  assign n45796 = ( x749 & n45794 ) | ( x749 & ~n45795 ) | ( n45794 & ~n45795 ) ;
  assign n45797 = x1130 & n45748 ;
  assign n45798 = x750 | n45748 ;
  assign n45799 = ( x966 & ~n45797 ) | ( x966 & n45798 ) | ( ~n45797 & n45798 ) ;
  assign n45800 = ~x966 & n45799 ;
  assign n45801 = x751 | n45748 ;
  assign n45802 = x1123 & n45748 ;
  assign n45803 = ( x966 & n45801 ) | ( x966 & ~n45802 ) | ( n45801 & ~n45802 ) ;
  assign n45804 = ~x966 & n45803 ;
  assign n45805 = x752 | n45748 ;
  assign n45806 = x1124 & n45748 ;
  assign n45807 = ( x966 & n45805 ) | ( x966 & ~n45806 ) | ( n45805 & ~n45806 ) ;
  assign n45808 = ~x966 & n45807 ;
  assign n45809 = x753 | n45748 ;
  assign n45810 = x1117 & n45748 ;
  assign n45811 = ( x966 & n45809 ) | ( x966 & ~n45810 ) | ( n45809 & ~n45810 ) ;
  assign n45812 = ~x966 & n45811 ;
  assign n45813 = x754 | n45748 ;
  assign n45814 = x1118 & n45748 ;
  assign n45815 = ( x966 & n45813 ) | ( x966 & ~n45814 ) | ( n45813 & ~n45814 ) ;
  assign n45816 = ~x966 & n45815 ;
  assign n45817 = x755 | n45748 ;
  assign n45818 = x1120 & n45748 ;
  assign n45819 = ( x966 & n45817 ) | ( x966 & ~n45818 ) | ( n45817 & ~n45818 ) ;
  assign n45820 = ~x966 & n45819 ;
  assign n45821 = x756 | n45748 ;
  assign n45822 = x1119 & n45748 ;
  assign n45823 = ( x966 & n45821 ) | ( x966 & ~n45822 ) | ( n45821 & ~n45822 ) ;
  assign n45824 = ~x966 & n45823 ;
  assign n45825 = x757 | n45748 ;
  assign n45826 = x1113 & n45748 ;
  assign n45827 = ( x966 & n45825 ) | ( x966 & ~n45826 ) | ( n45825 & ~n45826 ) ;
  assign n45828 = ~x966 & n45827 ;
  assign n45829 = x1101 & n45748 ;
  assign n45830 = x966 | n45829 ;
  assign n45831 = n45748 & ~n45830 ;
  assign n45832 = ( x758 & n45830 ) | ( x758 & ~n45831 ) | ( n45830 & ~n45831 ) ;
  assign n45833 = x759 | n45748 ;
  assign n45834 = n44078 & n45747 ;
  assign n45835 = ( x966 & n45833 ) | ( x966 & ~n45834 ) | ( n45833 & ~n45834 ) ;
  assign n45836 = n45835 ^ n45833 ^ 1'b0 ;
  assign n45837 = ( x966 & n45835 ) | ( x966 & ~n45836 ) | ( n45835 & ~n45836 ) ;
  assign n45838 = x760 | n45748 ;
  assign n45839 = x1115 & n45748 ;
  assign n45840 = ( x966 & n45838 ) | ( x966 & ~n45839 ) | ( n45838 & ~n45839 ) ;
  assign n45841 = ~x966 & n45840 ;
  assign n45842 = x761 | n45748 ;
  assign n45843 = x1121 & n45748 ;
  assign n45844 = ( x966 & n45842 ) | ( x966 & ~n45843 ) | ( n45842 & ~n45843 ) ;
  assign n45845 = ~x966 & n45844 ;
  assign n45846 = x1129 & n45748 ;
  assign n45847 = x762 | n45748 ;
  assign n45848 = ( x966 & ~n45846 ) | ( x966 & n45847 ) | ( ~n45846 & n45847 ) ;
  assign n45849 = ~x966 & n45848 ;
  assign n45850 = x1103 & n45748 ;
  assign n45851 = x966 | n45850 ;
  assign n45852 = n45748 & ~n45851 ;
  assign n45853 = ( x763 & n45851 ) | ( x763 & ~n45852 ) | ( n45851 & ~n45852 ) ;
  assign n45854 = x1107 & n45748 ;
  assign n45855 = x966 | n45854 ;
  assign n45856 = n45748 & ~n45855 ;
  assign n45857 = ( x764 & n45855 ) | ( x764 & ~n45856 ) | ( n45855 & ~n45856 ) ;
  assign n45858 = n45563 | n45779 ;
  assign n45859 = x765 & n45858 ;
  assign n45860 = n45679 ^ x731 ^ 1'b0 ;
  assign n45861 = x771 & x800 ;
  assign n45862 = x769 & x794 ;
  assign n45863 = ( x765 & ~n45861 ) | ( x765 & n45862 ) | ( ~n45861 & n45862 ) ;
  assign n45864 = n45861 | n45863 ;
  assign n45865 = ( ~n45550 & n45557 ) | ( ~n45550 & n45864 ) | ( n45557 & n45864 ) ;
  assign n45866 = ~n45550 & n45865 ;
  assign n45867 = n45551 | n45866 ;
  assign n45868 = ~n45562 & n45867 ;
  assign n45869 = x721 | n45868 ;
  assign n45870 = ~n45587 & n45869 ;
  assign n45871 = ~n45565 & n45567 ;
  assign n45872 = n45870 & ~n45871 ;
  assign n45873 = n45588 & ~n45677 ;
  assign n45874 = x765 | n45873 ;
  assign n45875 = ( ~x795 & n45872 ) | ( ~x795 & n45874 ) | ( n45872 & n45874 ) ;
  assign n45876 = ~x795 & n45875 ;
  assign n45877 = ( n45679 & ~n45860 ) | ( n45679 & n45876 ) | ( ~n45860 & n45876 ) ;
  assign n45878 = x731 | n45876 ;
  assign n45879 = x795 | n45878 ;
  assign n45880 = n45877 ^ x765 ^ 1'b0 ;
  assign n45881 = ( ~x765 & n45879 ) | ( ~x765 & n45880 ) | ( n45879 & n45880 ) ;
  assign n45882 = ( x765 & n45877 ) | ( x765 & n45881 ) | ( n45877 & n45881 ) ;
  assign n45883 = n45882 ^ x945 ^ 1'b0 ;
  assign n45884 = ( ~n45859 & n45882 ) | ( ~n45859 & n45883 ) | ( n45882 & n45883 ) ;
  assign n45885 = x1110 & n45748 ;
  assign n45886 = x966 | n45885 ;
  assign n45887 = n45748 & ~n45886 ;
  assign n45888 = ( x766 & n45886 ) | ( x766 & ~n45887 ) | ( n45886 & ~n45887 ) ;
  assign n45889 = x767 | n45748 ;
  assign n45890 = x1116 & n45748 ;
  assign n45891 = ( x966 & n45889 ) | ( x966 & ~n45890 ) | ( n45889 & ~n45890 ) ;
  assign n45892 = ~x966 & n45891 ;
  assign n45893 = x768 | n45748 ;
  assign n45894 = x1125 & n45748 ;
  assign n45895 = ( x966 & n45893 ) | ( x966 & ~n45894 ) | ( n45893 & ~n45894 ) ;
  assign n45896 = ~x966 & n45895 ;
  assign n45897 = x769 & ~n45582 ;
  assign n45898 = x775 & n45574 ;
  assign n45899 = n45898 ^ x769 ^ 1'b0 ;
  assign n45900 = x794 & ~n45552 ;
  assign n45901 = ~n45553 & n45900 ;
  assign n45902 = ( n45560 & ~n45669 ) | ( n45560 & n45901 ) | ( ~n45669 & n45901 ) ;
  assign n45903 = ~n45560 & n45902 ;
  assign n45904 = ~x775 & n45903 ;
  assign n45905 = n45873 | n45904 ;
  assign n45906 = x795 & n45905 ;
  assign n45907 = n45582 & ~n45906 ;
  assign n45908 = n45899 & n45907 ;
  assign n45909 = ~n45595 & n45903 ;
  assign n45910 = ~n45908 & n45909 ;
  assign n45911 = ( n45897 & n45908 ) | ( n45897 & ~n45910 ) | ( n45908 & ~n45910 ) ;
  assign n45912 = x770 | n45748 ;
  assign n45913 = x1126 & n45748 ;
  assign n45914 = ( x966 & n45912 ) | ( x966 & ~n45913 ) | ( n45912 & ~n45913 ) ;
  assign n45915 = ~x966 & n45914 ;
  assign n45916 = x771 & x945 ;
  assign n45917 = n45858 & n45916 ;
  assign n45918 = n45588 | n45870 ;
  assign n45919 = ~n45593 & n45918 ;
  assign n45920 = ( ~n45589 & n45594 ) | ( ~n45589 & n45919 ) | ( n45594 & n45919 ) ;
  assign n45921 = ( n45563 & ~n45668 ) | ( n45563 & n45920 ) | ( ~n45668 & n45920 ) ;
  assign n45922 = ~n45563 & n45921 ;
  assign n45923 = ~x945 & x987 ;
  assign n45924 = ( n45917 & ~n45922 ) | ( n45917 & n45923 ) | ( ~n45922 & n45923 ) ;
  assign n45925 = n45922 ^ n45917 ^ 1'b0 ;
  assign n45926 = ( n45917 & n45924 ) | ( n45917 & ~n45925 ) | ( n45924 & ~n45925 ) ;
  assign n45927 = x1102 & n45748 ;
  assign n45928 = x966 | n45927 ;
  assign n45929 = n45748 & ~n45928 ;
  assign n45930 = ( x772 & n45928 ) | ( x772 & ~n45929 ) | ( n45928 & ~n45929 ) ;
  assign n45931 = x801 | n45562 ;
  assign n45932 = n45922 & ~n45931 ;
  assign n45933 = n45581 & ~n45932 ;
  assign n45934 = ( n45563 & n45858 ) | ( n45563 & n45931 ) | ( n45858 & n45931 ) ;
  assign n45935 = x773 & n45934 ;
  assign n45936 = ( ~n45777 & n45933 ) | ( ~n45777 & n45935 ) | ( n45933 & n45935 ) ;
  assign n45937 = ~n45777 & n45936 ;
  assign n45938 = x774 | n45748 ;
  assign n45939 = x1127 & n45748 ;
  assign n45940 = ( x966 & n45938 ) | ( x966 & ~n45939 ) | ( n45938 & ~n45939 ) ;
  assign n45941 = ~x966 & n45940 ;
  assign n45942 = x775 & n45858 ;
  assign n45943 = x731 & ~x945 ;
  assign n45944 = n45943 ^ n45942 ^ 1'b0 ;
  assign n45945 = x765 & x771 ;
  assign n45946 = n45574 & n45945 ;
  assign n45947 = x795 & x800 ;
  assign n45948 = x801 & ~x816 ;
  assign n45949 = n45947 & n45948 ;
  assign n45950 = ( n45561 & ~n45668 ) | ( n45561 & n45949 ) | ( ~n45668 & n45949 ) ;
  assign n45951 = ~n45561 & n45950 ;
  assign n45952 = ( x775 & n45946 ) | ( x775 & ~n45951 ) | ( n45946 & ~n45951 ) ;
  assign n45953 = n45952 ^ n45946 ^ 1'b0 ;
  assign n45954 = ( x775 & n45952 ) | ( x775 & ~n45953 ) | ( n45952 & ~n45953 ) ;
  assign n45955 = ( n45943 & ~n45944 ) | ( n45943 & n45954 ) | ( ~n45944 & n45954 ) ;
  assign n45956 = ( n45942 & n45944 ) | ( n45942 & n45955 ) | ( n45944 & n45955 ) ;
  assign n45957 = n45679 | n45946 ;
  assign n45958 = x775 & n45943 ;
  assign n45959 = n45956 & ~n45958 ;
  assign n45960 = ( n45956 & ~n45957 ) | ( n45956 & n45959 ) | ( ~n45957 & n45959 ) ;
  assign n45961 = x1128 & n45748 ;
  assign n45962 = x776 | n45748 ;
  assign n45963 = ( x966 & ~n45961 ) | ( x966 & n45962 ) | ( ~n45961 & n45962 ) ;
  assign n45964 = ~x966 & n45963 ;
  assign n45965 = x777 | n45748 ;
  assign n45966 = x1122 & n45748 ;
  assign n45967 = ( x966 & n45965 ) | ( x966 & ~n45966 ) | ( n45965 & ~n45966 ) ;
  assign n45968 = ~x966 & n45967 ;
  assign n45969 = x1046 | x1083 ;
  assign n45970 = x832 & x956 ;
  assign n45971 = ( x1085 & n45969 ) | ( x1085 & n45970 ) | ( n45969 & n45970 ) ;
  assign n45972 = ~n45969 & n45971 ;
  assign n45973 = ~x968 & n45972 ;
  assign n45974 = n45973 ^ x1100 ^ 1'b0 ;
  assign n45975 = ( x778 & x1100 ) | ( x778 & ~n45974 ) | ( x1100 & ~n45974 ) ;
  assign n45976 = x779 & ~n44133 ;
  assign n45977 = x780 & ~n44044 ;
  assign n45978 = n45973 ^ x1101 ^ 1'b0 ;
  assign n45979 = ( x781 & x1101 ) | ( x781 & ~n45978 ) | ( x1101 & ~n45978 ) ;
  assign n45980 = n39971 & ~n44083 ;
  assign n45981 = n44043 & n45980 ;
  assign n45982 = n45973 ^ x1109 ^ 1'b0 ;
  assign n45983 = ( x783 & x1109 ) | ( x783 & ~n45982 ) | ( x1109 & ~n45982 ) ;
  assign n45984 = n45973 ^ x1110 ^ 1'b0 ;
  assign n45985 = ( x784 & x1110 ) | ( x784 & ~n45984 ) | ( x1110 & ~n45984 ) ;
  assign n45986 = n45973 ^ x1102 ^ 1'b0 ;
  assign n45987 = ( x785 & x1102 ) | ( x785 & ~n45986 ) | ( x1102 & ~n45986 ) ;
  assign n45988 = ( x24 & x786 ) | ( x24 & n6306 ) | ( x786 & n6306 ) ;
  assign n45989 = n45973 ^ x1104 ^ 1'b0 ;
  assign n45990 = ( x787 & x1104 ) | ( x787 & ~n45989 ) | ( x1104 & ~n45989 ) ;
  assign n45991 = n45973 ^ x1105 ^ 1'b0 ;
  assign n45992 = ( x788 & x1105 ) | ( x788 & ~n45991 ) | ( x1105 & ~n45991 ) ;
  assign n45993 = n45973 ^ x1106 ^ 1'b0 ;
  assign n45994 = ( x789 & x1106 ) | ( x789 & ~n45993 ) | ( x1106 & ~n45993 ) ;
  assign n45995 = n45973 ^ x1107 ^ 1'b0 ;
  assign n45996 = ( x790 & x1107 ) | ( x790 & ~n45995 ) | ( x1107 & ~n45995 ) ;
  assign n45997 = n45973 ^ x1108 ^ 1'b0 ;
  assign n45998 = ( x791 & x1108 ) | ( x791 & ~n45997 ) | ( x1108 & ~n45997 ) ;
  assign n45999 = n45973 ^ x1103 ^ 1'b0 ;
  assign n46000 = ( x792 & x1103 ) | ( x792 & ~n45999 ) | ( x1103 & ~n45999 ) ;
  assign n46001 = x968 & n45972 ;
  assign n46002 = n46001 ^ x1130 ^ 1'b0 ;
  assign n46003 = ( x794 & x1130 ) | ( x794 & ~n46002 ) | ( x1130 & ~n46002 ) ;
  assign n46004 = n46001 ^ x1128 ^ 1'b0 ;
  assign n46005 = ( x795 & x1128 ) | ( x795 & ~n46004 ) | ( x1128 & ~n46004 ) ;
  assign n46006 = x266 & ~x269 ;
  assign n46007 = x278 & x279 ;
  assign n46008 = ( x280 & n46006 ) | ( x280 & n46007 ) | ( n46006 & n46007 ) ;
  assign n46009 = ~x280 & n46008 ;
  assign n46010 = ~x281 & n46009 ;
  assign n46011 = ~n44322 & n46010 ;
  assign n46012 = n46011 ^ x264 ^ 1'b0 ;
  assign n46013 = n46001 ^ x1124 ^ 1'b0 ;
  assign n46014 = ( x798 & x1124 ) | ( x798 & ~n46013 ) | ( x1124 & ~n46013 ) ;
  assign n46015 = n46001 ^ x1107 ^ 1'b0 ;
  assign n46016 = ( x799 & ~x1107 ) | ( x799 & n46015 ) | ( ~x1107 & n46015 ) ;
  assign n46017 = n46001 ^ x1125 ^ 1'b0 ;
  assign n46018 = ( x800 & x1125 ) | ( x800 & ~n46017 ) | ( x1125 & ~n46017 ) ;
  assign n46019 = n46001 ^ x1126 ^ 1'b0 ;
  assign n46020 = ( x801 & x1126 ) | ( x801 & ~n46019 ) | ( x1126 & ~n46019 ) ;
  assign n46021 = ~x274 & n44325 ;
  assign n46022 = n46001 ^ x1106 ^ 1'b0 ;
  assign n46023 = ( x803 & ~x1106 ) | ( x803 & n46022 ) | ( ~x1106 & n46022 ) ;
  assign n46024 = n46001 ^ x1109 ^ 1'b0 ;
  assign n46025 = ( x804 & x1109 ) | ( x804 & ~n46024 ) | ( x1109 & ~n46024 ) ;
  assign n46026 = ~x282 & n44320 ;
  assign n46027 = n46026 ^ x270 ^ 1'b0 ;
  assign n46028 = n46001 ^ x1127 ^ 1'b0 ;
  assign n46029 = ( x807 & x1127 ) | ( x807 & ~n46028 ) | ( x1127 & ~n46028 ) ;
  assign n46030 = n46001 ^ x1101 ^ 1'b0 ;
  assign n46031 = ( x808 & x1101 ) | ( x808 & ~n46030 ) | ( x1101 & ~n46030 ) ;
  assign n46032 = n46001 ^ x1103 ^ 1'b0 ;
  assign n46033 = ( x809 & ~x1103 ) | ( x809 & n46032 ) | ( ~x1103 & n46032 ) ;
  assign n46034 = n46001 ^ x1108 ^ 1'b0 ;
  assign n46035 = ( x810 & x1108 ) | ( x810 & ~n46034 ) | ( x1108 & ~n46034 ) ;
  assign n46036 = n46001 ^ x1102 ^ 1'b0 ;
  assign n46037 = ( x811 & x1102 ) | ( x811 & ~n46036 ) | ( x1102 & ~n46036 ) ;
  assign n46038 = n46001 ^ x1104 ^ 1'b0 ;
  assign n46039 = ( x812 & ~x1104 ) | ( x812 & n46038 ) | ( ~x1104 & n46038 ) ;
  assign n46040 = n46001 ^ x1131 ^ 1'b0 ;
  assign n46041 = ( x813 & x1131 ) | ( x813 & ~n46040 ) | ( x1131 & ~n46040 ) ;
  assign n46042 = n46001 ^ x1105 ^ 1'b0 ;
  assign n46043 = ( x814 & ~x1105 ) | ( x814 & n46042 ) | ( ~x1105 & n46042 ) ;
  assign n46044 = n46001 ^ x1110 ^ 1'b0 ;
  assign n46045 = ( x815 & x1110 ) | ( x815 & ~n46044 ) | ( x1110 & ~n46044 ) ;
  assign n46046 = n46001 ^ x1129 ^ 1'b0 ;
  assign n46047 = ( x816 & x1129 ) | ( x816 & ~n46046 ) | ( x1129 & ~n46046 ) ;
  assign n46048 = n44318 ^ x269 ^ 1'b0 ;
  assign n46049 = ~n10841 & n12746 ;
  assign n46050 = n12545 | n46049 ;
  assign n46051 = n44324 ^ x265 ^ 1'b0 ;
  assign n46052 = ~x270 & n46026 ;
  assign n46053 = x277 & ~n46052 ;
  assign n46054 = n44323 | n46053 ;
  assign n46055 = x811 | x893 ;
  assign n46056 = n6489 & ~n10841 ;
  assign n46057 = x982 | n8671 ;
  assign n46058 = n5020 & ~n46057 ;
  assign n46059 = ( n5020 & n46056 ) | ( n5020 & n46058 ) | ( n46056 & n46058 ) ;
  assign n46060 = x1126 ^ x1125 ^ 1'b0 ;
  assign n46061 = n46060 ^ x1129 ^ x1128 ;
  assign n46062 = n46061 ^ x1130 ^ x1124 ;
  assign n46063 = x123 & ~n1360 ;
  assign n46064 = x1127 & ~n46063 ;
  assign n46065 = x1131 & n46064 ;
  assign n46066 = ~n46062 & n46065 ;
  assign n46068 = x1127 | x1131 ;
  assign n46069 = ~n46063 & n46068 ;
  assign n46067 = x825 & n46063 ;
  assign n46070 = n46069 ^ n46067 ^ n46063 ;
  assign n46071 = ( n46062 & ~n46066 ) | ( n46062 & n46070 ) | ( ~n46066 & n46070 ) ;
  assign n46072 = n46067 | n46069 ;
  assign n46073 = n46062 & ~n46065 ;
  assign n46074 = n46071 & ~n46073 ;
  assign n46075 = ( n46071 & ~n46072 ) | ( n46071 & n46074 ) | ( ~n46072 & n46074 ) ;
  assign n46076 = x1117 ^ x1116 ^ 1'b0 ;
  assign n46077 = n46076 ^ x1121 ^ x1120 ;
  assign n46078 = n46077 ^ x1119 ^ x1118 ;
  assign n46079 = x1122 & ~n46063 ;
  assign n46080 = x1123 & n46079 ;
  assign n46081 = ~n46078 & n46080 ;
  assign n46083 = x1122 | x1123 ;
  assign n46084 = ~n46063 & n46083 ;
  assign n46082 = x826 & n46063 ;
  assign n46085 = n46084 ^ n46082 ^ n46063 ;
  assign n46086 = ( n46078 & ~n46081 ) | ( n46078 & n46085 ) | ( ~n46081 & n46085 ) ;
  assign n46087 = n46082 | n46084 ;
  assign n46088 = n46078 & ~n46080 ;
  assign n46089 = n46086 & ~n46088 ;
  assign n46090 = ( n46086 & ~n46087 ) | ( n46086 & n46089 ) | ( ~n46087 & n46089 ) ;
  assign n46091 = x1106 ^ x1104 ^ 1'b0 ;
  assign n46092 = n46091 ^ x1102 ^ x1101 ;
  assign n46093 = n46092 ^ x1105 ^ x1103 ;
  assign n46094 = x1107 & ~n46063 ;
  assign n46095 = x1100 & n46094 ;
  assign n46096 = ~n46093 & n46095 ;
  assign n46098 = x1100 | x1107 ;
  assign n46099 = ~n46063 & n46098 ;
  assign n46097 = x827 & n46063 ;
  assign n46100 = n46099 ^ n46097 ^ n46063 ;
  assign n46101 = ( n46093 & ~n46096 ) | ( n46093 & n46100 ) | ( ~n46096 & n46100 ) ;
  assign n46102 = n46097 | n46099 ;
  assign n46103 = n46093 & ~n46095 ;
  assign n46104 = n46101 & ~n46103 ;
  assign n46105 = ( n46101 & ~n46102 ) | ( n46101 & n46104 ) | ( ~n46102 & n46104 ) ;
  assign n46106 = x1109 ^ x1108 ^ 1'b0 ;
  assign n46107 = n46106 ^ x1113 ^ x1112 ;
  assign n46108 = n46107 ^ x1111 ^ x1110 ;
  assign n46109 = x1114 & ~n46063 ;
  assign n46110 = x1115 & n46109 ;
  assign n46111 = ~n46108 & n46110 ;
  assign n46113 = x1114 | x1115 ;
  assign n46114 = ~n46063 & n46113 ;
  assign n46112 = x828 & n46063 ;
  assign n46115 = n46114 ^ n46112 ^ n46063 ;
  assign n46116 = ( n46108 & ~n46111 ) | ( n46108 & n46115 ) | ( ~n46111 & n46115 ) ;
  assign n46117 = n46112 | n46114 ;
  assign n46118 = n46108 & ~n46110 ;
  assign n46119 = n46116 & ~n46118 ;
  assign n46120 = ( n46116 & ~n46117 ) | ( n46116 & n46119 ) | ( ~n46117 & n46119 ) ;
  assign n46121 = n8670 & ~n10841 ;
  assign n46122 = x951 & ~n46121 ;
  assign n46123 = x1092 & ~n46122 ;
  assign n46124 = n46009 ^ x281 ^ 1'b0 ;
  assign n46125 = ~x832 & x1091 ;
  assign n46126 = ( ~x1162 & n7430 ) | ( ~x1162 & n46125 ) | ( n7430 & n46125 ) ;
  assign n46127 = x1162 & n46126 ;
  assign n46128 = x833 & ~n1611 ;
  assign n46129 = n15279 | n46128 ;
  assign n46130 = x946 & n1611 ;
  assign n46131 = n44320 ^ x282 ^ 1'b0 ;
  assign n46132 = x1049 ^ x955 ^ 1'b0 ;
  assign n46133 = ( x837 & x1049 ) | ( x837 & n46132 ) | ( x1049 & n46132 ) ;
  assign n46134 = x1047 ^ x955 ^ 1'b0 ;
  assign n46135 = ( x838 & x1047 ) | ( x838 & n46134 ) | ( x1047 & n46134 ) ;
  assign n46136 = x1074 ^ x955 ^ 1'b0 ;
  assign n46137 = ( x839 & x1074 ) | ( x839 & n46136 ) | ( x1074 & n46136 ) ;
  assign n46138 = n1611 ^ x1196 ^ 1'b0 ;
  assign n46139 = ( x840 & x1196 ) | ( x840 & ~n46138 ) | ( x1196 & ~n46138 ) ;
  assign n46140 = x33 | n8263 ;
  assign n46141 = x1035 ^ x955 ^ 1'b0 ;
  assign n46142 = ( x842 & x1035 ) | ( x842 & n46141 ) | ( x1035 & n46141 ) ;
  assign n46143 = x1079 ^ x955 ^ 1'b0 ;
  assign n46144 = ( x843 & x1079 ) | ( x843 & n46143 ) | ( x1079 & n46143 ) ;
  assign n46145 = x1078 ^ x955 ^ 1'b0 ;
  assign n46146 = ( x844 & x1078 ) | ( x844 & n46145 ) | ( x1078 & n46145 ) ;
  assign n46147 = x1043 ^ x955 ^ 1'b0 ;
  assign n46148 = ( x845 & x1043 ) | ( x845 & n46147 ) | ( x1043 & n46147 ) ;
  assign n46149 = n40529 ^ x1134 ^ 1'b0 ;
  assign n46150 = ( x846 & x1134 ) | ( x846 & ~n46149 ) | ( x1134 & ~n46149 ) ;
  assign n46151 = x1055 ^ x955 ^ 1'b0 ;
  assign n46152 = ( x847 & x1055 ) | ( x847 & n46151 ) | ( x1055 & n46151 ) ;
  assign n46153 = x1039 ^ x955 ^ 1'b0 ;
  assign n46154 = ( x848 & x1039 ) | ( x848 & n46153 ) | ( x1039 & n46153 ) ;
  assign n46155 = n1611 ^ x1198 ^ 1'b0 ;
  assign n46156 = ( x849 & x1198 ) | ( x849 & ~n46155 ) | ( x1198 & ~n46155 ) ;
  assign n46157 = x1048 ^ x955 ^ 1'b0 ;
  assign n46158 = ( x850 & x1048 ) | ( x850 & n46157 ) | ( x1048 & n46157 ) ;
  assign n46159 = x1045 ^ x955 ^ 1'b0 ;
  assign n46160 = ( x851 & x1045 ) | ( x851 & n46159 ) | ( x1045 & n46159 ) ;
  assign n46161 = x1062 ^ x955 ^ 1'b0 ;
  assign n46162 = ( x852 & x1062 ) | ( x852 & n46161 ) | ( x1062 & n46161 ) ;
  assign n46163 = x1080 ^ x955 ^ 1'b0 ;
  assign n46164 = ( x853 & x1080 ) | ( x853 & n46163 ) | ( x1080 & n46163 ) ;
  assign n46165 = x1051 ^ x955 ^ 1'b0 ;
  assign n46166 = ( x854 & x1051 ) | ( x854 & n46165 ) | ( x1051 & n46165 ) ;
  assign n46167 = x1065 ^ x955 ^ 1'b0 ;
  assign n46168 = ( x855 & x1065 ) | ( x855 & n46167 ) | ( x1065 & n46167 ) ;
  assign n46169 = x1067 ^ x955 ^ 1'b0 ;
  assign n46170 = ( x856 & x1067 ) | ( x856 & n46169 ) | ( x1067 & n46169 ) ;
  assign n46171 = x1058 ^ x955 ^ 1'b0 ;
  assign n46172 = ( x857 & x1058 ) | ( x857 & n46171 ) | ( x1058 & n46171 ) ;
  assign n46173 = x1087 ^ x955 ^ 1'b0 ;
  assign n46174 = ( x858 & x1087 ) | ( x858 & n46173 ) | ( x1087 & n46173 ) ;
  assign n46175 = x1070 ^ x955 ^ 1'b0 ;
  assign n46176 = ( x859 & x1070 ) | ( x859 & n46175 ) | ( x1070 & n46175 ) ;
  assign n46177 = x1076 ^ x955 ^ 1'b0 ;
  assign n46178 = ( x860 & x1076 ) | ( x860 & n46177 ) | ( x1076 & n46177 ) ;
  assign n46179 = x123 | x1141 ;
  assign n46180 = x123 & ~x861 ;
  assign n46181 = x228 & ~n46180 ;
  assign n46182 = n46179 & n46181 ;
  assign n46183 = x1093 ^ x861 ^ 1'b0 ;
  assign n46184 = ( x861 & x1141 ) | ( x861 & n46183 ) | ( x1141 & n46183 ) ;
  assign n46185 = ( ~x228 & n46182 ) | ( ~x228 & n46184 ) | ( n46182 & n46184 ) ;
  assign n46186 = n46182 ^ x228 ^ 1'b0 ;
  assign n46187 = ( n46182 & n46185 ) | ( n46182 & ~n46186 ) | ( n46185 & ~n46186 ) ;
  assign n46188 = n40529 ^ x1139 ^ 1'b0 ;
  assign n46189 = ( x862 & x1139 ) | ( x862 & ~n46188 ) | ( x1139 & ~n46188 ) ;
  assign n46190 = n1611 ^ x1199 ^ 1'b0 ;
  assign n46191 = ( x863 & x1199 ) | ( x863 & ~n46190 ) | ( x1199 & ~n46190 ) ;
  assign n46192 = n1611 ^ x1197 ^ 1'b0 ;
  assign n46193 = ( x864 & x1197 ) | ( x864 & ~n46192 ) | ( x1197 & ~n46192 ) ;
  assign n46194 = x1040 ^ x955 ^ 1'b0 ;
  assign n46195 = ( x865 & x1040 ) | ( x865 & n46194 ) | ( x1040 & n46194 ) ;
  assign n46196 = x1053 ^ x955 ^ 1'b0 ;
  assign n46197 = ( x866 & x1053 ) | ( x866 & n46196 ) | ( x1053 & n46196 ) ;
  assign n46198 = x1057 ^ x955 ^ 1'b0 ;
  assign n46199 = ( x867 & x1057 ) | ( x867 & n46198 ) | ( x1057 & n46198 ) ;
  assign n46200 = x1063 ^ x955 ^ 1'b0 ;
  assign n46201 = ( x868 & x1063 ) | ( x868 & n46200 ) | ( x1063 & n46200 ) ;
  assign n46202 = x123 | x1140 ;
  assign n46203 = x123 & ~x869 ;
  assign n46204 = x228 & ~n46203 ;
  assign n46205 = n46202 & n46204 ;
  assign n46206 = x1093 ^ x869 ^ 1'b0 ;
  assign n46207 = ( x869 & x1140 ) | ( x869 & n46206 ) | ( x1140 & n46206 ) ;
  assign n46208 = ( ~x228 & n46205 ) | ( ~x228 & n46207 ) | ( n46205 & n46207 ) ;
  assign n46209 = n46205 ^ x228 ^ 1'b0 ;
  assign n46210 = ( n46205 & n46208 ) | ( n46205 & ~n46209 ) | ( n46208 & ~n46209 ) ;
  assign n46211 = x1069 ^ x955 ^ 1'b0 ;
  assign n46212 = ( x870 & x1069 ) | ( x870 & n46211 ) | ( x1069 & n46211 ) ;
  assign n46213 = x1072 ^ x955 ^ 1'b0 ;
  assign n46214 = ( x871 & x1072 ) | ( x871 & n46213 ) | ( x1072 & n46213 ) ;
  assign n46215 = x1084 ^ x955 ^ 1'b0 ;
  assign n46216 = ( x872 & x1084 ) | ( x872 & n46215 ) | ( x1084 & n46215 ) ;
  assign n46217 = x1044 ^ x955 ^ 1'b0 ;
  assign n46218 = ( x873 & x1044 ) | ( x873 & n46217 ) | ( x1044 & n46217 ) ;
  assign n46219 = x1036 ^ x955 ^ 1'b0 ;
  assign n46220 = ( x874 & x1036 ) | ( x874 & n46219 ) | ( x1036 & n46219 ) ;
  assign n46221 = x123 & x875 ;
  assign n46222 = ~x123 & x1136 ;
  assign n46223 = ( x228 & n46221 ) | ( x228 & ~n46222 ) | ( n46221 & ~n46222 ) ;
  assign n46224 = ~n46221 & n46223 ;
  assign n46225 = x1093 ^ x875 ^ 1'b0 ;
  assign n46226 = ( x875 & x1136 ) | ( x875 & n46225 ) | ( x1136 & n46225 ) ;
  assign n46227 = ( x228 & ~n46224 ) | ( x228 & n46226 ) | ( ~n46224 & n46226 ) ;
  assign n46228 = ~n46224 & n46227 ;
  assign n46229 = x1037 ^ x955 ^ 1'b0 ;
  assign n46230 = ( x876 & x1037 ) | ( x876 & n46229 ) | ( x1037 & n46229 ) ;
  assign n46231 = x123 | x1138 ;
  assign n46232 = x123 & ~x877 ;
  assign n46233 = x228 & ~n46232 ;
  assign n46234 = n46231 & n46233 ;
  assign n46235 = x1093 ^ x877 ^ 1'b0 ;
  assign n46236 = ( x877 & x1138 ) | ( x877 & n46235 ) | ( x1138 & n46235 ) ;
  assign n46237 = ( ~x228 & n46234 ) | ( ~x228 & n46236 ) | ( n46234 & n46236 ) ;
  assign n46238 = n46234 ^ x228 ^ 1'b0 ;
  assign n46239 = ( n46234 & n46237 ) | ( n46234 & ~n46238 ) | ( n46237 & ~n46238 ) ;
  assign n46240 = x123 | x1137 ;
  assign n46241 = x123 & ~x878 ;
  assign n46242 = x228 & ~n46241 ;
  assign n46243 = n46240 & n46242 ;
  assign n46244 = x1093 ^ x878 ^ 1'b0 ;
  assign n46245 = ( x878 & x1137 ) | ( x878 & n46244 ) | ( x1137 & n46244 ) ;
  assign n46246 = ( ~x228 & n46243 ) | ( ~x228 & n46245 ) | ( n46243 & n46245 ) ;
  assign n46247 = n46243 ^ x228 ^ 1'b0 ;
  assign n46248 = ( n46243 & n46246 ) | ( n46243 & ~n46247 ) | ( n46246 & ~n46247 ) ;
  assign n46249 = x123 | x1135 ;
  assign n46250 = x123 & ~x879 ;
  assign n46251 = x228 & ~n46250 ;
  assign n46252 = n46249 & n46251 ;
  assign n46253 = x1093 ^ x879 ^ 1'b0 ;
  assign n46254 = ( x879 & x1135 ) | ( x879 & n46253 ) | ( x1135 & n46253 ) ;
  assign n46255 = ( ~x228 & n46252 ) | ( ~x228 & n46254 ) | ( n46252 & n46254 ) ;
  assign n46256 = n46252 ^ x228 ^ 1'b0 ;
  assign n46257 = ( n46252 & n46255 ) | ( n46252 & ~n46256 ) | ( n46255 & ~n46256 ) ;
  assign n46258 = x1081 ^ x955 ^ 1'b0 ;
  assign n46259 = ( x880 & x1081 ) | ( x880 & n46258 ) | ( x1081 & n46258 ) ;
  assign n46260 = x1059 ^ x955 ^ 1'b0 ;
  assign n46261 = ( x881 & x1059 ) | ( x881 & n46260 ) | ( x1059 & n46260 ) ;
  assign n46262 = ~x883 & n46063 ;
  assign n46263 = n46094 | n46262 ;
  assign n46264 = n46063 ^ x884 ^ 1'b0 ;
  assign n46265 = ( ~x884 & x1124 ) | ( ~x884 & n46264 ) | ( x1124 & n46264 ) ;
  assign n46266 = n46063 ^ x885 ^ 1'b0 ;
  assign n46267 = ( ~x885 & x1125 ) | ( ~x885 & n46266 ) | ( x1125 & n46266 ) ;
  assign n46268 = n46063 ^ x886 ^ 1'b0 ;
  assign n46269 = ( ~x886 & x1109 ) | ( ~x886 & n46268 ) | ( x1109 & n46268 ) ;
  assign n46270 = n46063 ^ x887 ^ 1'b0 ;
  assign n46271 = ( ~x887 & x1100 ) | ( ~x887 & n46270 ) | ( x1100 & n46270 ) ;
  assign n46272 = n46063 ^ x888 ^ 1'b0 ;
  assign n46273 = ( ~x888 & x1120 ) | ( ~x888 & n46272 ) | ( x1120 & n46272 ) ;
  assign n46274 = n46063 ^ x889 ^ 1'b0 ;
  assign n46275 = ( ~x889 & x1103 ) | ( ~x889 & n46274 ) | ( x1103 & n46274 ) ;
  assign n46276 = n46063 ^ x890 ^ 1'b0 ;
  assign n46277 = ( ~x890 & x1126 ) | ( ~x890 & n46276 ) | ( x1126 & n46276 ) ;
  assign n46278 = n46063 ^ x891 ^ 1'b0 ;
  assign n46279 = ( ~x891 & x1116 ) | ( ~x891 & n46278 ) | ( x1116 & n46278 ) ;
  assign n46280 = n46063 ^ x892 ^ 1'b0 ;
  assign n46281 = ( ~x892 & x1101 ) | ( ~x892 & n46280 ) | ( x1101 & n46280 ) ;
  assign n46282 = n46063 ^ x894 ^ 1'b0 ;
  assign n46283 = ( ~x894 & x1119 ) | ( ~x894 & n46282 ) | ( x1119 & n46282 ) ;
  assign n46284 = n46063 ^ x895 ^ 1'b0 ;
  assign n46285 = ( ~x895 & x1113 ) | ( ~x895 & n46284 ) | ( x1113 & n46284 ) ;
  assign n46286 = n46063 ^ x896 ^ 1'b0 ;
  assign n46287 = ( ~x896 & x1118 ) | ( ~x896 & n46286 ) | ( x1118 & n46286 ) ;
  assign n46288 = n46063 ^ x898 ^ 1'b0 ;
  assign n46289 = ( ~x898 & x1129 ) | ( ~x898 & n46288 ) | ( x1129 & n46288 ) ;
  assign n46290 = n46063 ^ x899 ^ 1'b0 ;
  assign n46291 = ( ~x899 & x1115 ) | ( ~x899 & n46290 ) | ( x1115 & n46290 ) ;
  assign n46292 = n46063 ^ x900 ^ 1'b0 ;
  assign n46293 = ( ~x900 & x1110 ) | ( ~x900 & n46292 ) | ( x1110 & n46292 ) ;
  assign n46294 = n46063 ^ x902 ^ 1'b0 ;
  assign n46295 = ( ~x902 & x1111 ) | ( ~x902 & n46294 ) | ( x1111 & n46294 ) ;
  assign n46296 = n46063 ^ x903 ^ 1'b0 ;
  assign n46297 = ( ~x903 & x1121 ) | ( ~x903 & n46296 ) | ( x1121 & n46296 ) ;
  assign n46298 = ~x904 & n46063 ;
  assign n46299 = n46064 | n46298 ;
  assign n46300 = n46063 ^ x905 ^ 1'b0 ;
  assign n46301 = ( ~x905 & x1131 ) | ( ~x905 & n46300 ) | ( x1131 & n46300 ) ;
  assign n46302 = n46063 ^ x906 ^ 1'b0 ;
  assign n46303 = ( ~x906 & x1128 ) | ( ~x906 & n46302 ) | ( x1128 & n46302 ) ;
  assign n46304 = x624 | x979 ;
  assign n46305 = ~x598 & x979 ;
  assign n46306 = x782 & ~n46305 ;
  assign n46307 = n46304 & n46306 ;
  assign n46308 = x782 | x907 ;
  assign n46309 = x979 ^ x615 ^ 1'b0 ;
  assign n46310 = ( x604 & ~x615 ) | ( x604 & n46309 ) | ( ~x615 & n46309 ) ;
  assign n46311 = x782 & ~n46310 ;
  assign n46312 = ( n46307 & n46308 ) | ( n46307 & ~n46311 ) | ( n46308 & ~n46311 ) ;
  assign n46313 = ~n46307 & n46312 ;
  assign n46314 = ~x908 & n46063 ;
  assign n46315 = n46079 | n46314 ;
  assign n46316 = n46063 ^ x909 ^ 1'b0 ;
  assign n46317 = ( ~x909 & x1105 ) | ( ~x909 & n46316 ) | ( x1105 & n46316 ) ;
  assign n46318 = n46063 ^ x910 ^ 1'b0 ;
  assign n46319 = ( ~x910 & x1117 ) | ( ~x910 & n46318 ) | ( x1117 & n46318 ) ;
  assign n46320 = n46063 ^ x911 ^ 1'b0 ;
  assign n46321 = ( ~x911 & x1130 ) | ( ~x911 & n46320 ) | ( x1130 & n46320 ) ;
  assign n46322 = ~x912 & n46063 ;
  assign n46323 = n46109 | n46322 ;
  assign n46324 = n46063 ^ x913 ^ 1'b0 ;
  assign n46325 = ( ~x913 & x1106 ) | ( ~x913 & n46324 ) | ( x1106 & n46324 ) ;
  assign n46326 = n44317 ^ x280 ^ 1'b0 ;
  assign n46327 = n46063 ^ x915 ^ 1'b0 ;
  assign n46328 = ( ~x915 & x1108 ) | ( ~x915 & n46327 ) | ( x1108 & n46327 ) ;
  assign n46329 = n46063 ^ x916 ^ 1'b0 ;
  assign n46330 = ( ~x916 & x1123 ) | ( ~x916 & n46329 ) | ( x1123 & n46329 ) ;
  assign n46331 = n46063 ^ x917 ^ 1'b0 ;
  assign n46332 = ( ~x917 & x1112 ) | ( ~x917 & n46331 ) | ( x1112 & n46331 ) ;
  assign n46333 = n46063 ^ x918 ^ 1'b0 ;
  assign n46334 = ( ~x918 & x1104 ) | ( ~x918 & n46333 ) | ( x1104 & n46333 ) ;
  assign n46335 = n46063 ^ x919 ^ 1'b0 ;
  assign n46336 = ( ~x919 & x1102 ) | ( ~x919 & n46335 ) | ( x1102 & n46335 ) ;
  assign n46337 = x1093 ^ x920 ^ 1'b0 ;
  assign n46338 = ( x920 & x1139 ) | ( x920 & n46337 ) | ( x1139 & n46337 ) ;
  assign n46339 = x1093 ^ x921 ^ 1'b0 ;
  assign n46340 = ( x921 & x1140 ) | ( x921 & n46339 ) | ( x1140 & n46339 ) ;
  assign n46341 = x1093 ^ x922 ^ 1'b0 ;
  assign n46342 = ( x922 & x1152 ) | ( x922 & n46341 ) | ( x1152 & n46341 ) ;
  assign n46343 = x1093 ^ x923 ^ 1'b0 ;
  assign n46344 = ( x923 & x1154 ) | ( x923 & n46343 ) | ( x1154 & n46343 ) ;
  assign n46345 = ~x300 & x301 ;
  assign n46346 = x311 & ~x312 ;
  assign n46347 = n46345 & n46346 ;
  assign n46348 = x1093 ^ x925 ^ 1'b0 ;
  assign n46349 = ( x925 & x1155 ) | ( x925 & n46348 ) | ( x1155 & n46348 ) ;
  assign n46350 = x1093 ^ x926 ^ 1'b0 ;
  assign n46351 = ( x926 & x1157 ) | ( x926 & n46350 ) | ( x1157 & n46350 ) ;
  assign n46352 = x1093 ^ x927 ^ 1'b0 ;
  assign n46353 = ( x927 & x1145 ) | ( x927 & n46352 ) | ( x1145 & n46352 ) ;
  assign n46354 = x1093 ^ x928 ^ 1'b0 ;
  assign n46355 = ( x928 & x1136 ) | ( x928 & n46354 ) | ( x1136 & n46354 ) ;
  assign n46356 = x1093 ^ x929 ^ 1'b0 ;
  assign n46357 = ( x929 & x1144 ) | ( x929 & n46356 ) | ( x1144 & n46356 ) ;
  assign n46358 = x1093 ^ x930 ^ 1'b0 ;
  assign n46359 = ( x930 & x1134 ) | ( x930 & n46358 ) | ( x1134 & n46358 ) ;
  assign n46360 = x1093 ^ x931 ^ 1'b0 ;
  assign n46361 = ( x931 & x1150 ) | ( x931 & n46360 ) | ( x1150 & n46360 ) ;
  assign n46362 = x932 & ~x1093 ;
  assign n46363 = n40522 | n46362 ;
  assign n46364 = x1093 ^ x933 ^ 1'b0 ;
  assign n46365 = ( x933 & x1137 ) | ( x933 & n46364 ) | ( x1137 & n46364 ) ;
  assign n46366 = x1093 ^ x934 ^ 1'b0 ;
  assign n46367 = ( x934 & x1147 ) | ( x934 & n46366 ) | ( x1147 & n46366 ) ;
  assign n46368 = x1093 ^ x935 ^ 1'b0 ;
  assign n46369 = ( x935 & x1141 ) | ( x935 & n46368 ) | ( x1141 & n46368 ) ;
  assign n46370 = x1093 ^ x936 ^ 1'b0 ;
  assign n46371 = ( x936 & x1149 ) | ( x936 & n46370 ) | ( x1149 & n46370 ) ;
  assign n46372 = x1093 ^ x937 ^ 1'b0 ;
  assign n46373 = ( x937 & x1148 ) | ( x937 & n46372 ) | ( x1148 & n46372 ) ;
  assign n46374 = x1093 ^ x938 ^ 1'b0 ;
  assign n46375 = ( x938 & x1135 ) | ( x938 & n46374 ) | ( x1135 & n46374 ) ;
  assign n46376 = x1093 ^ x939 ^ 1'b0 ;
  assign n46377 = ( x939 & x1146 ) | ( x939 & n46376 ) | ( x1146 & n46376 ) ;
  assign n46378 = x1093 ^ x940 ^ 1'b0 ;
  assign n46379 = ( x940 & x1138 ) | ( x940 & n46378 ) | ( x1138 & n46378 ) ;
  assign n46380 = x1093 ^ x941 ^ 1'b0 ;
  assign n46381 = ( x941 & x1153 ) | ( x941 & n46380 ) | ( x1153 & n46380 ) ;
  assign n46382 = x1093 ^ x942 ^ 1'b0 ;
  assign n46383 = ( x942 & x1156 ) | ( x942 & n46382 ) | ( x1156 & n46382 ) ;
  assign n46384 = x1093 ^ x943 ^ 1'b0 ;
  assign n46385 = ( x943 & x1151 ) | ( x943 & n46384 ) | ( x1151 & n46384 ) ;
  assign n46386 = x1093 ^ x944 ^ 1'b0 ;
  assign n46387 = ( x944 & x1143 ) | ( x944 & n46386 ) | ( x1143 & n46386 ) ;
  assign n46388 = x230 & n1611 ;
  assign n46389 = ~x782 & x947 ;
  assign n46390 = n46307 | n46389 ;
  assign n46391 = x992 ^ x266 ^ 1'b0 ;
  assign n46392 = ( x313 & ~x949 ) | ( x313 & n42288 ) | ( ~x949 & n42288 ) ;
  assign n46393 = ~n6489 & n12833 ;
  assign n46394 = x957 & x1092 ;
  assign n46395 = x31 | n46394 ;
  assign n46396 = ~x782 & x960 ;
  assign n46397 = ~x230 & x961 ;
  assign n46398 = ~x782 & x963 ;
  assign n46399 = ~x230 & x967 ;
  assign n46400 = ~x230 & x969 ;
  assign n46401 = ~x782 & x970 ;
  assign n46402 = ~x230 & x971 ;
  assign n46403 = ~x782 & x972 ;
  assign n46404 = ~x230 & x974 ;
  assign n46405 = ~x782 & x975 ;
  assign n46406 = ~x230 & x977 ;
  assign n46407 = ~x782 & x978 ;
  assign n46408 = ~x598 & x615 ;
  assign n46409 = x824 & x1092 ;
  assign n46410 = x604 | x624 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = n2119 ;
  assign y154 = n2359 ;
  assign y155 = n2535 ;
  assign y156 = ~n2779 ;
  assign y157 = ~n3007 ;
  assign y158 = n3239 ;
  assign y159 = n3471 ;
  assign y160 = n3711 ;
  assign y161 = n3944 ;
  assign y162 = n4177 ;
  assign y163 = n4413 ;
  assign y164 = n4650 ;
  assign y165 = n5002 ;
  assign y166 = ~1'b0 ;
  assign y167 = n5191 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n5489 ;
  assign y172 = ~n5622 ;
  assign y173 = ~n5754 ;
  assign y174 = ~n5854 ;
  assign y175 = ~n5953 ;
  assign y176 = ~n6052 ;
  assign y177 = ~n6151 ;
  assign y178 = ~n6247 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = n5191 ;
  assign y182 = n6307 ;
  assign y183 = n6357 ;
  assign y184 = ~n6362 ;
  assign y185 = ~n6364 ;
  assign y186 = ~n6366 ;
  assign y187 = ~n6368 ;
  assign y188 = x37 ;
  assign y189 = n7445 ;
  assign y190 = n7545 ;
  assign y191 = n8269 ;
  assign y192 = n8661 ;
  assign y193 = n8741 ;
  assign y194 = n8763 ;
  assign y195 = n6305 ;
  assign y196 = n8795 ;
  assign y197 = n8880 ;
  assign y198 = n8894 ;
  assign y199 = n9090 ;
  assign y200 = n9342 ;
  assign y201 = n9526 ;
  assign y202 = n9603 ;
  assign y203 = n9607 ;
  assign y204 = n9628 ;
  assign y205 = n9676 ;
  assign y206 = n9682 ;
  assign y207 = n9702 ;
  assign y208 = n9730 ;
  assign y209 = n9738 ;
  assign y210 = n9894 ;
  assign y211 = n9907 ;
  assign y212 = n9928 ;
  assign y213 = n9942 ;
  assign y214 = n9950 ;
  assign y215 = n9961 ;
  assign y216 = n9964 ;
  assign y217 = n9969 ;
  assign y218 = n9978 ;
  assign y219 = n9982 ;
  assign y220 = n9986 ;
  assign y221 = n9992 ;
  assign y222 = n10003 ;
  assign y223 = n10007 ;
  assign y224 = n10024 ;
  assign y225 = n10029 ;
  assign y226 = n10038 ;
  assign y227 = n10051 ;
  assign y228 = n10072 ;
  assign y229 = n10094 ;
  assign y230 = n10111 ;
  assign y231 = n10123 ;
  assign y232 = n10137 ;
  assign y233 = n10149 ;
  assign y234 = n10308 ;
  assign y235 = n10319 ;
  assign y236 = n10321 ;
  assign y237 = n10840 ;
  assign y238 = n11515 ;
  assign y239 = n11525 ;
  assign y240 = n11534 ;
  assign y241 = n11548 ;
  assign y242 = n11554 ;
  assign y243 = n11559 ;
  assign y244 = n11564 ;
  assign y245 = n11568 ;
  assign y246 = n11589 ;
  assign y247 = n11600 ;
  assign y248 = n11605 ;
  assign y249 = n11617 ;
  assign y250 = n11629 ;
  assign y251 = n11636 ;
  assign y252 = n11654 ;
  assign y253 = n11670 ;
  assign y254 = n11681 ;
  assign y255 = n11691 ;
  assign y256 = n11696 ;
  assign y257 = n11780 ;
  assign y258 = n11797 ;
  assign y259 = n11877 ;
  assign y260 = n11880 ;
  assign y261 = n11888 ;
  assign y262 = n11909 ;
  assign y263 = x117 ;
  assign y264 = n11920 ;
  assign y265 = n11922 ;
  assign y266 = n11940 ;
  assign y267 = n11942 ;
  assign y268 = n11953 ;
  assign y269 = n11959 ;
  assign y270 = ~n11960 ;
  assign y271 = n12010 ;
  assign y272 = n12052 ;
  assign y273 = n12094 ;
  assign y274 = n12145 ;
  assign y275 = n12165 ;
  assign y276 = n12485 ;
  assign y277 = n12543 ;
  assign y278 = n12958 ;
  assign y279 = n13386 ;
  assign y280 = n13394 ;
  assign y281 = ~n13453 ;
  assign y282 = n13871 ;
  assign y283 = n14194 ;
  assign y284 = n14289 ;
  assign y285 = x131 ;
  assign y286 = n14313 ;
  assign y287 = n14447 ;
  assign y288 = n14457 ;
  assign y289 = n14682 ;
  assign y290 = n14748 ;
  assign y291 = n14869 ;
  assign y292 = n15001 ;
  assign y293 = n15093 ;
  assign y294 = n15109 ;
  assign y295 = n15195 ;
  assign y296 = n15254 ;
  assign y297 = ~n16609 ;
  assign y298 = ~n17078 ;
  assign y299 = n17836 ;
  assign y300 = ~n18305 ;
  assign y301 = n18813 ;
  assign y302 = ~n19253 ;
  assign y303 = n19337 ;
  assign y304 = ~n19476 ;
  assign y305 = ~n19540 ;
  assign y306 = ~n19602 ;
  assign y307 = ~n19663 ;
  assign y308 = ~n19748 ;
  assign y309 = n19855 ;
  assign y310 = ~n19940 ;
  assign y311 = ~n19993 ;
  assign y312 = ~n20032 ;
  assign y313 = ~n20066 ;
  assign y314 = ~n20126 ;
  assign y315 = ~n20187 ;
  assign y316 = ~n20248 ;
  assign y317 = ~n20310 ;
  assign y318 = n20404 ;
  assign y319 = ~n20462 ;
  assign y320 = ~n20523 ;
  assign y321 = ~n20563 ;
  assign y322 = ~n20603 ;
  assign y323 = n20701 ;
  assign y324 = ~n20743 ;
  assign y325 = ~n20827 ;
  assign y326 = ~n20911 ;
  assign y327 = ~n20992 ;
  assign y328 = ~n21076 ;
  assign y329 = ~n21160 ;
  assign y330 = ~n21595 ;
  assign y331 = n22068 ;
  assign y332 = ~n22519 ;
  assign y333 = ~n22927 ;
  assign y334 = ~n23367 ;
  assign y335 = ~n23800 ;
  assign y336 = ~n24237 ;
  assign y337 = ~n24679 ;
  assign y338 = ~n25121 ;
  assign y339 = ~n25554 ;
  assign y340 = ~n25987 ;
  assign y341 = ~n26420 ;
  assign y342 = ~n26862 ;
  assign y343 = ~n27292 ;
  assign y344 = ~n27725 ;
  assign y345 = ~n28155 ;
  assign y346 = n28624 ;
  assign y347 = ~n29071 ;
  assign y348 = ~n29518 ;
  assign y349 = ~n29965 ;
  assign y350 = ~n30398 ;
  assign y351 = ~n30818 ;
  assign y352 = n30876 ;
  assign y353 = n30953 ;
  assign y354 = ~n31017 ;
  assign y355 = n31646 ;
  assign y356 = n31914 ;
  assign y357 = n32177 ;
  assign y358 = ~n32362 ;
  assign y359 = ~n32368 ;
  assign y360 = ~n32374 ;
  assign y361 = ~n32482 ;
  assign y362 = ~n32487 ;
  assign y363 = ~n32493 ;
  assign y364 = ~n32961 ;
  assign y365 = ~n33029 ;
  assign y366 = ~n33179 ;
  assign y367 = n33306 ;
  assign y368 = n33334 ;
  assign y369 = ~n33357 ;
  assign y370 = ~n33379 ;
  assign y371 = ~n33402 ;
  assign y372 = n33524 ;
  assign y373 = n33639 ;
  assign y374 = ~n33658 ;
  assign y375 = ~n33663 ;
  assign y376 = n33686 ;
  assign y377 = ~n33691 ;
  assign y378 = n33800 ;
  assign y379 = n34421 ;
  assign y380 = n35004 ;
  assign y381 = n35578 ;
  assign y382 = n35700 ;
  assign y383 = n35755 ;
  assign y384 = ~n35791 ;
  assign y385 = n35805 ;
  assign y386 = x232 ;
  assign y387 = n35896 ;
  assign y388 = x236 ;
  assign y389 = n35959 ;
  assign y390 = ~n36385 ;
  assign y391 = n36709 ;
  assign y392 = n36916 ;
  assign y393 = n36934 ;
  assign y394 = ~n37192 ;
  assign y395 = n37532 ;
  assign y396 = n37630 ;
  assign y397 = n38064 ;
  assign y398 = n38364 ;
  assign y399 = n38457 ;
  assign y400 = ~n38769 ;
  assign y401 = n38822 ;
  assign y402 = n39066 ;
  assign y403 = n39348 ;
  assign y404 = n39590 ;
  assign y405 = n39751 ;
  assign y406 = n39951 ;
  assign y407 = n39960 ;
  assign y408 = n39969 ;
  assign y409 = n40009 ;
  assign y410 = n40253 ;
  assign y411 = n40485 ;
  assign y412 = n40489 ;
  assign y413 = n40493 ;
  assign y414 = n40497 ;
  assign y415 = n40501 ;
  assign y416 = n40505 ;
  assign y417 = n40511 ;
  assign y418 = n40517 ;
  assign y419 = ~n40551 ;
  assign y420 = ~n40765 ;
  assign y421 = ~n40812 ;
  assign y422 = ~n40853 ;
  assign y423 = n40920 ;
  assign y424 = n41140 ;
  assign y425 = n41306 ;
  assign y426 = ~n41354 ;
  assign y427 = ~n41397 ;
  assign y428 = n41442 ;
  assign y429 = n41549 ;
  assign y430 = n41614 ;
  assign y431 = ~n41657 ;
  assign y432 = n41729 ;
  assign y433 = n41761 ;
  assign y434 = ~n41807 ;
  assign y435 = n41872 ;
  assign y436 = n41934 ;
  assign y437 = ~n41977 ;
  assign y438 = ~n42017 ;
  assign y439 = ~n42055 ;
  assign y440 = n42116 ;
  assign y441 = ~n42120 ;
  assign y442 = n42138 ;
  assign y443 = n42156 ;
  assign y444 = ~n42158 ;
  assign y445 = n42164 ;
  assign y446 = n42177 ;
  assign y447 = n42179 ;
  assign y448 = n42181 ;
  assign y449 = n42183 ;
  assign y450 = n42185 ;
  assign y451 = n42187 ;
  assign y452 = n42189 ;
  assign y453 = n42191 ;
  assign y454 = n42193 ;
  assign y455 = n42195 ;
  assign y456 = n42203 ;
  assign y457 = n42210 ;
  assign y458 = ~n42214 ;
  assign y459 = ~n42236 ;
  assign y460 = n42238 ;
  assign y461 = n42240 ;
  assign y462 = n42242 ;
  assign y463 = n42244 ;
  assign y464 = n42246 ;
  assign y465 = n42248 ;
  assign y466 = n42250 ;
  assign y467 = ~n42278 ;
  assign y468 = ~n42281 ;
  assign y469 = n42283 ;
  assign y470 = n42289 ;
  assign y471 = ~n42301 ;
  assign y472 = n42304 ;
  assign y473 = n42306 ;
  assign y474 = n42309 ;
  assign y475 = n42312 ;
  assign y476 = n42314 ;
  assign y477 = n42316 ;
  assign y478 = n42318 ;
  assign y479 = n42320 ;
  assign y480 = n42322 ;
  assign y481 = n42324 ;
  assign y482 = n42326 ;
  assign y483 = n42328 ;
  assign y484 = n42330 ;
  assign y485 = n42332 ;
  assign y486 = n42334 ;
  assign y487 = n42343 ;
  assign y488 = n42350 ;
  assign y489 = n42363 ;
  assign y490 = n42365 ;
  assign y491 = n42367 ;
  assign y492 = n42369 ;
  assign y493 = n42371 ;
  assign y494 = n42373 ;
  assign y495 = n42375 ;
  assign y496 = n42377 ;
  assign y497 = ~n42385 ;
  assign y498 = n42388 ;
  assign y499 = n42390 ;
  assign y500 = n42392 ;
  assign y501 = n42394 ;
  assign y502 = n42396 ;
  assign y503 = n42398 ;
  assign y504 = n42400 ;
  assign y505 = n42402 ;
  assign y506 = n42404 ;
  assign y507 = n42406 ;
  assign y508 = n42408 ;
  assign y509 = n42410 ;
  assign y510 = n42412 ;
  assign y511 = n42414 ;
  assign y512 = n42416 ;
  assign y513 = n42418 ;
  assign y514 = n42420 ;
  assign y515 = n42422 ;
  assign y516 = n42424 ;
  assign y517 = n42426 ;
  assign y518 = n42428 ;
  assign y519 = n42430 ;
  assign y520 = n42432 ;
  assign y521 = n42434 ;
  assign y522 = n42436 ;
  assign y523 = n42438 ;
  assign y524 = n42440 ;
  assign y525 = n42442 ;
  assign y526 = n42444 ;
  assign y527 = n42446 ;
  assign y528 = n42448 ;
  assign y529 = n42450 ;
  assign y530 = n42452 ;
  assign y531 = n42454 ;
  assign y532 = n42456 ;
  assign y533 = n42458 ;
  assign y534 = n42460 ;
  assign y535 = n42462 ;
  assign y536 = n42464 ;
  assign y537 = n42466 ;
  assign y538 = n42468 ;
  assign y539 = n42470 ;
  assign y540 = n42472 ;
  assign y541 = n42474 ;
  assign y542 = n42476 ;
  assign y543 = n42478 ;
  assign y544 = n42480 ;
  assign y545 = n42482 ;
  assign y546 = n42484 ;
  assign y547 = n42486 ;
  assign y548 = n42488 ;
  assign y549 = n42490 ;
  assign y550 = n42492 ;
  assign y551 = n42494 ;
  assign y552 = n42496 ;
  assign y553 = n42498 ;
  assign y554 = n42500 ;
  assign y555 = n42502 ;
  assign y556 = n42504 ;
  assign y557 = n42506 ;
  assign y558 = n42508 ;
  assign y559 = n42510 ;
  assign y560 = n42512 ;
  assign y561 = n42514 ;
  assign y562 = n42516 ;
  assign y563 = n42518 ;
  assign y564 = n42520 ;
  assign y565 = n42522 ;
  assign y566 = n42524 ;
  assign y567 = n42526 ;
  assign y568 = n42528 ;
  assign y569 = n42530 ;
  assign y570 = n42532 ;
  assign y571 = n42535 ;
  assign y572 = n42537 ;
  assign y573 = n42539 ;
  assign y574 = n42541 ;
  assign y575 = n42543 ;
  assign y576 = n42545 ;
  assign y577 = n42547 ;
  assign y578 = n42549 ;
  assign y579 = n42551 ;
  assign y580 = n42553 ;
  assign y581 = n42555 ;
  assign y582 = n42557 ;
  assign y583 = n42559 ;
  assign y584 = n42561 ;
  assign y585 = n42563 ;
  assign y586 = n42565 ;
  assign y587 = n42567 ;
  assign y588 = n42569 ;
  assign y589 = n42571 ;
  assign y590 = n42573 ;
  assign y591 = n42575 ;
  assign y592 = n42577 ;
  assign y593 = n42579 ;
  assign y594 = n42581 ;
  assign y595 = n42583 ;
  assign y596 = n42585 ;
  assign y597 = n42587 ;
  assign y598 = n42589 ;
  assign y599 = n42591 ;
  assign y600 = n42593 ;
  assign y601 = n42595 ;
  assign y602 = n42597 ;
  assign y603 = n42599 ;
  assign y604 = n42601 ;
  assign y605 = n42603 ;
  assign y606 = n42605 ;
  assign y607 = n42607 ;
  assign y608 = n42609 ;
  assign y609 = n42611 ;
  assign y610 = n42613 ;
  assign y611 = n42615 ;
  assign y612 = n42617 ;
  assign y613 = n42619 ;
  assign y614 = n42645 ;
  assign y615 = n42647 ;
  assign y616 = n42649 ;
  assign y617 = n42651 ;
  assign y618 = n42653 ;
  assign y619 = n42655 ;
  assign y620 = n42657 ;
  assign y621 = n42659 ;
  assign y622 = n42684 ;
  assign y623 = n42702 ;
  assign y624 = n42729 ;
  assign y625 = n42734 ;
  assign y626 = n42754 ;
  assign y627 = n42774 ;
  assign y628 = n42794 ;
  assign y629 = n42814 ;
  assign y630 = n42826 ;
  assign y631 = n42838 ;
  assign y632 = n42850 ;
  assign y633 = n42864 ;
  assign y634 = ~n42287 ;
  assign y635 = n42865 ;
  assign y636 = x583 ;
  assign y637 = n42128 ;
  assign y638 = n42867 ;
  assign y639 = n42869 ;
  assign y640 = n42871 ;
  assign y641 = n42873 ;
  assign y642 = n42875 ;
  assign y643 = n42877 ;
  assign y644 = n42879 ;
  assign y645 = ~n42881 ;
  assign y646 = n42883 ;
  assign y647 = n42885 ;
  assign y648 = n42887 ;
  assign y649 = n42889 ;
  assign y650 = n42891 ;
  assign y651 = ~n42893 ;
  assign y652 = n42895 ;
  assign y653 = n42897 ;
  assign y654 = ~n42899 ;
  assign y655 = n42901 ;
  assign y656 = n42903 ;
  assign y657 = n42905 ;
  assign y658 = n42907 ;
  assign y659 = n42909 ;
  assign y660 = n42911 ;
  assign y661 = n42913 ;
  assign y662 = n42922 ;
  assign y663 = n42924 ;
  assign y664 = n42926 ;
  assign y665 = n42928 ;
  assign y666 = n42930 ;
  assign y667 = n42932 ;
  assign y668 = n42938 ;
  assign y669 = n42940 ;
  assign y670 = n42942 ;
  assign y671 = n42944 ;
  assign y672 = n42946 ;
  assign y673 = n42948 ;
  assign y674 = n42950 ;
  assign y675 = n42956 ;
  assign y676 = ~n42958 ;
  assign y677 = n42960 ;
  assign y678 = n42962 ;
  assign y679 = n42964 ;
  assign y680 = n42969 ;
  assign y681 = ~n42971 ;
  assign y682 = n42973 ;
  assign y683 = n42975 ;
  assign y684 = n42977 ;
  assign y685 = n42979 ;
  assign y686 = n42981 ;
  assign y687 = n42983 ;
  assign y688 = n42985 ;
  assign y689 = n42987 ;
  assign y690 = n42989 ;
  assign y691 = ~n42991 ;
  assign y692 = n42993 ;
  assign y693 = n42995 ;
  assign y694 = n42997 ;
  assign y695 = n42999 ;
  assign y696 = n43001 ;
  assign y697 = n43003 ;
  assign y698 = n43005 ;
  assign y699 = n43007 ;
  assign y700 = n43009 ;
  assign y701 = n43014 ;
  assign y702 = n43016 ;
  assign y703 = n43018 ;
  assign y704 = n43020 ;
  assign y705 = n43022 ;
  assign y706 = n43024 ;
  assign y707 = ~n43026 ;
  assign y708 = n43028 ;
  assign y709 = n43030 ;
  assign y710 = n43032 ;
  assign y711 = n43034 ;
  assign y712 = n43036 ;
  assign y713 = n43038 ;
  assign y714 = n43043 ;
  assign y715 = n43045 ;
  assign y716 = n43047 ;
  assign y717 = n43049 ;
  assign y718 = n43051 ;
  assign y719 = n43053 ;
  assign y720 = n43055 ;
  assign y721 = n43057 ;
  assign y722 = n43059 ;
  assign y723 = n43061 ;
  assign y724 = n43177 ;
  assign y725 = n43179 ;
  assign y726 = ~n43181 ;
  assign y727 = n43186 ;
  assign y728 = n43188 ;
  assign y729 = n43190 ;
  assign y730 = n43192 ;
  assign y731 = n43194 ;
  assign y732 = n43196 ;
  assign y733 = n43198 ;
  assign y734 = n43200 ;
  assign y735 = n43202 ;
  assign y736 = n43204 ;
  assign y737 = n43206 ;
  assign y738 = n43208 ;
  assign y739 = n43210 ;
  assign y740 = n5023 ;
  assign y741 = n43212 ;
  assign y742 = n43214 ;
  assign y743 = n43216 ;
  assign y744 = n43224 ;
  assign y745 = n43229 ;
  assign y746 = n43249 ;
  assign y747 = ~n43253 ;
  assign y748 = n43257 ;
  assign y749 = n43261 ;
  assign y750 = n44019 ;
  assign y751 = n44026 ;
  assign y752 = n44032 ;
  assign y753 = n44037 ;
  assign y754 = n44040 ;
  assign y755 = n44046 ;
  assign y756 = n44050 ;
  assign y757 = n44053 ;
  assign y758 = n44057 ;
  assign y759 = n44069 ;
  assign y760 = n44082 ;
  assign y761 = n44088 ;
  assign y762 = ~n44091 ;
  assign y763 = n44095 ;
  assign y764 = n44099 ;
  assign y765 = n44103 ;
  assign y766 = n44107 ;
  assign y767 = n44111 ;
  assign y768 = n44115 ;
  assign y769 = n44119 ;
  assign y770 = n44123 ;
  assign y771 = n44130 ;
  assign y772 = ~n44135 ;
  assign y773 = n44142 ;
  assign y774 = n44146 ;
  assign y775 = n44150 ;
  assign y776 = n44154 ;
  assign y777 = n44158 ;
  assign y778 = n44162 ;
  assign y779 = n44166 ;
  assign y780 = n44170 ;
  assign y781 = n44175 ;
  assign y782 = n44184 ;
  assign y783 = n44188 ;
  assign y784 = n44192 ;
  assign y785 = n44196 ;
  assign y786 = n44200 ;
  assign y787 = n44204 ;
  assign y788 = ~n44208 ;
  assign y789 = ~n44212 ;
  assign y790 = n44216 ;
  assign y791 = n44220 ;
  assign y792 = ~n44224 ;
  assign y793 = n44228 ;
  assign y794 = n44232 ;
  assign y795 = n44236 ;
  assign y796 = n44240 ;
  assign y797 = n44244 ;
  assign y798 = n44248 ;
  assign y799 = n44252 ;
  assign y800 = n44256 ;
  assign y801 = n44260 ;
  assign y802 = n44264 ;
  assign y803 = ~n44268 ;
  assign y804 = n44272 ;
  assign y805 = n44276 ;
  assign y806 = ~n44280 ;
  assign y807 = ~n44284 ;
  assign y808 = n44288 ;
  assign y809 = n44292 ;
  assign y810 = n44296 ;
  assign y811 = ~n44300 ;
  assign y812 = ~n44304 ;
  assign y813 = n44308 ;
  assign y814 = ~n44312 ;
  assign y815 = n44316 ;
  assign y816 = ~n44326 ;
  assign y817 = n44330 ;
  assign y818 = n44334 ;
  assign y819 = n44338 ;
  assign y820 = n44388 ;
  assign y821 = n44432 ;
  assign y822 = n44436 ;
  assign y823 = n44474 ;
  assign y824 = n44513 ;
  assign y825 = n44550 ;
  assign y826 = ~n44554 ;
  assign y827 = n44587 ;
  assign y828 = n44619 ;
  assign y829 = n44656 ;
  assign y830 = n44693 ;
  assign y831 = n44732 ;
  assign y832 = n44770 ;
  assign y833 = n44807 ;
  assign y834 = n44839 ;
  assign y835 = n44871 ;
  assign y836 = n44908 ;
  assign y837 = n44912 ;
  assign y838 = n44916 ;
  assign y839 = n44948 ;
  assign y840 = n7451 ;
  assign y841 = ~n44953 ;
  assign y842 = n44993 ;
  assign y843 = ~n44997 ;
  assign y844 = n45001 ;
  assign y845 = ~n45005 ;
  assign y846 = n45041 ;
  assign y847 = n45045 ;
  assign y848 = n45049 ;
  assign y849 = n45087 ;
  assign y850 = ~n45091 ;
  assign y851 = ~n45095 ;
  assign y852 = ~n45099 ;
  assign y853 = n45103 ;
  assign y854 = ~n45107 ;
  assign y855 = ~n45111 ;
  assign y856 = n45115 ;
  assign y857 = n45119 ;
  assign y858 = ~n45123 ;
  assign y859 = ~n45127 ;
  assign y860 = n45131 ;
  assign y861 = ~n45135 ;
  assign y862 = n45139 ;
  assign y863 = n45143 ;
  assign y864 = n45179 ;
  assign y865 = n45219 ;
  assign y866 = ~n45223 ;
  assign y867 = n45227 ;
  assign y868 = n45259 ;
  assign y869 = n45296 ;
  assign y870 = n45329 ;
  assign y871 = n45367 ;
  assign y872 = n45371 ;
  assign y873 = n45407 ;
  assign y874 = n45441 ;
  assign y875 = n45477 ;
  assign y876 = n45511 ;
  assign y877 = n45549 ;
  assign y878 = n45599 ;
  assign y879 = n45635 ;
  assign y880 = ~n45639 ;
  assign y881 = ~n45643 ;
  assign y882 = ~n45647 ;
  assign y883 = n45651 ;
  assign y884 = n45655 ;
  assign y885 = ~n45659 ;
  assign y886 = n45663 ;
  assign y887 = n45667 ;
  assign y888 = n45685 ;
  assign y889 = ~n45689 ;
  assign y890 = n45725 ;
  assign y891 = ~n45729 ;
  assign y892 = n45733 ;
  assign y893 = n45737 ;
  assign y894 = ~n45741 ;
  assign y895 = ~n45745 ;
  assign y896 = n45752 ;
  assign y897 = n44074 ;
  assign y898 = ~n45756 ;
  assign y899 = ~n45760 ;
  assign y900 = n45764 ;
  assign y901 = ~n45768 ;
  assign y902 = ~n45772 ;
  assign y903 = n45776 ;
  assign y904 = n45788 ;
  assign y905 = n45792 ;
  assign y906 = n45796 ;
  assign y907 = ~n45800 ;
  assign y908 = ~n45804 ;
  assign y909 = ~n45808 ;
  assign y910 = ~n45812 ;
  assign y911 = ~n45816 ;
  assign y912 = ~n45820 ;
  assign y913 = ~n45824 ;
  assign y914 = ~n45828 ;
  assign y915 = n45832 ;
  assign y916 = n45837 ;
  assign y917 = ~n45841 ;
  assign y918 = ~n45845 ;
  assign y919 = ~n45849 ;
  assign y920 = n45853 ;
  assign y921 = n45857 ;
  assign y922 = ~n45884 ;
  assign y923 = n45888 ;
  assign y924 = ~n45892 ;
  assign y925 = ~n45896 ;
  assign y926 = n45911 ;
  assign y927 = ~n45915 ;
  assign y928 = n45926 ;
  assign y929 = n45930 ;
  assign y930 = n45937 ;
  assign y931 = ~n45941 ;
  assign y932 = n45960 ;
  assign y933 = ~n45964 ;
  assign y934 = ~n45968 ;
  assign y935 = n45975 ;
  assign y936 = ~n45976 ;
  assign y937 = ~n45977 ;
  assign y938 = n45979 ;
  assign y939 = ~n45981 ;
  assign y940 = n45983 ;
  assign y941 = n45985 ;
  assign y942 = n45987 ;
  assign y943 = ~n45988 ;
  assign y944 = n45990 ;
  assign y945 = n45992 ;
  assign y946 = n45994 ;
  assign y947 = n45996 ;
  assign y948 = n45998 ;
  assign y949 = n46000 ;
  assign y950 = ~n35897 ;
  assign y951 = n46003 ;
  assign y952 = n46005 ;
  assign y953 = ~n46012 ;
  assign y954 = n44180 ;
  assign y955 = n46014 ;
  assign y956 = ~n46016 ;
  assign y957 = n46018 ;
  assign y958 = n46020 ;
  assign y959 = n46021 ;
  assign y960 = ~n46023 ;
  assign y961 = n46025 ;
  assign y962 = ~n46027 ;
  assign y963 = n45922 ;
  assign y964 = n46029 ;
  assign y965 = n46031 ;
  assign y966 = ~n46033 ;
  assign y967 = n46035 ;
  assign y968 = n46037 ;
  assign y969 = ~n46039 ;
  assign y970 = n46041 ;
  assign y971 = ~n46043 ;
  assign y972 = n46045 ;
  assign y973 = n46047 ;
  assign y974 = ~n46048 ;
  assign y975 = n46050 ;
  assign y976 = ~n46051 ;
  assign y977 = ~n46054 ;
  assign y978 = ~n45858 ;
  assign y979 = ~n46055 ;
  assign y980 = n44949 ;
  assign y981 = n46059 ;
  assign y982 = n46075 ;
  assign y983 = n46090 ;
  assign y984 = n46105 ;
  assign y985 = n46120 ;
  assign y986 = n46123 ;
  assign y987 = ~n46124 ;
  assign y988 = n45748 ;
  assign y989 = n46127 ;
  assign y990 = n46129 ;
  assign y991 = n46130 ;
  assign y992 = ~n46131 ;
  assign y993 = n46133 ;
  assign y994 = n46135 ;
  assign y995 = n46137 ;
  assign y996 = n46139 ;
  assign y997 = ~n46140 ;
  assign y998 = n46142 ;
  assign y999 = n46144 ;
  assign y1000 = n46146 ;
  assign y1001 = n46148 ;
  assign y1002 = n46150 ;
  assign y1003 = n46152 ;
  assign y1004 = n46154 ;
  assign y1005 = n46156 ;
  assign y1006 = n46158 ;
  assign y1007 = n46160 ;
  assign y1008 = n46162 ;
  assign y1009 = n46164 ;
  assign y1010 = n46166 ;
  assign y1011 = n46168 ;
  assign y1012 = n46170 ;
  assign y1013 = n46172 ;
  assign y1014 = n46174 ;
  assign y1015 = n46176 ;
  assign y1016 = n46178 ;
  assign y1017 = n46187 ;
  assign y1018 = n46189 ;
  assign y1019 = n46191 ;
  assign y1020 = n46193 ;
  assign y1021 = n46195 ;
  assign y1022 = n46197 ;
  assign y1023 = n46199 ;
  assign y1024 = n46201 ;
  assign y1025 = n46210 ;
  assign y1026 = n46212 ;
  assign y1027 = n46214 ;
  assign y1028 = n46216 ;
  assign y1029 = n46218 ;
  assign y1030 = n46220 ;
  assign y1031 = n46228 ;
  assign y1032 = n46230 ;
  assign y1033 = n46239 ;
  assign y1034 = n46248 ;
  assign y1035 = n46257 ;
  assign y1036 = n46259 ;
  assign y1037 = n46261 ;
  assign y1038 = n7318 ;
  assign y1039 = n46263 ;
  assign y1040 = n46265 ;
  assign y1041 = n46267 ;
  assign y1042 = n46269 ;
  assign y1043 = n46271 ;
  assign y1044 = n46273 ;
  assign y1045 = n46275 ;
  assign y1046 = n46277 ;
  assign y1047 = n46279 ;
  assign y1048 = n46281 ;
  assign y1049 = n5225 ;
  assign y1050 = n46283 ;
  assign y1051 = n46285 ;
  assign y1052 = n46287 ;
  assign y1053 = x67 ;
  assign y1054 = n46289 ;
  assign y1055 = n46291 ;
  assign y1056 = n46293 ;
  assign y1057 = n5035 ;
  assign y1058 = n46295 ;
  assign y1059 = n46297 ;
  assign y1060 = n46299 ;
  assign y1061 = n46301 ;
  assign y1062 = n46303 ;
  assign y1063 = n46313 ;
  assign y1064 = n46315 ;
  assign y1065 = n46317 ;
  assign y1066 = n46319 ;
  assign y1067 = n46321 ;
  assign y1068 = n46323 ;
  assign y1069 = n46325 ;
  assign y1070 = ~n46326 ;
  assign y1071 = n46328 ;
  assign y1072 = n46330 ;
  assign y1073 = n46332 ;
  assign y1074 = n46334 ;
  assign y1075 = n46336 ;
  assign y1076 = n46338 ;
  assign y1077 = n46340 ;
  assign y1078 = n46342 ;
  assign y1079 = n46344 ;
  assign y1080 = n46347 ;
  assign y1081 = n46349 ;
  assign y1082 = n46351 ;
  assign y1083 = n46353 ;
  assign y1084 = n46355 ;
  assign y1085 = n46357 ;
  assign y1086 = n46359 ;
  assign y1087 = n46361 ;
  assign y1088 = n46363 ;
  assign y1089 = n46365 ;
  assign y1090 = n46367 ;
  assign y1091 = n46369 ;
  assign y1092 = n46371 ;
  assign y1093 = n46373 ;
  assign y1094 = n46375 ;
  assign y1095 = n46377 ;
  assign y1096 = n46379 ;
  assign y1097 = n46381 ;
  assign y1098 = n46383 ;
  assign y1099 = n46385 ;
  assign y1100 = n46387 ;
  assign y1101 = n5082 ;
  assign y1102 = n46388 ;
  assign y1103 = n46390 ;
  assign y1104 = n46391 ;
  assign y1105 = ~n46392 ;
  assign y1106 = n15280 ;
  assign y1107 = n46393 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n46395 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n46396 ;
  assign y1116 = n46397 ;
  assign y1117 = x1014 ;
  assign y1118 = n46398 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n46399 ;
  assign y1123 = x1135 ;
  assign y1124 = n46400 ;
  assign y1125 = n46401 ;
  assign y1126 = n46402 ;
  assign y1127 = n46403 ;
  assign y1128 = n46404 ;
  assign y1129 = n46405 ;
  assign y1130 = ~x278 ;
  assign y1131 = n46406 ;
  assign y1132 = n46407 ;
  assign y1133 = ~n46408 ;
  assign y1134 = x1064 ;
  assign y1135 = n46409 ;
  assign y1136 = x299 ;
  assign y1137 = n46410 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
