module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 ;
  assign n1105 = ~x127 ;
  assign n196 = x126 & n1105 ;
  assign n1106 = ~n196 ;
  assign n197 = x125 & n1106 ;
  assign n1107 = ~x125 ;
  assign n198 = n1107 & x127 ;
  assign n199 = n197 | n198 ;
  assign n200 = x124 & n199 ;
  assign n201 = x124 | n196 ;
  assign n1108 = ~n200 ;
  assign n202 = n1108 & n201 ;
  assign n1109 = ~n202 ;
  assign n203 = x123 & n1109 ;
  assign n1110 = ~x123 ;
  assign n204 = n1110 & n199 ;
  assign n205 = n203 | n204 ;
  assign n206 = x122 & n205 ;
  assign n207 = x122 | n202 ;
  assign n1111 = ~n206 ;
  assign n208 = n1111 & n207 ;
  assign n1112 = ~n208 ;
  assign n209 = x121 & n1112 ;
  assign n1113 = ~x121 ;
  assign n210 = n1113 & n205 ;
  assign n211 = n209 | n210 ;
  assign n212 = x120 & n211 ;
  assign n213 = x120 | n208 ;
  assign n1114 = ~n212 ;
  assign n214 = n1114 & n213 ;
  assign n1115 = ~n214 ;
  assign n215 = x119 & n1115 ;
  assign n1116 = ~x119 ;
  assign n216 = n1116 & n211 ;
  assign n217 = n215 | n216 ;
  assign n218 = x118 & n217 ;
  assign n219 = x118 | n214 ;
  assign n1117 = ~n218 ;
  assign n220 = n1117 & n219 ;
  assign n1118 = ~n220 ;
  assign n221 = x117 & n1118 ;
  assign n1119 = ~x117 ;
  assign n222 = n1119 & n217 ;
  assign n223 = n221 | n222 ;
  assign n224 = x116 & n223 ;
  assign n225 = x116 | n220 ;
  assign n1120 = ~n224 ;
  assign n226 = n1120 & n225 ;
  assign n1121 = ~n226 ;
  assign n227 = x115 & n1121 ;
  assign n1122 = ~x115 ;
  assign n228 = n1122 & n223 ;
  assign n229 = n227 | n228 ;
  assign n230 = x114 & n229 ;
  assign n231 = x114 | n226 ;
  assign n1123 = ~n230 ;
  assign n232 = n1123 & n231 ;
  assign n1124 = ~n232 ;
  assign n233 = x113 & n1124 ;
  assign n1125 = ~x113 ;
  assign n234 = n1125 & n229 ;
  assign n235 = n233 | n234 ;
  assign n236 = x112 & n235 ;
  assign n237 = x112 | n232 ;
  assign n1126 = ~n236 ;
  assign n238 = n1126 & n237 ;
  assign n1127 = ~n238 ;
  assign n239 = x111 & n1127 ;
  assign n1128 = ~x111 ;
  assign n240 = n1128 & n235 ;
  assign n241 = n239 | n240 ;
  assign n242 = x110 & n241 ;
  assign n243 = x110 | n238 ;
  assign n1129 = ~n242 ;
  assign n244 = n1129 & n243 ;
  assign n1130 = ~n244 ;
  assign n245 = x109 & n1130 ;
  assign n1131 = ~x109 ;
  assign n246 = n1131 & n241 ;
  assign n247 = n245 | n246 ;
  assign n248 = x108 & n247 ;
  assign n249 = x108 | n244 ;
  assign n1132 = ~n248 ;
  assign n250 = n1132 & n249 ;
  assign n1133 = ~n250 ;
  assign n251 = x107 & n1133 ;
  assign n1134 = ~x107 ;
  assign n252 = n1134 & n247 ;
  assign n253 = n251 | n252 ;
  assign n254 = x106 & n253 ;
  assign n255 = x106 | n250 ;
  assign n1135 = ~n254 ;
  assign n256 = n1135 & n255 ;
  assign n1136 = ~n256 ;
  assign n257 = x105 & n1136 ;
  assign n1137 = ~x105 ;
  assign n258 = n1137 & n253 ;
  assign n259 = n257 | n258 ;
  assign n260 = x104 & n259 ;
  assign n261 = x104 | n256 ;
  assign n1138 = ~n260 ;
  assign n262 = n1138 & n261 ;
  assign n1139 = ~n262 ;
  assign n263 = x103 & n1139 ;
  assign n1140 = ~x103 ;
  assign n264 = n1140 & n259 ;
  assign n265 = n263 | n264 ;
  assign n266 = x102 & n265 ;
  assign n267 = x102 | n262 ;
  assign n1141 = ~n266 ;
  assign n268 = n1141 & n267 ;
  assign n1142 = ~n268 ;
  assign n269 = x101 & n1142 ;
  assign n1143 = ~x101 ;
  assign n270 = n1143 & n265 ;
  assign n271 = n269 | n270 ;
  assign n272 = x100 & n271 ;
  assign n273 = x100 | n268 ;
  assign n1144 = ~n272 ;
  assign n274 = n1144 & n273 ;
  assign n1145 = ~n274 ;
  assign n275 = x99 & n1145 ;
  assign n1146 = ~x99 ;
  assign n276 = n1146 & n271 ;
  assign n277 = n275 | n276 ;
  assign n278 = x98 & n277 ;
  assign n279 = x98 | n274 ;
  assign n1147 = ~n278 ;
  assign n280 = n1147 & n279 ;
  assign n1148 = ~n280 ;
  assign n281 = x97 & n1148 ;
  assign n1149 = ~x97 ;
  assign n282 = n1149 & n277 ;
  assign n283 = n281 | n282 ;
  assign n284 = x96 & n283 ;
  assign n285 = x96 | n280 ;
  assign n1150 = ~n284 ;
  assign n286 = n1150 & n285 ;
  assign n1151 = ~n286 ;
  assign n287 = x95 & n1151 ;
  assign n1152 = ~x95 ;
  assign n288 = n1152 & n283 ;
  assign n289 = n287 | n288 ;
  assign n290 = x94 & n289 ;
  assign n291 = x94 | n286 ;
  assign n1153 = ~n290 ;
  assign n292 = n1153 & n291 ;
  assign n1154 = ~n292 ;
  assign n293 = x93 & n1154 ;
  assign n1155 = ~x93 ;
  assign n294 = n1155 & n289 ;
  assign n295 = n293 | n294 ;
  assign n296 = x92 & n295 ;
  assign n297 = x92 | n292 ;
  assign n1156 = ~n296 ;
  assign n298 = n1156 & n297 ;
  assign n1157 = ~n298 ;
  assign n299 = x91 & n1157 ;
  assign n1158 = ~x91 ;
  assign n300 = n1158 & n295 ;
  assign n301 = n299 | n300 ;
  assign n302 = x90 & n301 ;
  assign n303 = x90 | n298 ;
  assign n1159 = ~n302 ;
  assign n304 = n1159 & n303 ;
  assign n1160 = ~n304 ;
  assign n305 = x89 & n1160 ;
  assign n1161 = ~x89 ;
  assign n306 = n1161 & n301 ;
  assign n307 = n305 | n306 ;
  assign n308 = x88 & n307 ;
  assign n309 = x88 | n304 ;
  assign n1162 = ~n308 ;
  assign n310 = n1162 & n309 ;
  assign n1163 = ~n310 ;
  assign n311 = x87 & n1163 ;
  assign n1164 = ~x87 ;
  assign n312 = n1164 & n307 ;
  assign n313 = n311 | n312 ;
  assign n314 = x86 & n313 ;
  assign n315 = x86 | n310 ;
  assign n1165 = ~n314 ;
  assign n316 = n1165 & n315 ;
  assign n1166 = ~n316 ;
  assign n317 = x85 & n1166 ;
  assign n1167 = ~x85 ;
  assign n318 = n1167 & n313 ;
  assign n319 = n317 | n318 ;
  assign n320 = x84 & n319 ;
  assign n321 = x84 | n316 ;
  assign n1168 = ~n320 ;
  assign n322 = n1168 & n321 ;
  assign n1169 = ~n322 ;
  assign n323 = x83 & n1169 ;
  assign n1170 = ~x83 ;
  assign n324 = n1170 & n319 ;
  assign n325 = n323 | n324 ;
  assign n326 = x82 & n325 ;
  assign n327 = x82 | n322 ;
  assign n1171 = ~n326 ;
  assign n328 = n1171 & n327 ;
  assign n1172 = ~n328 ;
  assign n329 = x81 & n1172 ;
  assign n1173 = ~x81 ;
  assign n330 = n1173 & n325 ;
  assign n331 = n329 | n330 ;
  assign n332 = x80 & n331 ;
  assign n333 = x80 | n328 ;
  assign n1174 = ~n332 ;
  assign n334 = n1174 & n333 ;
  assign n1175 = ~n334 ;
  assign n335 = x79 & n1175 ;
  assign n1176 = ~x79 ;
  assign n336 = n1176 & n331 ;
  assign n337 = n335 | n336 ;
  assign n338 = x78 & n337 ;
  assign n339 = x78 | n334 ;
  assign n1177 = ~n338 ;
  assign n340 = n1177 & n339 ;
  assign n1178 = ~n340 ;
  assign n341 = x77 & n1178 ;
  assign n1179 = ~x77 ;
  assign n342 = n1179 & n337 ;
  assign n343 = n341 | n342 ;
  assign n344 = x76 & n343 ;
  assign n345 = x76 | n340 ;
  assign n1180 = ~n344 ;
  assign n346 = n1180 & n345 ;
  assign n1181 = ~n346 ;
  assign n347 = x75 & n1181 ;
  assign n1182 = ~x75 ;
  assign n348 = n1182 & n343 ;
  assign n349 = n347 | n348 ;
  assign n350 = x74 & n349 ;
  assign n351 = x74 | n346 ;
  assign n1183 = ~n350 ;
  assign n352 = n1183 & n351 ;
  assign n1184 = ~n352 ;
  assign n353 = x73 & n1184 ;
  assign n1185 = ~x73 ;
  assign n354 = n1185 & n349 ;
  assign n355 = n353 | n354 ;
  assign n356 = x72 & n355 ;
  assign n357 = x72 | n352 ;
  assign n1186 = ~n356 ;
  assign n358 = n1186 & n357 ;
  assign n1187 = ~n358 ;
  assign n359 = x71 & n1187 ;
  assign n1188 = ~x71 ;
  assign n360 = n1188 & n355 ;
  assign n361 = n359 | n360 ;
  assign n362 = x70 & n361 ;
  assign n363 = x70 | n358 ;
  assign n1189 = ~n362 ;
  assign n364 = n1189 & n363 ;
  assign n1190 = ~n364 ;
  assign n365 = x69 & n1190 ;
  assign n1191 = ~x69 ;
  assign n366 = n1191 & n361 ;
  assign n367 = n365 | n366 ;
  assign n368 = x68 & n367 ;
  assign n369 = x68 | n364 ;
  assign n1192 = ~n368 ;
  assign n370 = n1192 & n369 ;
  assign n1193 = ~n370 ;
  assign n371 = x67 & n1193 ;
  assign n1194 = ~x67 ;
  assign n372 = n1194 & n367 ;
  assign n373 = n371 | n372 ;
  assign n374 = x66 & n373 ;
  assign n375 = x66 | n370 ;
  assign n1195 = ~n374 ;
  assign n376 = n1195 & n375 ;
  assign n1196 = ~n376 ;
  assign n377 = x65 & n1196 ;
  assign n1197 = ~x65 ;
  assign n378 = n1197 & n373 ;
  assign n379 = n377 | n378 ;
  assign n380 = x64 & n379 ;
  assign n381 = x64 | n376 ;
  assign n1198 = ~n380 ;
  assign n382 = n1198 & n381 ;
  assign n1199 = ~n382 ;
  assign n383 = x63 & n1199 ;
  assign n1200 = ~x63 ;
  assign n384 = n1200 & n379 ;
  assign n385 = n383 | n384 ;
  assign n386 = x62 & n385 ;
  assign n387 = x62 | n382 ;
  assign n1201 = ~n386 ;
  assign n388 = n1201 & n387 ;
  assign n1202 = ~n388 ;
  assign n389 = x61 & n1202 ;
  assign n1203 = ~x61 ;
  assign n390 = n1203 & n385 ;
  assign n391 = n389 | n390 ;
  assign n392 = x60 & n391 ;
  assign n393 = x60 | n388 ;
  assign n1204 = ~n392 ;
  assign n394 = n1204 & n393 ;
  assign n1205 = ~n394 ;
  assign n395 = x59 & n1205 ;
  assign n1206 = ~x59 ;
  assign n396 = n1206 & n391 ;
  assign n397 = n395 | n396 ;
  assign n398 = x58 & n397 ;
  assign n399 = x58 | n394 ;
  assign n1207 = ~n398 ;
  assign n400 = n1207 & n399 ;
  assign n1208 = ~n400 ;
  assign n401 = x57 & n1208 ;
  assign n1209 = ~x57 ;
  assign n402 = n1209 & n397 ;
  assign n403 = n401 | n402 ;
  assign n404 = x56 & n403 ;
  assign n405 = x56 | n400 ;
  assign n1210 = ~n404 ;
  assign n406 = n1210 & n405 ;
  assign n1211 = ~n406 ;
  assign n407 = x55 & n1211 ;
  assign n1212 = ~x55 ;
  assign n408 = n1212 & n403 ;
  assign n409 = n407 | n408 ;
  assign n410 = x54 & n409 ;
  assign n411 = x54 | n406 ;
  assign n1213 = ~n410 ;
  assign n412 = n1213 & n411 ;
  assign n1214 = ~n412 ;
  assign n413 = x53 & n1214 ;
  assign n1215 = ~x53 ;
  assign n414 = n1215 & n409 ;
  assign n415 = n413 | n414 ;
  assign n416 = x52 & n415 ;
  assign n417 = x52 | n412 ;
  assign n1216 = ~n416 ;
  assign n418 = n1216 & n417 ;
  assign n1217 = ~n418 ;
  assign n419 = x51 & n1217 ;
  assign n1218 = ~x51 ;
  assign n420 = n1218 & n415 ;
  assign n421 = n419 | n420 ;
  assign n422 = x50 & n421 ;
  assign n423 = x50 | n418 ;
  assign n1219 = ~n422 ;
  assign n424 = n1219 & n423 ;
  assign n1220 = ~n424 ;
  assign n425 = x49 & n1220 ;
  assign n1221 = ~x49 ;
  assign n426 = n1221 & n421 ;
  assign n427 = n425 | n426 ;
  assign n428 = x48 & n427 ;
  assign n429 = x48 | n424 ;
  assign n1222 = ~n428 ;
  assign n430 = n1222 & n429 ;
  assign n1223 = ~n430 ;
  assign n431 = x47 & n1223 ;
  assign n1224 = ~x47 ;
  assign n432 = n1224 & n427 ;
  assign n433 = n431 | n432 ;
  assign n434 = x46 & n433 ;
  assign n435 = x46 | n430 ;
  assign n1225 = ~n434 ;
  assign n436 = n1225 & n435 ;
  assign n1226 = ~n436 ;
  assign n437 = x45 & n1226 ;
  assign n1227 = ~x45 ;
  assign n438 = n1227 & n433 ;
  assign n439 = n437 | n438 ;
  assign n440 = x44 & n439 ;
  assign n441 = x44 | n436 ;
  assign n1228 = ~n440 ;
  assign n442 = n1228 & n441 ;
  assign n1229 = ~n442 ;
  assign n443 = x43 & n1229 ;
  assign n1230 = ~x43 ;
  assign n444 = n1230 & n439 ;
  assign n445 = n443 | n444 ;
  assign n446 = x42 & n445 ;
  assign n447 = x42 | n442 ;
  assign n1231 = ~n446 ;
  assign n448 = n1231 & n447 ;
  assign n1232 = ~n448 ;
  assign n449 = x41 & n1232 ;
  assign n1233 = ~x41 ;
  assign n450 = n1233 & n445 ;
  assign n451 = n449 | n450 ;
  assign n452 = x40 & n451 ;
  assign n453 = x40 | n448 ;
  assign n1234 = ~n452 ;
  assign n454 = n1234 & n453 ;
  assign n1235 = ~n454 ;
  assign n455 = x39 & n1235 ;
  assign n1236 = ~x39 ;
  assign n456 = n1236 & n451 ;
  assign n457 = n455 | n456 ;
  assign n458 = x38 & n457 ;
  assign n459 = x38 | n454 ;
  assign n1237 = ~n458 ;
  assign n460 = n1237 & n459 ;
  assign n1238 = ~n460 ;
  assign n461 = x37 & n1238 ;
  assign n1239 = ~x37 ;
  assign n462 = n1239 & n457 ;
  assign n463 = n461 | n462 ;
  assign n464 = x36 & n463 ;
  assign n465 = x36 | n460 ;
  assign n1240 = ~n464 ;
  assign n466 = n1240 & n465 ;
  assign n1241 = ~n466 ;
  assign n467 = x35 & n1241 ;
  assign n1242 = ~x35 ;
  assign n468 = n1242 & n463 ;
  assign n469 = n467 | n468 ;
  assign n470 = x34 & n469 ;
  assign n471 = x34 | n466 ;
  assign n1243 = ~n470 ;
  assign n472 = n1243 & n471 ;
  assign n1244 = ~n472 ;
  assign n473 = x33 & n1244 ;
  assign n1245 = ~x33 ;
  assign n474 = n1245 & n469 ;
  assign n475 = n473 | n474 ;
  assign n476 = x32 & n475 ;
  assign n477 = x32 | n472 ;
  assign n1246 = ~n476 ;
  assign n478 = n1246 & n477 ;
  assign n1247 = ~n478 ;
  assign n479 = x31 & n1247 ;
  assign n1248 = ~x31 ;
  assign n480 = n1248 & n475 ;
  assign n481 = n479 | n480 ;
  assign n482 = x30 & n481 ;
  assign n483 = x30 | n478 ;
  assign n1249 = ~n482 ;
  assign n484 = n1249 & n483 ;
  assign n1250 = ~n484 ;
  assign n485 = x29 & n1250 ;
  assign n1251 = ~x29 ;
  assign n486 = n1251 & n481 ;
  assign n487 = n485 | n486 ;
  assign n488 = x28 & n487 ;
  assign n489 = x28 | n484 ;
  assign n1252 = ~n488 ;
  assign n490 = n1252 & n489 ;
  assign n1253 = ~n490 ;
  assign n491 = x27 & n1253 ;
  assign n1254 = ~x27 ;
  assign n492 = n1254 & n487 ;
  assign n493 = n491 | n492 ;
  assign n494 = x26 & n493 ;
  assign n495 = x26 | n490 ;
  assign n1255 = ~n494 ;
  assign n496 = n1255 & n495 ;
  assign n1256 = ~n496 ;
  assign n497 = x25 & n1256 ;
  assign n1257 = ~x25 ;
  assign n498 = n1257 & n493 ;
  assign n499 = n497 | n498 ;
  assign n500 = x24 & n499 ;
  assign n501 = x24 | n496 ;
  assign n1258 = ~n500 ;
  assign n502 = n1258 & n501 ;
  assign n1259 = ~n502 ;
  assign n503 = x23 & n1259 ;
  assign n1260 = ~x23 ;
  assign n504 = n1260 & n499 ;
  assign n505 = n503 | n504 ;
  assign n506 = x22 & n505 ;
  assign n507 = x22 | n502 ;
  assign n1261 = ~n506 ;
  assign n508 = n1261 & n507 ;
  assign n1262 = ~n508 ;
  assign n509 = x21 & n1262 ;
  assign n1263 = ~x21 ;
  assign n510 = n1263 & n505 ;
  assign n511 = n509 | n510 ;
  assign n512 = x20 & n511 ;
  assign n513 = x20 | n508 ;
  assign n1264 = ~n512 ;
  assign n514 = n1264 & n513 ;
  assign n1265 = ~n514 ;
  assign n515 = x19 & n1265 ;
  assign n1266 = ~x19 ;
  assign n516 = n1266 & n511 ;
  assign n517 = n515 | n516 ;
  assign n518 = x18 & n517 ;
  assign n519 = x18 | n514 ;
  assign n1267 = ~n518 ;
  assign n520 = n1267 & n519 ;
  assign n1268 = ~n520 ;
  assign n521 = x17 & n1268 ;
  assign n1269 = ~x17 ;
  assign n522 = n1269 & n517 ;
  assign n523 = n521 | n522 ;
  assign n524 = x16 & n523 ;
  assign n525 = x16 | n520 ;
  assign n1270 = ~n524 ;
  assign n526 = n1270 & n525 ;
  assign n1271 = ~n526 ;
  assign n527 = x15 & n1271 ;
  assign n1272 = ~x15 ;
  assign n528 = n1272 & n523 ;
  assign n529 = n527 | n528 ;
  assign n530 = x14 & n529 ;
  assign n531 = x14 | n526 ;
  assign n1273 = ~n530 ;
  assign n532 = n1273 & n531 ;
  assign n1274 = ~n532 ;
  assign n533 = x13 & n1274 ;
  assign n1275 = ~x13 ;
  assign n534 = n1275 & n529 ;
  assign n535 = n533 | n534 ;
  assign n536 = x12 & n535 ;
  assign n537 = x12 | n532 ;
  assign n1276 = ~n536 ;
  assign n538 = n1276 & n537 ;
  assign n1277 = ~n538 ;
  assign n539 = x11 & n1277 ;
  assign n1278 = ~x11 ;
  assign n540 = n1278 & n535 ;
  assign n541 = n539 | n540 ;
  assign n542 = x10 & n541 ;
  assign n543 = x10 | n538 ;
  assign n1279 = ~n542 ;
  assign n544 = n1279 & n543 ;
  assign n1280 = ~n544 ;
  assign n545 = x9 & n1280 ;
  assign n1281 = ~x9 ;
  assign n546 = n1281 & n541 ;
  assign n547 = n545 | n546 ;
  assign n548 = x8 & n547 ;
  assign n549 = x8 | n544 ;
  assign n1282 = ~n548 ;
  assign n550 = n1282 & n549 ;
  assign n1283 = ~n550 ;
  assign n551 = x7 & n1283 ;
  assign n1284 = ~x7 ;
  assign n552 = n1284 & n547 ;
  assign n553 = n551 | n552 ;
  assign n554 = x6 & n553 ;
  assign n555 = x6 | n550 ;
  assign n1285 = ~n554 ;
  assign n556 = n1285 & n555 ;
  assign n1286 = ~n556 ;
  assign n557 = x5 & n1286 ;
  assign n1287 = ~x5 ;
  assign n558 = n1287 & n553 ;
  assign n559 = n557 | n558 ;
  assign n560 = x4 & n559 ;
  assign n561 = x4 | n556 ;
  assign n1288 = ~n560 ;
  assign n562 = n1288 & n561 ;
  assign n1289 = ~x2 ;
  assign n566 = x1 & n1289 ;
  assign n1290 = ~n562 ;
  assign n567 = n1290 & n566 ;
  assign n563 = x3 & n1290 ;
  assign n1291 = ~x3 ;
  assign n564 = n1291 & n559 ;
  assign n565 = n563 | n564 ;
  assign n1292 = ~n566 ;
  assign n568 = n565 & n1292 ;
  assign n129 = n567 | n568 ;
  assign n163 = x78 | x79 ;
  assign n171 = x94 | x95 ;
  assign n146 = x102 | x103 ;
  assign n150 = x110 | x111 ;
  assign n137 = x114 | x115 ;
  assign n139 = x118 | x119 ;
  assign n195 = x126 | x127 ;
  assign n569 = x124 | x125 ;
  assign n942 = x122 | x123 ;
  assign n1293 = ~n569 ;
  assign n570 = n1293 & n942 ;
  assign n571 = n195 | n570 ;
  assign n1294 = ~n139 ;
  assign n573 = n1294 & n571 ;
  assign n572 = x120 & n571 ;
  assign n1295 = ~n942 ;
  assign n1024 = x121 & n1295 ;
  assign n574 = n569 | n1024 ;
  assign n1296 = ~n195 ;
  assign n575 = n1296 & n574 ;
  assign n576 = x120 | n575 ;
  assign n1297 = ~n572 ;
  assign n577 = n1297 & n576 ;
  assign n1298 = ~n577 ;
  assign n578 = n139 & n1298 ;
  assign n579 = n573 | n578 ;
  assign n1299 = ~n137 ;
  assign n580 = n1299 & n579 ;
  assign n581 = x116 | x117 ;
  assign n582 = n577 | n581 ;
  assign n583 = n579 & n581 ;
  assign n1300 = ~n583 ;
  assign n584 = n582 & n1300 ;
  assign n1301 = ~n584 ;
  assign n585 = n137 & n1301 ;
  assign n586 = n580 | n585 ;
  assign n1302 = ~n150 ;
  assign n587 = n1302 & n586 ;
  assign n588 = x112 | x113 ;
  assign n589 = n584 | n588 ;
  assign n590 = n586 & n588 ;
  assign n1303 = ~n590 ;
  assign n591 = n589 & n1303 ;
  assign n1304 = ~n591 ;
  assign n592 = n150 & n1304 ;
  assign n593 = n587 | n592 ;
  assign n598 = x106 | x107 ;
  assign n1305 = ~n598 ;
  assign n599 = n593 & n1305 ;
  assign n594 = x108 | x109 ;
  assign n595 = n591 | n594 ;
  assign n596 = n593 & n594 ;
  assign n1306 = ~n596 ;
  assign n597 = n595 & n1306 ;
  assign n1307 = ~n597 ;
  assign n600 = n1307 & n598 ;
  assign n601 = n599 | n600 ;
  assign n1308 = ~n146 ;
  assign n602 = n1308 & n601 ;
  assign n603 = x104 | x105 ;
  assign n604 = n597 | n603 ;
  assign n605 = n601 & n603 ;
  assign n1309 = ~n605 ;
  assign n606 = n604 & n1309 ;
  assign n1310 = ~n606 ;
  assign n607 = n146 & n1310 ;
  assign n608 = n602 | n607 ;
  assign n613 = x98 | x99 ;
  assign n1311 = ~n613 ;
  assign n614 = n608 & n1311 ;
  assign n609 = x100 | x101 ;
  assign n610 = n606 | n609 ;
  assign n611 = n608 & n609 ;
  assign n1312 = ~n611 ;
  assign n612 = n610 & n1312 ;
  assign n1313 = ~n612 ;
  assign n615 = n1313 & n613 ;
  assign n616 = n614 | n615 ;
  assign n1314 = ~n171 ;
  assign n617 = n1314 & n616 ;
  assign n618 = x96 | x97 ;
  assign n619 = n612 | n618 ;
  assign n620 = n616 & n618 ;
  assign n1315 = ~n620 ;
  assign n621 = n619 & n1315 ;
  assign n1316 = ~n621 ;
  assign n622 = n171 & n1316 ;
  assign n623 = n617 | n622 ;
  assign n628 = x90 | x91 ;
  assign n1317 = ~n628 ;
  assign n629 = n623 & n1317 ;
  assign n624 = x92 | x93 ;
  assign n625 = n621 | n624 ;
  assign n626 = n623 & n624 ;
  assign n1318 = ~n626 ;
  assign n627 = n625 & n1318 ;
  assign n1319 = ~n627 ;
  assign n630 = n1319 & n628 ;
  assign n631 = n629 | n630 ;
  assign n636 = x86 | x87 ;
  assign n1320 = ~n636 ;
  assign n637 = n631 & n1320 ;
  assign n632 = x88 | x89 ;
  assign n633 = n627 | n632 ;
  assign n634 = n631 & n632 ;
  assign n1321 = ~n634 ;
  assign n635 = n633 & n1321 ;
  assign n1322 = ~n635 ;
  assign n638 = n1322 & n636 ;
  assign n639 = n637 | n638 ;
  assign n644 = x82 | x83 ;
  assign n1323 = ~n644 ;
  assign n645 = n639 & n1323 ;
  assign n640 = x84 | x85 ;
  assign n641 = n635 | n640 ;
  assign n642 = n639 & n640 ;
  assign n1324 = ~n642 ;
  assign n643 = n641 & n1324 ;
  assign n1325 = ~n643 ;
  assign n646 = n1325 & n644 ;
  assign n647 = n645 | n646 ;
  assign n1326 = ~n163 ;
  assign n648 = n1326 & n647 ;
  assign n649 = x80 | x81 ;
  assign n650 = n643 | n649 ;
  assign n651 = n647 & n649 ;
  assign n1327 = ~n651 ;
  assign n652 = n650 & n1327 ;
  assign n1328 = ~n652 ;
  assign n653 = n163 & n1328 ;
  assign n654 = n648 | n653 ;
  assign n659 = x74 | x75 ;
  assign n1329 = ~n659 ;
  assign n660 = n654 & n1329 ;
  assign n655 = x76 | x77 ;
  assign n656 = n652 | n655 ;
  assign n657 = n654 & n655 ;
  assign n1330 = ~n657 ;
  assign n658 = n656 & n1330 ;
  assign n1331 = ~n658 ;
  assign n661 = n1331 & n659 ;
  assign n662 = n660 | n661 ;
  assign n667 = x70 | x71 ;
  assign n1332 = ~n667 ;
  assign n668 = n662 & n1332 ;
  assign n663 = x72 | x73 ;
  assign n664 = n658 | n663 ;
  assign n665 = n662 & n663 ;
  assign n1333 = ~n665 ;
  assign n666 = n664 & n1333 ;
  assign n1334 = ~n666 ;
  assign n669 = n1334 & n667 ;
  assign n670 = n668 | n669 ;
  assign n675 = x66 | x67 ;
  assign n1335 = ~n675 ;
  assign n676 = n670 & n1335 ;
  assign n671 = x68 | x69 ;
  assign n672 = n666 | n671 ;
  assign n673 = n670 & n671 ;
  assign n1336 = ~n673 ;
  assign n674 = n672 & n1336 ;
  assign n1337 = ~n674 ;
  assign n677 = n1337 & n675 ;
  assign n678 = n676 | n677 ;
  assign n683 = x62 | x63 ;
  assign n1338 = ~n683 ;
  assign n684 = n678 & n1338 ;
  assign n679 = x64 | x65 ;
  assign n680 = n674 | n679 ;
  assign n681 = n678 & n679 ;
  assign n1339 = ~n681 ;
  assign n682 = n680 & n1339 ;
  assign n1340 = ~n682 ;
  assign n685 = n1340 & n683 ;
  assign n686 = n684 | n685 ;
  assign n691 = x58 | x59 ;
  assign n1341 = ~n691 ;
  assign n692 = n686 & n1341 ;
  assign n687 = x60 | x61 ;
  assign n688 = n682 | n687 ;
  assign n689 = n686 & n687 ;
  assign n1342 = ~n689 ;
  assign n690 = n688 & n1342 ;
  assign n1343 = ~n690 ;
  assign n693 = n1343 & n691 ;
  assign n694 = n692 | n693 ;
  assign n699 = x54 | x55 ;
  assign n1344 = ~n699 ;
  assign n700 = n694 & n1344 ;
  assign n695 = x56 | x57 ;
  assign n696 = n690 | n695 ;
  assign n697 = n694 & n695 ;
  assign n1345 = ~n697 ;
  assign n698 = n696 & n1345 ;
  assign n1346 = ~n698 ;
  assign n701 = n1346 & n699 ;
  assign n702 = n700 | n701 ;
  assign n707 = x50 | x51 ;
  assign n1347 = ~n707 ;
  assign n708 = n702 & n1347 ;
  assign n703 = x52 | x53 ;
  assign n704 = n698 | n703 ;
  assign n705 = n702 & n703 ;
  assign n1348 = ~n705 ;
  assign n706 = n704 & n1348 ;
  assign n1349 = ~n706 ;
  assign n709 = n1349 & n707 ;
  assign n710 = n708 | n709 ;
  assign n715 = x46 | x47 ;
  assign n1350 = ~n715 ;
  assign n716 = n710 & n1350 ;
  assign n711 = x48 | x49 ;
  assign n712 = n706 | n711 ;
  assign n713 = n710 & n711 ;
  assign n1351 = ~n713 ;
  assign n714 = n712 & n1351 ;
  assign n1352 = ~n714 ;
  assign n717 = n1352 & n715 ;
  assign n718 = n716 | n717 ;
  assign n723 = x42 | x43 ;
  assign n1353 = ~n723 ;
  assign n724 = n718 & n1353 ;
  assign n719 = x44 | x45 ;
  assign n720 = n714 | n719 ;
  assign n721 = n718 & n719 ;
  assign n1354 = ~n721 ;
  assign n722 = n720 & n1354 ;
  assign n1355 = ~n722 ;
  assign n725 = n1355 & n723 ;
  assign n726 = n724 | n725 ;
  assign n731 = x38 | x39 ;
  assign n1356 = ~n731 ;
  assign n732 = n726 & n1356 ;
  assign n727 = x40 | x41 ;
  assign n728 = n722 | n727 ;
  assign n729 = n726 & n727 ;
  assign n1357 = ~n729 ;
  assign n730 = n728 & n1357 ;
  assign n1358 = ~n730 ;
  assign n733 = n1358 & n731 ;
  assign n734 = n732 | n733 ;
  assign n739 = x34 | x35 ;
  assign n1359 = ~n739 ;
  assign n740 = n734 & n1359 ;
  assign n735 = x36 | x37 ;
  assign n736 = n730 | n735 ;
  assign n737 = n734 & n735 ;
  assign n1360 = ~n737 ;
  assign n738 = n736 & n1360 ;
  assign n1361 = ~n738 ;
  assign n741 = n1361 & n739 ;
  assign n742 = n740 | n741 ;
  assign n747 = x30 | x31 ;
  assign n1362 = ~n747 ;
  assign n748 = n742 & n1362 ;
  assign n743 = x32 | x33 ;
  assign n744 = n738 | n743 ;
  assign n745 = n742 & n743 ;
  assign n1363 = ~n745 ;
  assign n746 = n744 & n1363 ;
  assign n1364 = ~n746 ;
  assign n749 = n1364 & n747 ;
  assign n750 = n748 | n749 ;
  assign n755 = x26 | x27 ;
  assign n1365 = ~n755 ;
  assign n756 = n750 & n1365 ;
  assign n751 = x28 | x29 ;
  assign n752 = n746 | n751 ;
  assign n753 = n750 & n751 ;
  assign n1366 = ~n753 ;
  assign n754 = n752 & n1366 ;
  assign n1367 = ~n754 ;
  assign n757 = n1367 & n755 ;
  assign n758 = n756 | n757 ;
  assign n763 = x22 | x23 ;
  assign n1368 = ~n763 ;
  assign n764 = n758 & n1368 ;
  assign n759 = x24 | x25 ;
  assign n760 = n754 | n759 ;
  assign n761 = n758 & n759 ;
  assign n1369 = ~n761 ;
  assign n762 = n760 & n1369 ;
  assign n1370 = ~n762 ;
  assign n765 = n1370 & n763 ;
  assign n766 = n764 | n765 ;
  assign n771 = x18 | x19 ;
  assign n1371 = ~n771 ;
  assign n772 = n766 & n1371 ;
  assign n767 = x20 | x21 ;
  assign n768 = n762 | n767 ;
  assign n769 = n766 & n767 ;
  assign n1372 = ~n769 ;
  assign n770 = n768 & n1372 ;
  assign n1373 = ~n770 ;
  assign n773 = n1373 & n771 ;
  assign n774 = n772 | n773 ;
  assign n779 = x14 | x15 ;
  assign n1374 = ~n779 ;
  assign n780 = n774 & n1374 ;
  assign n775 = x16 | x17 ;
  assign n776 = n770 | n775 ;
  assign n777 = n774 & n775 ;
  assign n1375 = ~n777 ;
  assign n778 = n776 & n1375 ;
  assign n1376 = ~n778 ;
  assign n781 = n1376 & n779 ;
  assign n782 = n780 | n781 ;
  assign n787 = x10 | x11 ;
  assign n1377 = ~n787 ;
  assign n788 = n782 & n1377 ;
  assign n783 = x12 | x13 ;
  assign n784 = n778 | n783 ;
  assign n785 = n782 & n783 ;
  assign n1378 = ~n785 ;
  assign n786 = n784 & n1378 ;
  assign n1379 = ~n786 ;
  assign n789 = n1379 & n787 ;
  assign n790 = n788 | n789 ;
  assign n795 = x6 | x7 ;
  assign n1380 = ~n795 ;
  assign n796 = n790 & n1380 ;
  assign n791 = x8 | x9 ;
  assign n792 = n786 | n791 ;
  assign n793 = n790 & n791 ;
  assign n1381 = ~n793 ;
  assign n794 = n792 & n1381 ;
  assign n1382 = ~n794 ;
  assign n797 = n1382 & n795 ;
  assign n798 = n796 | n797 ;
  assign n803 = x2 | x3 ;
  assign n1383 = ~n803 ;
  assign n804 = n798 & n1383 ;
  assign n799 = x4 | x5 ;
  assign n800 = n794 | n799 ;
  assign n801 = n798 & n799 ;
  assign n1384 = ~n801 ;
  assign n802 = n800 & n1384 ;
  assign n1385 = ~n802 ;
  assign n805 = n1385 & n803 ;
  assign n130 = n804 | n805 ;
  assign n164 = x77 | n163 ;
  assign n165 = x76 | n164 ;
  assign n172 = x93 | n171 ;
  assign n173 = x92 | n172 ;
  assign n147 = x101 | n146 ;
  assign n148 = x100 | n147 ;
  assign n151 = x109 | n150 ;
  assign n152 = x108 | n151 ;
  assign n806 = n195 | n569 ;
  assign n1078 = x120 | x121 ;
  assign n1098 = n942 | n1078 ;
  assign n140 = x117 | n139 ;
  assign n141 = x116 | n140 ;
  assign n1386 = ~n1098 ;
  assign n807 = n1386 & n141 ;
  assign n808 = n806 | n807 ;
  assign n1387 = ~n152 ;
  assign n809 = n1387 & n808 ;
  assign n810 = x113 | x114 ;
  assign n811 = x112 | n810 ;
  assign n812 = n808 & n811 ;
  assign n1388 = ~n141 ;
  assign n143 = x115 & n1388 ;
  assign n813 = n1098 | n143 ;
  assign n1389 = ~n806 ;
  assign n814 = n1389 & n813 ;
  assign n815 = n811 | n814 ;
  assign n1390 = ~n812 ;
  assign n816 = n1390 & n815 ;
  assign n1391 = ~n816 ;
  assign n817 = n152 & n1391 ;
  assign n818 = n809 | n817 ;
  assign n1392 = ~n148 ;
  assign n819 = n1392 & n818 ;
  assign n820 = x105 | n598 ;
  assign n821 = x104 | n820 ;
  assign n822 = n816 | n821 ;
  assign n823 = n818 & n821 ;
  assign n1393 = ~n823 ;
  assign n824 = n822 & n1393 ;
  assign n1394 = ~n824 ;
  assign n825 = n148 & n1394 ;
  assign n826 = n819 | n825 ;
  assign n1395 = ~n173 ;
  assign n827 = n1395 & n826 ;
  assign n828 = x97 | n613 ;
  assign n829 = x96 | n828 ;
  assign n830 = n824 | n829 ;
  assign n831 = n826 & n829 ;
  assign n1396 = ~n831 ;
  assign n832 = n830 & n1396 ;
  assign n1397 = ~n832 ;
  assign n833 = n173 & n1397 ;
  assign n834 = n827 | n833 ;
  assign n840 = x85 | n636 ;
  assign n841 = x84 | n840 ;
  assign n1398 = ~n841 ;
  assign n842 = n834 & n1398 ;
  assign n835 = x89 | n628 ;
  assign n836 = x88 | n835 ;
  assign n837 = n832 | n836 ;
  assign n838 = n834 & n836 ;
  assign n1399 = ~n838 ;
  assign n839 = n837 & n1399 ;
  assign n1400 = ~n839 ;
  assign n843 = n1400 & n841 ;
  assign n844 = n842 | n843 ;
  assign n1401 = ~n165 ;
  assign n845 = n1401 & n844 ;
  assign n846 = x81 | n644 ;
  assign n847 = x80 | n846 ;
  assign n848 = n839 | n847 ;
  assign n849 = n844 & n847 ;
  assign n1402 = ~n849 ;
  assign n850 = n848 & n1402 ;
  assign n1403 = ~n850 ;
  assign n851 = n165 & n1403 ;
  assign n852 = n845 | n851 ;
  assign n858 = x69 | n667 ;
  assign n859 = x68 | n858 ;
  assign n1404 = ~n859 ;
  assign n860 = n852 & n1404 ;
  assign n853 = x73 | n659 ;
  assign n854 = x72 | n853 ;
  assign n855 = n850 | n854 ;
  assign n856 = n852 & n854 ;
  assign n1405 = ~n856 ;
  assign n857 = n855 & n1405 ;
  assign n1406 = ~n857 ;
  assign n861 = n1406 & n859 ;
  assign n862 = n860 | n861 ;
  assign n868 = x61 | n683 ;
  assign n869 = x60 | n868 ;
  assign n1407 = ~n869 ;
  assign n870 = n862 & n1407 ;
  assign n863 = x65 | n675 ;
  assign n864 = x64 | n863 ;
  assign n865 = n857 | n864 ;
  assign n866 = n862 & n864 ;
  assign n1408 = ~n866 ;
  assign n867 = n865 & n1408 ;
  assign n1409 = ~n867 ;
  assign n871 = n1409 & n869 ;
  assign n872 = n870 | n871 ;
  assign n878 = x53 | n699 ;
  assign n879 = x52 | n878 ;
  assign n1410 = ~n879 ;
  assign n880 = n872 & n1410 ;
  assign n873 = x57 | n691 ;
  assign n874 = x56 | n873 ;
  assign n875 = n867 | n874 ;
  assign n876 = n872 & n874 ;
  assign n1411 = ~n876 ;
  assign n877 = n875 & n1411 ;
  assign n1412 = ~n877 ;
  assign n881 = n1412 & n879 ;
  assign n882 = n880 | n881 ;
  assign n888 = x45 | n715 ;
  assign n889 = x44 | n888 ;
  assign n1413 = ~n889 ;
  assign n890 = n882 & n1413 ;
  assign n883 = x49 | n707 ;
  assign n884 = x48 | n883 ;
  assign n885 = n877 | n884 ;
  assign n886 = n882 & n884 ;
  assign n1414 = ~n886 ;
  assign n887 = n885 & n1414 ;
  assign n1415 = ~n887 ;
  assign n891 = n1415 & n889 ;
  assign n892 = n890 | n891 ;
  assign n898 = x37 | n731 ;
  assign n899 = x36 | n898 ;
  assign n1416 = ~n899 ;
  assign n900 = n892 & n1416 ;
  assign n893 = x41 | n723 ;
  assign n894 = x40 | n893 ;
  assign n895 = n887 | n894 ;
  assign n896 = n892 & n894 ;
  assign n1417 = ~n896 ;
  assign n897 = n895 & n1417 ;
  assign n1418 = ~n897 ;
  assign n901 = n1418 & n899 ;
  assign n902 = n900 | n901 ;
  assign n908 = x29 | n747 ;
  assign n909 = x28 | n908 ;
  assign n1419 = ~n909 ;
  assign n910 = n902 & n1419 ;
  assign n903 = x33 | n739 ;
  assign n904 = x32 | n903 ;
  assign n905 = n897 | n904 ;
  assign n906 = n902 & n904 ;
  assign n1420 = ~n906 ;
  assign n907 = n905 & n1420 ;
  assign n1421 = ~n907 ;
  assign n911 = n1421 & n909 ;
  assign n912 = n910 | n911 ;
  assign n918 = x21 | n763 ;
  assign n919 = x20 | n918 ;
  assign n1422 = ~n919 ;
  assign n920 = n912 & n1422 ;
  assign n913 = x25 | n755 ;
  assign n914 = x24 | n913 ;
  assign n915 = n907 | n914 ;
  assign n916 = n912 & n914 ;
  assign n1423 = ~n916 ;
  assign n917 = n915 & n1423 ;
  assign n1424 = ~n917 ;
  assign n921 = n1424 & n919 ;
  assign n922 = n920 | n921 ;
  assign n928 = x13 | n779 ;
  assign n929 = x12 | n928 ;
  assign n1425 = ~n929 ;
  assign n930 = n922 & n1425 ;
  assign n923 = x17 | n771 ;
  assign n924 = x16 | n923 ;
  assign n925 = n917 | n924 ;
  assign n926 = n922 & n924 ;
  assign n1426 = ~n926 ;
  assign n927 = n925 & n1426 ;
  assign n1427 = ~n927 ;
  assign n931 = n1427 & n929 ;
  assign n932 = n930 | n931 ;
  assign n938 = x5 | n795 ;
  assign n939 = x4 | n938 ;
  assign n1428 = ~n939 ;
  assign n940 = n932 & n1428 ;
  assign n933 = x9 | n787 ;
  assign n934 = x8 | n933 ;
  assign n935 = n927 | n934 ;
  assign n936 = n932 & n934 ;
  assign n1429 = ~n936 ;
  assign n937 = n935 & n1429 ;
  assign n1430 = ~n937 ;
  assign n941 = n1430 & n939 ;
  assign n131 = n940 | n941 ;
  assign n166 = x75 | n165 ;
  assign n167 = x74 | n166 ;
  assign n168 = x73 | n167 ;
  assign n169 = x72 | n168 ;
  assign n174 = x91 | n173 ;
  assign n175 = x90 | n174 ;
  assign n176 = x89 | n175 ;
  assign n177 = x88 | n176 ;
  assign n1104 = n806 | n1098 ;
  assign n138 = x113 | n137 ;
  assign n142 = x112 | n141 ;
  assign n144 = n138 | n142 ;
  assign n153 = x107 | n152 ;
  assign n154 = x106 | n153 ;
  assign n155 = x105 | n154 ;
  assign n156 = x104 | n155 ;
  assign n1431 = ~n144 ;
  assign n943 = n1431 & n156 ;
  assign n944 = n1104 | n943 ;
  assign n1432 = ~n177 ;
  assign n945 = n1432 & n944 ;
  assign n946 = x101 | x102 ;
  assign n947 = x100 | n946 ;
  assign n948 = x99 | n947 ;
  assign n949 = x98 | n948 ;
  assign n950 = x97 | n949 ;
  assign n951 = x96 | n950 ;
  assign n952 = n944 & n951 ;
  assign n1433 = ~n156 ;
  assign n158 = x103 & n1433 ;
  assign n953 = n144 | n158 ;
  assign n1434 = ~n1104 ;
  assign n954 = n1434 & n953 ;
  assign n955 = n951 | n954 ;
  assign n1435 = ~n952 ;
  assign n956 = n1435 & n955 ;
  assign n1436 = ~n956 ;
  assign n957 = n177 & n1436 ;
  assign n958 = n945 | n957 ;
  assign n1437 = ~n169 ;
  assign n959 = n1437 & n958 ;
  assign n960 = x83 | n841 ;
  assign n961 = x82 | n960 ;
  assign n962 = x81 | n961 ;
  assign n963 = x80 | n962 ;
  assign n964 = n956 | n963 ;
  assign n965 = n958 & n963 ;
  assign n1438 = ~n965 ;
  assign n966 = n964 & n1438 ;
  assign n1439 = ~n966 ;
  assign n967 = n169 & n1439 ;
  assign n968 = n959 | n967 ;
  assign n976 = x59 | n869 ;
  assign n977 = x58 | n976 ;
  assign n978 = x57 | n977 ;
  assign n979 = x56 | n978 ;
  assign n1440 = ~n979 ;
  assign n980 = n968 & n1440 ;
  assign n969 = x67 | n859 ;
  assign n970 = x66 | n969 ;
  assign n971 = x65 | n970 ;
  assign n972 = x64 | n971 ;
  assign n973 = n966 | n972 ;
  assign n974 = n968 & n972 ;
  assign n1441 = ~n974 ;
  assign n975 = n973 & n1441 ;
  assign n1442 = ~n975 ;
  assign n981 = n1442 & n979 ;
  assign n982 = n980 | n981 ;
  assign n990 = x43 | n889 ;
  assign n991 = x42 | n990 ;
  assign n992 = x41 | n991 ;
  assign n993 = x40 | n992 ;
  assign n1443 = ~n993 ;
  assign n994 = n982 & n1443 ;
  assign n983 = x51 | n879 ;
  assign n984 = x50 | n983 ;
  assign n985 = x49 | n984 ;
  assign n986 = x48 | n985 ;
  assign n987 = n975 | n986 ;
  assign n988 = n982 & n986 ;
  assign n1444 = ~n988 ;
  assign n989 = n987 & n1444 ;
  assign n1445 = ~n989 ;
  assign n995 = n1445 & n993 ;
  assign n996 = n994 | n995 ;
  assign n1004 = x27 | n909 ;
  assign n1005 = x26 | n1004 ;
  assign n1006 = x25 | n1005 ;
  assign n1007 = x24 | n1006 ;
  assign n1446 = ~n1007 ;
  assign n1008 = n996 & n1446 ;
  assign n997 = x35 | n899 ;
  assign n998 = x34 | n997 ;
  assign n999 = x33 | n998 ;
  assign n1000 = x32 | n999 ;
  assign n1001 = n989 | n1000 ;
  assign n1002 = n996 & n1000 ;
  assign n1447 = ~n1002 ;
  assign n1003 = n1001 & n1447 ;
  assign n1448 = ~n1003 ;
  assign n1009 = n1448 & n1007 ;
  assign n1010 = n1008 | n1009 ;
  assign n1018 = x11 | n929 ;
  assign n1019 = x10 | n1018 ;
  assign n1020 = x9 | n1019 ;
  assign n1021 = x8 | n1020 ;
  assign n1449 = ~n1021 ;
  assign n1022 = n1010 & n1449 ;
  assign n1011 = x19 | n919 ;
  assign n1012 = x18 | n1011 ;
  assign n1013 = x17 | n1012 ;
  assign n1014 = x16 | n1013 ;
  assign n1015 = n1003 | n1014 ;
  assign n1016 = n1010 & n1014 ;
  assign n1450 = ~n1016 ;
  assign n1017 = n1015 & n1450 ;
  assign n1451 = ~n1017 ;
  assign n1023 = n1451 & n1021 ;
  assign n132 = n1022 | n1023 ;
  assign n145 = n1104 | n144 ;
  assign n149 = x99 | n148 ;
  assign n157 = x98 | n156 ;
  assign n159 = x97 | n157 ;
  assign n160 = x96 | n159 ;
  assign n161 = n149 | n160 ;
  assign n178 = x87 | n177 ;
  assign n179 = x86 | n178 ;
  assign n180 = x85 | n179 ;
  assign n181 = x84 | n180 ;
  assign n182 = x83 | n181 ;
  assign n183 = x82 | n182 ;
  assign n184 = x81 | n183 ;
  assign n185 = x80 | n184 ;
  assign n1452 = ~n161 ;
  assign n1025 = n1452 & n185 ;
  assign n1026 = n145 | n1025 ;
  assign n1046 = x55 | n979 ;
  assign n1047 = x54 | n1046 ;
  assign n1048 = x53 | n1047 ;
  assign n1049 = x52 | n1048 ;
  assign n1050 = x51 | n1049 ;
  assign n1051 = x50 | n1050 ;
  assign n1052 = x49 | n1051 ;
  assign n1053 = x48 | n1052 ;
  assign n1453 = ~n1053 ;
  assign n1054 = n1026 & n1453 ;
  assign n1027 = x77 | x78 ;
  assign n1028 = x76 | n1027 ;
  assign n1029 = x75 | n1028 ;
  assign n1030 = x74 | n1029 ;
  assign n1031 = x73 | n1030 ;
  assign n1032 = x72 | n1031 ;
  assign n1033 = x71 | n1032 ;
  assign n1034 = x70 | n1033 ;
  assign n1035 = x69 | n1034 ;
  assign n1036 = x68 | n1035 ;
  assign n1037 = x67 | n1036 ;
  assign n1038 = x66 | n1037 ;
  assign n1039 = x65 | n1038 ;
  assign n1040 = x64 | n1039 ;
  assign n1041 = n1026 & n1040 ;
  assign n1454 = ~n185 ;
  assign n187 = x79 & n1454 ;
  assign n1042 = n161 | n187 ;
  assign n1455 = ~n145 ;
  assign n1043 = n1455 & n1042 ;
  assign n1044 = n1040 | n1043 ;
  assign n1456 = ~n1041 ;
  assign n1045 = n1456 & n1044 ;
  assign n1457 = ~n1045 ;
  assign n1055 = n1457 & n1053 ;
  assign n1056 = n1054 | n1055 ;
  assign n1068 = x23 | n1007 ;
  assign n1069 = x22 | n1068 ;
  assign n1070 = x21 | n1069 ;
  assign n1071 = x20 | n1070 ;
  assign n1072 = x19 | n1071 ;
  assign n1073 = x18 | n1072 ;
  assign n1074 = x17 | n1073 ;
  assign n1075 = x16 | n1074 ;
  assign n1458 = ~n1075 ;
  assign n1076 = n1056 & n1458 ;
  assign n1057 = x39 | n993 ;
  assign n1058 = x38 | n1057 ;
  assign n1059 = x37 | n1058 ;
  assign n1060 = x36 | n1059 ;
  assign n1061 = x35 | n1060 ;
  assign n1062 = x34 | n1061 ;
  assign n1063 = x33 | n1062 ;
  assign n1064 = x32 | n1063 ;
  assign n1065 = n1045 | n1064 ;
  assign n1066 = n1056 & n1064 ;
  assign n1459 = ~n1066 ;
  assign n1067 = n1065 & n1459 ;
  assign n1460 = ~n1067 ;
  assign n1077 = n1460 & n1075 ;
  assign n133 = n1076 | n1077 ;
  assign n162 = n145 | n161 ;
  assign n170 = x71 | n169 ;
  assign n186 = x70 | n185 ;
  assign n188 = x69 | n186 ;
  assign n189 = x68 | n188 ;
  assign n190 = x67 | n189 ;
  assign n191 = x66 | n190 ;
  assign n192 = x65 | n191 ;
  assign n193 = x64 | n192 ;
  assign n194 = n170 | n193 ;
  assign n1079 = x47 | n1053 ;
  assign n1080 = x46 | n1079 ;
  assign n1081 = x45 | n1080 ;
  assign n1082 = x44 | n1081 ;
  assign n1083 = x43 | n1082 ;
  assign n1084 = x42 | n1083 ;
  assign n1085 = x41 | n1084 ;
  assign n1086 = x40 | n1085 ;
  assign n1087 = x39 | n1086 ;
  assign n1088 = x38 | n1087 ;
  assign n1089 = x37 | n1088 ;
  assign n1090 = x36 | n1089 ;
  assign n1091 = x35 | n1090 ;
  assign n1092 = x34 | n1091 ;
  assign n1093 = x33 | n1092 ;
  assign n1094 = x32 | n1093 ;
  assign n1461 = ~n194 ;
  assign n1097 = n1461 & n1094 ;
  assign n134 = n162 | n1097 ;
  assign n135 = n162 | n194 ;
  assign n1099 = x0 | n135 ;
  assign n1100 = n1021 | n1099 ;
  assign n1101 = x3 | n1100 ;
  assign n1102 = x2 | n1101 ;
  assign n1095 = n1075 | n1094 ;
  assign n1096 = n939 | n1095 ;
  assign n1103 = x1 | n1096 ;
  assign n136 = n1102 | n1103 ;
  assign y0 = n129 ;
  assign y1 = n130 ;
  assign y2 = n131 ;
  assign y3 = n132 ;
  assign y4 = n133 ;
  assign y5 = n134 ;
  assign y6 = n135 ;
  assign y7 = n136 ;
endmodule
