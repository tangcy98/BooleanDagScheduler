module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 ;
  assign n257 = x128 ^ x0 ^ 1'b0 ;
  assign n258 = x0 & x128 ;
  assign n259 = n258 ^ x129 ^ x1 ;
  assign n260 = ( x1 & x129 ) | ( x1 & n258 ) | ( x129 & n258 ) ;
  assign n261 = n260 ^ x130 ^ x2 ;
  assign n265 = ( x2 & x130 ) | ( x2 & n260 ) | ( x130 & n260 ) ;
  assign n262 = x3 | x131 ;
  assign n263 = x3 & x131 ;
  assign n264 = n262 & ~n263 ;
  assign n266 = n265 ^ n264 ^ 1'b0 ;
  assign n270 = ( x3 & x131 ) | ( x3 & n265 ) | ( x131 & n265 ) ;
  assign n267 = x4 | x132 ;
  assign n268 = x4 & x132 ;
  assign n269 = n267 & ~n268 ;
  assign n271 = n270 ^ n269 ^ 1'b0 ;
  assign n275 = ( x4 & x132 ) | ( x4 & n270 ) | ( x132 & n270 ) ;
  assign n272 = x5 | x133 ;
  assign n273 = x5 & x133 ;
  assign n274 = n272 & ~n273 ;
  assign n276 = n275 ^ n274 ^ 1'b0 ;
  assign n280 = ( x5 & x133 ) | ( x5 & n275 ) | ( x133 & n275 ) ;
  assign n277 = x6 | x134 ;
  assign n278 = x6 & x134 ;
  assign n279 = n277 & ~n278 ;
  assign n281 = n280 ^ n279 ^ 1'b0 ;
  assign n285 = ( x6 & x134 ) | ( x6 & n280 ) | ( x134 & n280 ) ;
  assign n282 = x7 | x135 ;
  assign n283 = x7 & x135 ;
  assign n284 = n282 & ~n283 ;
  assign n286 = n285 ^ n284 ^ 1'b0 ;
  assign n290 = ( x7 & x135 ) | ( x7 & n285 ) | ( x135 & n285 ) ;
  assign n287 = x8 | x136 ;
  assign n288 = x8 & x136 ;
  assign n289 = n287 & ~n288 ;
  assign n291 = n290 ^ n289 ^ 1'b0 ;
  assign n295 = ( x8 & x136 ) | ( x8 & n290 ) | ( x136 & n290 ) ;
  assign n292 = x9 | x137 ;
  assign n293 = x9 & x137 ;
  assign n294 = n292 & ~n293 ;
  assign n296 = n295 ^ n294 ^ 1'b0 ;
  assign n300 = ( x9 & x137 ) | ( x9 & n295 ) | ( x137 & n295 ) ;
  assign n297 = x10 | x138 ;
  assign n298 = x10 & x138 ;
  assign n299 = n297 & ~n298 ;
  assign n301 = n300 ^ n299 ^ 1'b0 ;
  assign n305 = ( x10 & x138 ) | ( x10 & n300 ) | ( x138 & n300 ) ;
  assign n302 = x11 | x139 ;
  assign n303 = x11 & x139 ;
  assign n304 = n302 & ~n303 ;
  assign n306 = n305 ^ n304 ^ 1'b0 ;
  assign n310 = ( x11 & x139 ) | ( x11 & n305 ) | ( x139 & n305 ) ;
  assign n307 = x12 | x140 ;
  assign n308 = x12 & x140 ;
  assign n309 = n307 & ~n308 ;
  assign n311 = n310 ^ n309 ^ 1'b0 ;
  assign n315 = ( x12 & x140 ) | ( x12 & n310 ) | ( x140 & n310 ) ;
  assign n312 = x13 | x141 ;
  assign n313 = x13 & x141 ;
  assign n314 = n312 & ~n313 ;
  assign n316 = n315 ^ n314 ^ 1'b0 ;
  assign n320 = ( x13 & x141 ) | ( x13 & n315 ) | ( x141 & n315 ) ;
  assign n317 = x14 | x142 ;
  assign n318 = x14 & x142 ;
  assign n319 = n317 & ~n318 ;
  assign n321 = n320 ^ n319 ^ 1'b0 ;
  assign n325 = ( x14 & x142 ) | ( x14 & n320 ) | ( x142 & n320 ) ;
  assign n322 = x15 | x143 ;
  assign n323 = x15 & x143 ;
  assign n324 = n322 & ~n323 ;
  assign n326 = n325 ^ n324 ^ 1'b0 ;
  assign n330 = ( x15 & x143 ) | ( x15 & n325 ) | ( x143 & n325 ) ;
  assign n327 = x16 | x144 ;
  assign n328 = x16 & x144 ;
  assign n329 = n327 & ~n328 ;
  assign n331 = n330 ^ n329 ^ 1'b0 ;
  assign n335 = ( x16 & x144 ) | ( x16 & n330 ) | ( x144 & n330 ) ;
  assign n332 = x17 | x145 ;
  assign n333 = x17 & x145 ;
  assign n334 = n332 & ~n333 ;
  assign n336 = n335 ^ n334 ^ 1'b0 ;
  assign n340 = ( x17 & x145 ) | ( x17 & n335 ) | ( x145 & n335 ) ;
  assign n337 = x18 | x146 ;
  assign n338 = x18 & x146 ;
  assign n339 = n337 & ~n338 ;
  assign n341 = n340 ^ n339 ^ 1'b0 ;
  assign n345 = ( x18 & x146 ) | ( x18 & n340 ) | ( x146 & n340 ) ;
  assign n342 = x19 | x147 ;
  assign n343 = x19 & x147 ;
  assign n344 = n342 & ~n343 ;
  assign n346 = n345 ^ n344 ^ 1'b0 ;
  assign n350 = ( x19 & x147 ) | ( x19 & n345 ) | ( x147 & n345 ) ;
  assign n347 = x20 | x148 ;
  assign n348 = x20 & x148 ;
  assign n349 = n347 & ~n348 ;
  assign n351 = n350 ^ n349 ^ 1'b0 ;
  assign n355 = ( x20 & x148 ) | ( x20 & n350 ) | ( x148 & n350 ) ;
  assign n352 = x21 | x149 ;
  assign n353 = x21 & x149 ;
  assign n354 = n352 & ~n353 ;
  assign n356 = n355 ^ n354 ^ 1'b0 ;
  assign n360 = ( x21 & x149 ) | ( x21 & n355 ) | ( x149 & n355 ) ;
  assign n357 = x22 | x150 ;
  assign n358 = x22 & x150 ;
  assign n359 = n357 & ~n358 ;
  assign n361 = n360 ^ n359 ^ 1'b0 ;
  assign n365 = ( x22 & x150 ) | ( x22 & n360 ) | ( x150 & n360 ) ;
  assign n362 = x23 | x151 ;
  assign n363 = x23 & x151 ;
  assign n364 = n362 & ~n363 ;
  assign n366 = n365 ^ n364 ^ 1'b0 ;
  assign n370 = ( x23 & x151 ) | ( x23 & n365 ) | ( x151 & n365 ) ;
  assign n367 = x24 | x152 ;
  assign n368 = x24 & x152 ;
  assign n369 = n367 & ~n368 ;
  assign n371 = n370 ^ n369 ^ 1'b0 ;
  assign n375 = ( x24 & x152 ) | ( x24 & n370 ) | ( x152 & n370 ) ;
  assign n372 = x25 | x153 ;
  assign n373 = x25 & x153 ;
  assign n374 = n372 & ~n373 ;
  assign n376 = n375 ^ n374 ^ 1'b0 ;
  assign n380 = ( x25 & x153 ) | ( x25 & n375 ) | ( x153 & n375 ) ;
  assign n377 = x26 | x154 ;
  assign n378 = x26 & x154 ;
  assign n379 = n377 & ~n378 ;
  assign n381 = n380 ^ n379 ^ 1'b0 ;
  assign n385 = ( x26 & x154 ) | ( x26 & n380 ) | ( x154 & n380 ) ;
  assign n382 = x27 | x155 ;
  assign n383 = x27 & x155 ;
  assign n384 = n382 & ~n383 ;
  assign n386 = n385 ^ n384 ^ 1'b0 ;
  assign n390 = ( x27 & x155 ) | ( x27 & n385 ) | ( x155 & n385 ) ;
  assign n387 = x28 | x156 ;
  assign n388 = x28 & x156 ;
  assign n389 = n387 & ~n388 ;
  assign n391 = n390 ^ n389 ^ 1'b0 ;
  assign n395 = ( x28 & x156 ) | ( x28 & n390 ) | ( x156 & n390 ) ;
  assign n392 = x29 | x157 ;
  assign n393 = x29 & x157 ;
  assign n394 = n392 & ~n393 ;
  assign n396 = n395 ^ n394 ^ 1'b0 ;
  assign n400 = ( x29 & x157 ) | ( x29 & n395 ) | ( x157 & n395 ) ;
  assign n397 = x30 | x158 ;
  assign n398 = x30 & x158 ;
  assign n399 = n397 & ~n398 ;
  assign n401 = n400 ^ n399 ^ 1'b0 ;
  assign n405 = ( x30 & x158 ) | ( x30 & n400 ) | ( x158 & n400 ) ;
  assign n402 = x31 | x159 ;
  assign n403 = x31 & x159 ;
  assign n404 = n402 & ~n403 ;
  assign n406 = n405 ^ n404 ^ 1'b0 ;
  assign n410 = ( x31 & x159 ) | ( x31 & n405 ) | ( x159 & n405 ) ;
  assign n407 = x32 | x160 ;
  assign n408 = x32 & x160 ;
  assign n409 = n407 & ~n408 ;
  assign n411 = n410 ^ n409 ^ 1'b0 ;
  assign n415 = ( x32 & x160 ) | ( x32 & n410 ) | ( x160 & n410 ) ;
  assign n412 = x33 | x161 ;
  assign n413 = x33 & x161 ;
  assign n414 = n412 & ~n413 ;
  assign n416 = n415 ^ n414 ^ 1'b0 ;
  assign n420 = ( x33 & x161 ) | ( x33 & n415 ) | ( x161 & n415 ) ;
  assign n417 = x34 | x162 ;
  assign n418 = x34 & x162 ;
  assign n419 = n417 & ~n418 ;
  assign n421 = n420 ^ n419 ^ 1'b0 ;
  assign n425 = ( x34 & x162 ) | ( x34 & n420 ) | ( x162 & n420 ) ;
  assign n422 = x35 | x163 ;
  assign n423 = x35 & x163 ;
  assign n424 = n422 & ~n423 ;
  assign n426 = n425 ^ n424 ^ 1'b0 ;
  assign n430 = ( x35 & x163 ) | ( x35 & n425 ) | ( x163 & n425 ) ;
  assign n427 = x36 | x164 ;
  assign n428 = x36 & x164 ;
  assign n429 = n427 & ~n428 ;
  assign n431 = n430 ^ n429 ^ 1'b0 ;
  assign n435 = ( x36 & x164 ) | ( x36 & n430 ) | ( x164 & n430 ) ;
  assign n432 = x37 | x165 ;
  assign n433 = x37 & x165 ;
  assign n434 = n432 & ~n433 ;
  assign n436 = n435 ^ n434 ^ 1'b0 ;
  assign n440 = ( x37 & x165 ) | ( x37 & n435 ) | ( x165 & n435 ) ;
  assign n437 = x38 | x166 ;
  assign n438 = x38 & x166 ;
  assign n439 = n437 & ~n438 ;
  assign n441 = n440 ^ n439 ^ 1'b0 ;
  assign n445 = ( x38 & x166 ) | ( x38 & n440 ) | ( x166 & n440 ) ;
  assign n442 = x39 | x167 ;
  assign n443 = x39 & x167 ;
  assign n444 = n442 & ~n443 ;
  assign n446 = n445 ^ n444 ^ 1'b0 ;
  assign n450 = ( x39 & x167 ) | ( x39 & n445 ) | ( x167 & n445 ) ;
  assign n447 = x40 | x168 ;
  assign n448 = x40 & x168 ;
  assign n449 = n447 & ~n448 ;
  assign n451 = n450 ^ n449 ^ 1'b0 ;
  assign n455 = ( x40 & x168 ) | ( x40 & n450 ) | ( x168 & n450 ) ;
  assign n452 = x41 | x169 ;
  assign n453 = x41 & x169 ;
  assign n454 = n452 & ~n453 ;
  assign n456 = n455 ^ n454 ^ 1'b0 ;
  assign n460 = ( x41 & x169 ) | ( x41 & n455 ) | ( x169 & n455 ) ;
  assign n457 = x42 | x170 ;
  assign n458 = x42 & x170 ;
  assign n459 = n457 & ~n458 ;
  assign n461 = n460 ^ n459 ^ 1'b0 ;
  assign n465 = ( x42 & x170 ) | ( x42 & n460 ) | ( x170 & n460 ) ;
  assign n462 = x43 | x171 ;
  assign n463 = x43 & x171 ;
  assign n464 = n462 & ~n463 ;
  assign n466 = n465 ^ n464 ^ 1'b0 ;
  assign n470 = ( x43 & x171 ) | ( x43 & n465 ) | ( x171 & n465 ) ;
  assign n467 = x44 | x172 ;
  assign n468 = x44 & x172 ;
  assign n469 = n467 & ~n468 ;
  assign n471 = n470 ^ n469 ^ 1'b0 ;
  assign n475 = ( x44 & x172 ) | ( x44 & n470 ) | ( x172 & n470 ) ;
  assign n472 = x45 | x173 ;
  assign n473 = x45 & x173 ;
  assign n474 = n472 & ~n473 ;
  assign n476 = n475 ^ n474 ^ 1'b0 ;
  assign n480 = ( x45 & x173 ) | ( x45 & n475 ) | ( x173 & n475 ) ;
  assign n477 = x46 | x174 ;
  assign n478 = x46 & x174 ;
  assign n479 = n477 & ~n478 ;
  assign n481 = n480 ^ n479 ^ 1'b0 ;
  assign n485 = ( x46 & x174 ) | ( x46 & n480 ) | ( x174 & n480 ) ;
  assign n482 = x47 | x175 ;
  assign n483 = x47 & x175 ;
  assign n484 = n482 & ~n483 ;
  assign n486 = n485 ^ n484 ^ 1'b0 ;
  assign n490 = ( x47 & x175 ) | ( x47 & n485 ) | ( x175 & n485 ) ;
  assign n487 = x48 | x176 ;
  assign n488 = x48 & x176 ;
  assign n489 = n487 & ~n488 ;
  assign n491 = n490 ^ n489 ^ 1'b0 ;
  assign n495 = ( x48 & x176 ) | ( x48 & n490 ) | ( x176 & n490 ) ;
  assign n492 = x49 | x177 ;
  assign n493 = x49 & x177 ;
  assign n494 = n492 & ~n493 ;
  assign n496 = n495 ^ n494 ^ 1'b0 ;
  assign n500 = ( x49 & x177 ) | ( x49 & n495 ) | ( x177 & n495 ) ;
  assign n497 = x50 | x178 ;
  assign n498 = x50 & x178 ;
  assign n499 = n497 & ~n498 ;
  assign n501 = n500 ^ n499 ^ 1'b0 ;
  assign n505 = ( x50 & x178 ) | ( x50 & n500 ) | ( x178 & n500 ) ;
  assign n502 = x51 | x179 ;
  assign n503 = x51 & x179 ;
  assign n504 = n502 & ~n503 ;
  assign n506 = n505 ^ n504 ^ 1'b0 ;
  assign n510 = ( x51 & x179 ) | ( x51 & n505 ) | ( x179 & n505 ) ;
  assign n507 = x52 | x180 ;
  assign n508 = x52 & x180 ;
  assign n509 = n507 & ~n508 ;
  assign n511 = n510 ^ n509 ^ 1'b0 ;
  assign n515 = ( x52 & x180 ) | ( x52 & n510 ) | ( x180 & n510 ) ;
  assign n512 = x53 | x181 ;
  assign n513 = x53 & x181 ;
  assign n514 = n512 & ~n513 ;
  assign n516 = n515 ^ n514 ^ 1'b0 ;
  assign n520 = ( x53 & x181 ) | ( x53 & n515 ) | ( x181 & n515 ) ;
  assign n517 = x54 | x182 ;
  assign n518 = x54 & x182 ;
  assign n519 = n517 & ~n518 ;
  assign n521 = n520 ^ n519 ^ 1'b0 ;
  assign n525 = ( x54 & x182 ) | ( x54 & n520 ) | ( x182 & n520 ) ;
  assign n522 = x55 | x183 ;
  assign n523 = x55 & x183 ;
  assign n524 = n522 & ~n523 ;
  assign n526 = n525 ^ n524 ^ 1'b0 ;
  assign n530 = ( x55 & x183 ) | ( x55 & n525 ) | ( x183 & n525 ) ;
  assign n527 = x56 | x184 ;
  assign n528 = x56 & x184 ;
  assign n529 = n527 & ~n528 ;
  assign n531 = n530 ^ n529 ^ 1'b0 ;
  assign n535 = ( x56 & x184 ) | ( x56 & n530 ) | ( x184 & n530 ) ;
  assign n532 = x57 | x185 ;
  assign n533 = x57 & x185 ;
  assign n534 = n532 & ~n533 ;
  assign n536 = n535 ^ n534 ^ 1'b0 ;
  assign n540 = ( x57 & x185 ) | ( x57 & n535 ) | ( x185 & n535 ) ;
  assign n537 = x58 | x186 ;
  assign n538 = x58 & x186 ;
  assign n539 = n537 & ~n538 ;
  assign n541 = n540 ^ n539 ^ 1'b0 ;
  assign n545 = ( x58 & x186 ) | ( x58 & n540 ) | ( x186 & n540 ) ;
  assign n542 = x59 | x187 ;
  assign n543 = x59 & x187 ;
  assign n544 = n542 & ~n543 ;
  assign n546 = n545 ^ n544 ^ 1'b0 ;
  assign n550 = ( x59 & x187 ) | ( x59 & n545 ) | ( x187 & n545 ) ;
  assign n547 = x60 | x188 ;
  assign n548 = x60 & x188 ;
  assign n549 = n547 & ~n548 ;
  assign n551 = n550 ^ n549 ^ 1'b0 ;
  assign n555 = ( x60 & x188 ) | ( x60 & n550 ) | ( x188 & n550 ) ;
  assign n552 = x61 | x189 ;
  assign n553 = x61 & x189 ;
  assign n554 = n552 & ~n553 ;
  assign n556 = n555 ^ n554 ^ 1'b0 ;
  assign n560 = ( x61 & x189 ) | ( x61 & n555 ) | ( x189 & n555 ) ;
  assign n557 = x62 | x190 ;
  assign n558 = x62 & x190 ;
  assign n559 = n557 & ~n558 ;
  assign n561 = n560 ^ n559 ^ 1'b0 ;
  assign n565 = ( x62 & x190 ) | ( x62 & n560 ) | ( x190 & n560 ) ;
  assign n562 = x63 | x191 ;
  assign n563 = x63 & x191 ;
  assign n564 = n562 & ~n563 ;
  assign n566 = n565 ^ n564 ^ 1'b0 ;
  assign n570 = ( x63 & x191 ) | ( x63 & n565 ) | ( x191 & n565 ) ;
  assign n567 = x64 | x192 ;
  assign n568 = x64 & x192 ;
  assign n569 = n567 & ~n568 ;
  assign n571 = n570 ^ n569 ^ 1'b0 ;
  assign n575 = ( x64 & x192 ) | ( x64 & n570 ) | ( x192 & n570 ) ;
  assign n572 = x65 | x193 ;
  assign n573 = x65 & x193 ;
  assign n574 = n572 & ~n573 ;
  assign n576 = n575 ^ n574 ^ 1'b0 ;
  assign n580 = ( x65 & x193 ) | ( x65 & n575 ) | ( x193 & n575 ) ;
  assign n577 = x66 | x194 ;
  assign n578 = x66 & x194 ;
  assign n579 = n577 & ~n578 ;
  assign n581 = n580 ^ n579 ^ 1'b0 ;
  assign n585 = ( x66 & x194 ) | ( x66 & n580 ) | ( x194 & n580 ) ;
  assign n582 = x67 | x195 ;
  assign n583 = x67 & x195 ;
  assign n584 = n582 & ~n583 ;
  assign n586 = n585 ^ n584 ^ 1'b0 ;
  assign n590 = ( x67 & x195 ) | ( x67 & n585 ) | ( x195 & n585 ) ;
  assign n587 = x68 | x196 ;
  assign n588 = x68 & x196 ;
  assign n589 = n587 & ~n588 ;
  assign n591 = n590 ^ n589 ^ 1'b0 ;
  assign n595 = ( x68 & x196 ) | ( x68 & n590 ) | ( x196 & n590 ) ;
  assign n592 = x69 | x197 ;
  assign n593 = x69 & x197 ;
  assign n594 = n592 & ~n593 ;
  assign n596 = n595 ^ n594 ^ 1'b0 ;
  assign n600 = ( x69 & x197 ) | ( x69 & n595 ) | ( x197 & n595 ) ;
  assign n597 = x70 | x198 ;
  assign n598 = x70 & x198 ;
  assign n599 = n597 & ~n598 ;
  assign n601 = n600 ^ n599 ^ 1'b0 ;
  assign n605 = ( x70 & x198 ) | ( x70 & n600 ) | ( x198 & n600 ) ;
  assign n602 = x71 | x199 ;
  assign n603 = x71 & x199 ;
  assign n604 = n602 & ~n603 ;
  assign n606 = n605 ^ n604 ^ 1'b0 ;
  assign n610 = ( x71 & x199 ) | ( x71 & n605 ) | ( x199 & n605 ) ;
  assign n607 = x72 | x200 ;
  assign n608 = x72 & x200 ;
  assign n609 = n607 & ~n608 ;
  assign n611 = n610 ^ n609 ^ 1'b0 ;
  assign n615 = ( x72 & x200 ) | ( x72 & n610 ) | ( x200 & n610 ) ;
  assign n612 = x73 | x201 ;
  assign n613 = x73 & x201 ;
  assign n614 = n612 & ~n613 ;
  assign n616 = n615 ^ n614 ^ 1'b0 ;
  assign n620 = ( x73 & x201 ) | ( x73 & n615 ) | ( x201 & n615 ) ;
  assign n617 = x74 | x202 ;
  assign n618 = x74 & x202 ;
  assign n619 = n617 & ~n618 ;
  assign n621 = n620 ^ n619 ^ 1'b0 ;
  assign n625 = ( x74 & x202 ) | ( x74 & n620 ) | ( x202 & n620 ) ;
  assign n622 = x75 | x203 ;
  assign n623 = x75 & x203 ;
  assign n624 = n622 & ~n623 ;
  assign n626 = n625 ^ n624 ^ 1'b0 ;
  assign n630 = ( x75 & x203 ) | ( x75 & n625 ) | ( x203 & n625 ) ;
  assign n627 = x76 | x204 ;
  assign n628 = x76 & x204 ;
  assign n629 = n627 & ~n628 ;
  assign n631 = n630 ^ n629 ^ 1'b0 ;
  assign n635 = ( x76 & x204 ) | ( x76 & n630 ) | ( x204 & n630 ) ;
  assign n632 = x77 | x205 ;
  assign n633 = x77 & x205 ;
  assign n634 = n632 & ~n633 ;
  assign n636 = n635 ^ n634 ^ 1'b0 ;
  assign n640 = ( x77 & x205 ) | ( x77 & n635 ) | ( x205 & n635 ) ;
  assign n637 = x78 | x206 ;
  assign n638 = x78 & x206 ;
  assign n639 = n637 & ~n638 ;
  assign n641 = n640 ^ n639 ^ 1'b0 ;
  assign n645 = ( x78 & x206 ) | ( x78 & n640 ) | ( x206 & n640 ) ;
  assign n642 = x79 | x207 ;
  assign n643 = x79 & x207 ;
  assign n644 = n642 & ~n643 ;
  assign n646 = n645 ^ n644 ^ 1'b0 ;
  assign n650 = ( x79 & x207 ) | ( x79 & n645 ) | ( x207 & n645 ) ;
  assign n647 = x80 | x208 ;
  assign n648 = x80 & x208 ;
  assign n649 = n647 & ~n648 ;
  assign n651 = n650 ^ n649 ^ 1'b0 ;
  assign n655 = ( x80 & x208 ) | ( x80 & n650 ) | ( x208 & n650 ) ;
  assign n652 = x81 | x209 ;
  assign n653 = x81 & x209 ;
  assign n654 = n652 & ~n653 ;
  assign n656 = n655 ^ n654 ^ 1'b0 ;
  assign n660 = ( x81 & x209 ) | ( x81 & n655 ) | ( x209 & n655 ) ;
  assign n657 = x82 | x210 ;
  assign n658 = x82 & x210 ;
  assign n659 = n657 & ~n658 ;
  assign n661 = n660 ^ n659 ^ 1'b0 ;
  assign n665 = ( x82 & x210 ) | ( x82 & n660 ) | ( x210 & n660 ) ;
  assign n662 = x83 | x211 ;
  assign n663 = x83 & x211 ;
  assign n664 = n662 & ~n663 ;
  assign n666 = n665 ^ n664 ^ 1'b0 ;
  assign n670 = ( x83 & x211 ) | ( x83 & n665 ) | ( x211 & n665 ) ;
  assign n667 = x84 | x212 ;
  assign n668 = x84 & x212 ;
  assign n669 = n667 & ~n668 ;
  assign n671 = n670 ^ n669 ^ 1'b0 ;
  assign n675 = ( x84 & x212 ) | ( x84 & n670 ) | ( x212 & n670 ) ;
  assign n672 = x85 | x213 ;
  assign n673 = x85 & x213 ;
  assign n674 = n672 & ~n673 ;
  assign n676 = n675 ^ n674 ^ 1'b0 ;
  assign n680 = ( x85 & x213 ) | ( x85 & n675 ) | ( x213 & n675 ) ;
  assign n677 = x86 | x214 ;
  assign n678 = x86 & x214 ;
  assign n679 = n677 & ~n678 ;
  assign n681 = n680 ^ n679 ^ 1'b0 ;
  assign n685 = ( x86 & x214 ) | ( x86 & n680 ) | ( x214 & n680 ) ;
  assign n682 = x87 | x215 ;
  assign n683 = x87 & x215 ;
  assign n684 = n682 & ~n683 ;
  assign n686 = n685 ^ n684 ^ 1'b0 ;
  assign n690 = ( x87 & x215 ) | ( x87 & n685 ) | ( x215 & n685 ) ;
  assign n687 = x88 | x216 ;
  assign n688 = x88 & x216 ;
  assign n689 = n687 & ~n688 ;
  assign n691 = n690 ^ n689 ^ 1'b0 ;
  assign n695 = ( x88 & x216 ) | ( x88 & n690 ) | ( x216 & n690 ) ;
  assign n692 = x89 | x217 ;
  assign n693 = x89 & x217 ;
  assign n694 = n692 & ~n693 ;
  assign n696 = n695 ^ n694 ^ 1'b0 ;
  assign n700 = ( x89 & x217 ) | ( x89 & n695 ) | ( x217 & n695 ) ;
  assign n697 = x90 | x218 ;
  assign n698 = x90 & x218 ;
  assign n699 = n697 & ~n698 ;
  assign n701 = n700 ^ n699 ^ 1'b0 ;
  assign n705 = ( x90 & x218 ) | ( x90 & n700 ) | ( x218 & n700 ) ;
  assign n702 = x91 | x219 ;
  assign n703 = x91 & x219 ;
  assign n704 = n702 & ~n703 ;
  assign n706 = n705 ^ n704 ^ 1'b0 ;
  assign n710 = ( x91 & x219 ) | ( x91 & n705 ) | ( x219 & n705 ) ;
  assign n707 = x92 | x220 ;
  assign n708 = x92 & x220 ;
  assign n709 = n707 & ~n708 ;
  assign n711 = n710 ^ n709 ^ 1'b0 ;
  assign n715 = ( x92 & x220 ) | ( x92 & n710 ) | ( x220 & n710 ) ;
  assign n712 = x93 | x221 ;
  assign n713 = x93 & x221 ;
  assign n714 = n712 & ~n713 ;
  assign n716 = n715 ^ n714 ^ 1'b0 ;
  assign n720 = ( x93 & x221 ) | ( x93 & n715 ) | ( x221 & n715 ) ;
  assign n717 = x94 | x222 ;
  assign n718 = x94 & x222 ;
  assign n719 = n717 & ~n718 ;
  assign n721 = n720 ^ n719 ^ 1'b0 ;
  assign n725 = ( x94 & x222 ) | ( x94 & n720 ) | ( x222 & n720 ) ;
  assign n722 = x95 | x223 ;
  assign n723 = x95 & x223 ;
  assign n724 = n722 & ~n723 ;
  assign n726 = n725 ^ n724 ^ 1'b0 ;
  assign n730 = ( x95 & x223 ) | ( x95 & n725 ) | ( x223 & n725 ) ;
  assign n727 = x96 | x224 ;
  assign n728 = x96 & x224 ;
  assign n729 = n727 & ~n728 ;
  assign n731 = n730 ^ n729 ^ 1'b0 ;
  assign n735 = ( x96 & x224 ) | ( x96 & n730 ) | ( x224 & n730 ) ;
  assign n732 = x97 | x225 ;
  assign n733 = x97 & x225 ;
  assign n734 = n732 & ~n733 ;
  assign n736 = n735 ^ n734 ^ 1'b0 ;
  assign n740 = ( x97 & x225 ) | ( x97 & n735 ) | ( x225 & n735 ) ;
  assign n737 = x98 | x226 ;
  assign n738 = x98 & x226 ;
  assign n739 = n737 & ~n738 ;
  assign n741 = n740 ^ n739 ^ 1'b0 ;
  assign n745 = ( x98 & x226 ) | ( x98 & n740 ) | ( x226 & n740 ) ;
  assign n742 = x99 | x227 ;
  assign n743 = x99 & x227 ;
  assign n744 = n742 & ~n743 ;
  assign n746 = n745 ^ n744 ^ 1'b0 ;
  assign n750 = ( x99 & x227 ) | ( x99 & n745 ) | ( x227 & n745 ) ;
  assign n747 = x100 | x228 ;
  assign n748 = x100 & x228 ;
  assign n749 = n747 & ~n748 ;
  assign n751 = n750 ^ n749 ^ 1'b0 ;
  assign n755 = ( x100 & x228 ) | ( x100 & n750 ) | ( x228 & n750 ) ;
  assign n752 = x101 | x229 ;
  assign n753 = x101 & x229 ;
  assign n754 = n752 & ~n753 ;
  assign n756 = n755 ^ n754 ^ 1'b0 ;
  assign n760 = ( x101 & x229 ) | ( x101 & n755 ) | ( x229 & n755 ) ;
  assign n757 = x102 | x230 ;
  assign n758 = x102 & x230 ;
  assign n759 = n757 & ~n758 ;
  assign n761 = n760 ^ n759 ^ 1'b0 ;
  assign n765 = ( x102 & x230 ) | ( x102 & n760 ) | ( x230 & n760 ) ;
  assign n762 = x103 | x231 ;
  assign n763 = x103 & x231 ;
  assign n764 = n762 & ~n763 ;
  assign n766 = n765 ^ n764 ^ 1'b0 ;
  assign n770 = ( x103 & x231 ) | ( x103 & n765 ) | ( x231 & n765 ) ;
  assign n767 = x104 | x232 ;
  assign n768 = x104 & x232 ;
  assign n769 = n767 & ~n768 ;
  assign n771 = n770 ^ n769 ^ 1'b0 ;
  assign n775 = ( x104 & x232 ) | ( x104 & n770 ) | ( x232 & n770 ) ;
  assign n772 = x105 | x233 ;
  assign n773 = x105 & x233 ;
  assign n774 = n772 & ~n773 ;
  assign n776 = n775 ^ n774 ^ 1'b0 ;
  assign n780 = ( x105 & x233 ) | ( x105 & n775 ) | ( x233 & n775 ) ;
  assign n777 = x106 | x234 ;
  assign n778 = x106 & x234 ;
  assign n779 = n777 & ~n778 ;
  assign n781 = n780 ^ n779 ^ 1'b0 ;
  assign n785 = ( x106 & x234 ) | ( x106 & n780 ) | ( x234 & n780 ) ;
  assign n782 = x107 | x235 ;
  assign n783 = x107 & x235 ;
  assign n784 = n782 & ~n783 ;
  assign n786 = n785 ^ n784 ^ 1'b0 ;
  assign n790 = ( x107 & x235 ) | ( x107 & n785 ) | ( x235 & n785 ) ;
  assign n787 = x108 | x236 ;
  assign n788 = x108 & x236 ;
  assign n789 = n787 & ~n788 ;
  assign n791 = n790 ^ n789 ^ 1'b0 ;
  assign n795 = ( x108 & x236 ) | ( x108 & n790 ) | ( x236 & n790 ) ;
  assign n792 = x109 | x237 ;
  assign n793 = x109 & x237 ;
  assign n794 = n792 & ~n793 ;
  assign n796 = n795 ^ n794 ^ 1'b0 ;
  assign n800 = ( x109 & x237 ) | ( x109 & n795 ) | ( x237 & n795 ) ;
  assign n797 = x110 | x238 ;
  assign n798 = x110 & x238 ;
  assign n799 = n797 & ~n798 ;
  assign n801 = n800 ^ n799 ^ 1'b0 ;
  assign n805 = ( x110 & x238 ) | ( x110 & n800 ) | ( x238 & n800 ) ;
  assign n802 = x111 | x239 ;
  assign n803 = x111 & x239 ;
  assign n804 = n802 & ~n803 ;
  assign n806 = n805 ^ n804 ^ 1'b0 ;
  assign n810 = ( x111 & x239 ) | ( x111 & n805 ) | ( x239 & n805 ) ;
  assign n807 = x112 | x240 ;
  assign n808 = x112 & x240 ;
  assign n809 = n807 & ~n808 ;
  assign n811 = n810 ^ n809 ^ 1'b0 ;
  assign n815 = ( x112 & x240 ) | ( x112 & n810 ) | ( x240 & n810 ) ;
  assign n812 = x113 | x241 ;
  assign n813 = x113 & x241 ;
  assign n814 = n812 & ~n813 ;
  assign n816 = n815 ^ n814 ^ 1'b0 ;
  assign n820 = ( x113 & x241 ) | ( x113 & n815 ) | ( x241 & n815 ) ;
  assign n817 = x114 | x242 ;
  assign n818 = x114 & x242 ;
  assign n819 = n817 & ~n818 ;
  assign n821 = n820 ^ n819 ^ 1'b0 ;
  assign n825 = ( x114 & x242 ) | ( x114 & n820 ) | ( x242 & n820 ) ;
  assign n822 = x115 | x243 ;
  assign n823 = x115 & x243 ;
  assign n824 = n822 & ~n823 ;
  assign n826 = n825 ^ n824 ^ 1'b0 ;
  assign n830 = ( x115 & x243 ) | ( x115 & n825 ) | ( x243 & n825 ) ;
  assign n827 = x116 | x244 ;
  assign n828 = x116 & x244 ;
  assign n829 = n827 & ~n828 ;
  assign n831 = n830 ^ n829 ^ 1'b0 ;
  assign n835 = ( x116 & x244 ) | ( x116 & n830 ) | ( x244 & n830 ) ;
  assign n832 = x117 | x245 ;
  assign n833 = x117 & x245 ;
  assign n834 = n832 & ~n833 ;
  assign n836 = n835 ^ n834 ^ 1'b0 ;
  assign n840 = ( x117 & x245 ) | ( x117 & n835 ) | ( x245 & n835 ) ;
  assign n837 = x118 | x246 ;
  assign n838 = x118 & x246 ;
  assign n839 = n837 & ~n838 ;
  assign n841 = n840 ^ n839 ^ 1'b0 ;
  assign n845 = ( x118 & x246 ) | ( x118 & n840 ) | ( x246 & n840 ) ;
  assign n842 = x119 | x247 ;
  assign n843 = x119 & x247 ;
  assign n844 = n842 & ~n843 ;
  assign n846 = n845 ^ n844 ^ 1'b0 ;
  assign n850 = ( x119 & x247 ) | ( x119 & n845 ) | ( x247 & n845 ) ;
  assign n847 = x120 | x248 ;
  assign n848 = x120 & x248 ;
  assign n849 = n847 & ~n848 ;
  assign n851 = n850 ^ n849 ^ 1'b0 ;
  assign n855 = ( x120 & x248 ) | ( x120 & n850 ) | ( x248 & n850 ) ;
  assign n852 = x121 | x249 ;
  assign n853 = x121 & x249 ;
  assign n854 = n852 & ~n853 ;
  assign n856 = n855 ^ n854 ^ 1'b0 ;
  assign n860 = ( x121 & x249 ) | ( x121 & n855 ) | ( x249 & n855 ) ;
  assign n857 = x122 | x250 ;
  assign n858 = x122 & x250 ;
  assign n859 = n857 & ~n858 ;
  assign n861 = n860 ^ n859 ^ 1'b0 ;
  assign n865 = ( x122 & x250 ) | ( x122 & n860 ) | ( x250 & n860 ) ;
  assign n862 = x123 | x251 ;
  assign n863 = x123 & x251 ;
  assign n864 = n862 & ~n863 ;
  assign n866 = n865 ^ n864 ^ 1'b0 ;
  assign n870 = ( x123 & x251 ) | ( x123 & n865 ) | ( x251 & n865 ) ;
  assign n867 = x124 | x252 ;
  assign n868 = x124 & x252 ;
  assign n869 = n867 & ~n868 ;
  assign n871 = n870 ^ n869 ^ 1'b0 ;
  assign n875 = ( x124 & x252 ) | ( x124 & n870 ) | ( x252 & n870 ) ;
  assign n872 = x125 | x253 ;
  assign n873 = x125 & x253 ;
  assign n874 = n872 & ~n873 ;
  assign n876 = n875 ^ n874 ^ 1'b0 ;
  assign n880 = ( x125 & x253 ) | ( x125 & n875 ) | ( x253 & n875 ) ;
  assign n877 = x126 | x254 ;
  assign n878 = x126 & x254 ;
  assign n879 = n877 & ~n878 ;
  assign n881 = n880 ^ n879 ^ 1'b0 ;
  assign n885 = ( x126 & x254 ) | ( x126 & n880 ) | ( x254 & n880 ) ;
  assign n882 = x127 | x255 ;
  assign n883 = x127 & x255 ;
  assign n884 = n882 & ~n883 ;
  assign n886 = n885 ^ n884 ^ 1'b0 ;
  assign n887 = ( x127 & x255 ) | ( x127 & n885 ) | ( x255 & n885 ) ;
  assign y0 = n257 ;
  assign y1 = n259 ;
  assign y2 = n261 ;
  assign y3 = n266 ;
  assign y4 = n271 ;
  assign y5 = n276 ;
  assign y6 = n281 ;
  assign y7 = n286 ;
  assign y8 = n291 ;
  assign y9 = n296 ;
  assign y10 = n301 ;
  assign y11 = n306 ;
  assign y12 = n311 ;
  assign y13 = n316 ;
  assign y14 = n321 ;
  assign y15 = n326 ;
  assign y16 = n331 ;
  assign y17 = n336 ;
  assign y18 = n341 ;
  assign y19 = n346 ;
  assign y20 = n351 ;
  assign y21 = n356 ;
  assign y22 = n361 ;
  assign y23 = n366 ;
  assign y24 = n371 ;
  assign y25 = n376 ;
  assign y26 = n381 ;
  assign y27 = n386 ;
  assign y28 = n391 ;
  assign y29 = n396 ;
  assign y30 = n401 ;
  assign y31 = n406 ;
  assign y32 = n411 ;
  assign y33 = n416 ;
  assign y34 = n421 ;
  assign y35 = n426 ;
  assign y36 = n431 ;
  assign y37 = n436 ;
  assign y38 = n441 ;
  assign y39 = n446 ;
  assign y40 = n451 ;
  assign y41 = n456 ;
  assign y42 = n461 ;
  assign y43 = n466 ;
  assign y44 = n471 ;
  assign y45 = n476 ;
  assign y46 = n481 ;
  assign y47 = n486 ;
  assign y48 = n491 ;
  assign y49 = n496 ;
  assign y50 = n501 ;
  assign y51 = n506 ;
  assign y52 = n511 ;
  assign y53 = n516 ;
  assign y54 = n521 ;
  assign y55 = n526 ;
  assign y56 = n531 ;
  assign y57 = n536 ;
  assign y58 = n541 ;
  assign y59 = n546 ;
  assign y60 = n551 ;
  assign y61 = n556 ;
  assign y62 = n561 ;
  assign y63 = n566 ;
  assign y64 = n571 ;
  assign y65 = n576 ;
  assign y66 = n581 ;
  assign y67 = n586 ;
  assign y68 = n591 ;
  assign y69 = n596 ;
  assign y70 = n601 ;
  assign y71 = n606 ;
  assign y72 = n611 ;
  assign y73 = n616 ;
  assign y74 = n621 ;
  assign y75 = n626 ;
  assign y76 = n631 ;
  assign y77 = n636 ;
  assign y78 = n641 ;
  assign y79 = n646 ;
  assign y80 = n651 ;
  assign y81 = n656 ;
  assign y82 = n661 ;
  assign y83 = n666 ;
  assign y84 = n671 ;
  assign y85 = n676 ;
  assign y86 = n681 ;
  assign y87 = n686 ;
  assign y88 = n691 ;
  assign y89 = n696 ;
  assign y90 = n701 ;
  assign y91 = n706 ;
  assign y92 = n711 ;
  assign y93 = n716 ;
  assign y94 = n721 ;
  assign y95 = n726 ;
  assign y96 = n731 ;
  assign y97 = n736 ;
  assign y98 = n741 ;
  assign y99 = n746 ;
  assign y100 = n751 ;
  assign y101 = n756 ;
  assign y102 = n761 ;
  assign y103 = n766 ;
  assign y104 = n771 ;
  assign y105 = n776 ;
  assign y106 = n781 ;
  assign y107 = n786 ;
  assign y108 = n791 ;
  assign y109 = n796 ;
  assign y110 = n801 ;
  assign y111 = n806 ;
  assign y112 = n811 ;
  assign y113 = n816 ;
  assign y114 = n821 ;
  assign y115 = n826 ;
  assign y116 = n831 ;
  assign y117 = n836 ;
  assign y118 = n841 ;
  assign y119 = n846 ;
  assign y120 = n851 ;
  assign y121 = n856 ;
  assign y122 = n861 ;
  assign y123 = n866 ;
  assign y124 = n871 ;
  assign y125 = n876 ;
  assign y126 = n881 ;
  assign y127 = n886 ;
  assign y128 = n887 ;
endmodule
