module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 ;
  assign n383 = x0 & x128 ;
  assign n397 = x0 | x128 ;
  assign n1276 = ~n383 ;
  assign n398 = n1276 & n397 ;
  assign n384 = x1 & x129 ;
  assign n399 = x1 | x129 ;
  assign n1277 = ~n384 ;
  assign n400 = n1277 & n399 ;
  assign n401 = n383 & n400 ;
  assign n402 = n383 | n400 ;
  assign n1278 = ~n401 ;
  assign n403 = n1278 & n402 ;
  assign n404 = n383 & n399 ;
  assign n405 = n384 | n404 ;
  assign n257 = x2 & x130 ;
  assign n406 = x2 | x130 ;
  assign n1279 = ~n257 ;
  assign n408 = n1279 & n406 ;
  assign n409 = n405 & n408 ;
  assign n410 = n405 | n408 ;
  assign n1280 = ~n409 ;
  assign n411 = n1280 & n410 ;
  assign n407 = n405 & n406 ;
  assign n412 = n257 | n407 ;
  assign n258 = x3 & x131 ;
  assign n413 = x3 | x131 ;
  assign n1281 = ~n258 ;
  assign n414 = n1281 & n413 ;
  assign n415 = n412 | n414 ;
  assign n416 = n412 & n414 ;
  assign n1282 = ~n416 ;
  assign n417 = n415 & n1282 ;
  assign n418 = n412 & n413 ;
  assign n419 = n258 | n418 ;
  assign n259 = x4 & x132 ;
  assign n420 = x4 | x132 ;
  assign n1283 = ~n259 ;
  assign n422 = n1283 & n420 ;
  assign n423 = n419 & n422 ;
  assign n424 = n419 | n422 ;
  assign n1284 = ~n423 ;
  assign n425 = n1284 & n424 ;
  assign n421 = n419 & n420 ;
  assign n426 = n259 | n421 ;
  assign n260 = x5 & x133 ;
  assign n427 = x5 | x133 ;
  assign n1285 = ~n260 ;
  assign n428 = n1285 & n427 ;
  assign n429 = n426 | n428 ;
  assign n430 = n426 & n428 ;
  assign n1286 = ~n430 ;
  assign n431 = n429 & n1286 ;
  assign n432 = n426 & n427 ;
  assign n433 = n260 | n432 ;
  assign n261 = x6 & x134 ;
  assign n434 = x6 | x134 ;
  assign n1287 = ~n261 ;
  assign n436 = n1287 & n434 ;
  assign n437 = n433 & n436 ;
  assign n438 = n433 | n436 ;
  assign n1288 = ~n437 ;
  assign n439 = n1288 & n438 ;
  assign n435 = n433 & n434 ;
  assign n440 = n261 | n435 ;
  assign n262 = x7 & x135 ;
  assign n441 = x7 | x135 ;
  assign n1289 = ~n262 ;
  assign n442 = n1289 & n441 ;
  assign n443 = n440 | n442 ;
  assign n444 = n440 & n442 ;
  assign n1290 = ~n444 ;
  assign n445 = n443 & n1290 ;
  assign n446 = n440 & n441 ;
  assign n447 = n262 | n446 ;
  assign n263 = x8 & x136 ;
  assign n448 = x8 | x136 ;
  assign n1291 = ~n263 ;
  assign n450 = n1291 & n448 ;
  assign n451 = n447 & n450 ;
  assign n452 = n447 | n450 ;
  assign n1292 = ~n451 ;
  assign n453 = n1292 & n452 ;
  assign n449 = n447 & n448 ;
  assign n454 = n263 | n449 ;
  assign n264 = x9 & x137 ;
  assign n455 = x9 | x137 ;
  assign n1293 = ~n264 ;
  assign n456 = n1293 & n455 ;
  assign n457 = n454 | n456 ;
  assign n458 = n454 & n456 ;
  assign n1294 = ~n458 ;
  assign n459 = n457 & n1294 ;
  assign n460 = n454 & n455 ;
  assign n461 = n264 | n460 ;
  assign n265 = x10 & x138 ;
  assign n462 = x10 | x138 ;
  assign n1295 = ~n265 ;
  assign n464 = n1295 & n462 ;
  assign n465 = n461 & n464 ;
  assign n466 = n461 | n464 ;
  assign n1296 = ~n465 ;
  assign n467 = n1296 & n466 ;
  assign n463 = n461 & n462 ;
  assign n468 = n265 | n463 ;
  assign n266 = x11 & x139 ;
  assign n469 = x11 | x139 ;
  assign n1297 = ~n266 ;
  assign n470 = n1297 & n469 ;
  assign n471 = n468 | n470 ;
  assign n472 = n468 & n470 ;
  assign n1298 = ~n472 ;
  assign n473 = n471 & n1298 ;
  assign n474 = n468 & n469 ;
  assign n475 = n266 | n474 ;
  assign n267 = x12 & x140 ;
  assign n476 = x12 | x140 ;
  assign n1299 = ~n267 ;
  assign n478 = n1299 & n476 ;
  assign n479 = n475 & n478 ;
  assign n480 = n475 | n478 ;
  assign n1300 = ~n479 ;
  assign n481 = n1300 & n480 ;
  assign n477 = n475 & n476 ;
  assign n482 = n267 | n477 ;
  assign n268 = x13 & x141 ;
  assign n483 = x13 | x141 ;
  assign n1301 = ~n268 ;
  assign n484 = n1301 & n483 ;
  assign n485 = n482 | n484 ;
  assign n486 = n482 & n484 ;
  assign n1302 = ~n486 ;
  assign n487 = n485 & n1302 ;
  assign n488 = n482 & n483 ;
  assign n489 = n268 | n488 ;
  assign n269 = x14 & x142 ;
  assign n490 = x14 | x142 ;
  assign n1303 = ~n269 ;
  assign n492 = n1303 & n490 ;
  assign n493 = n489 & n492 ;
  assign n494 = n489 | n492 ;
  assign n1304 = ~n493 ;
  assign n495 = n1304 & n494 ;
  assign n491 = n489 & n490 ;
  assign n496 = n269 | n491 ;
  assign n270 = x15 & x143 ;
  assign n497 = x15 | x143 ;
  assign n1305 = ~n270 ;
  assign n498 = n1305 & n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n496 & n498 ;
  assign n1306 = ~n500 ;
  assign n501 = n499 & n1306 ;
  assign n502 = n496 & n497 ;
  assign n503 = n270 | n502 ;
  assign n271 = x16 & x144 ;
  assign n504 = x16 | x144 ;
  assign n1307 = ~n271 ;
  assign n506 = n1307 & n504 ;
  assign n507 = n503 & n506 ;
  assign n508 = n503 | n506 ;
  assign n1308 = ~n507 ;
  assign n509 = n1308 & n508 ;
  assign n505 = n503 & n504 ;
  assign n510 = n271 | n505 ;
  assign n272 = x17 & x145 ;
  assign n511 = x17 | x145 ;
  assign n1309 = ~n272 ;
  assign n512 = n1309 & n511 ;
  assign n513 = n510 | n512 ;
  assign n514 = n510 & n512 ;
  assign n1310 = ~n514 ;
  assign n515 = n513 & n1310 ;
  assign n516 = n510 & n511 ;
  assign n517 = n272 | n516 ;
  assign n273 = x18 & x146 ;
  assign n518 = x18 | x146 ;
  assign n1311 = ~n273 ;
  assign n520 = n1311 & n518 ;
  assign n521 = n517 & n520 ;
  assign n522 = n517 | n520 ;
  assign n1312 = ~n521 ;
  assign n523 = n1312 & n522 ;
  assign n519 = n517 & n518 ;
  assign n524 = n273 | n519 ;
  assign n274 = x19 & x147 ;
  assign n525 = x19 | x147 ;
  assign n1313 = ~n274 ;
  assign n526 = n1313 & n525 ;
  assign n527 = n524 | n526 ;
  assign n528 = n524 & n526 ;
  assign n1314 = ~n528 ;
  assign n529 = n527 & n1314 ;
  assign n530 = n524 & n525 ;
  assign n531 = n274 | n530 ;
  assign n275 = x20 & x148 ;
  assign n532 = x20 | x148 ;
  assign n1315 = ~n275 ;
  assign n534 = n1315 & n532 ;
  assign n535 = n531 & n534 ;
  assign n536 = n531 | n534 ;
  assign n1316 = ~n535 ;
  assign n537 = n1316 & n536 ;
  assign n533 = n531 & n532 ;
  assign n538 = n275 | n533 ;
  assign n276 = x21 & x149 ;
  assign n539 = x21 | x149 ;
  assign n1317 = ~n276 ;
  assign n540 = n1317 & n539 ;
  assign n541 = n538 | n540 ;
  assign n542 = n538 & n540 ;
  assign n1318 = ~n542 ;
  assign n543 = n541 & n1318 ;
  assign n544 = n538 & n539 ;
  assign n545 = n276 | n544 ;
  assign n277 = x22 & x150 ;
  assign n546 = x22 | x150 ;
  assign n1319 = ~n277 ;
  assign n548 = n1319 & n546 ;
  assign n549 = n545 & n548 ;
  assign n550 = n545 | n548 ;
  assign n1320 = ~n549 ;
  assign n551 = n1320 & n550 ;
  assign n547 = n545 & n546 ;
  assign n552 = n277 | n547 ;
  assign n278 = x23 & x151 ;
  assign n553 = x23 | x151 ;
  assign n1321 = ~n278 ;
  assign n554 = n1321 & n553 ;
  assign n555 = n552 | n554 ;
  assign n556 = n552 & n554 ;
  assign n1322 = ~n556 ;
  assign n557 = n555 & n1322 ;
  assign n558 = n552 & n553 ;
  assign n559 = n278 | n558 ;
  assign n279 = x24 & x152 ;
  assign n560 = x24 | x152 ;
  assign n1323 = ~n279 ;
  assign n562 = n1323 & n560 ;
  assign n563 = n559 & n562 ;
  assign n564 = n559 | n562 ;
  assign n1324 = ~n563 ;
  assign n565 = n1324 & n564 ;
  assign n561 = n559 & n560 ;
  assign n566 = n279 | n561 ;
  assign n280 = x25 & x153 ;
  assign n567 = x25 | x153 ;
  assign n1325 = ~n280 ;
  assign n568 = n1325 & n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = n566 & n568 ;
  assign n1326 = ~n570 ;
  assign n571 = n569 & n1326 ;
  assign n572 = n566 & n567 ;
  assign n573 = n280 | n572 ;
  assign n281 = x26 & x154 ;
  assign n574 = x26 | x154 ;
  assign n1327 = ~n281 ;
  assign n576 = n1327 & n574 ;
  assign n577 = n573 & n576 ;
  assign n578 = n573 | n576 ;
  assign n1328 = ~n577 ;
  assign n579 = n1328 & n578 ;
  assign n575 = n573 & n574 ;
  assign n580 = n281 | n575 ;
  assign n282 = x27 & x155 ;
  assign n581 = x27 | x155 ;
  assign n1329 = ~n282 ;
  assign n582 = n1329 & n581 ;
  assign n583 = n580 | n582 ;
  assign n584 = n580 & n582 ;
  assign n1330 = ~n584 ;
  assign n585 = n583 & n1330 ;
  assign n586 = n580 & n581 ;
  assign n587 = n282 | n586 ;
  assign n283 = x28 & x156 ;
  assign n588 = x28 | x156 ;
  assign n1331 = ~n283 ;
  assign n590 = n1331 & n588 ;
  assign n591 = n587 & n590 ;
  assign n592 = n587 | n590 ;
  assign n1332 = ~n591 ;
  assign n593 = n1332 & n592 ;
  assign n589 = n587 & n588 ;
  assign n594 = n283 | n589 ;
  assign n284 = x29 & x157 ;
  assign n595 = x29 | x157 ;
  assign n1333 = ~n284 ;
  assign n596 = n1333 & n595 ;
  assign n597 = n594 | n596 ;
  assign n598 = n594 & n596 ;
  assign n1334 = ~n598 ;
  assign n599 = n597 & n1334 ;
  assign n600 = n594 & n595 ;
  assign n601 = n284 | n600 ;
  assign n285 = x30 & x158 ;
  assign n602 = x30 | x158 ;
  assign n1335 = ~n285 ;
  assign n604 = n1335 & n602 ;
  assign n605 = n601 & n604 ;
  assign n606 = n601 | n604 ;
  assign n1336 = ~n605 ;
  assign n607 = n1336 & n606 ;
  assign n603 = n601 & n602 ;
  assign n608 = n285 | n603 ;
  assign n286 = x31 & x159 ;
  assign n609 = x31 | x159 ;
  assign n1337 = ~n286 ;
  assign n610 = n1337 & n609 ;
  assign n611 = n608 | n610 ;
  assign n612 = n608 & n610 ;
  assign n1338 = ~n612 ;
  assign n613 = n611 & n1338 ;
  assign n614 = n608 & n609 ;
  assign n615 = n286 | n614 ;
  assign n287 = x32 & x160 ;
  assign n616 = x32 | x160 ;
  assign n1339 = ~n287 ;
  assign n618 = n1339 & n616 ;
  assign n619 = n615 & n618 ;
  assign n620 = n615 | n618 ;
  assign n1340 = ~n619 ;
  assign n621 = n1340 & n620 ;
  assign n617 = n615 & n616 ;
  assign n622 = n287 | n617 ;
  assign n288 = x33 & x161 ;
  assign n623 = x33 | x161 ;
  assign n1341 = ~n288 ;
  assign n624 = n1341 & n623 ;
  assign n625 = n622 | n624 ;
  assign n626 = n622 & n624 ;
  assign n1342 = ~n626 ;
  assign n627 = n625 & n1342 ;
  assign n628 = n622 & n623 ;
  assign n629 = n288 | n628 ;
  assign n289 = x34 & x162 ;
  assign n630 = x34 | x162 ;
  assign n1343 = ~n289 ;
  assign n632 = n1343 & n630 ;
  assign n633 = n629 & n632 ;
  assign n634 = n629 | n632 ;
  assign n1344 = ~n633 ;
  assign n635 = n1344 & n634 ;
  assign n631 = n629 & n630 ;
  assign n636 = n289 | n631 ;
  assign n290 = x35 & x163 ;
  assign n637 = x35 | x163 ;
  assign n1345 = ~n290 ;
  assign n638 = n1345 & n637 ;
  assign n639 = n636 | n638 ;
  assign n640 = n636 & n638 ;
  assign n1346 = ~n640 ;
  assign n641 = n639 & n1346 ;
  assign n642 = n636 & n637 ;
  assign n643 = n290 | n642 ;
  assign n291 = x36 & x164 ;
  assign n644 = x36 | x164 ;
  assign n1347 = ~n291 ;
  assign n646 = n1347 & n644 ;
  assign n647 = n643 & n646 ;
  assign n648 = n643 | n646 ;
  assign n1348 = ~n647 ;
  assign n649 = n1348 & n648 ;
  assign n645 = n643 & n644 ;
  assign n650 = n291 | n645 ;
  assign n292 = x37 & x165 ;
  assign n651 = x37 | x165 ;
  assign n1349 = ~n292 ;
  assign n652 = n1349 & n651 ;
  assign n653 = n650 | n652 ;
  assign n654 = n650 & n652 ;
  assign n1350 = ~n654 ;
  assign n655 = n653 & n1350 ;
  assign n656 = n650 & n651 ;
  assign n657 = n292 | n656 ;
  assign n293 = x38 & x166 ;
  assign n658 = x38 | x166 ;
  assign n1351 = ~n293 ;
  assign n660 = n1351 & n658 ;
  assign n661 = n657 & n660 ;
  assign n662 = n657 | n660 ;
  assign n1352 = ~n661 ;
  assign n663 = n1352 & n662 ;
  assign n659 = n657 & n658 ;
  assign n664 = n293 | n659 ;
  assign n294 = x39 & x167 ;
  assign n665 = x39 | x167 ;
  assign n1353 = ~n294 ;
  assign n666 = n1353 & n665 ;
  assign n667 = n664 | n666 ;
  assign n668 = n664 & n666 ;
  assign n1354 = ~n668 ;
  assign n669 = n667 & n1354 ;
  assign n670 = n664 & n665 ;
  assign n671 = n294 | n670 ;
  assign n295 = x40 & x168 ;
  assign n672 = x40 | x168 ;
  assign n1355 = ~n295 ;
  assign n674 = n1355 & n672 ;
  assign n675 = n671 & n674 ;
  assign n676 = n671 | n674 ;
  assign n1356 = ~n675 ;
  assign n677 = n1356 & n676 ;
  assign n673 = n671 & n672 ;
  assign n678 = n295 | n673 ;
  assign n296 = x41 & x169 ;
  assign n679 = x41 | x169 ;
  assign n1357 = ~n296 ;
  assign n680 = n1357 & n679 ;
  assign n681 = n678 | n680 ;
  assign n682 = n678 & n680 ;
  assign n1358 = ~n682 ;
  assign n683 = n681 & n1358 ;
  assign n684 = n678 & n679 ;
  assign n685 = n296 | n684 ;
  assign n297 = x42 & x170 ;
  assign n686 = x42 | x170 ;
  assign n1359 = ~n297 ;
  assign n688 = n1359 & n686 ;
  assign n689 = n685 & n688 ;
  assign n690 = n685 | n688 ;
  assign n1360 = ~n689 ;
  assign n691 = n1360 & n690 ;
  assign n687 = n685 & n686 ;
  assign n692 = n297 | n687 ;
  assign n298 = x43 & x171 ;
  assign n693 = x43 | x171 ;
  assign n1361 = ~n298 ;
  assign n694 = n1361 & n693 ;
  assign n695 = n692 | n694 ;
  assign n696 = n692 & n694 ;
  assign n1362 = ~n696 ;
  assign n697 = n695 & n1362 ;
  assign n698 = n692 & n693 ;
  assign n699 = n298 | n698 ;
  assign n299 = x44 & x172 ;
  assign n700 = x44 | x172 ;
  assign n1363 = ~n299 ;
  assign n702 = n1363 & n700 ;
  assign n703 = n699 & n702 ;
  assign n704 = n699 | n702 ;
  assign n1364 = ~n703 ;
  assign n705 = n1364 & n704 ;
  assign n701 = n699 & n700 ;
  assign n706 = n299 | n701 ;
  assign n300 = x45 & x173 ;
  assign n707 = x45 | x173 ;
  assign n1365 = ~n300 ;
  assign n708 = n1365 & n707 ;
  assign n709 = n706 | n708 ;
  assign n710 = n706 & n708 ;
  assign n1366 = ~n710 ;
  assign n711 = n709 & n1366 ;
  assign n712 = n706 & n707 ;
  assign n713 = n300 | n712 ;
  assign n301 = x46 & x174 ;
  assign n714 = x46 | x174 ;
  assign n1367 = ~n301 ;
  assign n716 = n1367 & n714 ;
  assign n717 = n713 & n716 ;
  assign n718 = n713 | n716 ;
  assign n1368 = ~n717 ;
  assign n719 = n1368 & n718 ;
  assign n715 = n713 & n714 ;
  assign n720 = n301 | n715 ;
  assign n302 = x47 & x175 ;
  assign n721 = x47 | x175 ;
  assign n1369 = ~n302 ;
  assign n722 = n1369 & n721 ;
  assign n723 = n720 | n722 ;
  assign n724 = n720 & n722 ;
  assign n1370 = ~n724 ;
  assign n725 = n723 & n1370 ;
  assign n726 = n720 & n721 ;
  assign n727 = n302 | n726 ;
  assign n303 = x48 & x176 ;
  assign n728 = x48 | x176 ;
  assign n1371 = ~n303 ;
  assign n730 = n1371 & n728 ;
  assign n731 = n727 & n730 ;
  assign n732 = n727 | n730 ;
  assign n1372 = ~n731 ;
  assign n733 = n1372 & n732 ;
  assign n729 = n727 & n728 ;
  assign n734 = n303 | n729 ;
  assign n304 = x49 & x177 ;
  assign n735 = x49 | x177 ;
  assign n1373 = ~n304 ;
  assign n736 = n1373 & n735 ;
  assign n737 = n734 | n736 ;
  assign n738 = n734 & n736 ;
  assign n1374 = ~n738 ;
  assign n739 = n737 & n1374 ;
  assign n740 = n734 & n735 ;
  assign n741 = n304 | n740 ;
  assign n305 = x50 & x178 ;
  assign n742 = x50 | x178 ;
  assign n1375 = ~n305 ;
  assign n744 = n1375 & n742 ;
  assign n745 = n741 & n744 ;
  assign n746 = n741 | n744 ;
  assign n1376 = ~n745 ;
  assign n747 = n1376 & n746 ;
  assign n743 = n741 & n742 ;
  assign n748 = n305 | n743 ;
  assign n306 = x51 & x179 ;
  assign n749 = x51 | x179 ;
  assign n1377 = ~n306 ;
  assign n750 = n1377 & n749 ;
  assign n751 = n748 | n750 ;
  assign n752 = n748 & n750 ;
  assign n1378 = ~n752 ;
  assign n753 = n751 & n1378 ;
  assign n754 = n748 & n749 ;
  assign n755 = n306 | n754 ;
  assign n307 = x52 & x180 ;
  assign n756 = x52 | x180 ;
  assign n1379 = ~n307 ;
  assign n758 = n1379 & n756 ;
  assign n759 = n755 & n758 ;
  assign n760 = n755 | n758 ;
  assign n1380 = ~n759 ;
  assign n761 = n1380 & n760 ;
  assign n757 = n755 & n756 ;
  assign n762 = n307 | n757 ;
  assign n308 = x53 & x181 ;
  assign n763 = x53 | x181 ;
  assign n1381 = ~n308 ;
  assign n764 = n1381 & n763 ;
  assign n765 = n762 | n764 ;
  assign n766 = n762 & n764 ;
  assign n1382 = ~n766 ;
  assign n767 = n765 & n1382 ;
  assign n768 = n762 & n763 ;
  assign n769 = n308 | n768 ;
  assign n309 = x54 & x182 ;
  assign n770 = x54 | x182 ;
  assign n1383 = ~n309 ;
  assign n772 = n1383 & n770 ;
  assign n773 = n769 & n772 ;
  assign n774 = n769 | n772 ;
  assign n1384 = ~n773 ;
  assign n775 = n1384 & n774 ;
  assign n771 = n769 & n770 ;
  assign n776 = n309 | n771 ;
  assign n310 = x55 & x183 ;
  assign n777 = x55 | x183 ;
  assign n1385 = ~n310 ;
  assign n778 = n1385 & n777 ;
  assign n779 = n776 | n778 ;
  assign n780 = n776 & n778 ;
  assign n1386 = ~n780 ;
  assign n781 = n779 & n1386 ;
  assign n782 = n776 & n777 ;
  assign n783 = n310 | n782 ;
  assign n311 = x56 & x184 ;
  assign n784 = x56 | x184 ;
  assign n1387 = ~n311 ;
  assign n786 = n1387 & n784 ;
  assign n787 = n783 & n786 ;
  assign n788 = n783 | n786 ;
  assign n1388 = ~n787 ;
  assign n789 = n1388 & n788 ;
  assign n785 = n783 & n784 ;
  assign n790 = n311 | n785 ;
  assign n312 = x57 & x185 ;
  assign n791 = x57 | x185 ;
  assign n1389 = ~n312 ;
  assign n792 = n1389 & n791 ;
  assign n793 = n790 | n792 ;
  assign n794 = n790 & n792 ;
  assign n1390 = ~n794 ;
  assign n795 = n793 & n1390 ;
  assign n796 = n790 & n791 ;
  assign n797 = n312 | n796 ;
  assign n313 = x58 & x186 ;
  assign n798 = x58 | x186 ;
  assign n1391 = ~n313 ;
  assign n800 = n1391 & n798 ;
  assign n801 = n797 & n800 ;
  assign n802 = n797 | n800 ;
  assign n1392 = ~n801 ;
  assign n803 = n1392 & n802 ;
  assign n799 = n797 & n798 ;
  assign n804 = n313 | n799 ;
  assign n314 = x59 & x187 ;
  assign n805 = x59 | x187 ;
  assign n1393 = ~n314 ;
  assign n806 = n1393 & n805 ;
  assign n807 = n804 | n806 ;
  assign n808 = n804 & n806 ;
  assign n1394 = ~n808 ;
  assign n809 = n807 & n1394 ;
  assign n810 = n804 & n805 ;
  assign n811 = n314 | n810 ;
  assign n315 = x60 & x188 ;
  assign n812 = x60 | x188 ;
  assign n1395 = ~n315 ;
  assign n814 = n1395 & n812 ;
  assign n815 = n811 & n814 ;
  assign n816 = n811 | n814 ;
  assign n1396 = ~n815 ;
  assign n817 = n1396 & n816 ;
  assign n813 = n811 & n812 ;
  assign n818 = n315 | n813 ;
  assign n316 = x61 & x189 ;
  assign n819 = x61 | x189 ;
  assign n1397 = ~n316 ;
  assign n820 = n1397 & n819 ;
  assign n821 = n818 | n820 ;
  assign n822 = n818 & n820 ;
  assign n1398 = ~n822 ;
  assign n823 = n821 & n1398 ;
  assign n824 = n818 & n819 ;
  assign n825 = n316 | n824 ;
  assign n317 = x62 & x190 ;
  assign n826 = x62 | x190 ;
  assign n1399 = ~n317 ;
  assign n828 = n1399 & n826 ;
  assign n829 = n825 & n828 ;
  assign n830 = n825 | n828 ;
  assign n1400 = ~n829 ;
  assign n831 = n1400 & n830 ;
  assign n827 = n825 & n826 ;
  assign n832 = n317 | n827 ;
  assign n318 = x63 & x191 ;
  assign n833 = x63 | x191 ;
  assign n1401 = ~n318 ;
  assign n834 = n1401 & n833 ;
  assign n835 = n832 | n834 ;
  assign n836 = n832 & n834 ;
  assign n1402 = ~n836 ;
  assign n837 = n835 & n1402 ;
  assign n838 = n832 & n833 ;
  assign n839 = n318 | n838 ;
  assign n319 = x64 & x192 ;
  assign n840 = x64 | x192 ;
  assign n1403 = ~n319 ;
  assign n842 = n1403 & n840 ;
  assign n843 = n839 & n842 ;
  assign n844 = n839 | n842 ;
  assign n1404 = ~n843 ;
  assign n845 = n1404 & n844 ;
  assign n841 = n839 & n840 ;
  assign n846 = n319 | n841 ;
  assign n320 = x65 & x193 ;
  assign n847 = x65 | x193 ;
  assign n1405 = ~n320 ;
  assign n848 = n1405 & n847 ;
  assign n849 = n846 | n848 ;
  assign n850 = n846 & n848 ;
  assign n1406 = ~n850 ;
  assign n851 = n849 & n1406 ;
  assign n852 = n846 & n847 ;
  assign n853 = n320 | n852 ;
  assign n321 = x66 & x194 ;
  assign n854 = x66 | x194 ;
  assign n1407 = ~n321 ;
  assign n856 = n1407 & n854 ;
  assign n857 = n853 & n856 ;
  assign n858 = n853 | n856 ;
  assign n1408 = ~n857 ;
  assign n859 = n1408 & n858 ;
  assign n855 = n853 & n854 ;
  assign n860 = n321 | n855 ;
  assign n322 = x67 & x195 ;
  assign n861 = x67 | x195 ;
  assign n1409 = ~n322 ;
  assign n862 = n1409 & n861 ;
  assign n863 = n860 | n862 ;
  assign n864 = n860 & n862 ;
  assign n1410 = ~n864 ;
  assign n865 = n863 & n1410 ;
  assign n866 = n860 & n861 ;
  assign n867 = n322 | n866 ;
  assign n323 = x68 & x196 ;
  assign n868 = x68 | x196 ;
  assign n1411 = ~n323 ;
  assign n870 = n1411 & n868 ;
  assign n871 = n867 & n870 ;
  assign n872 = n867 | n870 ;
  assign n1412 = ~n871 ;
  assign n873 = n1412 & n872 ;
  assign n869 = n867 & n868 ;
  assign n874 = n323 | n869 ;
  assign n324 = x69 & x197 ;
  assign n875 = x69 | x197 ;
  assign n1413 = ~n324 ;
  assign n876 = n1413 & n875 ;
  assign n877 = n874 | n876 ;
  assign n878 = n874 & n876 ;
  assign n1414 = ~n878 ;
  assign n879 = n877 & n1414 ;
  assign n880 = n874 & n875 ;
  assign n881 = n324 | n880 ;
  assign n325 = x70 & x198 ;
  assign n882 = x70 | x198 ;
  assign n1415 = ~n325 ;
  assign n884 = n1415 & n882 ;
  assign n885 = n881 & n884 ;
  assign n886 = n881 | n884 ;
  assign n1416 = ~n885 ;
  assign n887 = n1416 & n886 ;
  assign n883 = n881 & n882 ;
  assign n888 = n325 | n883 ;
  assign n326 = x71 & x199 ;
  assign n889 = x71 | x199 ;
  assign n1417 = ~n326 ;
  assign n890 = n1417 & n889 ;
  assign n891 = n888 | n890 ;
  assign n892 = n888 & n890 ;
  assign n1418 = ~n892 ;
  assign n893 = n891 & n1418 ;
  assign n894 = n888 & n889 ;
  assign n895 = n326 | n894 ;
  assign n327 = x72 & x200 ;
  assign n896 = x72 | x200 ;
  assign n1419 = ~n327 ;
  assign n898 = n1419 & n896 ;
  assign n899 = n895 & n898 ;
  assign n900 = n895 | n898 ;
  assign n1420 = ~n899 ;
  assign n901 = n1420 & n900 ;
  assign n897 = n895 & n896 ;
  assign n902 = n327 | n897 ;
  assign n328 = x73 & x201 ;
  assign n903 = x73 | x201 ;
  assign n1421 = ~n328 ;
  assign n904 = n1421 & n903 ;
  assign n905 = n902 | n904 ;
  assign n906 = n902 & n904 ;
  assign n1422 = ~n906 ;
  assign n907 = n905 & n1422 ;
  assign n908 = n902 & n903 ;
  assign n909 = n328 | n908 ;
  assign n329 = x74 & x202 ;
  assign n910 = x74 | x202 ;
  assign n1423 = ~n329 ;
  assign n912 = n1423 & n910 ;
  assign n913 = n909 & n912 ;
  assign n914 = n909 | n912 ;
  assign n1424 = ~n913 ;
  assign n915 = n1424 & n914 ;
  assign n911 = n909 & n910 ;
  assign n916 = n329 | n911 ;
  assign n330 = x75 & x203 ;
  assign n917 = x75 | x203 ;
  assign n1425 = ~n330 ;
  assign n918 = n1425 & n917 ;
  assign n919 = n916 | n918 ;
  assign n920 = n916 & n918 ;
  assign n1426 = ~n920 ;
  assign n921 = n919 & n1426 ;
  assign n922 = n916 & n917 ;
  assign n923 = n330 | n922 ;
  assign n331 = x76 & x204 ;
  assign n924 = x76 | x204 ;
  assign n1427 = ~n331 ;
  assign n926 = n1427 & n924 ;
  assign n927 = n923 & n926 ;
  assign n928 = n923 | n926 ;
  assign n1428 = ~n927 ;
  assign n929 = n1428 & n928 ;
  assign n925 = n923 & n924 ;
  assign n930 = n331 | n925 ;
  assign n332 = x77 & x205 ;
  assign n931 = x77 | x205 ;
  assign n1429 = ~n332 ;
  assign n932 = n1429 & n931 ;
  assign n933 = n930 | n932 ;
  assign n934 = n930 & n932 ;
  assign n1430 = ~n934 ;
  assign n935 = n933 & n1430 ;
  assign n936 = n930 & n931 ;
  assign n937 = n332 | n936 ;
  assign n333 = x78 & x206 ;
  assign n938 = x78 | x206 ;
  assign n1431 = ~n333 ;
  assign n940 = n1431 & n938 ;
  assign n941 = n937 & n940 ;
  assign n942 = n937 | n940 ;
  assign n1432 = ~n941 ;
  assign n943 = n1432 & n942 ;
  assign n939 = n937 & n938 ;
  assign n944 = n333 | n939 ;
  assign n334 = x79 & x207 ;
  assign n945 = x79 | x207 ;
  assign n1433 = ~n334 ;
  assign n946 = n1433 & n945 ;
  assign n947 = n944 | n946 ;
  assign n948 = n944 & n946 ;
  assign n1434 = ~n948 ;
  assign n949 = n947 & n1434 ;
  assign n950 = n944 & n945 ;
  assign n951 = n334 | n950 ;
  assign n335 = x80 & x208 ;
  assign n952 = x80 | x208 ;
  assign n1435 = ~n335 ;
  assign n954 = n1435 & n952 ;
  assign n955 = n951 & n954 ;
  assign n956 = n951 | n954 ;
  assign n1436 = ~n955 ;
  assign n957 = n1436 & n956 ;
  assign n953 = n951 & n952 ;
  assign n958 = n335 | n953 ;
  assign n336 = x81 & x209 ;
  assign n959 = x81 | x209 ;
  assign n1437 = ~n336 ;
  assign n960 = n1437 & n959 ;
  assign n961 = n958 | n960 ;
  assign n962 = n958 & n960 ;
  assign n1438 = ~n962 ;
  assign n963 = n961 & n1438 ;
  assign n964 = n958 & n959 ;
  assign n965 = n336 | n964 ;
  assign n337 = x82 & x210 ;
  assign n966 = x82 | x210 ;
  assign n1439 = ~n337 ;
  assign n968 = n1439 & n966 ;
  assign n969 = n965 & n968 ;
  assign n970 = n965 | n968 ;
  assign n1440 = ~n969 ;
  assign n971 = n1440 & n970 ;
  assign n967 = n965 & n966 ;
  assign n972 = n337 | n967 ;
  assign n338 = x83 & x211 ;
  assign n973 = x83 | x211 ;
  assign n1441 = ~n338 ;
  assign n974 = n1441 & n973 ;
  assign n975 = n972 | n974 ;
  assign n976 = n972 & n974 ;
  assign n1442 = ~n976 ;
  assign n977 = n975 & n1442 ;
  assign n978 = n972 & n973 ;
  assign n979 = n338 | n978 ;
  assign n339 = x84 & x212 ;
  assign n980 = x84 | x212 ;
  assign n1443 = ~n339 ;
  assign n982 = n1443 & n980 ;
  assign n983 = n979 & n982 ;
  assign n984 = n979 | n982 ;
  assign n1444 = ~n983 ;
  assign n985 = n1444 & n984 ;
  assign n981 = n979 & n980 ;
  assign n986 = n339 | n981 ;
  assign n340 = x85 & x213 ;
  assign n987 = x85 | x213 ;
  assign n1445 = ~n340 ;
  assign n988 = n1445 & n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = n986 & n988 ;
  assign n1446 = ~n990 ;
  assign n991 = n989 & n1446 ;
  assign n992 = n986 & n987 ;
  assign n993 = n340 | n992 ;
  assign n341 = x86 & x214 ;
  assign n994 = x86 | x214 ;
  assign n1447 = ~n341 ;
  assign n996 = n1447 & n994 ;
  assign n997 = n993 & n996 ;
  assign n998 = n993 | n996 ;
  assign n1448 = ~n997 ;
  assign n999 = n1448 & n998 ;
  assign n995 = n993 & n994 ;
  assign n1000 = n341 | n995 ;
  assign n342 = x87 & x215 ;
  assign n1001 = x87 | x215 ;
  assign n1449 = ~n342 ;
  assign n1002 = n1449 & n1001 ;
  assign n1003 = n1000 | n1002 ;
  assign n1004 = n1000 & n1002 ;
  assign n1450 = ~n1004 ;
  assign n1005 = n1003 & n1450 ;
  assign n1006 = n1000 & n1001 ;
  assign n1007 = n342 | n1006 ;
  assign n343 = x88 & x216 ;
  assign n1008 = x88 | x216 ;
  assign n1451 = ~n343 ;
  assign n1010 = n1451 & n1008 ;
  assign n1011 = n1007 & n1010 ;
  assign n1012 = n1007 | n1010 ;
  assign n1452 = ~n1011 ;
  assign n1013 = n1452 & n1012 ;
  assign n1009 = n1007 & n1008 ;
  assign n1014 = n343 | n1009 ;
  assign n344 = x89 & x217 ;
  assign n1015 = x89 | x217 ;
  assign n1453 = ~n344 ;
  assign n1016 = n1453 & n1015 ;
  assign n1017 = n1014 | n1016 ;
  assign n1018 = n1014 & n1016 ;
  assign n1454 = ~n1018 ;
  assign n1019 = n1017 & n1454 ;
  assign n1020 = n1014 & n1015 ;
  assign n1021 = n344 | n1020 ;
  assign n345 = x90 & x218 ;
  assign n1022 = x90 | x218 ;
  assign n1455 = ~n345 ;
  assign n1024 = n1455 & n1022 ;
  assign n1025 = n1021 & n1024 ;
  assign n1026 = n1021 | n1024 ;
  assign n1456 = ~n1025 ;
  assign n1027 = n1456 & n1026 ;
  assign n1023 = n1021 & n1022 ;
  assign n1028 = n345 | n1023 ;
  assign n346 = x91 & x219 ;
  assign n1029 = x91 | x219 ;
  assign n1457 = ~n346 ;
  assign n1030 = n1457 & n1029 ;
  assign n1031 = n1028 | n1030 ;
  assign n1032 = n1028 & n1030 ;
  assign n1458 = ~n1032 ;
  assign n1033 = n1031 & n1458 ;
  assign n1034 = n1028 & n1029 ;
  assign n1035 = n346 | n1034 ;
  assign n347 = x92 & x220 ;
  assign n1036 = x92 | x220 ;
  assign n1459 = ~n347 ;
  assign n1038 = n1459 & n1036 ;
  assign n1039 = n1035 & n1038 ;
  assign n1040 = n1035 | n1038 ;
  assign n1460 = ~n1039 ;
  assign n1041 = n1460 & n1040 ;
  assign n1037 = n1035 & n1036 ;
  assign n1042 = n347 | n1037 ;
  assign n348 = x93 & x221 ;
  assign n1043 = x93 | x221 ;
  assign n1461 = ~n348 ;
  assign n1044 = n1461 & n1043 ;
  assign n1045 = n1042 | n1044 ;
  assign n1046 = n1042 & n1044 ;
  assign n1462 = ~n1046 ;
  assign n1047 = n1045 & n1462 ;
  assign n1048 = n1042 & n1043 ;
  assign n1049 = n348 | n1048 ;
  assign n349 = x94 & x222 ;
  assign n1050 = x94 | x222 ;
  assign n1463 = ~n349 ;
  assign n1052 = n1463 & n1050 ;
  assign n1053 = n1049 & n1052 ;
  assign n1054 = n1049 | n1052 ;
  assign n1464 = ~n1053 ;
  assign n1055 = n1464 & n1054 ;
  assign n1051 = n1049 & n1050 ;
  assign n1056 = n349 | n1051 ;
  assign n350 = x95 & x223 ;
  assign n1057 = x95 | x223 ;
  assign n1465 = ~n350 ;
  assign n1058 = n1465 & n1057 ;
  assign n1059 = n1056 | n1058 ;
  assign n1060 = n1056 & n1058 ;
  assign n1466 = ~n1060 ;
  assign n1061 = n1059 & n1466 ;
  assign n1062 = n1056 & n1057 ;
  assign n1063 = n350 | n1062 ;
  assign n351 = x96 & x224 ;
  assign n1064 = x96 | x224 ;
  assign n1467 = ~n351 ;
  assign n1066 = n1467 & n1064 ;
  assign n1067 = n1063 & n1066 ;
  assign n1068 = n1063 | n1066 ;
  assign n1468 = ~n1067 ;
  assign n1069 = n1468 & n1068 ;
  assign n1065 = n1063 & n1064 ;
  assign n1070 = n351 | n1065 ;
  assign n352 = x97 & x225 ;
  assign n1071 = x97 | x225 ;
  assign n1469 = ~n352 ;
  assign n1072 = n1469 & n1071 ;
  assign n1073 = n1070 | n1072 ;
  assign n1074 = n1070 & n1072 ;
  assign n1470 = ~n1074 ;
  assign n1075 = n1073 & n1470 ;
  assign n1076 = n1070 & n1071 ;
  assign n1077 = n352 | n1076 ;
  assign n353 = x98 & x226 ;
  assign n1078 = x98 | x226 ;
  assign n1471 = ~n353 ;
  assign n1080 = n1471 & n1078 ;
  assign n1081 = n1077 & n1080 ;
  assign n1082 = n1077 | n1080 ;
  assign n1472 = ~n1081 ;
  assign n1083 = n1472 & n1082 ;
  assign n1079 = n1077 & n1078 ;
  assign n1084 = n353 | n1079 ;
  assign n354 = x99 & x227 ;
  assign n1085 = x99 | x227 ;
  assign n1473 = ~n354 ;
  assign n1086 = n1473 & n1085 ;
  assign n1087 = n1084 | n1086 ;
  assign n1088 = n1084 & n1086 ;
  assign n1474 = ~n1088 ;
  assign n1089 = n1087 & n1474 ;
  assign n1090 = n1084 & n1085 ;
  assign n1091 = n354 | n1090 ;
  assign n355 = x100 & x228 ;
  assign n1092 = x100 | x228 ;
  assign n1475 = ~n355 ;
  assign n1094 = n1475 & n1092 ;
  assign n1095 = n1091 & n1094 ;
  assign n1096 = n1091 | n1094 ;
  assign n1476 = ~n1095 ;
  assign n1097 = n1476 & n1096 ;
  assign n1093 = n1091 & n1092 ;
  assign n1098 = n355 | n1093 ;
  assign n356 = x101 & x229 ;
  assign n1099 = x101 | x229 ;
  assign n1477 = ~n356 ;
  assign n1100 = n1477 & n1099 ;
  assign n1101 = n1098 | n1100 ;
  assign n1102 = n1098 & n1100 ;
  assign n1478 = ~n1102 ;
  assign n1103 = n1101 & n1478 ;
  assign n1104 = n1098 & n1099 ;
  assign n1105 = n356 | n1104 ;
  assign n357 = x102 & x230 ;
  assign n1106 = x102 | x230 ;
  assign n1479 = ~n357 ;
  assign n1108 = n1479 & n1106 ;
  assign n1109 = n1105 & n1108 ;
  assign n1110 = n1105 | n1108 ;
  assign n1480 = ~n1109 ;
  assign n1111 = n1480 & n1110 ;
  assign n1107 = n1105 & n1106 ;
  assign n1112 = n357 | n1107 ;
  assign n358 = x103 & x231 ;
  assign n1113 = x103 | x231 ;
  assign n1481 = ~n358 ;
  assign n1114 = n1481 & n1113 ;
  assign n1115 = n1112 | n1114 ;
  assign n1116 = n1112 & n1114 ;
  assign n1482 = ~n1116 ;
  assign n1117 = n1115 & n1482 ;
  assign n1118 = n1112 & n1113 ;
  assign n1119 = n358 | n1118 ;
  assign n359 = x104 & x232 ;
  assign n1120 = x104 | x232 ;
  assign n1483 = ~n359 ;
  assign n1122 = n1483 & n1120 ;
  assign n1123 = n1119 & n1122 ;
  assign n1124 = n1119 | n1122 ;
  assign n1484 = ~n1123 ;
  assign n1125 = n1484 & n1124 ;
  assign n1121 = n1119 & n1120 ;
  assign n1126 = n359 | n1121 ;
  assign n360 = x105 & x233 ;
  assign n1127 = x105 | x233 ;
  assign n1485 = ~n360 ;
  assign n1128 = n1485 & n1127 ;
  assign n1129 = n1126 | n1128 ;
  assign n1130 = n1126 & n1128 ;
  assign n1486 = ~n1130 ;
  assign n1131 = n1129 & n1486 ;
  assign n1132 = n1126 & n1127 ;
  assign n1133 = n360 | n1132 ;
  assign n361 = x106 & x234 ;
  assign n1134 = x106 | x234 ;
  assign n1487 = ~n361 ;
  assign n1136 = n1487 & n1134 ;
  assign n1137 = n1133 & n1136 ;
  assign n1138 = n1133 | n1136 ;
  assign n1488 = ~n1137 ;
  assign n1139 = n1488 & n1138 ;
  assign n1135 = n1133 & n1134 ;
  assign n1140 = n361 | n1135 ;
  assign n362 = x107 & x235 ;
  assign n1141 = x107 | x235 ;
  assign n1489 = ~n362 ;
  assign n1142 = n1489 & n1141 ;
  assign n1143 = n1140 | n1142 ;
  assign n1144 = n1140 & n1142 ;
  assign n1490 = ~n1144 ;
  assign n1145 = n1143 & n1490 ;
  assign n1146 = n1140 & n1141 ;
  assign n1147 = n362 | n1146 ;
  assign n363 = x108 & x236 ;
  assign n1148 = x108 | x236 ;
  assign n1491 = ~n363 ;
  assign n1150 = n1491 & n1148 ;
  assign n1151 = n1147 & n1150 ;
  assign n1152 = n1147 | n1150 ;
  assign n1492 = ~n1151 ;
  assign n1153 = n1492 & n1152 ;
  assign n1149 = n1147 & n1148 ;
  assign n1154 = n363 | n1149 ;
  assign n364 = x109 & x237 ;
  assign n1155 = x109 | x237 ;
  assign n1493 = ~n364 ;
  assign n1156 = n1493 & n1155 ;
  assign n1157 = n1154 | n1156 ;
  assign n1158 = n1154 & n1156 ;
  assign n1494 = ~n1158 ;
  assign n1159 = n1157 & n1494 ;
  assign n1160 = n1154 & n1155 ;
  assign n1161 = n364 | n1160 ;
  assign n365 = x110 & x238 ;
  assign n1162 = x110 | x238 ;
  assign n1495 = ~n365 ;
  assign n1164 = n1495 & n1162 ;
  assign n1165 = n1161 & n1164 ;
  assign n1166 = n1161 | n1164 ;
  assign n1496 = ~n1165 ;
  assign n1167 = n1496 & n1166 ;
  assign n1163 = n1161 & n1162 ;
  assign n1168 = n365 | n1163 ;
  assign n366 = x111 & x239 ;
  assign n1169 = x111 | x239 ;
  assign n1497 = ~n366 ;
  assign n1170 = n1497 & n1169 ;
  assign n1171 = n1168 | n1170 ;
  assign n1172 = n1168 & n1170 ;
  assign n1498 = ~n1172 ;
  assign n1173 = n1171 & n1498 ;
  assign n1174 = n1168 & n1169 ;
  assign n1175 = n366 | n1174 ;
  assign n367 = x112 & x240 ;
  assign n1176 = x112 | x240 ;
  assign n1499 = ~n367 ;
  assign n1178 = n1499 & n1176 ;
  assign n1179 = n1175 & n1178 ;
  assign n1180 = n1175 | n1178 ;
  assign n1500 = ~n1179 ;
  assign n1181 = n1500 & n1180 ;
  assign n1177 = n1175 & n1176 ;
  assign n1182 = n367 | n1177 ;
  assign n368 = x113 & x241 ;
  assign n1183 = x113 | x241 ;
  assign n1501 = ~n368 ;
  assign n1184 = n1501 & n1183 ;
  assign n1185 = n1182 | n1184 ;
  assign n1186 = n1182 & n1184 ;
  assign n1502 = ~n1186 ;
  assign n1187 = n1185 & n1502 ;
  assign n1188 = n1182 & n1183 ;
  assign n1189 = n368 | n1188 ;
  assign n369 = x114 & x242 ;
  assign n1190 = x114 | x242 ;
  assign n1503 = ~n369 ;
  assign n1192 = n1503 & n1190 ;
  assign n1193 = n1189 & n1192 ;
  assign n1194 = n1189 | n1192 ;
  assign n1504 = ~n1193 ;
  assign n1195 = n1504 & n1194 ;
  assign n1191 = n1189 & n1190 ;
  assign n1196 = n369 | n1191 ;
  assign n370 = x115 & x243 ;
  assign n1197 = x115 | x243 ;
  assign n1505 = ~n370 ;
  assign n1198 = n1505 & n1197 ;
  assign n1199 = n1196 | n1198 ;
  assign n1200 = n1196 & n1198 ;
  assign n1506 = ~n1200 ;
  assign n1201 = n1199 & n1506 ;
  assign n1202 = n1196 & n1197 ;
  assign n1203 = n370 | n1202 ;
  assign n371 = x116 & x244 ;
  assign n1204 = x116 | x244 ;
  assign n1507 = ~n371 ;
  assign n1206 = n1507 & n1204 ;
  assign n1207 = n1203 & n1206 ;
  assign n1208 = n1203 | n1206 ;
  assign n1508 = ~n1207 ;
  assign n1209 = n1508 & n1208 ;
  assign n1205 = n1203 & n1204 ;
  assign n1210 = n371 | n1205 ;
  assign n372 = x117 & x245 ;
  assign n1211 = x117 | x245 ;
  assign n1509 = ~n372 ;
  assign n1212 = n1509 & n1211 ;
  assign n1213 = n1210 | n1212 ;
  assign n1214 = n1210 & n1212 ;
  assign n1510 = ~n1214 ;
  assign n1215 = n1213 & n1510 ;
  assign n1216 = n1210 & n1211 ;
  assign n1217 = n372 | n1216 ;
  assign n373 = x118 & x246 ;
  assign n1218 = x118 | x246 ;
  assign n1511 = ~n373 ;
  assign n1220 = n1511 & n1218 ;
  assign n1221 = n1217 & n1220 ;
  assign n1222 = n1217 | n1220 ;
  assign n1512 = ~n1221 ;
  assign n1223 = n1512 & n1222 ;
  assign n1219 = n1217 & n1218 ;
  assign n1224 = n373 | n1219 ;
  assign n374 = x119 & x247 ;
  assign n1225 = x119 | x247 ;
  assign n1513 = ~n374 ;
  assign n1226 = n1513 & n1225 ;
  assign n1227 = n1224 | n1226 ;
  assign n1228 = n1224 & n1226 ;
  assign n1514 = ~n1228 ;
  assign n1229 = n1227 & n1514 ;
  assign n1230 = n1224 & n1225 ;
  assign n1231 = n374 | n1230 ;
  assign n375 = x120 & x248 ;
  assign n1232 = x120 | x248 ;
  assign n1515 = ~n375 ;
  assign n1234 = n1515 & n1232 ;
  assign n1235 = n1231 & n1234 ;
  assign n1236 = n1231 | n1234 ;
  assign n1516 = ~n1235 ;
  assign n1237 = n1516 & n1236 ;
  assign n1233 = n1231 & n1232 ;
  assign n1238 = n375 | n1233 ;
  assign n376 = x121 & x249 ;
  assign n1239 = x121 | x249 ;
  assign n1517 = ~n376 ;
  assign n1240 = n1517 & n1239 ;
  assign n1241 = n1238 | n1240 ;
  assign n1242 = n1238 & n1240 ;
  assign n1518 = ~n1242 ;
  assign n1243 = n1241 & n1518 ;
  assign n377 = x122 & x250 ;
  assign n385 = x122 | x250 ;
  assign n1519 = ~n377 ;
  assign n386 = n1519 & n385 ;
  assign n1244 = n1238 & n1239 ;
  assign n1245 = n376 | n1244 ;
  assign n1246 = n386 & n1245 ;
  assign n1274 = n386 | n1245 ;
  assign n1520 = ~n1246 ;
  assign n1275 = n1520 & n1274 ;
  assign n378 = x123 & x251 ;
  assign n387 = x123 | x251 ;
  assign n1521 = ~n378 ;
  assign n388 = n1521 & n387 ;
  assign n1247 = n385 & n1245 ;
  assign n1248 = n377 | n1247 ;
  assign n1249 = n388 | n1248 ;
  assign n1250 = n388 & n1248 ;
  assign n1522 = ~n1250 ;
  assign n1251 = n1249 & n1522 ;
  assign n379 = x124 & x252 ;
  assign n389 = x124 | x252 ;
  assign n1523 = ~n379 ;
  assign n390 = n1523 & n389 ;
  assign n1252 = n387 & n1248 ;
  assign n1253 = n378 | n1252 ;
  assign n1254 = n390 & n1253 ;
  assign n1272 = n390 | n1253 ;
  assign n1524 = ~n1254 ;
  assign n1273 = n1524 & n1272 ;
  assign n380 = x125 & x253 ;
  assign n391 = x125 | x253 ;
  assign n1525 = ~n380 ;
  assign n392 = n1525 & n391 ;
  assign n1255 = n389 & n1253 ;
  assign n1256 = n379 | n1255 ;
  assign n1257 = n392 | n1256 ;
  assign n1258 = n392 & n1256 ;
  assign n1526 = ~n1258 ;
  assign n1259 = n1257 & n1526 ;
  assign n381 = x126 & x254 ;
  assign n393 = x126 | x254 ;
  assign n1527 = ~n381 ;
  assign n394 = n1527 & n393 ;
  assign n1260 = n391 & n1256 ;
  assign n1261 = n380 | n1260 ;
  assign n1262 = n394 & n1261 ;
  assign n1263 = n394 | n1261 ;
  assign n1528 = ~n1262 ;
  assign n1264 = n1528 & n1263 ;
  assign n382 = x127 & x255 ;
  assign n395 = x127 | x255 ;
  assign n1529 = ~n382 ;
  assign n396 = n1529 & n395 ;
  assign n1265 = n393 & n1261 ;
  assign n1266 = n381 | n1265 ;
  assign n1267 = n396 | n1266 ;
  assign n1268 = n396 & n1266 ;
  assign n1530 = ~n1268 ;
  assign n1269 = n1267 & n1530 ;
  assign n1270 = n395 & n1266 ;
  assign n1271 = n382 | n1270 ;
  assign y0 = n398 ;
  assign y1 = n403 ;
  assign y2 = n411 ;
  assign y3 = n417 ;
  assign y4 = n425 ;
  assign y5 = n431 ;
  assign y6 = n439 ;
  assign y7 = n445 ;
  assign y8 = n453 ;
  assign y9 = n459 ;
  assign y10 = n467 ;
  assign y11 = n473 ;
  assign y12 = n481 ;
  assign y13 = n487 ;
  assign y14 = n495 ;
  assign y15 = n501 ;
  assign y16 = n509 ;
  assign y17 = n515 ;
  assign y18 = n523 ;
  assign y19 = n529 ;
  assign y20 = n537 ;
  assign y21 = n543 ;
  assign y22 = n551 ;
  assign y23 = n557 ;
  assign y24 = n565 ;
  assign y25 = n571 ;
  assign y26 = n579 ;
  assign y27 = n585 ;
  assign y28 = n593 ;
  assign y29 = n599 ;
  assign y30 = n607 ;
  assign y31 = n613 ;
  assign y32 = n621 ;
  assign y33 = n627 ;
  assign y34 = n635 ;
  assign y35 = n641 ;
  assign y36 = n649 ;
  assign y37 = n655 ;
  assign y38 = n663 ;
  assign y39 = n669 ;
  assign y40 = n677 ;
  assign y41 = n683 ;
  assign y42 = n691 ;
  assign y43 = n697 ;
  assign y44 = n705 ;
  assign y45 = n711 ;
  assign y46 = n719 ;
  assign y47 = n725 ;
  assign y48 = n733 ;
  assign y49 = n739 ;
  assign y50 = n747 ;
  assign y51 = n753 ;
  assign y52 = n761 ;
  assign y53 = n767 ;
  assign y54 = n775 ;
  assign y55 = n781 ;
  assign y56 = n789 ;
  assign y57 = n795 ;
  assign y58 = n803 ;
  assign y59 = n809 ;
  assign y60 = n817 ;
  assign y61 = n823 ;
  assign y62 = n831 ;
  assign y63 = n837 ;
  assign y64 = n845 ;
  assign y65 = n851 ;
  assign y66 = n859 ;
  assign y67 = n865 ;
  assign y68 = n873 ;
  assign y69 = n879 ;
  assign y70 = n887 ;
  assign y71 = n893 ;
  assign y72 = n901 ;
  assign y73 = n907 ;
  assign y74 = n915 ;
  assign y75 = n921 ;
  assign y76 = n929 ;
  assign y77 = n935 ;
  assign y78 = n943 ;
  assign y79 = n949 ;
  assign y80 = n957 ;
  assign y81 = n963 ;
  assign y82 = n971 ;
  assign y83 = n977 ;
  assign y84 = n985 ;
  assign y85 = n991 ;
  assign y86 = n999 ;
  assign y87 = n1005 ;
  assign y88 = n1013 ;
  assign y89 = n1019 ;
  assign y90 = n1027 ;
  assign y91 = n1033 ;
  assign y92 = n1041 ;
  assign y93 = n1047 ;
  assign y94 = n1055 ;
  assign y95 = n1061 ;
  assign y96 = n1069 ;
  assign y97 = n1075 ;
  assign y98 = n1083 ;
  assign y99 = n1089 ;
  assign y100 = n1097 ;
  assign y101 = n1103 ;
  assign y102 = n1111 ;
  assign y103 = n1117 ;
  assign y104 = n1125 ;
  assign y105 = n1131 ;
  assign y106 = n1139 ;
  assign y107 = n1145 ;
  assign y108 = n1153 ;
  assign y109 = n1159 ;
  assign y110 = n1167 ;
  assign y111 = n1173 ;
  assign y112 = n1181 ;
  assign y113 = n1187 ;
  assign y114 = n1195 ;
  assign y115 = n1201 ;
  assign y116 = n1209 ;
  assign y117 = n1215 ;
  assign y118 = n1223 ;
  assign y119 = n1229 ;
  assign y120 = n1237 ;
  assign y121 = n1243 ;
  assign y122 = n1275 ;
  assign y123 = n1251 ;
  assign y124 = n1273 ;
  assign y125 = n1259 ;
  assign y126 = n1264 ;
  assign y127 = n1269 ;
  assign y128 = n1271 ;
endmodule
