module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 ;
  assign n513 = ~x119 & x247 ;
  assign n514 = ~x118 & x246 ;
  assign n515 = n513 | n514 ;
  assign n516 = ~x112 & x240 ;
  assign n517 = ~x114 & x242 ;
  assign n518 = ~x115 & x243 ;
  assign n519 = n517 | n518 ;
  assign n520 = ~x111 & x239 ;
  assign n521 = x238 | n520 ;
  assign n522 = x110 & ~n521 ;
  assign n523 = ~x110 & x238 ;
  assign n524 = x108 & ~x236 ;
  assign n525 = ( x109 & ~x237 ) | ( x109 & n524 ) | ( ~x237 & n524 ) ;
  assign n526 = ( n520 & ~n523 ) | ( n520 & n525 ) | ( ~n523 & n525 ) ;
  assign n527 = ~n520 & n526 ;
  assign n528 = n520 | n523 ;
  assign n529 = ~x103 & x231 ;
  assign n530 = x230 | n529 ;
  assign n531 = x102 & ~n530 ;
  assign n532 = ~x102 & x230 ;
  assign n533 = x100 & ~x228 ;
  assign n534 = ( x101 & ~x229 ) | ( x101 & n533 ) | ( ~x229 & n533 ) ;
  assign n535 = ( n529 & ~n532 ) | ( n529 & n534 ) | ( ~n532 & n534 ) ;
  assign n536 = ~n529 & n535 ;
  assign n537 = n529 | n532 ;
  assign n538 = ~x96 & x224 ;
  assign n539 = ~x98 & x226 ;
  assign n540 = ~x99 & x227 ;
  assign n541 = n539 | n540 ;
  assign n542 = ~x97 & x225 ;
  assign n543 = x95 & ~x223 ;
  assign n544 = ~x95 & x223 ;
  assign n545 = x222 | n544 ;
  assign n546 = x94 & ~n545 ;
  assign n547 = ~x94 & x222 ;
  assign n548 = x92 & ~x220 ;
  assign n549 = ( x93 & ~x221 ) | ( x93 & n548 ) | ( ~x221 & n548 ) ;
  assign n550 = ( n544 & ~n547 ) | ( n544 & n549 ) | ( ~n547 & n549 ) ;
  assign n551 = ~n544 & n550 ;
  assign n552 = n544 | n547 ;
  assign n553 = ~x87 & x215 ;
  assign n554 = x214 | n553 ;
  assign n555 = x86 & ~n554 ;
  assign n556 = ~x86 & x214 ;
  assign n557 = x84 & ~x212 ;
  assign n558 = ( x85 & ~x213 ) | ( x85 & n557 ) | ( ~x213 & n557 ) ;
  assign n559 = ( n553 & ~n556 ) | ( n553 & n558 ) | ( ~n556 & n558 ) ;
  assign n560 = ~n553 & n559 ;
  assign n561 = n553 | n556 ;
  assign n562 = ~x80 & x208 ;
  assign n563 = ~x82 & x210 ;
  assign n564 = ~x83 & x211 ;
  assign n565 = n563 | n564 ;
  assign n566 = ~x81 & x209 ;
  assign n567 = x79 & ~x207 ;
  assign n568 = ~x79 & x207 ;
  assign n569 = x206 | n568 ;
  assign n570 = x78 & ~n569 ;
  assign n571 = ~x78 & x206 ;
  assign n572 = x76 & ~x204 ;
  assign n573 = ( x77 & ~x205 ) | ( x77 & n572 ) | ( ~x205 & n572 ) ;
  assign n574 = ( n568 & ~n571 ) | ( n568 & n573 ) | ( ~n571 & n573 ) ;
  assign n575 = ~n568 & n574 ;
  assign n576 = n568 | n571 ;
  assign n577 = ~x71 & x199 ;
  assign n578 = x198 | n577 ;
  assign n579 = x70 & ~n578 ;
  assign n580 = ~x70 & x198 ;
  assign n581 = x68 & ~x196 ;
  assign n582 = ( x69 & ~x197 ) | ( x69 & n581 ) | ( ~x197 & n581 ) ;
  assign n583 = ( n577 & ~n580 ) | ( n577 & n582 ) | ( ~n580 & n582 ) ;
  assign n584 = ~n577 & n583 ;
  assign n585 = n577 | n580 ;
  assign n586 = ~x66 & x194 ;
  assign n587 = ~x67 & x195 ;
  assign n588 = ~x65 & x193 ;
  assign n589 = ~x64 & x192 ;
  assign n590 = ~x63 & x191 ;
  assign n591 = ~x62 & x190 ;
  assign n592 = n590 | n591 ;
  assign n593 = ~x60 & x188 ;
  assign n594 = ~x61 & x189 ;
  assign n595 = n593 | n594 ;
  assign n596 = n592 | n595 ;
  assign n597 = x59 & ~x187 ;
  assign n598 = ~x59 & x187 ;
  assign n599 = ~x58 & x186 ;
  assign n600 = x56 & ~x184 ;
  assign n601 = ( x57 & ~x185 ) | ( x57 & n600 ) | ( ~x185 & n600 ) ;
  assign n602 = x186 & ~n601 ;
  assign n603 = ( x58 & n601 ) | ( x58 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = ( n598 & ~n599 ) | ( n598 & n603 ) | ( ~n599 & n603 ) ;
  assign n605 = ~n598 & n604 ;
  assign n606 = ( ~n596 & n597 ) | ( ~n596 & n605 ) | ( n597 & n605 ) ;
  assign n607 = ~n596 & n606 ;
  assign n608 = n598 | n599 ;
  assign n609 = ~x47 & x175 ;
  assign n610 = ~x46 & x174 ;
  assign n611 = n609 | n610 ;
  assign n612 = ~x44 & x172 ;
  assign n613 = ~x45 & x173 ;
  assign n614 = n612 | n613 ;
  assign n615 = n611 | n614 ;
  assign n616 = ~x42 & x170 ;
  assign n617 = ~x43 & x171 ;
  assign n618 = x40 & ~x168 ;
  assign n619 = ( x41 & ~x169 ) | ( x41 & n618 ) | ( ~x169 & n618 ) ;
  assign n620 = x170 & ~n619 ;
  assign n621 = ( x42 & n619 ) | ( x42 & ~n620 ) | ( n619 & ~n620 ) ;
  assign n622 = ( n616 & ~n617 ) | ( n616 & n621 ) | ( ~n617 & n621 ) ;
  assign n623 = ~n616 & n622 ;
  assign n624 = x43 & ~x171 ;
  assign n625 = ( ~n615 & n623 ) | ( ~n615 & n624 ) | ( n623 & n624 ) ;
  assign n626 = ~n615 & n625 ;
  assign n627 = x44 & ~x172 ;
  assign n628 = ( x45 & ~x173 ) | ( x45 & n627 ) | ( ~x173 & n627 ) ;
  assign n629 = ( n609 & ~n610 ) | ( n609 & n628 ) | ( ~n610 & n628 ) ;
  assign n630 = ~n609 & n629 ;
  assign n631 = ~x32 & x160 ;
  assign n632 = ~x2 & x130 ;
  assign n633 = x0 & ~x128 ;
  assign n634 = x1 & ~x129 ;
  assign n635 = n633 | n634 ;
  assign n636 = ~x1 & x129 ;
  assign n637 = ( n632 & n635 ) | ( n632 & ~n636 ) | ( n635 & ~n636 ) ;
  assign n638 = ~n632 & n637 ;
  assign n639 = x130 & ~n638 ;
  assign n640 = ( x2 & n638 ) | ( x2 & ~n639 ) | ( n638 & ~n639 ) ;
  assign n641 = ( x3 & ~x131 ) | ( x3 & n640 ) | ( ~x131 & n640 ) ;
  assign n642 = ( x4 & ~x132 ) | ( x4 & n641 ) | ( ~x132 & n641 ) ;
  assign n643 = ( x5 & ~x133 ) | ( x5 & n642 ) | ( ~x133 & n642 ) ;
  assign n644 = ( x6 & ~x134 ) | ( x6 & n643 ) | ( ~x134 & n643 ) ;
  assign n645 = ( x7 & ~x135 ) | ( x7 & n644 ) | ( ~x135 & n644 ) ;
  assign n646 = ( x8 & ~x136 ) | ( x8 & n645 ) | ( ~x136 & n645 ) ;
  assign n647 = ( x9 & ~x137 ) | ( x9 & n646 ) | ( ~x137 & n646 ) ;
  assign n648 = ( x10 & ~x138 ) | ( x10 & n647 ) | ( ~x138 & n647 ) ;
  assign n649 = ( x11 & ~x139 ) | ( x11 & n648 ) | ( ~x139 & n648 ) ;
  assign n650 = ( x12 & ~x140 ) | ( x12 & n649 ) | ( ~x140 & n649 ) ;
  assign n651 = ( x13 & ~x141 ) | ( x13 & n650 ) | ( ~x141 & n650 ) ;
  assign n652 = ( x14 & ~x142 ) | ( x14 & n651 ) | ( ~x142 & n651 ) ;
  assign n653 = ( x15 & ~x143 ) | ( x15 & n652 ) | ( ~x143 & n652 ) ;
  assign n654 = ( x16 & ~x144 ) | ( x16 & n653 ) | ( ~x144 & n653 ) ;
  assign n655 = ( x17 & ~x145 ) | ( x17 & n654 ) | ( ~x145 & n654 ) ;
  assign n656 = ( x18 & ~x146 ) | ( x18 & n655 ) | ( ~x146 & n655 ) ;
  assign n657 = ( x19 & ~x147 ) | ( x19 & n656 ) | ( ~x147 & n656 ) ;
  assign n658 = ( x20 & ~x148 ) | ( x20 & n657 ) | ( ~x148 & n657 ) ;
  assign n659 = ( x21 & ~x149 ) | ( x21 & n658 ) | ( ~x149 & n658 ) ;
  assign n660 = ( x22 & ~x150 ) | ( x22 & n659 ) | ( ~x150 & n659 ) ;
  assign n661 = ( x23 & ~x151 ) | ( x23 & n660 ) | ( ~x151 & n660 ) ;
  assign n662 = ( x24 & ~x152 ) | ( x24 & n661 ) | ( ~x152 & n661 ) ;
  assign n663 = ( x25 & ~x153 ) | ( x25 & n662 ) | ( ~x153 & n662 ) ;
  assign n664 = ( x26 & ~x154 ) | ( x26 & n663 ) | ( ~x154 & n663 ) ;
  assign n665 = ( x27 & ~x155 ) | ( x27 & n664 ) | ( ~x155 & n664 ) ;
  assign n666 = ( x28 & ~x156 ) | ( x28 & n665 ) | ( ~x156 & n665 ) ;
  assign n667 = ( x29 & ~x157 ) | ( x29 & n666 ) | ( ~x157 & n666 ) ;
  assign n668 = ( x30 & ~x158 ) | ( x30 & n667 ) | ( ~x158 & n667 ) ;
  assign n669 = ( x31 & ~x159 ) | ( x31 & n668 ) | ( ~x159 & n668 ) ;
  assign n670 = ~x39 & x167 ;
  assign n671 = ~x38 & x166 ;
  assign n672 = n670 | n671 ;
  assign n673 = ~x36 & x164 ;
  assign n674 = ~x37 & x165 ;
  assign n675 = n673 | n674 ;
  assign n676 = n672 | n675 ;
  assign n677 = ~x33 & x161 ;
  assign n678 = ~x35 & x163 ;
  assign n679 = ~x34 & x162 ;
  assign n680 = n678 | n679 ;
  assign n681 = n677 | n680 ;
  assign n682 = n676 | n681 ;
  assign n683 = ( n631 & n669 ) | ( n631 & ~n682 ) | ( n669 & ~n682 ) ;
  assign n684 = ~n631 & n683 ;
  assign n685 = x39 & ~x167 ;
  assign n686 = x166 | n670 ;
  assign n687 = x38 & ~n686 ;
  assign n688 = x36 & ~x164 ;
  assign n689 = ( x37 & ~x165 ) | ( x37 & n688 ) | ( ~x165 & n688 ) ;
  assign n690 = ( n670 & ~n671 ) | ( n670 & n689 ) | ( ~n671 & n689 ) ;
  assign n691 = ~n670 & n690 ;
  assign n692 = x35 & ~x163 ;
  assign n693 = x33 & ~x161 ;
  assign n694 = x160 | n677 ;
  assign n695 = ~n693 & n694 ;
  assign n696 = ( x32 & n693 ) | ( x32 & ~n695 ) | ( n693 & ~n695 ) ;
  assign n697 = x34 & ~x162 ;
  assign n698 = ( ~n680 & n696 ) | ( ~n680 & n697 ) | ( n696 & n697 ) ;
  assign n699 = ~n680 & n698 ;
  assign n700 = ( ~n676 & n692 ) | ( ~n676 & n699 ) | ( n692 & n699 ) ;
  assign n701 = ~n676 & n700 ;
  assign n702 = ( ~n687 & n691 ) | ( ~n687 & n701 ) | ( n691 & n701 ) ;
  assign n703 = n687 | n702 ;
  assign n704 = ( ~n684 & n685 ) | ( ~n684 & n703 ) | ( n685 & n703 ) ;
  assign n705 = n684 | n704 ;
  assign n706 = n616 | n617 ;
  assign n707 = ~x41 & x169 ;
  assign n708 = ~x40 & x168 ;
  assign n709 = n707 | n708 ;
  assign n710 = n706 | n709 ;
  assign n711 = ( n615 & n705 ) | ( n615 & ~n710 ) | ( n705 & ~n710 ) ;
  assign n712 = ~n615 & n711 ;
  assign n713 = x174 | n609 ;
  assign n714 = ~n712 & n713 ;
  assign n715 = ( x46 & n712 ) | ( x46 & ~n714 ) | ( n712 & ~n714 ) ;
  assign n716 = ( ~n626 & n630 ) | ( ~n626 & n715 ) | ( n630 & n715 ) ;
  assign n717 = n626 | n716 ;
  assign n718 = x175 & ~n717 ;
  assign n719 = ( x47 & n717 ) | ( x47 & ~n718 ) | ( n717 & ~n718 ) ;
  assign n720 = ~x54 & x182 ;
  assign n721 = ~x55 & x183 ;
  assign n722 = n720 | n721 ;
  assign n723 = x52 & ~x180 ;
  assign n724 = ( x53 & ~x181 ) | ( x53 & n723 ) | ( ~x181 & n723 ) ;
  assign n725 = x54 & ~x182 ;
  assign n726 = ( ~n722 & n724 ) | ( ~n722 & n725 ) | ( n724 & n725 ) ;
  assign n727 = ~n722 & n726 ;
  assign n728 = ~x53 & x181 ;
  assign n729 = ~x52 & x180 ;
  assign n730 = n728 | n729 ;
  assign n731 = n722 | n730 ;
  assign n732 = ~x51 & x179 ;
  assign n733 = ~x50 & x178 ;
  assign n734 = n732 | n733 ;
  assign n735 = x49 & ~x177 ;
  assign n736 = ~x49 & x177 ;
  assign n737 = x176 | n736 ;
  assign n738 = ~n735 & n737 ;
  assign n739 = ( x48 & n735 ) | ( x48 & ~n738 ) | ( n735 & ~n738 ) ;
  assign n740 = x50 & ~x178 ;
  assign n741 = ( ~n734 & n739 ) | ( ~n734 & n740 ) | ( n739 & n740 ) ;
  assign n742 = ~n734 & n741 ;
  assign n743 = x179 & ~n742 ;
  assign n744 = ( x51 & n742 ) | ( x51 & ~n743 ) | ( n742 & ~n743 ) ;
  assign n745 = ( n727 & ~n731 ) | ( n727 & n744 ) | ( ~n731 & n744 ) ;
  assign n746 = n731 ^ n727 ^ 1'b0 ;
  assign n747 = ( n727 & n745 ) | ( n727 & ~n746 ) | ( n745 & ~n746 ) ;
  assign n748 = x183 & ~n747 ;
  assign n749 = ( x55 & n747 ) | ( x55 & ~n748 ) | ( n747 & ~n748 ) ;
  assign n750 = ~x48 & x176 ;
  assign n751 = n734 | n736 ;
  assign n752 = ( n731 & ~n750 ) | ( n731 & n751 ) | ( ~n750 & n751 ) ;
  assign n753 = n750 | n752 ;
  assign n754 = ~n749 & n753 ;
  assign n755 = ( n719 & n749 ) | ( n719 & ~n754 ) | ( n749 & ~n754 ) ;
  assign n756 = ~x57 & x185 ;
  assign n757 = ~x56 & x184 ;
  assign n758 = n756 | n757 ;
  assign n759 = n596 | n758 ;
  assign n760 = ( n608 & n755 ) | ( n608 & ~n759 ) | ( n755 & ~n759 ) ;
  assign n761 = ~n608 & n760 ;
  assign n762 = x190 | n590 ;
  assign n763 = ~n761 & n762 ;
  assign n764 = ( x62 & n761 ) | ( x62 & ~n763 ) | ( n761 & ~n763 ) ;
  assign n765 = x60 & ~x188 ;
  assign n766 = ( x61 & ~x189 ) | ( x61 & n765 ) | ( ~x189 & n765 ) ;
  assign n767 = ( n590 & ~n591 ) | ( n590 & n766 ) | ( ~n591 & n766 ) ;
  assign n768 = ~n590 & n767 ;
  assign n769 = ( ~n607 & n764 ) | ( ~n607 & n768 ) | ( n764 & n768 ) ;
  assign n770 = n607 | n769 ;
  assign n771 = x191 & ~n770 ;
  assign n772 = ( x63 & n770 ) | ( x63 & ~n771 ) | ( n770 & ~n771 ) ;
  assign n773 = ( n588 & ~n589 ) | ( n588 & n772 ) | ( ~n589 & n772 ) ;
  assign n774 = ~n588 & n773 ;
  assign n775 = ( n586 & ~n587 ) | ( n586 & n774 ) | ( ~n587 & n774 ) ;
  assign n776 = ~n586 & n775 ;
  assign n777 = x64 & ~x192 ;
  assign n778 = ( x65 & ~x193 ) | ( x65 & n777 ) | ( ~x193 & n777 ) ;
  assign n779 = x194 & ~n778 ;
  assign n780 = ( x66 & n778 ) | ( x66 & ~n779 ) | ( n778 & ~n779 ) ;
  assign n781 = ( n586 & ~n587 ) | ( n586 & n780 ) | ( ~n587 & n780 ) ;
  assign n782 = ~n586 & n781 ;
  assign n783 = x67 & ~x195 ;
  assign n784 = ( ~n776 & n782 ) | ( ~n776 & n783 ) | ( n782 & n783 ) ;
  assign n785 = n776 | n784 ;
  assign n786 = ~x69 & x197 ;
  assign n787 = ~x68 & x196 ;
  assign n788 = n786 | n787 ;
  assign n789 = ( n585 & n785 ) | ( n585 & ~n788 ) | ( n785 & ~n788 ) ;
  assign n790 = ~n585 & n789 ;
  assign n791 = ( ~n579 & n584 ) | ( ~n579 & n790 ) | ( n584 & n790 ) ;
  assign n792 = n579 | n791 ;
  assign n793 = x199 & ~n792 ;
  assign n794 = ( x71 & n792 ) | ( x71 & ~n793 ) | ( n792 & ~n793 ) ;
  assign n795 = ~x74 & x202 ;
  assign n796 = ~x75 & x203 ;
  assign n797 = n795 | n796 ;
  assign n798 = x72 & ~x200 ;
  assign n799 = ( x73 & ~x201 ) | ( x73 & n798 ) | ( ~x201 & n798 ) ;
  assign n800 = x74 & ~x202 ;
  assign n801 = ( ~n797 & n799 ) | ( ~n797 & n800 ) | ( n799 & n800 ) ;
  assign n802 = ~n797 & n801 ;
  assign n803 = x203 & ~n802 ;
  assign n804 = ( x75 & n802 ) | ( x75 & ~n803 ) | ( n802 & ~n803 ) ;
  assign n805 = ~x73 & x201 ;
  assign n806 = ~x72 & x200 ;
  assign n807 = n805 | n806 ;
  assign n808 = n797 | n807 ;
  assign n809 = ~n804 & n808 ;
  assign n810 = ( n794 & n804 ) | ( n794 & ~n809 ) | ( n804 & ~n809 ) ;
  assign n811 = ~x77 & x205 ;
  assign n812 = ~x76 & x204 ;
  assign n813 = n811 | n812 ;
  assign n814 = ( n576 & n810 ) | ( n576 & ~n813 ) | ( n810 & ~n813 ) ;
  assign n815 = ~n576 & n814 ;
  assign n816 = ( ~n570 & n575 ) | ( ~n570 & n815 ) | ( n575 & n815 ) ;
  assign n817 = n570 | n816 ;
  assign n818 = ( ~n566 & n567 ) | ( ~n566 & n817 ) | ( n567 & n817 ) ;
  assign n819 = ~n566 & n818 ;
  assign n820 = ( n562 & ~n565 ) | ( n562 & n819 ) | ( ~n565 & n819 ) ;
  assign n821 = ~n562 & n820 ;
  assign n822 = x81 & ~x209 ;
  assign n823 = x208 | n566 ;
  assign n824 = ~n822 & n823 ;
  assign n825 = ( x80 & n822 ) | ( x80 & ~n824 ) | ( n822 & ~n824 ) ;
  assign n826 = x210 & ~n825 ;
  assign n827 = ( x82 & n825 ) | ( x82 & ~n826 ) | ( n825 & ~n826 ) ;
  assign n828 = ( n563 & ~n564 ) | ( n563 & n827 ) | ( ~n564 & n827 ) ;
  assign n829 = ~n563 & n828 ;
  assign n830 = x83 & ~x211 ;
  assign n831 = ( ~n821 & n829 ) | ( ~n821 & n830 ) | ( n829 & n830 ) ;
  assign n832 = n821 | n831 ;
  assign n833 = ~x85 & x213 ;
  assign n834 = ~x84 & x212 ;
  assign n835 = n833 | n834 ;
  assign n836 = ( n561 & n832 ) | ( n561 & ~n835 ) | ( n832 & ~n835 ) ;
  assign n837 = ~n561 & n836 ;
  assign n838 = ( ~n555 & n560 ) | ( ~n555 & n837 ) | ( n560 & n837 ) ;
  assign n839 = n555 | n838 ;
  assign n840 = x215 & ~n839 ;
  assign n841 = ( x87 & n839 ) | ( x87 & ~n840 ) | ( n839 & ~n840 ) ;
  assign n842 = ~x90 & x218 ;
  assign n843 = ~x91 & x219 ;
  assign n844 = n842 | n843 ;
  assign n845 = x88 & ~x216 ;
  assign n846 = ( x89 & ~x217 ) | ( x89 & n845 ) | ( ~x217 & n845 ) ;
  assign n847 = x90 & ~x218 ;
  assign n848 = ( ~n844 & n846 ) | ( ~n844 & n847 ) | ( n846 & n847 ) ;
  assign n849 = ~n844 & n848 ;
  assign n850 = x219 & ~n849 ;
  assign n851 = ( x91 & n849 ) | ( x91 & ~n850 ) | ( n849 & ~n850 ) ;
  assign n852 = ~x89 & x217 ;
  assign n853 = ~x88 & x216 ;
  assign n854 = n852 | n853 ;
  assign n855 = n844 | n854 ;
  assign n856 = ~n851 & n855 ;
  assign n857 = ( n841 & n851 ) | ( n841 & ~n856 ) | ( n851 & ~n856 ) ;
  assign n858 = ~x93 & x221 ;
  assign n859 = ~x92 & x220 ;
  assign n860 = n858 | n859 ;
  assign n861 = ( n552 & n857 ) | ( n552 & ~n860 ) | ( n857 & ~n860 ) ;
  assign n862 = ~n552 & n861 ;
  assign n863 = ( ~n546 & n551 ) | ( ~n546 & n862 ) | ( n551 & n862 ) ;
  assign n864 = n546 | n863 ;
  assign n865 = ( ~n542 & n543 ) | ( ~n542 & n864 ) | ( n543 & n864 ) ;
  assign n866 = ~n542 & n865 ;
  assign n867 = ( n538 & ~n541 ) | ( n538 & n866 ) | ( ~n541 & n866 ) ;
  assign n868 = ~n538 & n867 ;
  assign n869 = x97 & ~x225 ;
  assign n870 = x224 | n542 ;
  assign n871 = ~n869 & n870 ;
  assign n872 = ( x96 & n869 ) | ( x96 & ~n871 ) | ( n869 & ~n871 ) ;
  assign n873 = x226 & ~n872 ;
  assign n874 = ( x98 & n872 ) | ( x98 & ~n873 ) | ( n872 & ~n873 ) ;
  assign n875 = ( n539 & ~n540 ) | ( n539 & n874 ) | ( ~n540 & n874 ) ;
  assign n876 = ~n539 & n875 ;
  assign n877 = x99 & ~x227 ;
  assign n878 = ( ~n868 & n876 ) | ( ~n868 & n877 ) | ( n876 & n877 ) ;
  assign n879 = n868 | n878 ;
  assign n880 = ~x101 & x229 ;
  assign n881 = ~x100 & x228 ;
  assign n882 = n880 | n881 ;
  assign n883 = ( n537 & n879 ) | ( n537 & ~n882 ) | ( n879 & ~n882 ) ;
  assign n884 = ~n537 & n883 ;
  assign n885 = ( ~n531 & n536 ) | ( ~n531 & n884 ) | ( n536 & n884 ) ;
  assign n886 = n531 | n885 ;
  assign n887 = x231 & ~n886 ;
  assign n888 = ( x103 & n886 ) | ( x103 & ~n887 ) | ( n886 & ~n887 ) ;
  assign n889 = ~x106 & x234 ;
  assign n890 = ~x107 & x235 ;
  assign n891 = n889 | n890 ;
  assign n892 = x104 & ~x232 ;
  assign n893 = ( x105 & ~x233 ) | ( x105 & n892 ) | ( ~x233 & n892 ) ;
  assign n894 = x106 & ~x234 ;
  assign n895 = ( ~n891 & n893 ) | ( ~n891 & n894 ) | ( n893 & n894 ) ;
  assign n896 = ~n891 & n895 ;
  assign n897 = x235 & ~n896 ;
  assign n898 = ( x107 & n896 ) | ( x107 & ~n897 ) | ( n896 & ~n897 ) ;
  assign n899 = ~x105 & x233 ;
  assign n900 = ~x104 & x232 ;
  assign n901 = n899 | n900 ;
  assign n902 = n891 | n901 ;
  assign n903 = ~n898 & n902 ;
  assign n904 = ( n888 & n898 ) | ( n888 & ~n903 ) | ( n898 & ~n903 ) ;
  assign n905 = ~x109 & x237 ;
  assign n906 = ~x108 & x236 ;
  assign n907 = n905 | n906 ;
  assign n908 = ( n528 & n904 ) | ( n528 & ~n907 ) | ( n904 & ~n907 ) ;
  assign n909 = ~n528 & n908 ;
  assign n910 = ( ~n522 & n527 ) | ( ~n522 & n909 ) | ( n527 & n909 ) ;
  assign n911 = n522 | n910 ;
  assign n912 = x239 & ~n911 ;
  assign n913 = ( x111 & n911 ) | ( x111 & ~n912 ) | ( n911 & ~n912 ) ;
  assign n914 = n913 ^ x113 ^ 1'b0 ;
  assign n915 = ( x113 & ~x241 ) | ( x113 & n914 ) | ( ~x241 & n914 ) ;
  assign n916 = ( n913 & ~n914 ) | ( n913 & n915 ) | ( ~n914 & n915 ) ;
  assign n917 = ( n516 & ~n519 ) | ( n516 & n916 ) | ( ~n519 & n916 ) ;
  assign n918 = ~n516 & n917 ;
  assign n919 = ~x113 & x241 ;
  assign n920 = x240 | n919 ;
  assign n921 = x112 & ~n920 ;
  assign n922 = x241 & ~n921 ;
  assign n923 = ( x113 & n921 ) | ( x113 & ~n922 ) | ( n921 & ~n922 ) ;
  assign n924 = x242 & ~n923 ;
  assign n925 = ( x114 & n923 ) | ( x114 & ~n924 ) | ( n923 & ~n924 ) ;
  assign n926 = ( n517 & ~n518 ) | ( n517 & n925 ) | ( ~n518 & n925 ) ;
  assign n927 = ~n517 & n926 ;
  assign n928 = x115 & ~x243 ;
  assign n929 = ( ~n918 & n927 ) | ( ~n918 & n928 ) | ( n927 & n928 ) ;
  assign n930 = n918 | n929 ;
  assign n931 = ~x117 & x245 ;
  assign n932 = ~x116 & x244 ;
  assign n933 = n931 | n932 ;
  assign n934 = ( n515 & n930 ) | ( n515 & ~n933 ) | ( n930 & ~n933 ) ;
  assign n935 = ~n515 & n934 ;
  assign n936 = x116 & ~x244 ;
  assign n937 = ( x117 & ~x245 ) | ( x117 & n936 ) | ( ~x245 & n936 ) ;
  assign n938 = ( n513 & ~n514 ) | ( n513 & n937 ) | ( ~n514 & n937 ) ;
  assign n939 = ~n513 & n938 ;
  assign n940 = x246 | n513 ;
  assign n941 = x118 & ~n940 ;
  assign n942 = ( ~n935 & n939 ) | ( ~n935 & n941 ) | ( n939 & n941 ) ;
  assign n943 = n935 | n942 ;
  assign n944 = x247 & ~n943 ;
  assign n945 = ( x119 & n943 ) | ( x119 & ~n944 ) | ( n943 & ~n944 ) ;
  assign n946 = ~x122 & x250 ;
  assign n947 = ~x123 & x251 ;
  assign n948 = n946 | n947 ;
  assign n949 = x120 & ~x248 ;
  assign n950 = ( x121 & ~x249 ) | ( x121 & n949 ) | ( ~x249 & n949 ) ;
  assign n951 = x122 & ~x250 ;
  assign n952 = ( ~n948 & n950 ) | ( ~n948 & n951 ) | ( n950 & n951 ) ;
  assign n953 = ~n948 & n952 ;
  assign n954 = x251 & ~n953 ;
  assign n955 = ( x123 & n953 ) | ( x123 & ~n954 ) | ( n953 & ~n954 ) ;
  assign n956 = ~x121 & x249 ;
  assign n957 = ~x120 & x248 ;
  assign n958 = n956 | n957 ;
  assign n959 = n948 | n958 ;
  assign n960 = ~n955 & n959 ;
  assign n961 = ( n945 & n955 ) | ( n945 & ~n960 ) | ( n955 & ~n960 ) ;
  assign n962 = x127 & ~x255 ;
  assign n963 = ~x126 & x254 ;
  assign n964 = ~x125 & x253 ;
  assign n965 = n963 | n964 ;
  assign n966 = x125 & ~x253 ;
  assign n967 = x124 & ~x252 ;
  assign n968 = ( ~n965 & n966 ) | ( ~n965 & n967 ) | ( n966 & n967 ) ;
  assign n969 = ~n965 & n968 ;
  assign n970 = x126 & ~x254 ;
  assign n971 = ( ~n962 & n969 ) | ( ~n962 & n970 ) | ( n969 & n970 ) ;
  assign n972 = ~n962 & n971 ;
  assign n973 = n962 | n965 ;
  assign n974 = ~x124 & x252 ;
  assign n975 = n973 | n974 ;
  assign n976 = ~n972 & n975 ;
  assign n977 = ( n961 & n972 ) | ( n961 & ~n976 ) | ( n972 & ~n976 ) ;
  assign n978 = ~x127 & x255 ;
  assign n979 = n977 | n978 ;
  assign n980 = n979 ^ x0 ^ 1'b0 ;
  assign n981 = ( x0 & x128 ) | ( x0 & ~n980 ) | ( x128 & ~n980 ) ;
  assign n982 = ~x375 & x503 ;
  assign n983 = ~x374 & x502 ;
  assign n984 = n982 | n983 ;
  assign n985 = ~x368 & x496 ;
  assign n986 = ~x370 & x498 ;
  assign n987 = ~x371 & x499 ;
  assign n988 = n986 | n987 ;
  assign n989 = ~x367 & x495 ;
  assign n990 = x494 | n989 ;
  assign n991 = x366 & ~n990 ;
  assign n992 = ~x366 & x494 ;
  assign n993 = x364 & ~x492 ;
  assign n994 = ( x365 & ~x493 ) | ( x365 & n993 ) | ( ~x493 & n993 ) ;
  assign n995 = ( n989 & ~n992 ) | ( n989 & n994 ) | ( ~n992 & n994 ) ;
  assign n996 = ~n989 & n995 ;
  assign n997 = n989 | n992 ;
  assign n998 = ~x359 & x487 ;
  assign n999 = x486 | n998 ;
  assign n1000 = x358 & ~n999 ;
  assign n1001 = ~x358 & x486 ;
  assign n1002 = x356 & ~x484 ;
  assign n1003 = ( x357 & ~x485 ) | ( x357 & n1002 ) | ( ~x485 & n1002 ) ;
  assign n1004 = ( n998 & ~n1001 ) | ( n998 & n1003 ) | ( ~n1001 & n1003 ) ;
  assign n1005 = ~n998 & n1004 ;
  assign n1006 = n998 | n1001 ;
  assign n1007 = ~x352 & x480 ;
  assign n1008 = ~x354 & x482 ;
  assign n1009 = ~x355 & x483 ;
  assign n1010 = n1008 | n1009 ;
  assign n1011 = ~x351 & x479 ;
  assign n1012 = x478 | n1011 ;
  assign n1013 = x350 & ~n1012 ;
  assign n1014 = ~x350 & x478 ;
  assign n1015 = x348 & ~x476 ;
  assign n1016 = ( x349 & ~x477 ) | ( x349 & n1015 ) | ( ~x477 & n1015 ) ;
  assign n1017 = ( n1011 & ~n1014 ) | ( n1011 & n1016 ) | ( ~n1014 & n1016 ) ;
  assign n1018 = ~n1011 & n1017 ;
  assign n1019 = n1011 | n1014 ;
  assign n1020 = ~x343 & x471 ;
  assign n1021 = x470 | n1020 ;
  assign n1022 = x342 & ~n1021 ;
  assign n1023 = ~x342 & x470 ;
  assign n1024 = x340 & ~x468 ;
  assign n1025 = ( x341 & ~x469 ) | ( x341 & n1024 ) | ( ~x469 & n1024 ) ;
  assign n1026 = ( n1020 & ~n1023 ) | ( n1020 & n1025 ) | ( ~n1023 & n1025 ) ;
  assign n1027 = ~n1020 & n1026 ;
  assign n1028 = n1020 | n1023 ;
  assign n1029 = ~x336 & x464 ;
  assign n1030 = ~x338 & x466 ;
  assign n1031 = ~x339 & x467 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = ~x335 & x463 ;
  assign n1034 = x462 | n1033 ;
  assign n1035 = x334 & ~n1034 ;
  assign n1036 = ~x334 & x462 ;
  assign n1037 = x332 & ~x460 ;
  assign n1038 = ( x333 & ~x461 ) | ( x333 & n1037 ) | ( ~x461 & n1037 ) ;
  assign n1039 = ( n1033 & ~n1036 ) | ( n1033 & n1038 ) | ( ~n1036 & n1038 ) ;
  assign n1040 = ~n1033 & n1039 ;
  assign n1041 = n1033 | n1036 ;
  assign n1042 = ~x327 & x455 ;
  assign n1043 = x454 | n1042 ;
  assign n1044 = x326 & ~n1043 ;
  assign n1045 = ~x326 & x454 ;
  assign n1046 = x324 & ~x452 ;
  assign n1047 = ( x325 & ~x453 ) | ( x325 & n1046 ) | ( ~x453 & n1046 ) ;
  assign n1048 = ( n1042 & ~n1045 ) | ( n1042 & n1047 ) | ( ~n1045 & n1047 ) ;
  assign n1049 = ~n1042 & n1048 ;
  assign n1050 = n1042 | n1045 ;
  assign n1051 = ~x322 & x450 ;
  assign n1052 = ~x323 & x451 ;
  assign n1053 = ~x321 & x449 ;
  assign n1054 = ~x320 & x448 ;
  assign n1055 = ~x319 & x447 ;
  assign n1056 = ~x318 & x446 ;
  assign n1057 = n1055 | n1056 ;
  assign n1058 = ~x316 & x444 ;
  assign n1059 = ~x317 & x445 ;
  assign n1060 = n1058 | n1059 ;
  assign n1061 = n1057 | n1060 ;
  assign n1062 = ~x314 & x442 ;
  assign n1063 = ~x315 & x443 ;
  assign n1064 = x312 & ~x440 ;
  assign n1065 = ( x313 & ~x441 ) | ( x313 & n1064 ) | ( ~x441 & n1064 ) ;
  assign n1066 = x442 & ~n1065 ;
  assign n1067 = ( x314 & n1065 ) | ( x314 & ~n1066 ) | ( n1065 & ~n1066 ) ;
  assign n1068 = ( n1062 & ~n1063 ) | ( n1062 & n1067 ) | ( ~n1063 & n1067 ) ;
  assign n1069 = ~n1062 & n1068 ;
  assign n1070 = x315 & ~x443 ;
  assign n1071 = ( ~n1061 & n1069 ) | ( ~n1061 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1072 = ~n1061 & n1071 ;
  assign n1073 = n1062 | n1063 ;
  assign n1074 = ~x303 & x431 ;
  assign n1075 = ~x302 & x430 ;
  assign n1076 = n1074 | n1075 ;
  assign n1077 = ~x300 & x428 ;
  assign n1078 = ~x301 & x429 ;
  assign n1079 = n1077 | n1078 ;
  assign n1080 = n1076 | n1079 ;
  assign n1081 = ~x298 & x426 ;
  assign n1082 = ~x299 & x427 ;
  assign n1083 = x296 & ~x424 ;
  assign n1084 = ( x297 & ~x425 ) | ( x297 & n1083 ) | ( ~x425 & n1083 ) ;
  assign n1085 = x426 & ~n1084 ;
  assign n1086 = ( x298 & n1084 ) | ( x298 & ~n1085 ) | ( n1084 & ~n1085 ) ;
  assign n1087 = ( n1081 & ~n1082 ) | ( n1081 & n1086 ) | ( ~n1082 & n1086 ) ;
  assign n1088 = ~n1081 & n1087 ;
  assign n1089 = x299 & ~x427 ;
  assign n1090 = ( ~n1080 & n1088 ) | ( ~n1080 & n1089 ) | ( n1088 & n1089 ) ;
  assign n1091 = ~n1080 & n1090 ;
  assign n1092 = x300 & ~x428 ;
  assign n1093 = ( x301 & ~x429 ) | ( x301 & n1092 ) | ( ~x429 & n1092 ) ;
  assign n1094 = ( n1074 & ~n1075 ) | ( n1074 & n1093 ) | ( ~n1075 & n1093 ) ;
  assign n1095 = ~n1074 & n1094 ;
  assign n1096 = ~x288 & x416 ;
  assign n1097 = x256 & ~x384 ;
  assign n1098 = x257 & n1097 ;
  assign n1099 = x385 & ~n1098 ;
  assign n1100 = x257 | n1097 ;
  assign n1101 = ~x258 & x386 ;
  assign n1102 = ( n1099 & n1100 ) | ( n1099 & ~n1101 ) | ( n1100 & ~n1101 ) ;
  assign n1103 = ~n1099 & n1102 ;
  assign n1104 = x386 & ~n1103 ;
  assign n1105 = ( x258 & n1103 ) | ( x258 & ~n1104 ) | ( n1103 & ~n1104 ) ;
  assign n1106 = ( x259 & ~x387 ) | ( x259 & n1105 ) | ( ~x387 & n1105 ) ;
  assign n1107 = ( x260 & ~x388 ) | ( x260 & n1106 ) | ( ~x388 & n1106 ) ;
  assign n1108 = ( x261 & ~x389 ) | ( x261 & n1107 ) | ( ~x389 & n1107 ) ;
  assign n1109 = ( x262 & ~x390 ) | ( x262 & n1108 ) | ( ~x390 & n1108 ) ;
  assign n1110 = ( x263 & ~x391 ) | ( x263 & n1109 ) | ( ~x391 & n1109 ) ;
  assign n1111 = ( x264 & ~x392 ) | ( x264 & n1110 ) | ( ~x392 & n1110 ) ;
  assign n1112 = ( x265 & ~x393 ) | ( x265 & n1111 ) | ( ~x393 & n1111 ) ;
  assign n1113 = ( x266 & ~x394 ) | ( x266 & n1112 ) | ( ~x394 & n1112 ) ;
  assign n1114 = ( x267 & ~x395 ) | ( x267 & n1113 ) | ( ~x395 & n1113 ) ;
  assign n1115 = ( x268 & ~x396 ) | ( x268 & n1114 ) | ( ~x396 & n1114 ) ;
  assign n1116 = ( x269 & ~x397 ) | ( x269 & n1115 ) | ( ~x397 & n1115 ) ;
  assign n1117 = ( x270 & ~x398 ) | ( x270 & n1116 ) | ( ~x398 & n1116 ) ;
  assign n1118 = ( x271 & ~x399 ) | ( x271 & n1117 ) | ( ~x399 & n1117 ) ;
  assign n1119 = ( x272 & ~x400 ) | ( x272 & n1118 ) | ( ~x400 & n1118 ) ;
  assign n1120 = ( x273 & ~x401 ) | ( x273 & n1119 ) | ( ~x401 & n1119 ) ;
  assign n1121 = ( x274 & ~x402 ) | ( x274 & n1120 ) | ( ~x402 & n1120 ) ;
  assign n1122 = ( x275 & ~x403 ) | ( x275 & n1121 ) | ( ~x403 & n1121 ) ;
  assign n1123 = ( x276 & ~x404 ) | ( x276 & n1122 ) | ( ~x404 & n1122 ) ;
  assign n1124 = ( x277 & ~x405 ) | ( x277 & n1123 ) | ( ~x405 & n1123 ) ;
  assign n1125 = ( x278 & ~x406 ) | ( x278 & n1124 ) | ( ~x406 & n1124 ) ;
  assign n1126 = ( x279 & ~x407 ) | ( x279 & n1125 ) | ( ~x407 & n1125 ) ;
  assign n1127 = ( x280 & ~x408 ) | ( x280 & n1126 ) | ( ~x408 & n1126 ) ;
  assign n1128 = ( x281 & ~x409 ) | ( x281 & n1127 ) | ( ~x409 & n1127 ) ;
  assign n1129 = ( x282 & ~x410 ) | ( x282 & n1128 ) | ( ~x410 & n1128 ) ;
  assign n1130 = ( x283 & ~x411 ) | ( x283 & n1129 ) | ( ~x411 & n1129 ) ;
  assign n1131 = ( x284 & ~x412 ) | ( x284 & n1130 ) | ( ~x412 & n1130 ) ;
  assign n1132 = ( x285 & ~x413 ) | ( x285 & n1131 ) | ( ~x413 & n1131 ) ;
  assign n1133 = ( x286 & ~x414 ) | ( x286 & n1132 ) | ( ~x414 & n1132 ) ;
  assign n1134 = ( x287 & ~x415 ) | ( x287 & n1133 ) | ( ~x415 & n1133 ) ;
  assign n1135 = ~x295 & x423 ;
  assign n1136 = ~x294 & x422 ;
  assign n1137 = n1135 | n1136 ;
  assign n1138 = ~x292 & x420 ;
  assign n1139 = ~x293 & x421 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = n1137 | n1140 ;
  assign n1142 = ~x289 & x417 ;
  assign n1143 = ~x290 & x418 ;
  assign n1144 = ~x291 & x419 ;
  assign n1145 = n1143 | n1144 ;
  assign n1146 = n1142 | n1145 ;
  assign n1147 = n1141 | n1146 ;
  assign n1148 = ( n1096 & n1134 ) | ( n1096 & ~n1147 ) | ( n1134 & ~n1147 ) ;
  assign n1149 = ~n1096 & n1148 ;
  assign n1150 = x295 & ~x423 ;
  assign n1151 = x422 | n1135 ;
  assign n1152 = x294 & ~n1151 ;
  assign n1153 = x292 & ~x420 ;
  assign n1154 = ( x293 & ~x421 ) | ( x293 & n1153 ) | ( ~x421 & n1153 ) ;
  assign n1155 = ( n1135 & ~n1136 ) | ( n1135 & n1154 ) | ( ~n1136 & n1154 ) ;
  assign n1156 = ~n1135 & n1155 ;
  assign n1157 = x289 & ~x417 ;
  assign n1158 = x416 | n1142 ;
  assign n1159 = ~n1157 & n1158 ;
  assign n1160 = ( x288 & n1157 ) | ( x288 & ~n1159 ) | ( n1157 & ~n1159 ) ;
  assign n1161 = x290 & ~x418 ;
  assign n1162 = ( ~n1145 & n1160 ) | ( ~n1145 & n1161 ) | ( n1160 & n1161 ) ;
  assign n1163 = ~n1145 & n1162 ;
  assign n1164 = x291 & ~x419 ;
  assign n1165 = ( ~n1141 & n1163 ) | ( ~n1141 & n1164 ) | ( n1163 & n1164 ) ;
  assign n1166 = ~n1141 & n1165 ;
  assign n1167 = ( ~n1152 & n1156 ) | ( ~n1152 & n1166 ) | ( n1156 & n1166 ) ;
  assign n1168 = n1152 | n1167 ;
  assign n1169 = ( ~n1149 & n1150 ) | ( ~n1149 & n1168 ) | ( n1150 & n1168 ) ;
  assign n1170 = n1149 | n1169 ;
  assign n1171 = n1081 | n1082 ;
  assign n1172 = ~x297 & x425 ;
  assign n1173 = ~x296 & x424 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = n1171 | n1174 ;
  assign n1176 = ( n1080 & n1170 ) | ( n1080 & ~n1175 ) | ( n1170 & ~n1175 ) ;
  assign n1177 = ~n1080 & n1176 ;
  assign n1178 = x430 | n1074 ;
  assign n1179 = ~n1177 & n1178 ;
  assign n1180 = ( x302 & n1177 ) | ( x302 & ~n1179 ) | ( n1177 & ~n1179 ) ;
  assign n1181 = ( ~n1091 & n1095 ) | ( ~n1091 & n1180 ) | ( n1095 & n1180 ) ;
  assign n1182 = n1091 | n1181 ;
  assign n1183 = x431 & ~n1182 ;
  assign n1184 = ( x303 & n1182 ) | ( x303 & ~n1183 ) | ( n1182 & ~n1183 ) ;
  assign n1185 = ~x310 & x438 ;
  assign n1186 = ~x311 & x439 ;
  assign n1187 = n1185 | n1186 ;
  assign n1188 = x308 & ~x436 ;
  assign n1189 = ( x309 & ~x437 ) | ( x309 & n1188 ) | ( ~x437 & n1188 ) ;
  assign n1190 = x310 & ~x438 ;
  assign n1191 = ( ~n1187 & n1189 ) | ( ~n1187 & n1190 ) | ( n1189 & n1190 ) ;
  assign n1192 = ~n1187 & n1191 ;
  assign n1193 = ~x309 & x437 ;
  assign n1194 = ~x308 & x436 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = n1187 | n1195 ;
  assign n1197 = ~x306 & x434 ;
  assign n1198 = ~x307 & x435 ;
  assign n1199 = n1197 | n1198 ;
  assign n1200 = x305 & ~x433 ;
  assign n1201 = ~x305 & x433 ;
  assign n1202 = x432 | n1201 ;
  assign n1203 = ~n1200 & n1202 ;
  assign n1204 = ( x304 & n1200 ) | ( x304 & ~n1203 ) | ( n1200 & ~n1203 ) ;
  assign n1205 = x306 & ~x434 ;
  assign n1206 = ( ~n1199 & n1204 ) | ( ~n1199 & n1205 ) | ( n1204 & n1205 ) ;
  assign n1207 = ~n1199 & n1206 ;
  assign n1208 = x435 & ~n1207 ;
  assign n1209 = ( x307 & n1207 ) | ( x307 & ~n1208 ) | ( n1207 & ~n1208 ) ;
  assign n1210 = ( n1192 & ~n1196 ) | ( n1192 & n1209 ) | ( ~n1196 & n1209 ) ;
  assign n1211 = n1196 ^ n1192 ^ 1'b0 ;
  assign n1212 = ( n1192 & n1210 ) | ( n1192 & ~n1211 ) | ( n1210 & ~n1211 ) ;
  assign n1213 = x439 & ~n1212 ;
  assign n1214 = ( x311 & n1212 ) | ( x311 & ~n1213 ) | ( n1212 & ~n1213 ) ;
  assign n1215 = ~x304 & x432 ;
  assign n1216 = n1199 | n1201 ;
  assign n1217 = ( n1196 & ~n1215 ) | ( n1196 & n1216 ) | ( ~n1215 & n1216 ) ;
  assign n1218 = n1215 | n1217 ;
  assign n1219 = ~n1214 & n1218 ;
  assign n1220 = ( n1184 & n1214 ) | ( n1184 & ~n1219 ) | ( n1214 & ~n1219 ) ;
  assign n1221 = ~x313 & x441 ;
  assign n1222 = ~x312 & x440 ;
  assign n1223 = n1221 | n1222 ;
  assign n1224 = n1061 | n1223 ;
  assign n1225 = ( n1073 & n1220 ) | ( n1073 & ~n1224 ) | ( n1220 & ~n1224 ) ;
  assign n1226 = ~n1073 & n1225 ;
  assign n1227 = x446 | n1055 ;
  assign n1228 = ~n1226 & n1227 ;
  assign n1229 = ( x318 & n1226 ) | ( x318 & ~n1228 ) | ( n1226 & ~n1228 ) ;
  assign n1230 = x316 & ~x444 ;
  assign n1231 = ( x317 & ~x445 ) | ( x317 & n1230 ) | ( ~x445 & n1230 ) ;
  assign n1232 = ( n1055 & ~n1056 ) | ( n1055 & n1231 ) | ( ~n1056 & n1231 ) ;
  assign n1233 = ~n1055 & n1232 ;
  assign n1234 = ( ~n1072 & n1229 ) | ( ~n1072 & n1233 ) | ( n1229 & n1233 ) ;
  assign n1235 = n1072 | n1234 ;
  assign n1236 = x447 & ~n1235 ;
  assign n1237 = ( x319 & n1235 ) | ( x319 & ~n1236 ) | ( n1235 & ~n1236 ) ;
  assign n1238 = ( n1053 & ~n1054 ) | ( n1053 & n1237 ) | ( ~n1054 & n1237 ) ;
  assign n1239 = ~n1053 & n1238 ;
  assign n1240 = ( n1051 & ~n1052 ) | ( n1051 & n1239 ) | ( ~n1052 & n1239 ) ;
  assign n1241 = ~n1051 & n1240 ;
  assign n1242 = x320 & ~x448 ;
  assign n1243 = ( x321 & ~x449 ) | ( x321 & n1242 ) | ( ~x449 & n1242 ) ;
  assign n1244 = x450 & ~n1243 ;
  assign n1245 = ( x322 & n1243 ) | ( x322 & ~n1244 ) | ( n1243 & ~n1244 ) ;
  assign n1246 = ( n1051 & ~n1052 ) | ( n1051 & n1245 ) | ( ~n1052 & n1245 ) ;
  assign n1247 = ~n1051 & n1246 ;
  assign n1248 = x323 & ~x451 ;
  assign n1249 = ( ~n1241 & n1247 ) | ( ~n1241 & n1248 ) | ( n1247 & n1248 ) ;
  assign n1250 = n1241 | n1249 ;
  assign n1251 = ~x325 & x453 ;
  assign n1252 = ~x324 & x452 ;
  assign n1253 = n1251 | n1252 ;
  assign n1254 = ( n1050 & n1250 ) | ( n1050 & ~n1253 ) | ( n1250 & ~n1253 ) ;
  assign n1255 = ~n1050 & n1254 ;
  assign n1256 = ( ~n1044 & n1049 ) | ( ~n1044 & n1255 ) | ( n1049 & n1255 ) ;
  assign n1257 = n1044 | n1256 ;
  assign n1258 = x455 & ~n1257 ;
  assign n1259 = ( x327 & n1257 ) | ( x327 & ~n1258 ) | ( n1257 & ~n1258 ) ;
  assign n1260 = ~x330 & x458 ;
  assign n1261 = ~x331 & x459 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = x328 & ~x456 ;
  assign n1264 = ( x329 & ~x457 ) | ( x329 & n1263 ) | ( ~x457 & n1263 ) ;
  assign n1265 = x330 & ~x458 ;
  assign n1266 = ( ~n1262 & n1264 ) | ( ~n1262 & n1265 ) | ( n1264 & n1265 ) ;
  assign n1267 = ~n1262 & n1266 ;
  assign n1268 = x459 & ~n1267 ;
  assign n1269 = ( x331 & n1267 ) | ( x331 & ~n1268 ) | ( n1267 & ~n1268 ) ;
  assign n1270 = ~x329 & x457 ;
  assign n1271 = ~x328 & x456 ;
  assign n1272 = n1270 | n1271 ;
  assign n1273 = n1262 | n1272 ;
  assign n1274 = ~n1269 & n1273 ;
  assign n1275 = ( n1259 & n1269 ) | ( n1259 & ~n1274 ) | ( n1269 & ~n1274 ) ;
  assign n1276 = ~x333 & x461 ;
  assign n1277 = ~x332 & x460 ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = ( n1041 & n1275 ) | ( n1041 & ~n1278 ) | ( n1275 & ~n1278 ) ;
  assign n1280 = ~n1041 & n1279 ;
  assign n1281 = ( ~n1035 & n1040 ) | ( ~n1035 & n1280 ) | ( n1040 & n1280 ) ;
  assign n1282 = n1035 | n1281 ;
  assign n1283 = x463 & ~n1282 ;
  assign n1284 = ( x335 & n1282 ) | ( x335 & ~n1283 ) | ( n1282 & ~n1283 ) ;
  assign n1285 = n1284 ^ x337 ^ 1'b0 ;
  assign n1286 = ( x337 & ~x465 ) | ( x337 & n1285 ) | ( ~x465 & n1285 ) ;
  assign n1287 = ( n1284 & ~n1285 ) | ( n1284 & n1286 ) | ( ~n1285 & n1286 ) ;
  assign n1288 = ( n1029 & ~n1032 ) | ( n1029 & n1287 ) | ( ~n1032 & n1287 ) ;
  assign n1289 = ~n1029 & n1288 ;
  assign n1290 = ~x337 & x465 ;
  assign n1291 = x464 | n1290 ;
  assign n1292 = x336 & ~n1291 ;
  assign n1293 = x465 & ~n1292 ;
  assign n1294 = ( x337 & n1292 ) | ( x337 & ~n1293 ) | ( n1292 & ~n1293 ) ;
  assign n1295 = x466 & ~n1294 ;
  assign n1296 = ( x338 & n1294 ) | ( x338 & ~n1295 ) | ( n1294 & ~n1295 ) ;
  assign n1297 = ( n1030 & ~n1031 ) | ( n1030 & n1296 ) | ( ~n1031 & n1296 ) ;
  assign n1298 = ~n1030 & n1297 ;
  assign n1299 = x339 & ~x467 ;
  assign n1300 = ( ~n1289 & n1298 ) | ( ~n1289 & n1299 ) | ( n1298 & n1299 ) ;
  assign n1301 = n1289 | n1300 ;
  assign n1302 = ~x341 & x469 ;
  assign n1303 = ~x340 & x468 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = ( n1028 & n1301 ) | ( n1028 & ~n1304 ) | ( n1301 & ~n1304 ) ;
  assign n1306 = ~n1028 & n1305 ;
  assign n1307 = ( ~n1022 & n1027 ) | ( ~n1022 & n1306 ) | ( n1027 & n1306 ) ;
  assign n1308 = n1022 | n1307 ;
  assign n1309 = x471 & ~n1308 ;
  assign n1310 = ( x343 & n1308 ) | ( x343 & ~n1309 ) | ( n1308 & ~n1309 ) ;
  assign n1311 = ~x346 & x474 ;
  assign n1312 = ~x347 & x475 ;
  assign n1313 = n1311 | n1312 ;
  assign n1314 = x344 & ~x472 ;
  assign n1315 = ( x345 & ~x473 ) | ( x345 & n1314 ) | ( ~x473 & n1314 ) ;
  assign n1316 = x346 & ~x474 ;
  assign n1317 = ( ~n1313 & n1315 ) | ( ~n1313 & n1316 ) | ( n1315 & n1316 ) ;
  assign n1318 = ~n1313 & n1317 ;
  assign n1319 = x475 & ~n1318 ;
  assign n1320 = ( x347 & n1318 ) | ( x347 & ~n1319 ) | ( n1318 & ~n1319 ) ;
  assign n1321 = ~x345 & x473 ;
  assign n1322 = ~x344 & x472 ;
  assign n1323 = n1321 | n1322 ;
  assign n1324 = n1313 | n1323 ;
  assign n1325 = ~n1320 & n1324 ;
  assign n1326 = ( n1310 & n1320 ) | ( n1310 & ~n1325 ) | ( n1320 & ~n1325 ) ;
  assign n1327 = ~x349 & x477 ;
  assign n1328 = ~x348 & x476 ;
  assign n1329 = n1327 | n1328 ;
  assign n1330 = ( n1019 & n1326 ) | ( n1019 & ~n1329 ) | ( n1326 & ~n1329 ) ;
  assign n1331 = ~n1019 & n1330 ;
  assign n1332 = ( ~n1013 & n1018 ) | ( ~n1013 & n1331 ) | ( n1018 & n1331 ) ;
  assign n1333 = n1013 | n1332 ;
  assign n1334 = x479 & ~n1333 ;
  assign n1335 = ( x351 & n1333 ) | ( x351 & ~n1334 ) | ( n1333 & ~n1334 ) ;
  assign n1336 = n1335 ^ x353 ^ 1'b0 ;
  assign n1337 = ( x353 & ~x481 ) | ( x353 & n1336 ) | ( ~x481 & n1336 ) ;
  assign n1338 = ( n1335 & ~n1336 ) | ( n1335 & n1337 ) | ( ~n1336 & n1337 ) ;
  assign n1339 = ( n1007 & ~n1010 ) | ( n1007 & n1338 ) | ( ~n1010 & n1338 ) ;
  assign n1340 = ~n1007 & n1339 ;
  assign n1341 = ~x353 & x481 ;
  assign n1342 = x480 | n1341 ;
  assign n1343 = x352 & ~n1342 ;
  assign n1344 = x481 & ~n1343 ;
  assign n1345 = ( x353 & n1343 ) | ( x353 & ~n1344 ) | ( n1343 & ~n1344 ) ;
  assign n1346 = x482 & ~n1345 ;
  assign n1347 = ( x354 & n1345 ) | ( x354 & ~n1346 ) | ( n1345 & ~n1346 ) ;
  assign n1348 = ( n1008 & ~n1009 ) | ( n1008 & n1347 ) | ( ~n1009 & n1347 ) ;
  assign n1349 = ~n1008 & n1348 ;
  assign n1350 = x355 & ~x483 ;
  assign n1351 = ( ~n1340 & n1349 ) | ( ~n1340 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1352 = n1340 | n1351 ;
  assign n1353 = ~x357 & x485 ;
  assign n1354 = ~x356 & x484 ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = ( n1006 & n1352 ) | ( n1006 & ~n1355 ) | ( n1352 & ~n1355 ) ;
  assign n1357 = ~n1006 & n1356 ;
  assign n1358 = ( ~n1000 & n1005 ) | ( ~n1000 & n1357 ) | ( n1005 & n1357 ) ;
  assign n1359 = n1000 | n1358 ;
  assign n1360 = x487 & ~n1359 ;
  assign n1361 = ( x359 & n1359 ) | ( x359 & ~n1360 ) | ( n1359 & ~n1360 ) ;
  assign n1362 = ~x362 & x490 ;
  assign n1363 = ~x363 & x491 ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = x360 & ~x488 ;
  assign n1366 = ( x361 & ~x489 ) | ( x361 & n1365 ) | ( ~x489 & n1365 ) ;
  assign n1367 = x362 & ~x490 ;
  assign n1368 = ( ~n1364 & n1366 ) | ( ~n1364 & n1367 ) | ( n1366 & n1367 ) ;
  assign n1369 = ~n1364 & n1368 ;
  assign n1370 = x491 & ~n1369 ;
  assign n1371 = ( x363 & n1369 ) | ( x363 & ~n1370 ) | ( n1369 & ~n1370 ) ;
  assign n1372 = ~x361 & x489 ;
  assign n1373 = ~x360 & x488 ;
  assign n1374 = n1372 | n1373 ;
  assign n1375 = n1364 | n1374 ;
  assign n1376 = ~n1371 & n1375 ;
  assign n1377 = ( n1361 & n1371 ) | ( n1361 & ~n1376 ) | ( n1371 & ~n1376 ) ;
  assign n1378 = ~x365 & x493 ;
  assign n1379 = ~x364 & x492 ;
  assign n1380 = n1378 | n1379 ;
  assign n1381 = ( n997 & n1377 ) | ( n997 & ~n1380 ) | ( n1377 & ~n1380 ) ;
  assign n1382 = ~n997 & n1381 ;
  assign n1383 = ( ~n991 & n996 ) | ( ~n991 & n1382 ) | ( n996 & n1382 ) ;
  assign n1384 = n991 | n1383 ;
  assign n1385 = x495 & ~n1384 ;
  assign n1386 = ( x367 & n1384 ) | ( x367 & ~n1385 ) | ( n1384 & ~n1385 ) ;
  assign n1387 = n1386 ^ x369 ^ 1'b0 ;
  assign n1388 = ( x369 & ~x497 ) | ( x369 & n1387 ) | ( ~x497 & n1387 ) ;
  assign n1389 = ( n1386 & ~n1387 ) | ( n1386 & n1388 ) | ( ~n1387 & n1388 ) ;
  assign n1390 = ( n985 & ~n988 ) | ( n985 & n1389 ) | ( ~n988 & n1389 ) ;
  assign n1391 = ~n985 & n1390 ;
  assign n1392 = ~x369 & x497 ;
  assign n1393 = x496 | n1392 ;
  assign n1394 = x368 & ~n1393 ;
  assign n1395 = x497 & ~n1394 ;
  assign n1396 = ( x369 & n1394 ) | ( x369 & ~n1395 ) | ( n1394 & ~n1395 ) ;
  assign n1397 = x498 & ~n1396 ;
  assign n1398 = ( x370 & n1396 ) | ( x370 & ~n1397 ) | ( n1396 & ~n1397 ) ;
  assign n1399 = ( n986 & ~n987 ) | ( n986 & n1398 ) | ( ~n987 & n1398 ) ;
  assign n1400 = ~n986 & n1399 ;
  assign n1401 = x371 & ~x499 ;
  assign n1402 = ( ~n1391 & n1400 ) | ( ~n1391 & n1401 ) | ( n1400 & n1401 ) ;
  assign n1403 = n1391 | n1402 ;
  assign n1404 = ~x373 & x501 ;
  assign n1405 = ~x372 & x500 ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = ( n984 & n1403 ) | ( n984 & ~n1406 ) | ( n1403 & ~n1406 ) ;
  assign n1408 = ~n984 & n1407 ;
  assign n1409 = x372 & ~x500 ;
  assign n1410 = ( x373 & ~x501 ) | ( x373 & n1409 ) | ( ~x501 & n1409 ) ;
  assign n1411 = ( n982 & ~n983 ) | ( n982 & n1410 ) | ( ~n983 & n1410 ) ;
  assign n1412 = ~n982 & n1411 ;
  assign n1413 = x502 | n982 ;
  assign n1414 = x374 & ~n1413 ;
  assign n1415 = ( ~n1408 & n1412 ) | ( ~n1408 & n1414 ) | ( n1412 & n1414 ) ;
  assign n1416 = n1408 | n1415 ;
  assign n1417 = x503 & ~n1416 ;
  assign n1418 = ( x375 & n1416 ) | ( x375 & ~n1417 ) | ( n1416 & ~n1417 ) ;
  assign n1419 = ~x378 & x506 ;
  assign n1420 = ~x379 & x507 ;
  assign n1421 = n1419 | n1420 ;
  assign n1422 = x376 & ~x504 ;
  assign n1423 = ( x377 & ~x505 ) | ( x377 & n1422 ) | ( ~x505 & n1422 ) ;
  assign n1424 = x378 & ~x506 ;
  assign n1425 = ( ~n1421 & n1423 ) | ( ~n1421 & n1424 ) | ( n1423 & n1424 ) ;
  assign n1426 = ~n1421 & n1425 ;
  assign n1427 = x507 & ~n1426 ;
  assign n1428 = ( x379 & n1426 ) | ( x379 & ~n1427 ) | ( n1426 & ~n1427 ) ;
  assign n1429 = ~x377 & x505 ;
  assign n1430 = ~x376 & x504 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = n1421 | n1431 ;
  assign n1433 = ~n1428 & n1432 ;
  assign n1434 = ( n1418 & n1428 ) | ( n1418 & ~n1433 ) | ( n1428 & ~n1433 ) ;
  assign n1435 = x383 & ~x511 ;
  assign n1436 = ~x382 & x510 ;
  assign n1437 = ~x381 & x509 ;
  assign n1438 = n1436 | n1437 ;
  assign n1439 = x381 & ~x509 ;
  assign n1440 = x380 & ~x508 ;
  assign n1441 = ( ~n1438 & n1439 ) | ( ~n1438 & n1440 ) | ( n1439 & n1440 ) ;
  assign n1442 = ~n1438 & n1441 ;
  assign n1443 = x382 & ~x510 ;
  assign n1444 = ( ~n1435 & n1442 ) | ( ~n1435 & n1443 ) | ( n1442 & n1443 ) ;
  assign n1445 = ~n1435 & n1444 ;
  assign n1446 = n1435 | n1438 ;
  assign n1447 = ~x380 & x508 ;
  assign n1448 = n1446 | n1447 ;
  assign n1449 = ~n1445 & n1448 ;
  assign n1450 = ( n1434 & n1445 ) | ( n1434 & ~n1449 ) | ( n1445 & ~n1449 ) ;
  assign n1451 = ~x383 & x511 ;
  assign n1452 = n1450 | n1451 ;
  assign n1453 = n1452 ^ x256 ^ 1'b0 ;
  assign n1454 = ( x256 & x384 ) | ( x256 & ~n1453 ) | ( x384 & ~n1453 ) ;
  assign n1455 = x511 | n1450 ;
  assign n1456 = x383 & n1455 ;
  assign n1457 = x255 | n977 ;
  assign n1458 = x127 & n1457 ;
  assign n1459 = n1456 & ~n1458 ;
  assign n1460 = n979 ^ x123 ^ 1'b0 ;
  assign n1461 = ( x123 & x251 ) | ( x123 & ~n1460 ) | ( x251 & ~n1460 ) ;
  assign n1462 = n1452 ^ x379 ^ 1'b0 ;
  assign n1463 = ( x379 & x507 ) | ( x379 & ~n1462 ) | ( x507 & ~n1462 ) ;
  assign n1464 = n1461 & ~n1463 ;
  assign n1465 = n1452 ^ x378 ^ 1'b0 ;
  assign n1466 = ( x378 & x506 ) | ( x378 & ~n1465 ) | ( x506 & ~n1465 ) ;
  assign n1467 = n979 ^ x122 ^ 1'b0 ;
  assign n1468 = ( x122 & x250 ) | ( x122 & ~n1467 ) | ( x250 & ~n1467 ) ;
  assign n1469 = n1466 & ~n1468 ;
  assign n1470 = ~n1461 & n1463 ;
  assign n1471 = n1469 | n1470 ;
  assign n1472 = n979 ^ x121 ^ 1'b0 ;
  assign n1473 = ( x121 & x249 ) | ( x121 & ~n1472 ) | ( x249 & ~n1472 ) ;
  assign n1474 = n1452 ^ x377 ^ 1'b0 ;
  assign n1475 = ( x377 & x505 ) | ( x377 & ~n1474 ) | ( x505 & ~n1474 ) ;
  assign n1476 = ~n1473 & n1475 ;
  assign n1477 = n1452 ^ x376 ^ 1'b0 ;
  assign n1478 = ( x376 & x504 ) | ( x376 & ~n1477 ) | ( x504 & ~n1477 ) ;
  assign n1479 = n979 ^ x120 ^ 1'b0 ;
  assign n1480 = ( x120 & x248 ) | ( x120 & ~n1479 ) | ( x248 & ~n1479 ) ;
  assign n1481 = n1478 & ~n1480 ;
  assign n1482 = n1476 | n1481 ;
  assign n1483 = n979 ^ x119 ^ 1'b0 ;
  assign n1484 = ( x119 & x247 ) | ( x119 & ~n1483 ) | ( x247 & ~n1483 ) ;
  assign n1485 = n1452 ^ x375 ^ 1'b0 ;
  assign n1486 = ( x375 & x503 ) | ( x375 & ~n1485 ) | ( x503 & ~n1485 ) ;
  assign n1487 = ~n1484 & n1486 ;
  assign n1488 = n1452 ^ x374 ^ 1'b0 ;
  assign n1489 = ( x374 & x502 ) | ( x374 & ~n1488 ) | ( x502 & ~n1488 ) ;
  assign n1490 = n979 ^ x118 ^ 1'b0 ;
  assign n1491 = ( x118 & x246 ) | ( x118 & ~n1490 ) | ( x246 & ~n1490 ) ;
  assign n1492 = n1489 & ~n1491 ;
  assign n1493 = n1487 | n1492 ;
  assign n1494 = n979 ^ x117 ^ 1'b0 ;
  assign n1495 = ( x117 & x245 ) | ( x117 & ~n1494 ) | ( x245 & ~n1494 ) ;
  assign n1496 = n1452 ^ x373 ^ 1'b0 ;
  assign n1497 = ( x373 & x501 ) | ( x373 & ~n1496 ) | ( x501 & ~n1496 ) ;
  assign n1498 = n1495 & ~n1497 ;
  assign n1499 = n979 ^ x116 ^ 1'b0 ;
  assign n1500 = ( x116 & x244 ) | ( x116 & ~n1499 ) | ( x244 & ~n1499 ) ;
  assign n1501 = ~n1495 & n1497 ;
  assign n1502 = n1452 ^ x372 ^ 1'b0 ;
  assign n1503 = ( x372 & x500 ) | ( x372 & ~n1502 ) | ( x500 & ~n1502 ) ;
  assign n1504 = n1501 | n1503 ;
  assign n1505 = n1500 & ~n1504 ;
  assign n1506 = ( ~n1493 & n1498 ) | ( ~n1493 & n1505 ) | ( n1498 & n1505 ) ;
  assign n1507 = ~n1493 & n1506 ;
  assign n1508 = n1452 ^ x368 ^ 1'b0 ;
  assign n1509 = ( x368 & x496 ) | ( x368 & ~n1508 ) | ( x496 & ~n1508 ) ;
  assign n1510 = n979 ^ x112 ^ 1'b0 ;
  assign n1511 = ( x112 & x240 ) | ( x112 & ~n1510 ) | ( x240 & ~n1510 ) ;
  assign n1512 = n1509 & ~n1511 ;
  assign n1513 = n1452 ^ x370 ^ 1'b0 ;
  assign n1514 = ( x370 & x498 ) | ( x370 & ~n1513 ) | ( x498 & ~n1513 ) ;
  assign n1515 = n979 ^ x114 ^ 1'b0 ;
  assign n1516 = ( x114 & x242 ) | ( x114 & ~n1515 ) | ( x242 & ~n1515 ) ;
  assign n1517 = n1514 & ~n1516 ;
  assign n1518 = n979 ^ x115 ^ 1'b0 ;
  assign n1519 = ( x115 & x243 ) | ( x115 & ~n1518 ) | ( x243 & ~n1518 ) ;
  assign n1520 = n1452 ^ x371 ^ 1'b0 ;
  assign n1521 = ( x371 & x499 ) | ( x371 & ~n1520 ) | ( x499 & ~n1520 ) ;
  assign n1522 = ~n1519 & n1521 ;
  assign n1523 = n1517 | n1522 ;
  assign n1524 = n979 ^ x113 ^ 1'b0 ;
  assign n1525 = ( x113 & x241 ) | ( x113 & ~n1524 ) | ( x241 & ~n1524 ) ;
  assign n1526 = n1452 ^ x369 ^ 1'b0 ;
  assign n1527 = ( x369 & x497 ) | ( x369 & ~n1526 ) | ( x497 & ~n1526 ) ;
  assign n1528 = ~n1525 & n1527 ;
  assign n1529 = n979 ^ x111 ^ 1'b0 ;
  assign n1530 = ( x111 & x239 ) | ( x111 & ~n1529 ) | ( x239 & ~n1529 ) ;
  assign n1531 = n1452 ^ x367 ^ 1'b0 ;
  assign n1532 = ( x367 & x495 ) | ( x367 & ~n1531 ) | ( x495 & ~n1531 ) ;
  assign n1533 = n1530 & ~n1532 ;
  assign n1534 = ~n1530 & n1532 ;
  assign n1535 = n1452 ^ x366 ^ 1'b0 ;
  assign n1536 = ( x366 & x494 ) | ( x366 & ~n1535 ) | ( x494 & ~n1535 ) ;
  assign n1537 = n979 ^ x110 ^ 1'b0 ;
  assign n1538 = ( x110 & x238 ) | ( x110 & ~n1537 ) | ( x238 & ~n1537 ) ;
  assign n1539 = n1536 & ~n1538 ;
  assign n1540 = n1534 | n1539 ;
  assign n1541 = n979 ^ x103 ^ 1'b0 ;
  assign n1542 = ( x103 & x231 ) | ( x103 & ~n1541 ) | ( x231 & ~n1541 ) ;
  assign n1543 = n1452 ^ x359 ^ 1'b0 ;
  assign n1544 = ( x359 & x487 ) | ( x359 & ~n1543 ) | ( x487 & ~n1543 ) ;
  assign n1545 = ~n1542 & n1544 ;
  assign n1546 = n1452 ^ x358 ^ 1'b0 ;
  assign n1547 = ( x358 & x486 ) | ( x358 & ~n1546 ) | ( x486 & ~n1546 ) ;
  assign n1548 = n979 ^ x102 ^ 1'b0 ;
  assign n1549 = ( x102 & x230 ) | ( x102 & ~n1548 ) | ( x230 & ~n1548 ) ;
  assign n1550 = n1547 & ~n1549 ;
  assign n1551 = n1545 | n1550 ;
  assign n1552 = n1452 ^ x352 ^ 1'b0 ;
  assign n1553 = ( x352 & x480 ) | ( x352 & ~n1552 ) | ( x480 & ~n1552 ) ;
  assign n1554 = n979 ^ x96 ^ 1'b0 ;
  assign n1555 = ( x96 & x224 ) | ( x96 & ~n1554 ) | ( x224 & ~n1554 ) ;
  assign n1556 = n1553 & ~n1555 ;
  assign n1557 = n1452 ^ x354 ^ 1'b0 ;
  assign n1558 = ( x354 & x482 ) | ( x354 & ~n1557 ) | ( x482 & ~n1557 ) ;
  assign n1559 = n979 ^ x98 ^ 1'b0 ;
  assign n1560 = ( x98 & x226 ) | ( x98 & ~n1559 ) | ( x226 & ~n1559 ) ;
  assign n1561 = n1558 & ~n1560 ;
  assign n1562 = n979 ^ x99 ^ 1'b0 ;
  assign n1563 = ( x99 & x227 ) | ( x99 & ~n1562 ) | ( x227 & ~n1562 ) ;
  assign n1564 = n1452 ^ x355 ^ 1'b0 ;
  assign n1565 = ( x355 & x483 ) | ( x355 & ~n1564 ) | ( x483 & ~n1564 ) ;
  assign n1566 = ~n1563 & n1565 ;
  assign n1567 = n1561 | n1566 ;
  assign n1568 = n979 ^ x97 ^ 1'b0 ;
  assign n1569 = ( x97 & x225 ) | ( x97 & ~n1568 ) | ( x225 & ~n1568 ) ;
  assign n1570 = n1452 ^ x353 ^ 1'b0 ;
  assign n1571 = ( x353 & x481 ) | ( x353 & ~n1570 ) | ( x481 & ~n1570 ) ;
  assign n1572 = ~n1569 & n1571 ;
  assign n1573 = n979 ^ x95 ^ 1'b0 ;
  assign n1574 = ( x95 & x223 ) | ( x95 & ~n1573 ) | ( x223 & ~n1573 ) ;
  assign n1575 = n1452 ^ x351 ^ 1'b0 ;
  assign n1576 = ( x351 & x479 ) | ( x351 & ~n1575 ) | ( x479 & ~n1575 ) ;
  assign n1577 = n1574 & ~n1576 ;
  assign n1578 = ~n1574 & n1576 ;
  assign n1579 = n1452 ^ x350 ^ 1'b0 ;
  assign n1580 = ( x350 & x478 ) | ( x350 & ~n1579 ) | ( x478 & ~n1579 ) ;
  assign n1581 = n979 ^ x94 ^ 1'b0 ;
  assign n1582 = ( x94 & x222 ) | ( x94 & ~n1581 ) | ( x222 & ~n1581 ) ;
  assign n1583 = n1580 & ~n1582 ;
  assign n1584 = n1578 | n1583 ;
  assign n1585 = n979 ^ x87 ^ 1'b0 ;
  assign n1586 = ( x87 & x215 ) | ( x87 & ~n1585 ) | ( x215 & ~n1585 ) ;
  assign n1587 = n1452 ^ x343 ^ 1'b0 ;
  assign n1588 = ( x343 & x471 ) | ( x343 & ~n1587 ) | ( x471 & ~n1587 ) ;
  assign n1589 = ~n1586 & n1588 ;
  assign n1590 = n1452 ^ x342 ^ 1'b0 ;
  assign n1591 = ( x342 & x470 ) | ( x342 & ~n1590 ) | ( x470 & ~n1590 ) ;
  assign n1592 = n979 ^ x86 ^ 1'b0 ;
  assign n1593 = ( x86 & x214 ) | ( x86 & ~n1592 ) | ( x214 & ~n1592 ) ;
  assign n1594 = n1591 & ~n1593 ;
  assign n1595 = n1589 | n1594 ;
  assign n1596 = n1452 ^ x336 ^ 1'b0 ;
  assign n1597 = ( x336 & x464 ) | ( x336 & ~n1596 ) | ( x464 & ~n1596 ) ;
  assign n1598 = n979 ^ x80 ^ 1'b0 ;
  assign n1599 = ( x80 & x208 ) | ( x80 & ~n1598 ) | ( x208 & ~n1598 ) ;
  assign n1600 = n1597 & ~n1599 ;
  assign n1601 = n1452 ^ x338 ^ 1'b0 ;
  assign n1602 = ( x338 & x466 ) | ( x338 & ~n1601 ) | ( x466 & ~n1601 ) ;
  assign n1603 = n979 ^ x82 ^ 1'b0 ;
  assign n1604 = ( x82 & x210 ) | ( x82 & ~n1603 ) | ( x210 & ~n1603 ) ;
  assign n1605 = n1602 & ~n1604 ;
  assign n1606 = n979 ^ x83 ^ 1'b0 ;
  assign n1607 = ( x83 & x211 ) | ( x83 & ~n1606 ) | ( x211 & ~n1606 ) ;
  assign n1608 = n1452 ^ x339 ^ 1'b0 ;
  assign n1609 = ( x339 & x467 ) | ( x339 & ~n1608 ) | ( x467 & ~n1608 ) ;
  assign n1610 = ~n1607 & n1609 ;
  assign n1611 = n1605 | n1610 ;
  assign n1612 = n979 ^ x81 ^ 1'b0 ;
  assign n1613 = ( x81 & x209 ) | ( x81 & ~n1612 ) | ( x209 & ~n1612 ) ;
  assign n1614 = n1452 ^ x337 ^ 1'b0 ;
  assign n1615 = ( x337 & x465 ) | ( x337 & ~n1614 ) | ( x465 & ~n1614 ) ;
  assign n1616 = ~n1613 & n1615 ;
  assign n1617 = n979 ^ x79 ^ 1'b0 ;
  assign n1618 = ( x79 & x207 ) | ( x79 & ~n1617 ) | ( x207 & ~n1617 ) ;
  assign n1619 = n1452 ^ x335 ^ 1'b0 ;
  assign n1620 = ( x335 & x463 ) | ( x335 & ~n1619 ) | ( x463 & ~n1619 ) ;
  assign n1621 = n1618 & ~n1620 ;
  assign n1622 = ~n1618 & n1620 ;
  assign n1623 = n1452 ^ x334 ^ 1'b0 ;
  assign n1624 = ( x334 & x462 ) | ( x334 & ~n1623 ) | ( x462 & ~n1623 ) ;
  assign n1625 = n979 ^ x78 ^ 1'b0 ;
  assign n1626 = ( x78 & x206 ) | ( x78 & ~n1625 ) | ( x206 & ~n1625 ) ;
  assign n1627 = n1624 & ~n1626 ;
  assign n1628 = n1622 | n1627 ;
  assign n1629 = n979 ^ x71 ^ 1'b0 ;
  assign n1630 = ( x71 & x199 ) | ( x71 & ~n1629 ) | ( x199 & ~n1629 ) ;
  assign n1631 = n1452 ^ x327 ^ 1'b0 ;
  assign n1632 = ( x327 & x455 ) | ( x327 & ~n1631 ) | ( x455 & ~n1631 ) ;
  assign n1633 = ~n1630 & n1632 ;
  assign n1634 = n1452 ^ x326 ^ 1'b0 ;
  assign n1635 = ( x326 & x454 ) | ( x326 & ~n1634 ) | ( x454 & ~n1634 ) ;
  assign n1636 = n979 ^ x70 ^ 1'b0 ;
  assign n1637 = ( x70 & x198 ) | ( x70 & ~n1636 ) | ( x198 & ~n1636 ) ;
  assign n1638 = n1635 & ~n1637 ;
  assign n1639 = n1633 | n1638 ;
  assign n1640 = n979 ^ x67 ^ 1'b0 ;
  assign n1641 = ( x67 & x195 ) | ( x67 & ~n1640 ) | ( x195 & ~n1640 ) ;
  assign n1642 = n1452 ^ x323 ^ 1'b0 ;
  assign n1643 = ( x323 & x451 ) | ( x323 & ~n1642 ) | ( x451 & ~n1642 ) ;
  assign n1644 = ~n1641 & n1643 ;
  assign n1645 = n1452 ^ x322 ^ 1'b0 ;
  assign n1646 = ( x322 & x450 ) | ( x322 & ~n1645 ) | ( x450 & ~n1645 ) ;
  assign n1647 = n979 ^ x66 ^ 1'b0 ;
  assign n1648 = ( x66 & x194 ) | ( x66 & ~n1647 ) | ( x194 & ~n1647 ) ;
  assign n1649 = n1646 & ~n1648 ;
  assign n1650 = n1452 ^ x320 ^ 1'b0 ;
  assign n1651 = ( x320 & x448 ) | ( x320 & ~n1650 ) | ( x448 & ~n1650 ) ;
  assign n1652 = n979 ^ x64 ^ 1'b0 ;
  assign n1653 = ( x64 & x192 ) | ( x64 & ~n1652 ) | ( x192 & ~n1652 ) ;
  assign n1654 = n1651 & ~n1653 ;
  assign n1655 = n979 ^ x65 ^ 1'b0 ;
  assign n1656 = ( x65 & x193 ) | ( x65 & ~n1655 ) | ( x193 & ~n1655 ) ;
  assign n1657 = n1452 ^ x321 ^ 1'b0 ;
  assign n1658 = ( x321 & x449 ) | ( x321 & ~n1657 ) | ( x449 & ~n1657 ) ;
  assign n1659 = ~n1656 & n1658 ;
  assign n1660 = n979 ^ x63 ^ 1'b0 ;
  assign n1661 = ( x63 & x191 ) | ( x63 & ~n1660 ) | ( x191 & ~n1660 ) ;
  assign n1662 = n1452 ^ x319 ^ 1'b0 ;
  assign n1663 = ( x319 & x447 ) | ( x319 & ~n1662 ) | ( x447 & ~n1662 ) ;
  assign n1664 = ~n1661 & n1663 ;
  assign n1665 = n1452 ^ x318 ^ 1'b0 ;
  assign n1666 = ( x318 & x446 ) | ( x318 & ~n1665 ) | ( x446 & ~n1665 ) ;
  assign n1667 = n979 ^ x62 ^ 1'b0 ;
  assign n1668 = ( x62 & x190 ) | ( x62 & ~n1667 ) | ( x190 & ~n1667 ) ;
  assign n1669 = n1666 & ~n1668 ;
  assign n1670 = n1664 | n1669 ;
  assign n1671 = n979 ^ x60 ^ 1'b0 ;
  assign n1672 = ( x60 & x188 ) | ( x60 & ~n1671 ) | ( x188 & ~n1671 ) ;
  assign n1673 = n1452 ^ x316 ^ 1'b0 ;
  assign n1674 = ( x316 & x444 ) | ( x316 & ~n1673 ) | ( x444 & ~n1673 ) ;
  assign n1675 = ~n1672 & n1674 ;
  assign n1676 = n979 ^ x61 ^ 1'b0 ;
  assign n1677 = ( x61 & x189 ) | ( x61 & ~n1676 ) | ( x189 & ~n1676 ) ;
  assign n1678 = n1452 ^ x317 ^ 1'b0 ;
  assign n1679 = ( x317 & x445 ) | ( x317 & ~n1678 ) | ( x445 & ~n1678 ) ;
  assign n1680 = ~n1677 & n1679 ;
  assign n1681 = n1675 | n1680 ;
  assign n1682 = n1670 | n1681 ;
  assign n1683 = n979 ^ x59 ^ 1'b0 ;
  assign n1684 = ( x59 & x187 ) | ( x59 & ~n1683 ) | ( x187 & ~n1683 ) ;
  assign n1685 = n1452 ^ x315 ^ 1'b0 ;
  assign n1686 = ( x315 & x443 ) | ( x315 & ~n1685 ) | ( x443 & ~n1685 ) ;
  assign n1687 = n1684 & ~n1686 ;
  assign n1688 = n979 ^ x58 ^ 1'b0 ;
  assign n1689 = ( x58 & x186 ) | ( x58 & ~n1688 ) | ( x186 & ~n1688 ) ;
  assign n1690 = n1452 ^ x314 ^ 1'b0 ;
  assign n1691 = ( x314 & x442 ) | ( x314 & ~n1690 ) | ( x442 & ~n1690 ) ;
  assign n1692 = ~n1689 & n1691 ;
  assign n1693 = ~n1684 & n1686 ;
  assign n1694 = n979 ^ x57 ^ 1'b0 ;
  assign n1695 = ( x57 & x185 ) | ( x57 & ~n1694 ) | ( x185 & ~n1694 ) ;
  assign n1696 = n1452 ^ x313 ^ 1'b0 ;
  assign n1697 = ( x313 & x441 ) | ( x313 & ~n1696 ) | ( x441 & ~n1696 ) ;
  assign n1698 = n979 ^ x56 ^ 1'b0 ;
  assign n1699 = ( x56 & x184 ) | ( x56 & ~n1698 ) | ( x184 & ~n1698 ) ;
  assign n1700 = n1452 ^ x312 ^ 1'b0 ;
  assign n1701 = ( x312 & x440 ) | ( x312 & ~n1700 ) | ( x440 & ~n1700 ) ;
  assign n1702 = n1699 & ~n1701 ;
  assign n1703 = ( n1695 & ~n1697 ) | ( n1695 & n1702 ) | ( ~n1697 & n1702 ) ;
  assign n1704 = n1691 & ~n1703 ;
  assign n1705 = ( n1689 & n1703 ) | ( n1689 & ~n1704 ) | ( n1703 & ~n1704 ) ;
  assign n1706 = ( n1692 & ~n1693 ) | ( n1692 & n1705 ) | ( ~n1693 & n1705 ) ;
  assign n1707 = ~n1692 & n1706 ;
  assign n1708 = ( ~n1682 & n1687 ) | ( ~n1682 & n1707 ) | ( n1687 & n1707 ) ;
  assign n1709 = ~n1682 & n1708 ;
  assign n1710 = n1692 | n1693 ;
  assign n1711 = n979 ^ x47 ^ 1'b0 ;
  assign n1712 = ( x47 & x175 ) | ( x47 & ~n1711 ) | ( x175 & ~n1711 ) ;
  assign n1713 = n1452 ^ x303 ^ 1'b0 ;
  assign n1714 = ( x303 & x431 ) | ( x303 & ~n1713 ) | ( x431 & ~n1713 ) ;
  assign n1715 = ~n1712 & n1714 ;
  assign n1716 = n1452 ^ x302 ^ 1'b0 ;
  assign n1717 = ( x302 & x430 ) | ( x302 & ~n1716 ) | ( x430 & ~n1716 ) ;
  assign n1718 = n979 ^ x46 ^ 1'b0 ;
  assign n1719 = ( x46 & x174 ) | ( x46 & ~n1718 ) | ( x174 & ~n1718 ) ;
  assign n1720 = n1717 & ~n1719 ;
  assign n1721 = n1715 | n1720 ;
  assign n1722 = n979 ^ x44 ^ 1'b0 ;
  assign n1723 = ( x44 & x172 ) | ( x44 & ~n1722 ) | ( x172 & ~n1722 ) ;
  assign n1724 = n1452 ^ x300 ^ 1'b0 ;
  assign n1725 = ( x300 & x428 ) | ( x300 & ~n1724 ) | ( x428 & ~n1724 ) ;
  assign n1726 = ~n1723 & n1725 ;
  assign n1727 = n979 ^ x45 ^ 1'b0 ;
  assign n1728 = ( x45 & x173 ) | ( x45 & ~n1727 ) | ( x173 & ~n1727 ) ;
  assign n1729 = n1452 ^ x301 ^ 1'b0 ;
  assign n1730 = ( x301 & x429 ) | ( x301 & ~n1729 ) | ( x429 & ~n1729 ) ;
  assign n1731 = ~n1728 & n1730 ;
  assign n1732 = n1726 | n1731 ;
  assign n1733 = n1721 | n1732 ;
  assign n1734 = n979 ^ x42 ^ 1'b0 ;
  assign n1735 = ( x42 & x170 ) | ( x42 & ~n1734 ) | ( x170 & ~n1734 ) ;
  assign n1736 = n1452 ^ x298 ^ 1'b0 ;
  assign n1737 = ( x298 & x426 ) | ( x298 & ~n1736 ) | ( x426 & ~n1736 ) ;
  assign n1738 = ~n1735 & n1737 ;
  assign n1739 = n979 ^ x43 ^ 1'b0 ;
  assign n1740 = ( x43 & x171 ) | ( x43 & ~n1739 ) | ( x171 & ~n1739 ) ;
  assign n1741 = n1452 ^ x299 ^ 1'b0 ;
  assign n1742 = ( x299 & x427 ) | ( x299 & ~n1741 ) | ( x427 & ~n1741 ) ;
  assign n1743 = ~n1740 & n1742 ;
  assign n1744 = n979 ^ x41 ^ 1'b0 ;
  assign n1745 = ( x41 & x169 ) | ( x41 & ~n1744 ) | ( x169 & ~n1744 ) ;
  assign n1746 = n1452 ^ x297 ^ 1'b0 ;
  assign n1747 = ( x297 & x425 ) | ( x297 & ~n1746 ) | ( x425 & ~n1746 ) ;
  assign n1748 = n979 ^ x40 ^ 1'b0 ;
  assign n1749 = ( x40 & x168 ) | ( x40 & ~n1748 ) | ( x168 & ~n1748 ) ;
  assign n1750 = n1452 ^ x296 ^ 1'b0 ;
  assign n1751 = ( x296 & x424 ) | ( x296 & ~n1750 ) | ( x424 & ~n1750 ) ;
  assign n1752 = n1749 & ~n1751 ;
  assign n1753 = ( n1745 & ~n1747 ) | ( n1745 & n1752 ) | ( ~n1747 & n1752 ) ;
  assign n1754 = n1737 & ~n1753 ;
  assign n1755 = ( n1735 & n1753 ) | ( n1735 & ~n1754 ) | ( n1753 & ~n1754 ) ;
  assign n1756 = ( n1738 & ~n1743 ) | ( n1738 & n1755 ) | ( ~n1743 & n1755 ) ;
  assign n1757 = ~n1738 & n1756 ;
  assign n1758 = n1740 & ~n1742 ;
  assign n1759 = ( ~n1733 & n1757 ) | ( ~n1733 & n1758 ) | ( n1757 & n1758 ) ;
  assign n1760 = ~n1733 & n1759 ;
  assign n1761 = n1452 ^ x288 ^ 1'b0 ;
  assign n1762 = ( x288 & x416 ) | ( x288 & ~n1761 ) | ( x416 & ~n1761 ) ;
  assign n1763 = n979 ^ x32 ^ 1'b0 ;
  assign n1764 = ( x32 & x160 ) | ( x32 & ~n1763 ) | ( x160 & ~n1763 ) ;
  assign n1765 = n1762 & ~n1764 ;
  assign n1766 = n979 ^ x31 ^ 1'b0 ;
  assign n1767 = ( x31 & x159 ) | ( x31 & ~n1766 ) | ( x159 & ~n1766 ) ;
  assign n1768 = n1452 ^ x287 ^ 1'b0 ;
  assign n1769 = ( x287 & x415 ) | ( x287 & ~n1768 ) | ( x415 & ~n1768 ) ;
  assign n1770 = n979 ^ x30 ^ 1'b0 ;
  assign n1771 = ( x30 & x158 ) | ( x30 & ~n1770 ) | ( x158 & ~n1770 ) ;
  assign n1772 = n1452 ^ x286 ^ 1'b0 ;
  assign n1773 = ( x286 & x414 ) | ( x286 & ~n1772 ) | ( x414 & ~n1772 ) ;
  assign n1774 = n979 ^ x29 ^ 1'b0 ;
  assign n1775 = ( x29 & x157 ) | ( x29 & ~n1774 ) | ( x157 & ~n1774 ) ;
  assign n1776 = n1452 ^ x285 ^ 1'b0 ;
  assign n1777 = ( x285 & x413 ) | ( x285 & ~n1776 ) | ( x413 & ~n1776 ) ;
  assign n1778 = n979 ^ x28 ^ 1'b0 ;
  assign n1779 = ( x28 & x156 ) | ( x28 & ~n1778 ) | ( x156 & ~n1778 ) ;
  assign n1780 = n1452 ^ x284 ^ 1'b0 ;
  assign n1781 = ( x284 & x412 ) | ( x284 & ~n1780 ) | ( x412 & ~n1780 ) ;
  assign n1782 = n979 ^ x27 ^ 1'b0 ;
  assign n1783 = ( x27 & x155 ) | ( x27 & ~n1782 ) | ( x155 & ~n1782 ) ;
  assign n1784 = n1452 ^ x283 ^ 1'b0 ;
  assign n1785 = ( x283 & x411 ) | ( x283 & ~n1784 ) | ( x411 & ~n1784 ) ;
  assign n1786 = n979 ^ x26 ^ 1'b0 ;
  assign n1787 = ( x26 & x154 ) | ( x26 & ~n1786 ) | ( x154 & ~n1786 ) ;
  assign n1788 = n1452 ^ x282 ^ 1'b0 ;
  assign n1789 = ( x282 & x410 ) | ( x282 & ~n1788 ) | ( x410 & ~n1788 ) ;
  assign n1790 = n1452 ^ x281 ^ 1'b0 ;
  assign n1791 = ( x281 & x409 ) | ( x281 & ~n1790 ) | ( x409 & ~n1790 ) ;
  assign n1792 = n1452 ^ x280 ^ 1'b0 ;
  assign n1793 = ( x280 & x408 ) | ( x280 & ~n1792 ) | ( x408 & ~n1792 ) ;
  assign n1794 = n979 ^ x23 ^ 1'b0 ;
  assign n1795 = ( x23 & x151 ) | ( x23 & ~n1794 ) | ( x151 & ~n1794 ) ;
  assign n1796 = n1452 ^ x279 ^ 1'b0 ;
  assign n1797 = ( x279 & x407 ) | ( x279 & ~n1796 ) | ( x407 & ~n1796 ) ;
  assign n1798 = n979 ^ x22 ^ 1'b0 ;
  assign n1799 = ( x22 & x150 ) | ( x22 & ~n1798 ) | ( x150 & ~n1798 ) ;
  assign n1800 = n1452 ^ x278 ^ 1'b0 ;
  assign n1801 = ( x278 & x406 ) | ( x278 & ~n1800 ) | ( x406 & ~n1800 ) ;
  assign n1802 = n979 ^ x21 ^ 1'b0 ;
  assign n1803 = ( x21 & x149 ) | ( x21 & ~n1802 ) | ( x149 & ~n1802 ) ;
  assign n1804 = n1452 ^ x277 ^ 1'b0 ;
  assign n1805 = ( x277 & x405 ) | ( x277 & ~n1804 ) | ( x405 & ~n1804 ) ;
  assign n1806 = n979 ^ x20 ^ 1'b0 ;
  assign n1807 = ( x20 & x148 ) | ( x20 & ~n1806 ) | ( x148 & ~n1806 ) ;
  assign n1808 = n1452 ^ x276 ^ 1'b0 ;
  assign n1809 = ( x276 & x404 ) | ( x276 & ~n1808 ) | ( x404 & ~n1808 ) ;
  assign n1810 = n979 ^ x19 ^ 1'b0 ;
  assign n1811 = ( x19 & x147 ) | ( x19 & ~n1810 ) | ( x147 & ~n1810 ) ;
  assign n1812 = n1452 ^ x275 ^ 1'b0 ;
  assign n1813 = ( x275 & x403 ) | ( x275 & ~n1812 ) | ( x403 & ~n1812 ) ;
  assign n1814 = n979 ^ x18 ^ 1'b0 ;
  assign n1815 = ( x18 & x146 ) | ( x18 & ~n1814 ) | ( x146 & ~n1814 ) ;
  assign n1816 = n1452 ^ x274 ^ 1'b0 ;
  assign n1817 = ( x274 & x402 ) | ( x274 & ~n1816 ) | ( x402 & ~n1816 ) ;
  assign n1818 = n1452 ^ x273 ^ 1'b0 ;
  assign n1819 = ( x273 & x401 ) | ( x273 & ~n1818 ) | ( x401 & ~n1818 ) ;
  assign n1820 = n1452 ^ x272 ^ 1'b0 ;
  assign n1821 = ( x272 & x400 ) | ( x272 & ~n1820 ) | ( x400 & ~n1820 ) ;
  assign n1822 = n979 ^ x15 ^ 1'b0 ;
  assign n1823 = ( x15 & x143 ) | ( x15 & ~n1822 ) | ( x143 & ~n1822 ) ;
  assign n1824 = n1452 ^ x271 ^ 1'b0 ;
  assign n1825 = ( x271 & x399 ) | ( x271 & ~n1824 ) | ( x399 & ~n1824 ) ;
  assign n1826 = n979 ^ x14 ^ 1'b0 ;
  assign n1827 = ( x14 & x142 ) | ( x14 & ~n1826 ) | ( x142 & ~n1826 ) ;
  assign n1828 = n1452 ^ x270 ^ 1'b0 ;
  assign n1829 = ( x270 & x398 ) | ( x270 & ~n1828 ) | ( x398 & ~n1828 ) ;
  assign n1830 = n979 ^ x13 ^ 1'b0 ;
  assign n1831 = ( x13 & x141 ) | ( x13 & ~n1830 ) | ( x141 & ~n1830 ) ;
  assign n1832 = n1452 ^ x269 ^ 1'b0 ;
  assign n1833 = ( x269 & x397 ) | ( x269 & ~n1832 ) | ( x397 & ~n1832 ) ;
  assign n1834 = n979 ^ x12 ^ 1'b0 ;
  assign n1835 = ( x12 & x140 ) | ( x12 & ~n1834 ) | ( x140 & ~n1834 ) ;
  assign n1836 = n1452 ^ x268 ^ 1'b0 ;
  assign n1837 = ( x268 & x396 ) | ( x268 & ~n1836 ) | ( x396 & ~n1836 ) ;
  assign n1838 = n979 ^ x11 ^ 1'b0 ;
  assign n1839 = ( x11 & x139 ) | ( x11 & ~n1838 ) | ( x139 & ~n1838 ) ;
  assign n1840 = n1452 ^ x267 ^ 1'b0 ;
  assign n1841 = ( x267 & x395 ) | ( x267 & ~n1840 ) | ( x395 & ~n1840 ) ;
  assign n1842 = n979 ^ x10 ^ 1'b0 ;
  assign n1843 = ( x10 & x138 ) | ( x10 & ~n1842 ) | ( x138 & ~n1842 ) ;
  assign n1844 = n1452 ^ x266 ^ 1'b0 ;
  assign n1845 = ( x266 & x394 ) | ( x266 & ~n1844 ) | ( x394 & ~n1844 ) ;
  assign n1846 = n1452 ^ x265 ^ 1'b0 ;
  assign n1847 = ( x265 & x393 ) | ( x265 & ~n1846 ) | ( x393 & ~n1846 ) ;
  assign n1848 = n1452 ^ x264 ^ 1'b0 ;
  assign n1849 = ( x264 & x392 ) | ( x264 & ~n1848 ) | ( x392 & ~n1848 ) ;
  assign n1850 = n979 ^ x7 ^ 1'b0 ;
  assign n1851 = ( x7 & x135 ) | ( x7 & ~n1850 ) | ( x135 & ~n1850 ) ;
  assign n1852 = n1452 ^ x263 ^ 1'b0 ;
  assign n1853 = ( x263 & x391 ) | ( x263 & ~n1852 ) | ( x391 & ~n1852 ) ;
  assign n1854 = n1452 ^ x262 ^ 1'b0 ;
  assign n1855 = ( x262 & x390 ) | ( x262 & ~n1854 ) | ( x390 & ~n1854 ) ;
  assign n1856 = n979 ^ x6 ^ 1'b0 ;
  assign n1857 = ( x6 & x134 ) | ( x6 & ~n1856 ) | ( x134 & ~n1856 ) ;
  assign n1858 = n1452 ^ x261 ^ 1'b0 ;
  assign n1859 = ( x261 & x389 ) | ( x261 & ~n1858 ) | ( x389 & ~n1858 ) ;
  assign n1860 = n979 ^ x5 ^ 1'b0 ;
  assign n1861 = ( x5 & x133 ) | ( x5 & ~n1860 ) | ( x133 & ~n1860 ) ;
  assign n1862 = n1452 ^ x260 ^ 1'b0 ;
  assign n1863 = ( x260 & x388 ) | ( x260 & ~n1862 ) | ( x388 & ~n1862 ) ;
  assign n1864 = n979 ^ x4 ^ 1'b0 ;
  assign n1865 = ( x4 & x132 ) | ( x4 & ~n1864 ) | ( x132 & ~n1864 ) ;
  assign n1866 = n979 ^ x3 ^ 1'b0 ;
  assign n1867 = ( x3 & x131 ) | ( x3 & ~n1866 ) | ( x131 & ~n1866 ) ;
  assign n1868 = n1452 ^ x259 ^ 1'b0 ;
  assign n1869 = ( x259 & x387 ) | ( x259 & ~n1868 ) | ( x387 & ~n1868 ) ;
  assign n1870 = n979 ^ x2 ^ 1'b0 ;
  assign n1871 = ( x2 & x130 ) | ( x2 & ~n1870 ) | ( x130 & ~n1870 ) ;
  assign n1872 = n1452 ^ x258 ^ 1'b0 ;
  assign n1873 = ( x258 & x386 ) | ( x258 & ~n1872 ) | ( x386 & ~n1872 ) ;
  assign n1874 = ~n1871 & n1873 ;
  assign n1875 = n979 ^ x1 ^ 1'b0 ;
  assign n1876 = ( x1 & x129 ) | ( x1 & ~n1875 ) | ( x129 & ~n1875 ) ;
  assign n1877 = n1452 ^ x257 ^ 1'b0 ;
  assign n1878 = ( x257 & x385 ) | ( x257 & ~n1877 ) | ( x385 & ~n1877 ) ;
  assign n1879 = n981 & ~n1454 ;
  assign n1880 = ~n1878 & n1879 ;
  assign n1881 = n1876 | n1880 ;
  assign n1882 = n1878 & ~n1879 ;
  assign n1883 = ( n1874 & n1881 ) | ( n1874 & ~n1882 ) | ( n1881 & ~n1882 ) ;
  assign n1884 = ~n1874 & n1883 ;
  assign n1885 = n1873 & ~n1884 ;
  assign n1886 = ( n1871 & n1884 ) | ( n1871 & ~n1885 ) | ( n1884 & ~n1885 ) ;
  assign n1887 = ( n1867 & ~n1869 ) | ( n1867 & n1886 ) | ( ~n1869 & n1886 ) ;
  assign n1888 = ( ~n1863 & n1865 ) | ( ~n1863 & n1887 ) | ( n1865 & n1887 ) ;
  assign n1889 = ( ~n1859 & n1861 ) | ( ~n1859 & n1888 ) | ( n1861 & n1888 ) ;
  assign n1890 = ( ~n1855 & n1857 ) | ( ~n1855 & n1889 ) | ( n1857 & n1889 ) ;
  assign n1891 = ( n1851 & ~n1853 ) | ( n1851 & n1890 ) | ( ~n1853 & n1890 ) ;
  assign n1892 = n979 ^ x8 ^ 1'b0 ;
  assign n1893 = ( x8 & x136 ) | ( x8 & ~n1892 ) | ( x136 & ~n1892 ) ;
  assign n1894 = ( ~n1849 & n1891 ) | ( ~n1849 & n1893 ) | ( n1891 & n1893 ) ;
  assign n1895 = n979 ^ x9 ^ 1'b0 ;
  assign n1896 = ( x9 & x137 ) | ( x9 & ~n1895 ) | ( x137 & ~n1895 ) ;
  assign n1897 = ( ~n1847 & n1894 ) | ( ~n1847 & n1896 ) | ( n1894 & n1896 ) ;
  assign n1898 = ( n1843 & ~n1845 ) | ( n1843 & n1897 ) | ( ~n1845 & n1897 ) ;
  assign n1899 = ( n1839 & ~n1841 ) | ( n1839 & n1898 ) | ( ~n1841 & n1898 ) ;
  assign n1900 = ( n1835 & ~n1837 ) | ( n1835 & n1899 ) | ( ~n1837 & n1899 ) ;
  assign n1901 = ( n1831 & ~n1833 ) | ( n1831 & n1900 ) | ( ~n1833 & n1900 ) ;
  assign n1902 = ( n1827 & ~n1829 ) | ( n1827 & n1901 ) | ( ~n1829 & n1901 ) ;
  assign n1903 = ( n1823 & ~n1825 ) | ( n1823 & n1902 ) | ( ~n1825 & n1902 ) ;
  assign n1904 = n979 ^ x16 ^ 1'b0 ;
  assign n1905 = ( x16 & x144 ) | ( x16 & ~n1904 ) | ( x144 & ~n1904 ) ;
  assign n1906 = ( ~n1821 & n1903 ) | ( ~n1821 & n1905 ) | ( n1903 & n1905 ) ;
  assign n1907 = n979 ^ x17 ^ 1'b0 ;
  assign n1908 = ( x17 & x145 ) | ( x17 & ~n1907 ) | ( x145 & ~n1907 ) ;
  assign n1909 = ( ~n1819 & n1906 ) | ( ~n1819 & n1908 ) | ( n1906 & n1908 ) ;
  assign n1910 = ( n1815 & ~n1817 ) | ( n1815 & n1909 ) | ( ~n1817 & n1909 ) ;
  assign n1911 = ( n1811 & ~n1813 ) | ( n1811 & n1910 ) | ( ~n1813 & n1910 ) ;
  assign n1912 = ( n1807 & ~n1809 ) | ( n1807 & n1911 ) | ( ~n1809 & n1911 ) ;
  assign n1913 = ( n1803 & ~n1805 ) | ( n1803 & n1912 ) | ( ~n1805 & n1912 ) ;
  assign n1914 = ( n1799 & ~n1801 ) | ( n1799 & n1913 ) | ( ~n1801 & n1913 ) ;
  assign n1915 = ( n1795 & ~n1797 ) | ( n1795 & n1914 ) | ( ~n1797 & n1914 ) ;
  assign n1916 = n979 ^ x24 ^ 1'b0 ;
  assign n1917 = ( x24 & x152 ) | ( x24 & ~n1916 ) | ( x152 & ~n1916 ) ;
  assign n1918 = ( ~n1793 & n1915 ) | ( ~n1793 & n1917 ) | ( n1915 & n1917 ) ;
  assign n1919 = n979 ^ x25 ^ 1'b0 ;
  assign n1920 = ( x25 & x153 ) | ( x25 & ~n1919 ) | ( x153 & ~n1919 ) ;
  assign n1921 = ( ~n1791 & n1918 ) | ( ~n1791 & n1920 ) | ( n1918 & n1920 ) ;
  assign n1922 = ( n1787 & ~n1789 ) | ( n1787 & n1921 ) | ( ~n1789 & n1921 ) ;
  assign n1923 = ( n1783 & ~n1785 ) | ( n1783 & n1922 ) | ( ~n1785 & n1922 ) ;
  assign n1924 = ( n1779 & ~n1781 ) | ( n1779 & n1923 ) | ( ~n1781 & n1923 ) ;
  assign n1925 = ( n1775 & ~n1777 ) | ( n1775 & n1924 ) | ( ~n1777 & n1924 ) ;
  assign n1926 = ( n1771 & ~n1773 ) | ( n1771 & n1925 ) | ( ~n1773 & n1925 ) ;
  assign n1927 = ( n1767 & ~n1769 ) | ( n1767 & n1926 ) | ( ~n1769 & n1926 ) ;
  assign n1928 = n979 ^ x39 ^ 1'b0 ;
  assign n1929 = ( x39 & x167 ) | ( x39 & ~n1928 ) | ( x167 & ~n1928 ) ;
  assign n1930 = n1452 ^ x295 ^ 1'b0 ;
  assign n1931 = ( x295 & x423 ) | ( x295 & ~n1930 ) | ( x423 & ~n1930 ) ;
  assign n1932 = ~n1929 & n1931 ;
  assign n1933 = n1452 ^ x294 ^ 1'b0 ;
  assign n1934 = ( x294 & x422 ) | ( x294 & ~n1933 ) | ( x422 & ~n1933 ) ;
  assign n1935 = n979 ^ x38 ^ 1'b0 ;
  assign n1936 = ( x38 & x166 ) | ( x38 & ~n1935 ) | ( x166 & ~n1935 ) ;
  assign n1937 = n1934 & ~n1936 ;
  assign n1938 = n1932 | n1937 ;
  assign n1939 = n979 ^ x36 ^ 1'b0 ;
  assign n1940 = ( x36 & x164 ) | ( x36 & ~n1939 ) | ( x164 & ~n1939 ) ;
  assign n1941 = n1452 ^ x292 ^ 1'b0 ;
  assign n1942 = ( x292 & x420 ) | ( x292 & ~n1941 ) | ( x420 & ~n1941 ) ;
  assign n1943 = ~n1940 & n1942 ;
  assign n1944 = n979 ^ x37 ^ 1'b0 ;
  assign n1945 = ( x37 & x165 ) | ( x37 & ~n1944 ) | ( x165 & ~n1944 ) ;
  assign n1946 = n1452 ^ x293 ^ 1'b0 ;
  assign n1947 = ( x293 & x421 ) | ( x293 & ~n1946 ) | ( x421 & ~n1946 ) ;
  assign n1948 = ~n1945 & n1947 ;
  assign n1949 = n1943 | n1948 ;
  assign n1950 = n1938 | n1949 ;
  assign n1951 = n979 ^ x33 ^ 1'b0 ;
  assign n1952 = ( x33 & x161 ) | ( x33 & ~n1951 ) | ( x161 & ~n1951 ) ;
  assign n1953 = n1452 ^ x289 ^ 1'b0 ;
  assign n1954 = ( x289 & x417 ) | ( x289 & ~n1953 ) | ( x417 & ~n1953 ) ;
  assign n1955 = ~n1952 & n1954 ;
  assign n1956 = n979 ^ x35 ^ 1'b0 ;
  assign n1957 = ( x35 & x163 ) | ( x35 & ~n1956 ) | ( x163 & ~n1956 ) ;
  assign n1958 = n1452 ^ x291 ^ 1'b0 ;
  assign n1959 = ( x291 & x419 ) | ( x291 & ~n1958 ) | ( x419 & ~n1958 ) ;
  assign n1960 = ~n1957 & n1959 ;
  assign n1961 = n1452 ^ x290 ^ 1'b0 ;
  assign n1962 = ( x290 & x418 ) | ( x290 & ~n1961 ) | ( x418 & ~n1961 ) ;
  assign n1963 = n979 ^ x34 ^ 1'b0 ;
  assign n1964 = ( x34 & x162 ) | ( x34 & ~n1963 ) | ( x162 & ~n1963 ) ;
  assign n1965 = n1962 & ~n1964 ;
  assign n1966 = ( ~n1955 & n1960 ) | ( ~n1955 & n1965 ) | ( n1960 & n1965 ) ;
  assign n1967 = n1955 | n1966 ;
  assign n1968 = n1950 | n1967 ;
  assign n1969 = ( n1765 & n1927 ) | ( n1765 & ~n1968 ) | ( n1927 & ~n1968 ) ;
  assign n1970 = ~n1765 & n1969 ;
  assign n1971 = n1929 & ~n1931 ;
  assign n1972 = ~n1762 & n1764 ;
  assign n1973 = n1952 & ~n1954 ;
  assign n1974 = ( ~n1967 & n1972 ) | ( ~n1967 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1975 = ~n1967 & n1974 ;
  assign n1976 = n1960 | n1962 ;
  assign n1977 = ~n1975 & n1976 ;
  assign n1978 = ( n1964 & n1975 ) | ( n1964 & ~n1977 ) | ( n1975 & ~n1977 ) ;
  assign n1979 = n1957 & ~n1959 ;
  assign n1980 = ( ~n1950 & n1978 ) | ( ~n1950 & n1979 ) | ( n1978 & n1979 ) ;
  assign n1981 = ~n1950 & n1980 ;
  assign n1982 = n1932 | n1934 ;
  assign n1983 = ~n1981 & n1982 ;
  assign n1984 = ( n1936 & n1981 ) | ( n1936 & ~n1983 ) | ( n1981 & ~n1983 ) ;
  assign n1985 = n1940 & ~n1942 ;
  assign n1986 = ( n1945 & ~n1947 ) | ( n1945 & n1985 ) | ( ~n1947 & n1985 ) ;
  assign n1987 = ( ~n1938 & n1984 ) | ( ~n1938 & n1986 ) | ( n1984 & n1986 ) ;
  assign n1988 = n1984 ^ n1938 ^ 1'b0 ;
  assign n1989 = ( n1984 & n1987 ) | ( n1984 & ~n1988 ) | ( n1987 & ~n1988 ) ;
  assign n1990 = ( ~n1970 & n1971 ) | ( ~n1970 & n1989 ) | ( n1971 & n1989 ) ;
  assign n1991 = n1970 | n1990 ;
  assign n1992 = n1738 | n1743 ;
  assign n1993 = ~n1745 & n1747 ;
  assign n1994 = ~n1749 & n1751 ;
  assign n1995 = n1993 | n1994 ;
  assign n1996 = n1992 | n1995 ;
  assign n1997 = ( n1733 & n1991 ) | ( n1733 & ~n1996 ) | ( n1991 & ~n1996 ) ;
  assign n1998 = ~n1733 & n1997 ;
  assign n1999 = ~n1717 & n1719 ;
  assign n2000 = ( ~n1715 & n1998 ) | ( ~n1715 & n1999 ) | ( n1998 & n1999 ) ;
  assign n2001 = n1998 ^ n1715 ^ 1'b0 ;
  assign n2002 = ( n1998 & n2000 ) | ( n1998 & ~n2001 ) | ( n2000 & ~n2001 ) ;
  assign n2003 = n1723 & ~n1725 ;
  assign n2004 = ( n1728 & ~n1730 ) | ( n1728 & n2003 ) | ( ~n1730 & n2003 ) ;
  assign n2005 = ( n1715 & ~n1720 ) | ( n1715 & n2004 ) | ( ~n1720 & n2004 ) ;
  assign n2006 = ~n1715 & n2005 ;
  assign n2007 = ( ~n1760 & n2002 ) | ( ~n1760 & n2006 ) | ( n2002 & n2006 ) ;
  assign n2008 = n1760 | n2007 ;
  assign n2009 = n1714 & ~n2008 ;
  assign n2010 = ( n1712 & n2008 ) | ( n1712 & ~n2009 ) | ( n2008 & ~n2009 ) ;
  assign n2011 = n979 ^ x55 ^ 1'b0 ;
  assign n2012 = ( x55 & x183 ) | ( x55 & ~n2011 ) | ( x183 & ~n2011 ) ;
  assign n2013 = n1452 ^ x310 ^ 1'b0 ;
  assign n2014 = ( x310 & x438 ) | ( x310 & ~n2013 ) | ( x438 & ~n2013 ) ;
  assign n2015 = n979 ^ x54 ^ 1'b0 ;
  assign n2016 = ( x54 & x182 ) | ( x54 & ~n2015 ) | ( x182 & ~n2015 ) ;
  assign n2017 = n2014 & ~n2016 ;
  assign n2018 = n1452 ^ x311 ^ 1'b0 ;
  assign n2019 = ( x311 & x439 ) | ( x311 & ~n2018 ) | ( x439 & ~n2018 ) ;
  assign n2020 = ~n2012 & n2019 ;
  assign n2021 = n2017 | n2020 ;
  assign n2022 = n979 ^ x53 ^ 1'b0 ;
  assign n2023 = ( x53 & x181 ) | ( x53 & ~n2022 ) | ( x181 & ~n2022 ) ;
  assign n2024 = n1452 ^ x309 ^ 1'b0 ;
  assign n2025 = ( x309 & x437 ) | ( x309 & ~n2024 ) | ( x437 & ~n2024 ) ;
  assign n2026 = n1452 ^ x308 ^ 1'b0 ;
  assign n2027 = ( x308 & x436 ) | ( x308 & ~n2026 ) | ( x436 & ~n2026 ) ;
  assign n2028 = n979 ^ x52 ^ 1'b0 ;
  assign n2029 = ( x52 & x180 ) | ( x52 & ~n2028 ) | ( x180 & ~n2028 ) ;
  assign n2030 = ~n2027 & n2029 ;
  assign n2031 = ( n2023 & ~n2025 ) | ( n2023 & n2030 ) | ( ~n2025 & n2030 ) ;
  assign n2032 = ~n2014 & n2016 ;
  assign n2033 = ( ~n2021 & n2031 ) | ( ~n2021 & n2032 ) | ( n2031 & n2032 ) ;
  assign n2034 = ~n2021 & n2033 ;
  assign n2035 = ~n2023 & n2025 ;
  assign n2036 = n2027 & ~n2029 ;
  assign n2037 = n2035 | n2036 ;
  assign n2038 = n2021 | n2037 ;
  assign n2039 = n979 ^ x51 ^ 1'b0 ;
  assign n2040 = ( x51 & x179 ) | ( x51 & ~n2039 ) | ( x179 & ~n2039 ) ;
  assign n2041 = n979 ^ x50 ^ 1'b0 ;
  assign n2042 = ( x50 & x178 ) | ( x50 & ~n2041 ) | ( x178 & ~n2041 ) ;
  assign n2043 = n979 ^ x49 ^ 1'b0 ;
  assign n2044 = ( x49 & x177 ) | ( x49 & ~n2043 ) | ( x177 & ~n2043 ) ;
  assign n2045 = n1452 ^ x305 ^ 1'b0 ;
  assign n2046 = ( x305 & x433 ) | ( x305 & ~n2045 ) | ( x433 & ~n2045 ) ;
  assign n2047 = ~n2044 & n2046 ;
  assign n2048 = n1452 ^ x307 ^ 1'b0 ;
  assign n2049 = ( x307 & x435 ) | ( x307 & ~n2048 ) | ( x435 & ~n2048 ) ;
  assign n2050 = ~n2040 & n2049 ;
  assign n2051 = n1452 ^ x306 ^ 1'b0 ;
  assign n2052 = ( x306 & x434 ) | ( x306 & ~n2051 ) | ( x434 & ~n2051 ) ;
  assign n2053 = ~n2042 & n2052 ;
  assign n2054 = ( ~n2047 & n2050 ) | ( ~n2047 & n2053 ) | ( n2050 & n2053 ) ;
  assign n2055 = n2047 | n2054 ;
  assign n2056 = n2044 & ~n2046 ;
  assign n2057 = n1452 ^ x304 ^ 1'b0 ;
  assign n2058 = ( x304 & x432 ) | ( x304 & ~n2057 ) | ( x432 & ~n2057 ) ;
  assign n2059 = n979 ^ x48 ^ 1'b0 ;
  assign n2060 = ( x48 & x176 ) | ( x48 & ~n2059 ) | ( x176 & ~n2059 ) ;
  assign n2061 = ~n2058 & n2060 ;
  assign n2062 = ( ~n2055 & n2056 ) | ( ~n2055 & n2061 ) | ( n2056 & n2061 ) ;
  assign n2063 = ~n2055 & n2062 ;
  assign n2064 = n2050 | n2052 ;
  assign n2065 = ~n2063 & n2064 ;
  assign n2066 = ( n2042 & n2063 ) | ( n2042 & ~n2065 ) | ( n2063 & ~n2065 ) ;
  assign n2067 = n2049 & ~n2066 ;
  assign n2068 = ( n2040 & n2066 ) | ( n2040 & ~n2067 ) | ( n2066 & ~n2067 ) ;
  assign n2069 = ( n2034 & ~n2038 ) | ( n2034 & n2068 ) | ( ~n2038 & n2068 ) ;
  assign n2070 = n2038 ^ n2034 ^ 1'b0 ;
  assign n2071 = ( n2034 & n2069 ) | ( n2034 & ~n2070 ) | ( n2069 & ~n2070 ) ;
  assign n2072 = n2019 & ~n2071 ;
  assign n2073 = ( n2012 & n2071 ) | ( n2012 & ~n2072 ) | ( n2071 & ~n2072 ) ;
  assign n2074 = n2038 | n2055 ;
  assign n2075 = n2058 & ~n2060 ;
  assign n2076 = n2074 | n2075 ;
  assign n2077 = ~n2073 & n2076 ;
  assign n2078 = ( n2010 & n2073 ) | ( n2010 & ~n2077 ) | ( n2073 & ~n2077 ) ;
  assign n2079 = ~n1695 & n1697 ;
  assign n2080 = ~n1699 & n1701 ;
  assign n2081 = n2079 | n2080 ;
  assign n2082 = n1682 | n2081 ;
  assign n2083 = ( n1710 & n2078 ) | ( n1710 & ~n2082 ) | ( n2078 & ~n2082 ) ;
  assign n2084 = ~n1710 & n2083 ;
  assign n2085 = ~n1666 & n1668 ;
  assign n2086 = ( ~n1664 & n2084 ) | ( ~n1664 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2087 = n2084 ^ n1664 ^ 1'b0 ;
  assign n2088 = ( n2084 & n2086 ) | ( n2084 & ~n2087 ) | ( n2086 & ~n2087 ) ;
  assign n2089 = n1672 & ~n1674 ;
  assign n2090 = ( n1677 & ~n1679 ) | ( n1677 & n2089 ) | ( ~n1679 & n2089 ) ;
  assign n2091 = ( n1664 & ~n1669 ) | ( n1664 & n2090 ) | ( ~n1669 & n2090 ) ;
  assign n2092 = ~n1664 & n2091 ;
  assign n2093 = ( ~n1709 & n2088 ) | ( ~n1709 & n2092 ) | ( n2088 & n2092 ) ;
  assign n2094 = n1709 | n2093 ;
  assign n2095 = n1663 & ~n2094 ;
  assign n2096 = ( n1661 & n2094 ) | ( n1661 & ~n2095 ) | ( n2094 & ~n2095 ) ;
  assign n2097 = ( n1654 & ~n1659 ) | ( n1654 & n2096 ) | ( ~n1659 & n2096 ) ;
  assign n2098 = ~n1654 & n2097 ;
  assign n2099 = ( n1644 & ~n1649 ) | ( n1644 & n2098 ) | ( ~n1649 & n2098 ) ;
  assign n2100 = ~n1644 & n2099 ;
  assign n2101 = n1656 & ~n1658 ;
  assign n2102 = n1651 | n1659 ;
  assign n2103 = ~n2101 & n2102 ;
  assign n2104 = ( n1653 & n2101 ) | ( n1653 & ~n2103 ) | ( n2101 & ~n2103 ) ;
  assign n2105 = ( ~n1646 & n1648 ) | ( ~n1646 & n2104 ) | ( n1648 & n2104 ) ;
  assign n2106 = n2104 ^ n1646 ^ 1'b0 ;
  assign n2107 = ( n2104 & n2105 ) | ( n2104 & ~n2106 ) | ( n2105 & ~n2106 ) ;
  assign n2108 = ( n1644 & ~n1649 ) | ( n1644 & n2107 ) | ( ~n1649 & n2107 ) ;
  assign n2109 = ~n1644 & n2108 ;
  assign n2110 = n1641 & ~n1643 ;
  assign n2111 = ( ~n2100 & n2109 ) | ( ~n2100 & n2110 ) | ( n2109 & n2110 ) ;
  assign n2112 = n2100 | n2111 ;
  assign n2113 = n979 ^ x69 ^ 1'b0 ;
  assign n2114 = ( x69 & x197 ) | ( x69 & ~n2113 ) | ( x197 & ~n2113 ) ;
  assign n2115 = n1452 ^ x325 ^ 1'b0 ;
  assign n2116 = ( x325 & x453 ) | ( x325 & ~n2115 ) | ( x453 & ~n2115 ) ;
  assign n2117 = ~n2114 & n2116 ;
  assign n2118 = n979 ^ x68 ^ 1'b0 ;
  assign n2119 = ( x68 & x196 ) | ( x68 & ~n2118 ) | ( x196 & ~n2118 ) ;
  assign n2120 = n1452 ^ x324 ^ 1'b0 ;
  assign n2121 = ( x324 & x452 ) | ( x324 & ~n2120 ) | ( x452 & ~n2120 ) ;
  assign n2122 = ~n2119 & n2121 ;
  assign n2123 = n2117 | n2122 ;
  assign n2124 = ( n1639 & n2112 ) | ( n1639 & ~n2123 ) | ( n2112 & ~n2123 ) ;
  assign n2125 = ~n1639 & n2124 ;
  assign n2126 = ~n1635 & n1637 ;
  assign n2127 = ( ~n1633 & n2125 ) | ( ~n1633 & n2126 ) | ( n2125 & n2126 ) ;
  assign n2128 = n2125 ^ n1633 ^ 1'b0 ;
  assign n2129 = ( n2125 & n2127 ) | ( n2125 & ~n2128 ) | ( n2127 & ~n2128 ) ;
  assign n2130 = n2119 & ~n2121 ;
  assign n2131 = ( n2114 & ~n2116 ) | ( n2114 & n2130 ) | ( ~n2116 & n2130 ) ;
  assign n2132 = ( ~n1639 & n2129 ) | ( ~n1639 & n2131 ) | ( n2129 & n2131 ) ;
  assign n2133 = n2129 ^ n1639 ^ 1'b0 ;
  assign n2134 = ( n2129 & n2132 ) | ( n2129 & ~n2133 ) | ( n2132 & ~n2133 ) ;
  assign n2135 = n1632 & ~n2134 ;
  assign n2136 = ( n1630 & n2134 ) | ( n1630 & ~n2135 ) | ( n2134 & ~n2135 ) ;
  assign n2137 = n979 ^ x75 ^ 1'b0 ;
  assign n2138 = ( x75 & x203 ) | ( x75 & ~n2137 ) | ( x203 & ~n2137 ) ;
  assign n2139 = n1452 ^ x330 ^ 1'b0 ;
  assign n2140 = ( x330 & x458 ) | ( x330 & ~n2139 ) | ( x458 & ~n2139 ) ;
  assign n2141 = n979 ^ x74 ^ 1'b0 ;
  assign n2142 = ( x74 & x202 ) | ( x74 & ~n2141 ) | ( x202 & ~n2141 ) ;
  assign n2143 = n2140 & ~n2142 ;
  assign n2144 = n1452 ^ x331 ^ 1'b0 ;
  assign n2145 = ( x331 & x459 ) | ( x331 & ~n2144 ) | ( x459 & ~n2144 ) ;
  assign n2146 = ~n2138 & n2145 ;
  assign n2147 = n2143 | n2146 ;
  assign n2148 = n979 ^ x73 ^ 1'b0 ;
  assign n2149 = ( x73 & x201 ) | ( x73 & ~n2148 ) | ( x201 & ~n2148 ) ;
  assign n2150 = n1452 ^ x329 ^ 1'b0 ;
  assign n2151 = ( x329 & x457 ) | ( x329 & ~n2150 ) | ( x457 & ~n2150 ) ;
  assign n2152 = n1452 ^ x328 ^ 1'b0 ;
  assign n2153 = ( x328 & x456 ) | ( x328 & ~n2152 ) | ( x456 & ~n2152 ) ;
  assign n2154 = n979 ^ x72 ^ 1'b0 ;
  assign n2155 = ( x72 & x200 ) | ( x72 & ~n2154 ) | ( x200 & ~n2154 ) ;
  assign n2156 = ~n2153 & n2155 ;
  assign n2157 = ( n2149 & ~n2151 ) | ( n2149 & n2156 ) | ( ~n2151 & n2156 ) ;
  assign n2158 = ~n2140 & n2142 ;
  assign n2159 = ( ~n2147 & n2157 ) | ( ~n2147 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = ~n2147 & n2159 ;
  assign n2161 = n2145 & ~n2160 ;
  assign n2162 = ( n2138 & n2160 ) | ( n2138 & ~n2161 ) | ( n2160 & ~n2161 ) ;
  assign n2163 = ~n2149 & n2151 ;
  assign n2164 = n2153 & ~n2155 ;
  assign n2165 = n2163 | n2164 ;
  assign n2166 = n2147 | n2165 ;
  assign n2167 = ~n2162 & n2166 ;
  assign n2168 = ( n2136 & n2162 ) | ( n2136 & ~n2167 ) | ( n2162 & ~n2167 ) ;
  assign n2169 = n979 ^ x77 ^ 1'b0 ;
  assign n2170 = ( x77 & x205 ) | ( x77 & ~n2169 ) | ( x205 & ~n2169 ) ;
  assign n2171 = n1452 ^ x333 ^ 1'b0 ;
  assign n2172 = ( x333 & x461 ) | ( x333 & ~n2171 ) | ( x461 & ~n2171 ) ;
  assign n2173 = ~n2170 & n2172 ;
  assign n2174 = n979 ^ x76 ^ 1'b0 ;
  assign n2175 = ( x76 & x204 ) | ( x76 & ~n2174 ) | ( x204 & ~n2174 ) ;
  assign n2176 = n1452 ^ x332 ^ 1'b0 ;
  assign n2177 = ( x332 & x460 ) | ( x332 & ~n2176 ) | ( x460 & ~n2176 ) ;
  assign n2178 = ~n2175 & n2177 ;
  assign n2179 = n2173 | n2178 ;
  assign n2180 = ( n1628 & n2168 ) | ( n1628 & ~n2179 ) | ( n2168 & ~n2179 ) ;
  assign n2181 = ~n1628 & n2180 ;
  assign n2182 = ~n1624 & n1626 ;
  assign n2183 = ( ~n1622 & n2181 ) | ( ~n1622 & n2182 ) | ( n2181 & n2182 ) ;
  assign n2184 = n2181 ^ n1622 ^ 1'b0 ;
  assign n2185 = ( n2181 & n2183 ) | ( n2181 & ~n2184 ) | ( n2183 & ~n2184 ) ;
  assign n2186 = n2175 & ~n2177 ;
  assign n2187 = ( n2170 & ~n2172 ) | ( n2170 & n2186 ) | ( ~n2172 & n2186 ) ;
  assign n2188 = ( ~n1628 & n2185 ) | ( ~n1628 & n2187 ) | ( n2185 & n2187 ) ;
  assign n2189 = n2185 ^ n1628 ^ 1'b0 ;
  assign n2190 = ( n2185 & n2188 ) | ( n2185 & ~n2189 ) | ( n2188 & ~n2189 ) ;
  assign n2191 = ( ~n1616 & n1621 ) | ( ~n1616 & n2190 ) | ( n1621 & n2190 ) ;
  assign n2192 = ~n1616 & n2191 ;
  assign n2193 = ( n1600 & ~n1611 ) | ( n1600 & n2192 ) | ( ~n1611 & n2192 ) ;
  assign n2194 = ~n1600 & n2193 ;
  assign n2195 = n1597 | n1616 ;
  assign n2196 = n1599 & ~n2195 ;
  assign n2197 = n1615 & ~n2196 ;
  assign n2198 = ( n1613 & n2196 ) | ( n1613 & ~n2197 ) | ( n2196 & ~n2197 ) ;
  assign n2199 = ( ~n1602 & n1604 ) | ( ~n1602 & n2198 ) | ( n1604 & n2198 ) ;
  assign n2200 = n2198 ^ n1602 ^ 1'b0 ;
  assign n2201 = ( n2198 & n2199 ) | ( n2198 & ~n2200 ) | ( n2199 & ~n2200 ) ;
  assign n2202 = ( n1605 & ~n1610 ) | ( n1605 & n2201 ) | ( ~n1610 & n2201 ) ;
  assign n2203 = ~n1605 & n2202 ;
  assign n2204 = n1607 & ~n1609 ;
  assign n2205 = ( ~n2194 & n2203 ) | ( ~n2194 & n2204 ) | ( n2203 & n2204 ) ;
  assign n2206 = n2194 | n2205 ;
  assign n2207 = n979 ^ x85 ^ 1'b0 ;
  assign n2208 = ( x85 & x213 ) | ( x85 & ~n2207 ) | ( x213 & ~n2207 ) ;
  assign n2209 = n1452 ^ x341 ^ 1'b0 ;
  assign n2210 = ( x341 & x469 ) | ( x341 & ~n2209 ) | ( x469 & ~n2209 ) ;
  assign n2211 = ~n2208 & n2210 ;
  assign n2212 = n979 ^ x84 ^ 1'b0 ;
  assign n2213 = ( x84 & x212 ) | ( x84 & ~n2212 ) | ( x212 & ~n2212 ) ;
  assign n2214 = n1452 ^ x340 ^ 1'b0 ;
  assign n2215 = ( x340 & x468 ) | ( x340 & ~n2214 ) | ( x468 & ~n2214 ) ;
  assign n2216 = ~n2213 & n2215 ;
  assign n2217 = n2211 | n2216 ;
  assign n2218 = ( n1595 & n2206 ) | ( n1595 & ~n2217 ) | ( n2206 & ~n2217 ) ;
  assign n2219 = ~n1595 & n2218 ;
  assign n2220 = ~n1591 & n1593 ;
  assign n2221 = ( ~n1589 & n2219 ) | ( ~n1589 & n2220 ) | ( n2219 & n2220 ) ;
  assign n2222 = n2219 ^ n1589 ^ 1'b0 ;
  assign n2223 = ( n2219 & n2221 ) | ( n2219 & ~n2222 ) | ( n2221 & ~n2222 ) ;
  assign n2224 = n2213 & ~n2215 ;
  assign n2225 = ( n2208 & ~n2210 ) | ( n2208 & n2224 ) | ( ~n2210 & n2224 ) ;
  assign n2226 = ( ~n1595 & n2223 ) | ( ~n1595 & n2225 ) | ( n2223 & n2225 ) ;
  assign n2227 = n2223 ^ n1595 ^ 1'b0 ;
  assign n2228 = ( n2223 & n2226 ) | ( n2223 & ~n2227 ) | ( n2226 & ~n2227 ) ;
  assign n2229 = n1588 & ~n2228 ;
  assign n2230 = ( n1586 & n2228 ) | ( n1586 & ~n2229 ) | ( n2228 & ~n2229 ) ;
  assign n2231 = n979 ^ x91 ^ 1'b0 ;
  assign n2232 = ( x91 & x219 ) | ( x91 & ~n2231 ) | ( x219 & ~n2231 ) ;
  assign n2233 = n1452 ^ x346 ^ 1'b0 ;
  assign n2234 = ( x346 & x474 ) | ( x346 & ~n2233 ) | ( x474 & ~n2233 ) ;
  assign n2235 = n979 ^ x90 ^ 1'b0 ;
  assign n2236 = ( x90 & x218 ) | ( x90 & ~n2235 ) | ( x218 & ~n2235 ) ;
  assign n2237 = n2234 & ~n2236 ;
  assign n2238 = n1452 ^ x347 ^ 1'b0 ;
  assign n2239 = ( x347 & x475 ) | ( x347 & ~n2238 ) | ( x475 & ~n2238 ) ;
  assign n2240 = ~n2232 & n2239 ;
  assign n2241 = n2237 | n2240 ;
  assign n2242 = n979 ^ x89 ^ 1'b0 ;
  assign n2243 = ( x89 & x217 ) | ( x89 & ~n2242 ) | ( x217 & ~n2242 ) ;
  assign n2244 = n1452 ^ x345 ^ 1'b0 ;
  assign n2245 = ( x345 & x473 ) | ( x345 & ~n2244 ) | ( x473 & ~n2244 ) ;
  assign n2246 = n1452 ^ x344 ^ 1'b0 ;
  assign n2247 = ( x344 & x472 ) | ( x344 & ~n2246 ) | ( x472 & ~n2246 ) ;
  assign n2248 = n979 ^ x88 ^ 1'b0 ;
  assign n2249 = ( x88 & x216 ) | ( x88 & ~n2248 ) | ( x216 & ~n2248 ) ;
  assign n2250 = ~n2247 & n2249 ;
  assign n2251 = ( n2243 & ~n2245 ) | ( n2243 & n2250 ) | ( ~n2245 & n2250 ) ;
  assign n2252 = ~n2234 & n2236 ;
  assign n2253 = ( ~n2241 & n2251 ) | ( ~n2241 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2254 = ~n2241 & n2253 ;
  assign n2255 = n2239 & ~n2254 ;
  assign n2256 = ( n2232 & n2254 ) | ( n2232 & ~n2255 ) | ( n2254 & ~n2255 ) ;
  assign n2257 = ~n2243 & n2245 ;
  assign n2258 = n2247 & ~n2249 ;
  assign n2259 = n2257 | n2258 ;
  assign n2260 = n2241 | n2259 ;
  assign n2261 = ~n2256 & n2260 ;
  assign n2262 = ( n2230 & n2256 ) | ( n2230 & ~n2261 ) | ( n2256 & ~n2261 ) ;
  assign n2263 = n979 ^ x93 ^ 1'b0 ;
  assign n2264 = ( x93 & x221 ) | ( x93 & ~n2263 ) | ( x221 & ~n2263 ) ;
  assign n2265 = n1452 ^ x349 ^ 1'b0 ;
  assign n2266 = ( x349 & x477 ) | ( x349 & ~n2265 ) | ( x477 & ~n2265 ) ;
  assign n2267 = ~n2264 & n2266 ;
  assign n2268 = n979 ^ x92 ^ 1'b0 ;
  assign n2269 = ( x92 & x220 ) | ( x92 & ~n2268 ) | ( x220 & ~n2268 ) ;
  assign n2270 = n1452 ^ x348 ^ 1'b0 ;
  assign n2271 = ( x348 & x476 ) | ( x348 & ~n2270 ) | ( x476 & ~n2270 ) ;
  assign n2272 = ~n2269 & n2271 ;
  assign n2273 = n2267 | n2272 ;
  assign n2274 = ( n1584 & n2262 ) | ( n1584 & ~n2273 ) | ( n2262 & ~n2273 ) ;
  assign n2275 = ~n1584 & n2274 ;
  assign n2276 = ~n1580 & n1582 ;
  assign n2277 = ( ~n1578 & n2275 ) | ( ~n1578 & n2276 ) | ( n2275 & n2276 ) ;
  assign n2278 = n2275 ^ n1578 ^ 1'b0 ;
  assign n2279 = ( n2275 & n2277 ) | ( n2275 & ~n2278 ) | ( n2277 & ~n2278 ) ;
  assign n2280 = n2269 & ~n2271 ;
  assign n2281 = ( n2264 & ~n2266 ) | ( n2264 & n2280 ) | ( ~n2266 & n2280 ) ;
  assign n2282 = ( ~n1584 & n2279 ) | ( ~n1584 & n2281 ) | ( n2279 & n2281 ) ;
  assign n2283 = n2279 ^ n1584 ^ 1'b0 ;
  assign n2284 = ( n2279 & n2282 ) | ( n2279 & ~n2283 ) | ( n2282 & ~n2283 ) ;
  assign n2285 = ( ~n1572 & n1577 ) | ( ~n1572 & n2284 ) | ( n1577 & n2284 ) ;
  assign n2286 = ~n1572 & n2285 ;
  assign n2287 = ( n1556 & ~n1567 ) | ( n1556 & n2286 ) | ( ~n1567 & n2286 ) ;
  assign n2288 = ~n1556 & n2287 ;
  assign n2289 = n1553 | n1572 ;
  assign n2290 = n1555 & ~n2289 ;
  assign n2291 = n1571 & ~n2290 ;
  assign n2292 = ( n1569 & n2290 ) | ( n1569 & ~n2291 ) | ( n2290 & ~n2291 ) ;
  assign n2293 = ( ~n1558 & n1560 ) | ( ~n1558 & n2292 ) | ( n1560 & n2292 ) ;
  assign n2294 = n2292 ^ n1558 ^ 1'b0 ;
  assign n2295 = ( n2292 & n2293 ) | ( n2292 & ~n2294 ) | ( n2293 & ~n2294 ) ;
  assign n2296 = ( n1561 & ~n1566 ) | ( n1561 & n2295 ) | ( ~n1566 & n2295 ) ;
  assign n2297 = ~n1561 & n2296 ;
  assign n2298 = n1563 & ~n1565 ;
  assign n2299 = ( ~n2288 & n2297 ) | ( ~n2288 & n2298 ) | ( n2297 & n2298 ) ;
  assign n2300 = n2288 | n2299 ;
  assign n2301 = n979 ^ x101 ^ 1'b0 ;
  assign n2302 = ( x101 & x229 ) | ( x101 & ~n2301 ) | ( x229 & ~n2301 ) ;
  assign n2303 = n1452 ^ x357 ^ 1'b0 ;
  assign n2304 = ( x357 & x485 ) | ( x357 & ~n2303 ) | ( x485 & ~n2303 ) ;
  assign n2305 = ~n2302 & n2304 ;
  assign n2306 = n979 ^ x100 ^ 1'b0 ;
  assign n2307 = ( x100 & x228 ) | ( x100 & ~n2306 ) | ( x228 & ~n2306 ) ;
  assign n2308 = n1452 ^ x356 ^ 1'b0 ;
  assign n2309 = ( x356 & x484 ) | ( x356 & ~n2308 ) | ( x484 & ~n2308 ) ;
  assign n2310 = ~n2307 & n2309 ;
  assign n2311 = n2305 | n2310 ;
  assign n2312 = ( n1551 & n2300 ) | ( n1551 & ~n2311 ) | ( n2300 & ~n2311 ) ;
  assign n2313 = ~n1551 & n2312 ;
  assign n2314 = ~n1547 & n1549 ;
  assign n2315 = ( ~n1545 & n2313 ) | ( ~n1545 & n2314 ) | ( n2313 & n2314 ) ;
  assign n2316 = n2313 ^ n1545 ^ 1'b0 ;
  assign n2317 = ( n2313 & n2315 ) | ( n2313 & ~n2316 ) | ( n2315 & ~n2316 ) ;
  assign n2318 = n2307 & ~n2309 ;
  assign n2319 = ( n2302 & ~n2304 ) | ( n2302 & n2318 ) | ( ~n2304 & n2318 ) ;
  assign n2320 = ( ~n1551 & n2317 ) | ( ~n1551 & n2319 ) | ( n2317 & n2319 ) ;
  assign n2321 = n2317 ^ n1551 ^ 1'b0 ;
  assign n2322 = ( n2317 & n2320 ) | ( n2317 & ~n2321 ) | ( n2320 & ~n2321 ) ;
  assign n2323 = n1544 & ~n2322 ;
  assign n2324 = ( n1542 & n2322 ) | ( n1542 & ~n2323 ) | ( n2322 & ~n2323 ) ;
  assign n2325 = n979 ^ x107 ^ 1'b0 ;
  assign n2326 = ( x107 & x235 ) | ( x107 & ~n2325 ) | ( x235 & ~n2325 ) ;
  assign n2327 = n1452 ^ x362 ^ 1'b0 ;
  assign n2328 = ( x362 & x490 ) | ( x362 & ~n2327 ) | ( x490 & ~n2327 ) ;
  assign n2329 = n979 ^ x106 ^ 1'b0 ;
  assign n2330 = ( x106 & x234 ) | ( x106 & ~n2329 ) | ( x234 & ~n2329 ) ;
  assign n2331 = n2328 & ~n2330 ;
  assign n2332 = n1452 ^ x363 ^ 1'b0 ;
  assign n2333 = ( x363 & x491 ) | ( x363 & ~n2332 ) | ( x491 & ~n2332 ) ;
  assign n2334 = ~n2326 & n2333 ;
  assign n2335 = n2331 | n2334 ;
  assign n2336 = n979 ^ x105 ^ 1'b0 ;
  assign n2337 = ( x105 & x233 ) | ( x105 & ~n2336 ) | ( x233 & ~n2336 ) ;
  assign n2338 = n1452 ^ x361 ^ 1'b0 ;
  assign n2339 = ( x361 & x489 ) | ( x361 & ~n2338 ) | ( x489 & ~n2338 ) ;
  assign n2340 = n1452 ^ x360 ^ 1'b0 ;
  assign n2341 = ( x360 & x488 ) | ( x360 & ~n2340 ) | ( x488 & ~n2340 ) ;
  assign n2342 = n979 ^ x104 ^ 1'b0 ;
  assign n2343 = ( x104 & x232 ) | ( x104 & ~n2342 ) | ( x232 & ~n2342 ) ;
  assign n2344 = ~n2341 & n2343 ;
  assign n2345 = ( n2337 & ~n2339 ) | ( n2337 & n2344 ) | ( ~n2339 & n2344 ) ;
  assign n2346 = ~n2328 & n2330 ;
  assign n2347 = ( ~n2335 & n2345 ) | ( ~n2335 & n2346 ) | ( n2345 & n2346 ) ;
  assign n2348 = ~n2335 & n2347 ;
  assign n2349 = n2333 & ~n2348 ;
  assign n2350 = ( n2326 & n2348 ) | ( n2326 & ~n2349 ) | ( n2348 & ~n2349 ) ;
  assign n2351 = ~n2337 & n2339 ;
  assign n2352 = n2341 & ~n2343 ;
  assign n2353 = n2351 | n2352 ;
  assign n2354 = n2335 | n2353 ;
  assign n2355 = ~n2350 & n2354 ;
  assign n2356 = ( n2324 & n2350 ) | ( n2324 & ~n2355 ) | ( n2350 & ~n2355 ) ;
  assign n2357 = n979 ^ x109 ^ 1'b0 ;
  assign n2358 = ( x109 & x237 ) | ( x109 & ~n2357 ) | ( x237 & ~n2357 ) ;
  assign n2359 = n1452 ^ x365 ^ 1'b0 ;
  assign n2360 = ( x365 & x493 ) | ( x365 & ~n2359 ) | ( x493 & ~n2359 ) ;
  assign n2361 = ~n2358 & n2360 ;
  assign n2362 = n979 ^ x108 ^ 1'b0 ;
  assign n2363 = ( x108 & x236 ) | ( x108 & ~n2362 ) | ( x236 & ~n2362 ) ;
  assign n2364 = n1452 ^ x364 ^ 1'b0 ;
  assign n2365 = ( x364 & x492 ) | ( x364 & ~n2364 ) | ( x492 & ~n2364 ) ;
  assign n2366 = ~n2363 & n2365 ;
  assign n2367 = n2361 | n2366 ;
  assign n2368 = ( n1540 & n2356 ) | ( n1540 & ~n2367 ) | ( n2356 & ~n2367 ) ;
  assign n2369 = ~n1540 & n2368 ;
  assign n2370 = ~n1536 & n1538 ;
  assign n2371 = ( ~n1534 & n2369 ) | ( ~n1534 & n2370 ) | ( n2369 & n2370 ) ;
  assign n2372 = n2369 ^ n1534 ^ 1'b0 ;
  assign n2373 = ( n2369 & n2371 ) | ( n2369 & ~n2372 ) | ( n2371 & ~n2372 ) ;
  assign n2374 = n2363 & ~n2365 ;
  assign n2375 = ( n2358 & ~n2360 ) | ( n2358 & n2374 ) | ( ~n2360 & n2374 ) ;
  assign n2376 = ( ~n1540 & n2373 ) | ( ~n1540 & n2375 ) | ( n2373 & n2375 ) ;
  assign n2377 = n2373 ^ n1540 ^ 1'b0 ;
  assign n2378 = ( n2373 & n2376 ) | ( n2373 & ~n2377 ) | ( n2376 & ~n2377 ) ;
  assign n2379 = ( ~n1528 & n1533 ) | ( ~n1528 & n2378 ) | ( n1533 & n2378 ) ;
  assign n2380 = ~n1528 & n2379 ;
  assign n2381 = ( n1512 & ~n1523 ) | ( n1512 & n2380 ) | ( ~n1523 & n2380 ) ;
  assign n2382 = ~n1512 & n2381 ;
  assign n2383 = n1525 & ~n1527 ;
  assign n2384 = n1509 | n1528 ;
  assign n2385 = ~n2383 & n2384 ;
  assign n2386 = ( n1511 & n2383 ) | ( n1511 & ~n2385 ) | ( n2383 & ~n2385 ) ;
  assign n2387 = ( ~n1514 & n1516 ) | ( ~n1514 & n2386 ) | ( n1516 & n2386 ) ;
  assign n2388 = n2386 ^ n1514 ^ 1'b0 ;
  assign n2389 = ( n2386 & n2387 ) | ( n2386 & ~n2388 ) | ( n2387 & ~n2388 ) ;
  assign n2390 = ( n1517 & ~n1522 ) | ( n1517 & n2389 ) | ( ~n1522 & n2389 ) ;
  assign n2391 = ~n1517 & n2390 ;
  assign n2392 = n1519 & ~n1521 ;
  assign n2393 = ( ~n2382 & n2391 ) | ( ~n2382 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2394 = n2382 | n2393 ;
  assign n2395 = ~n1500 & n1503 ;
  assign n2396 = n1501 | n2395 ;
  assign n2397 = ( n1493 & n2394 ) | ( n1493 & ~n2396 ) | ( n2394 & ~n2396 ) ;
  assign n2398 = ~n1493 & n2397 ;
  assign n2399 = ~n1489 & n1491 ;
  assign n2400 = ~n1487 & n2399 ;
  assign n2401 = ( ~n1507 & n2398 ) | ( ~n1507 & n2400 ) | ( n2398 & n2400 ) ;
  assign n2402 = n1507 | n2401 ;
  assign n2403 = n1486 & ~n2402 ;
  assign n2404 = ( n1484 & n2402 ) | ( n1484 & ~n2403 ) | ( n2402 & ~n2403 ) ;
  assign n2405 = ( n1471 & ~n1482 ) | ( n1471 & n2404 ) | ( ~n1482 & n2404 ) ;
  assign n2406 = ~n1471 & n2405 ;
  assign n2407 = n1473 & ~n1475 ;
  assign n2408 = n1476 | n1478 ;
  assign n2409 = ~n2407 & n2408 ;
  assign n2410 = ( n1480 & n2407 ) | ( n1480 & ~n2409 ) | ( n2407 & ~n2409 ) ;
  assign n2411 = ~n1466 & n1468 ;
  assign n2412 = ( ~n1471 & n2410 ) | ( ~n1471 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = ~n1471 & n2412 ;
  assign n2414 = ( ~n1464 & n2406 ) | ( ~n1464 & n2413 ) | ( n2406 & n2413 ) ;
  assign n2415 = n1464 | n2414 ;
  assign n2416 = ~n1456 & n1458 ;
  assign n2417 = n979 ^ x126 ^ 1'b0 ;
  assign n2418 = ( x126 & x254 ) | ( x126 & ~n2417 ) | ( x254 & ~n2417 ) ;
  assign n2419 = n1452 ^ x382 ^ 1'b0 ;
  assign n2420 = ( x382 & x510 ) | ( x382 & ~n2419 ) | ( x510 & ~n2419 ) ;
  assign n2421 = n2418 & ~n2420 ;
  assign n2422 = ~n2418 & n2420 ;
  assign n2423 = n979 ^ x125 ^ 1'b0 ;
  assign n2424 = ( x125 & x253 ) | ( x125 & ~n2423 ) | ( x253 & ~n2423 ) ;
  assign n2425 = n1452 ^ x381 ^ 1'b0 ;
  assign n2426 = ( x381 & x509 ) | ( x381 & ~n2425 ) | ( x509 & ~n2425 ) ;
  assign n2427 = ~n2424 & n2426 ;
  assign n2428 = n2422 | n2427 ;
  assign n2429 = n2424 & ~n2426 ;
  assign n2430 = n979 ^ x124 ^ 1'b0 ;
  assign n2431 = ( x124 & x252 ) | ( x124 & ~n2430 ) | ( x252 & ~n2430 ) ;
  assign n2432 = n1452 ^ x380 ^ 1'b0 ;
  assign n2433 = ( x380 & x508 ) | ( x380 & ~n2432 ) | ( x508 & ~n2432 ) ;
  assign n2434 = n2431 & ~n2433 ;
  assign n2435 = ( ~n2428 & n2429 ) | ( ~n2428 & n2434 ) | ( n2429 & n2434 ) ;
  assign n2436 = ~n2428 & n2435 ;
  assign n2437 = ( ~n2416 & n2421 ) | ( ~n2416 & n2436 ) | ( n2421 & n2436 ) ;
  assign n2438 = ~n2416 & n2437 ;
  assign n2439 = n2416 | n2428 ;
  assign n2440 = ~n2431 & n2433 ;
  assign n2441 = n2439 | n2440 ;
  assign n2442 = ~n2438 & n2441 ;
  assign n2443 = ( n2415 & n2438 ) | ( n2415 & ~n2442 ) | ( n2438 & ~n2442 ) ;
  assign n2444 = n1459 | n2443 ;
  assign n2445 = n2444 ^ n981 ^ 1'b0 ;
  assign n2446 = ( n981 & n1454 ) | ( n981 & ~n2445 ) | ( n1454 & ~n2445 ) ;
  assign n2447 = n2444 ^ n1876 ^ 1'b0 ;
  assign n2448 = ( n1876 & n1878 ) | ( n1876 & ~n2447 ) | ( n1878 & ~n2447 ) ;
  assign n2449 = n2444 ^ n1871 ^ 1'b0 ;
  assign n2450 = ( n1871 & n1873 ) | ( n1871 & ~n2449 ) | ( n1873 & ~n2449 ) ;
  assign n2451 = n2444 ^ n1867 ^ 1'b0 ;
  assign n2452 = ( n1867 & n1869 ) | ( n1867 & ~n2451 ) | ( n1869 & ~n2451 ) ;
  assign n2453 = n2444 ^ n1865 ^ 1'b0 ;
  assign n2454 = ( n1863 & n1865 ) | ( n1863 & ~n2453 ) | ( n1865 & ~n2453 ) ;
  assign n2455 = n2444 ^ n1861 ^ 1'b0 ;
  assign n2456 = ( n1859 & n1861 ) | ( n1859 & ~n2455 ) | ( n1861 & ~n2455 ) ;
  assign n2457 = n2444 ^ n1857 ^ 1'b0 ;
  assign n2458 = ( n1855 & n1857 ) | ( n1855 & ~n2457 ) | ( n1857 & ~n2457 ) ;
  assign n2459 = n2444 ^ n1851 ^ 1'b0 ;
  assign n2460 = ( n1851 & n1853 ) | ( n1851 & ~n2459 ) | ( n1853 & ~n2459 ) ;
  assign n2461 = n2444 ^ n1893 ^ 1'b0 ;
  assign n2462 = ( n1849 & n1893 ) | ( n1849 & ~n2461 ) | ( n1893 & ~n2461 ) ;
  assign n2463 = n2444 ^ n1896 ^ 1'b0 ;
  assign n2464 = ( n1847 & n1896 ) | ( n1847 & ~n2463 ) | ( n1896 & ~n2463 ) ;
  assign n2465 = n2444 ^ n1843 ^ 1'b0 ;
  assign n2466 = ( n1843 & n1845 ) | ( n1843 & ~n2465 ) | ( n1845 & ~n2465 ) ;
  assign n2467 = n2444 ^ n1839 ^ 1'b0 ;
  assign n2468 = ( n1839 & n1841 ) | ( n1839 & ~n2467 ) | ( n1841 & ~n2467 ) ;
  assign n2469 = n2444 ^ n1835 ^ 1'b0 ;
  assign n2470 = ( n1835 & n1837 ) | ( n1835 & ~n2469 ) | ( n1837 & ~n2469 ) ;
  assign n2471 = n2444 ^ n1831 ^ 1'b0 ;
  assign n2472 = ( n1831 & n1833 ) | ( n1831 & ~n2471 ) | ( n1833 & ~n2471 ) ;
  assign n2473 = n2444 ^ n1827 ^ 1'b0 ;
  assign n2474 = ( n1827 & n1829 ) | ( n1827 & ~n2473 ) | ( n1829 & ~n2473 ) ;
  assign n2475 = n2444 ^ n1823 ^ 1'b0 ;
  assign n2476 = ( n1823 & n1825 ) | ( n1823 & ~n2475 ) | ( n1825 & ~n2475 ) ;
  assign n2477 = n2444 ^ n1905 ^ 1'b0 ;
  assign n2478 = ( n1821 & n1905 ) | ( n1821 & ~n2477 ) | ( n1905 & ~n2477 ) ;
  assign n2479 = n2444 ^ n1908 ^ 1'b0 ;
  assign n2480 = ( n1819 & n1908 ) | ( n1819 & ~n2479 ) | ( n1908 & ~n2479 ) ;
  assign n2481 = n2444 ^ n1815 ^ 1'b0 ;
  assign n2482 = ( n1815 & n1817 ) | ( n1815 & ~n2481 ) | ( n1817 & ~n2481 ) ;
  assign n2483 = n2444 ^ n1811 ^ 1'b0 ;
  assign n2484 = ( n1811 & n1813 ) | ( n1811 & ~n2483 ) | ( n1813 & ~n2483 ) ;
  assign n2485 = n2444 ^ n1807 ^ 1'b0 ;
  assign n2486 = ( n1807 & n1809 ) | ( n1807 & ~n2485 ) | ( n1809 & ~n2485 ) ;
  assign n2487 = n2444 ^ n1803 ^ 1'b0 ;
  assign n2488 = ( n1803 & n1805 ) | ( n1803 & ~n2487 ) | ( n1805 & ~n2487 ) ;
  assign n2489 = n2444 ^ n1799 ^ 1'b0 ;
  assign n2490 = ( n1799 & n1801 ) | ( n1799 & ~n2489 ) | ( n1801 & ~n2489 ) ;
  assign n2491 = n2444 ^ n1795 ^ 1'b0 ;
  assign n2492 = ( n1795 & n1797 ) | ( n1795 & ~n2491 ) | ( n1797 & ~n2491 ) ;
  assign n2493 = n2444 ^ n1917 ^ 1'b0 ;
  assign n2494 = ( n1793 & n1917 ) | ( n1793 & ~n2493 ) | ( n1917 & ~n2493 ) ;
  assign n2495 = n2444 ^ n1920 ^ 1'b0 ;
  assign n2496 = ( n1791 & n1920 ) | ( n1791 & ~n2495 ) | ( n1920 & ~n2495 ) ;
  assign n2497 = n2444 ^ n1787 ^ 1'b0 ;
  assign n2498 = ( n1787 & n1789 ) | ( n1787 & ~n2497 ) | ( n1789 & ~n2497 ) ;
  assign n2499 = n2444 ^ n1783 ^ 1'b0 ;
  assign n2500 = ( n1783 & n1785 ) | ( n1783 & ~n2499 ) | ( n1785 & ~n2499 ) ;
  assign n2501 = n2444 ^ n1779 ^ 1'b0 ;
  assign n2502 = ( n1779 & n1781 ) | ( n1779 & ~n2501 ) | ( n1781 & ~n2501 ) ;
  assign n2503 = n2444 ^ n1775 ^ 1'b0 ;
  assign n2504 = ( n1775 & n1777 ) | ( n1775 & ~n2503 ) | ( n1777 & ~n2503 ) ;
  assign n2505 = n2444 ^ n1771 ^ 1'b0 ;
  assign n2506 = ( n1771 & n1773 ) | ( n1771 & ~n2505 ) | ( n1773 & ~n2505 ) ;
  assign n2507 = n2444 ^ n1767 ^ 1'b0 ;
  assign n2508 = ( n1767 & n1769 ) | ( n1767 & ~n2507 ) | ( n1769 & ~n2507 ) ;
  assign n2509 = n2444 ^ n1764 ^ 1'b0 ;
  assign n2510 = ( n1762 & n1764 ) | ( n1762 & ~n2509 ) | ( n1764 & ~n2509 ) ;
  assign n2511 = n2444 ^ n1952 ^ 1'b0 ;
  assign n2512 = ( n1952 & n1954 ) | ( n1952 & ~n2511 ) | ( n1954 & ~n2511 ) ;
  assign n2513 = n2444 ^ n1964 ^ 1'b0 ;
  assign n2514 = ( n1962 & n1964 ) | ( n1962 & ~n2513 ) | ( n1964 & ~n2513 ) ;
  assign n2515 = n2444 ^ n1957 ^ 1'b0 ;
  assign n2516 = ( n1957 & n1959 ) | ( n1957 & ~n2515 ) | ( n1959 & ~n2515 ) ;
  assign n2517 = n2444 ^ n1940 ^ 1'b0 ;
  assign n2518 = ( n1940 & n1942 ) | ( n1940 & ~n2517 ) | ( n1942 & ~n2517 ) ;
  assign n2519 = n2444 ^ n1945 ^ 1'b0 ;
  assign n2520 = ( n1945 & n1947 ) | ( n1945 & ~n2519 ) | ( n1947 & ~n2519 ) ;
  assign n2521 = n2444 ^ n1936 ^ 1'b0 ;
  assign n2522 = ( n1934 & n1936 ) | ( n1934 & ~n2521 ) | ( n1936 & ~n2521 ) ;
  assign n2523 = n2444 ^ n1929 ^ 1'b0 ;
  assign n2524 = ( n1929 & n1931 ) | ( n1929 & ~n2523 ) | ( n1931 & ~n2523 ) ;
  assign n2525 = n2444 ^ n1749 ^ 1'b0 ;
  assign n2526 = ( n1749 & n1751 ) | ( n1749 & ~n2525 ) | ( n1751 & ~n2525 ) ;
  assign n2527 = n2444 ^ n1745 ^ 1'b0 ;
  assign n2528 = ( n1745 & n1747 ) | ( n1745 & ~n2527 ) | ( n1747 & ~n2527 ) ;
  assign n2529 = n2444 ^ n1735 ^ 1'b0 ;
  assign n2530 = ( n1735 & n1737 ) | ( n1735 & ~n2529 ) | ( n1737 & ~n2529 ) ;
  assign n2531 = n2444 ^ n1740 ^ 1'b0 ;
  assign n2532 = ( n1740 & n1742 ) | ( n1740 & ~n2531 ) | ( n1742 & ~n2531 ) ;
  assign n2533 = n2444 ^ n1723 ^ 1'b0 ;
  assign n2534 = ( n1723 & n1725 ) | ( n1723 & ~n2533 ) | ( n1725 & ~n2533 ) ;
  assign n2535 = n2444 ^ n1728 ^ 1'b0 ;
  assign n2536 = ( n1728 & n1730 ) | ( n1728 & ~n2535 ) | ( n1730 & ~n2535 ) ;
  assign n2537 = n2444 ^ n1719 ^ 1'b0 ;
  assign n2538 = ( n1717 & n1719 ) | ( n1717 & ~n2537 ) | ( n1719 & ~n2537 ) ;
  assign n2539 = n2444 ^ n1712 ^ 1'b0 ;
  assign n2540 = ( n1712 & n1714 ) | ( n1712 & ~n2539 ) | ( n1714 & ~n2539 ) ;
  assign n2541 = n2444 ^ n2060 ^ 1'b0 ;
  assign n2542 = ( n2058 & n2060 ) | ( n2058 & ~n2541 ) | ( n2060 & ~n2541 ) ;
  assign n2543 = n2444 ^ n2044 ^ 1'b0 ;
  assign n2544 = ( n2044 & n2046 ) | ( n2044 & ~n2543 ) | ( n2046 & ~n2543 ) ;
  assign n2545 = n2444 ^ n2042 ^ 1'b0 ;
  assign n2546 = ( n2042 & n2052 ) | ( n2042 & ~n2545 ) | ( n2052 & ~n2545 ) ;
  assign n2547 = n2444 ^ n2040 ^ 1'b0 ;
  assign n2548 = ( n2040 & n2049 ) | ( n2040 & ~n2547 ) | ( n2049 & ~n2547 ) ;
  assign n2549 = n2444 ^ n2029 ^ 1'b0 ;
  assign n2550 = ( n2027 & n2029 ) | ( n2027 & ~n2549 ) | ( n2029 & ~n2549 ) ;
  assign n2551 = n2444 ^ n2023 ^ 1'b0 ;
  assign n2552 = ( n2023 & n2025 ) | ( n2023 & ~n2551 ) | ( n2025 & ~n2551 ) ;
  assign n2553 = n2444 ^ n2016 ^ 1'b0 ;
  assign n2554 = ( n2014 & n2016 ) | ( n2014 & ~n2553 ) | ( n2016 & ~n2553 ) ;
  assign n2555 = n2444 ^ n2012 ^ 1'b0 ;
  assign n2556 = ( n2012 & n2019 ) | ( n2012 & ~n2555 ) | ( n2019 & ~n2555 ) ;
  assign n2557 = n2444 ^ n1699 ^ 1'b0 ;
  assign n2558 = ( n1699 & n1701 ) | ( n1699 & ~n2557 ) | ( n1701 & ~n2557 ) ;
  assign n2559 = n2444 ^ n1695 ^ 1'b0 ;
  assign n2560 = ( n1695 & n1697 ) | ( n1695 & ~n2559 ) | ( n1697 & ~n2559 ) ;
  assign n2561 = n2444 ^ n1689 ^ 1'b0 ;
  assign n2562 = ( n1689 & n1691 ) | ( n1689 & ~n2561 ) | ( n1691 & ~n2561 ) ;
  assign n2563 = n2444 ^ n1684 ^ 1'b0 ;
  assign n2564 = ( n1684 & n1686 ) | ( n1684 & ~n2563 ) | ( n1686 & ~n2563 ) ;
  assign n2565 = n2444 ^ n1672 ^ 1'b0 ;
  assign n2566 = ( n1672 & n1674 ) | ( n1672 & ~n2565 ) | ( n1674 & ~n2565 ) ;
  assign n2567 = n2444 ^ n1677 ^ 1'b0 ;
  assign n2568 = ( n1677 & n1679 ) | ( n1677 & ~n2567 ) | ( n1679 & ~n2567 ) ;
  assign n2569 = n2444 ^ n1668 ^ 1'b0 ;
  assign n2570 = ( n1666 & n1668 ) | ( n1666 & ~n2569 ) | ( n1668 & ~n2569 ) ;
  assign n2571 = n2444 ^ n1661 ^ 1'b0 ;
  assign n2572 = ( n1661 & n1663 ) | ( n1661 & ~n2571 ) | ( n1663 & ~n2571 ) ;
  assign n2573 = n2444 ^ n1653 ^ 1'b0 ;
  assign n2574 = ( n1651 & n1653 ) | ( n1651 & ~n2573 ) | ( n1653 & ~n2573 ) ;
  assign n2575 = n2444 ^ n1656 ^ 1'b0 ;
  assign n2576 = ( n1656 & n1658 ) | ( n1656 & ~n2575 ) | ( n1658 & ~n2575 ) ;
  assign n2577 = n2444 ^ n1648 ^ 1'b0 ;
  assign n2578 = ( n1646 & n1648 ) | ( n1646 & ~n2577 ) | ( n1648 & ~n2577 ) ;
  assign n2579 = n2444 ^ n1641 ^ 1'b0 ;
  assign n2580 = ( n1641 & n1643 ) | ( n1641 & ~n2579 ) | ( n1643 & ~n2579 ) ;
  assign n2581 = n2444 ^ n2119 ^ 1'b0 ;
  assign n2582 = ( n2119 & n2121 ) | ( n2119 & ~n2581 ) | ( n2121 & ~n2581 ) ;
  assign n2583 = n2444 ^ n2114 ^ 1'b0 ;
  assign n2584 = ( n2114 & n2116 ) | ( n2114 & ~n2583 ) | ( n2116 & ~n2583 ) ;
  assign n2585 = n2444 ^ n1637 ^ 1'b0 ;
  assign n2586 = ( n1635 & n1637 ) | ( n1635 & ~n2585 ) | ( n1637 & ~n2585 ) ;
  assign n2587 = n2444 ^ n1630 ^ 1'b0 ;
  assign n2588 = ( n1630 & n1632 ) | ( n1630 & ~n2587 ) | ( n1632 & ~n2587 ) ;
  assign n2589 = n2444 ^ n2155 ^ 1'b0 ;
  assign n2590 = ( n2153 & n2155 ) | ( n2153 & ~n2589 ) | ( n2155 & ~n2589 ) ;
  assign n2591 = n2444 ^ n2149 ^ 1'b0 ;
  assign n2592 = ( n2149 & n2151 ) | ( n2149 & ~n2591 ) | ( n2151 & ~n2591 ) ;
  assign n2593 = n2444 ^ n2142 ^ 1'b0 ;
  assign n2594 = ( n2140 & n2142 ) | ( n2140 & ~n2593 ) | ( n2142 & ~n2593 ) ;
  assign n2595 = n2444 ^ n2138 ^ 1'b0 ;
  assign n2596 = ( n2138 & n2145 ) | ( n2138 & ~n2595 ) | ( n2145 & ~n2595 ) ;
  assign n2597 = n2444 ^ n2175 ^ 1'b0 ;
  assign n2598 = ( n2175 & n2177 ) | ( n2175 & ~n2597 ) | ( n2177 & ~n2597 ) ;
  assign n2599 = n2444 ^ n2170 ^ 1'b0 ;
  assign n2600 = ( n2170 & n2172 ) | ( n2170 & ~n2599 ) | ( n2172 & ~n2599 ) ;
  assign n2601 = n2444 ^ n1626 ^ 1'b0 ;
  assign n2602 = ( n1624 & n1626 ) | ( n1624 & ~n2601 ) | ( n1626 & ~n2601 ) ;
  assign n2603 = n2444 ^ n1618 ^ 1'b0 ;
  assign n2604 = ( n1618 & n1620 ) | ( n1618 & ~n2603 ) | ( n1620 & ~n2603 ) ;
  assign n2605 = n2444 ^ n1599 ^ 1'b0 ;
  assign n2606 = ( n1597 & n1599 ) | ( n1597 & ~n2605 ) | ( n1599 & ~n2605 ) ;
  assign n2607 = n2444 ^ n1613 ^ 1'b0 ;
  assign n2608 = ( n1613 & n1615 ) | ( n1613 & ~n2607 ) | ( n1615 & ~n2607 ) ;
  assign n2609 = n2444 ^ n1604 ^ 1'b0 ;
  assign n2610 = ( n1602 & n1604 ) | ( n1602 & ~n2609 ) | ( n1604 & ~n2609 ) ;
  assign n2611 = n2444 ^ n1607 ^ 1'b0 ;
  assign n2612 = ( n1607 & n1609 ) | ( n1607 & ~n2611 ) | ( n1609 & ~n2611 ) ;
  assign n2613 = n2444 ^ n2213 ^ 1'b0 ;
  assign n2614 = ( n2213 & n2215 ) | ( n2213 & ~n2613 ) | ( n2215 & ~n2613 ) ;
  assign n2615 = n2444 ^ n2208 ^ 1'b0 ;
  assign n2616 = ( n2208 & n2210 ) | ( n2208 & ~n2615 ) | ( n2210 & ~n2615 ) ;
  assign n2617 = n2444 ^ n1593 ^ 1'b0 ;
  assign n2618 = ( n1591 & n1593 ) | ( n1591 & ~n2617 ) | ( n1593 & ~n2617 ) ;
  assign n2619 = n2444 ^ n1586 ^ 1'b0 ;
  assign n2620 = ( n1586 & n1588 ) | ( n1586 & ~n2619 ) | ( n1588 & ~n2619 ) ;
  assign n2621 = n2444 ^ n2249 ^ 1'b0 ;
  assign n2622 = ( n2247 & n2249 ) | ( n2247 & ~n2621 ) | ( n2249 & ~n2621 ) ;
  assign n2623 = n2444 ^ n2243 ^ 1'b0 ;
  assign n2624 = ( n2243 & n2245 ) | ( n2243 & ~n2623 ) | ( n2245 & ~n2623 ) ;
  assign n2625 = n2444 ^ n2236 ^ 1'b0 ;
  assign n2626 = ( n2234 & n2236 ) | ( n2234 & ~n2625 ) | ( n2236 & ~n2625 ) ;
  assign n2627 = n2444 ^ n2232 ^ 1'b0 ;
  assign n2628 = ( n2232 & n2239 ) | ( n2232 & ~n2627 ) | ( n2239 & ~n2627 ) ;
  assign n2629 = n2444 ^ n2269 ^ 1'b0 ;
  assign n2630 = ( n2269 & n2271 ) | ( n2269 & ~n2629 ) | ( n2271 & ~n2629 ) ;
  assign n2631 = n2444 ^ n2264 ^ 1'b0 ;
  assign n2632 = ( n2264 & n2266 ) | ( n2264 & ~n2631 ) | ( n2266 & ~n2631 ) ;
  assign n2633 = n2444 ^ n1582 ^ 1'b0 ;
  assign n2634 = ( n1580 & n1582 ) | ( n1580 & ~n2633 ) | ( n1582 & ~n2633 ) ;
  assign n2635 = n2444 ^ n1574 ^ 1'b0 ;
  assign n2636 = ( n1574 & n1576 ) | ( n1574 & ~n2635 ) | ( n1576 & ~n2635 ) ;
  assign n2637 = n2444 ^ n1555 ^ 1'b0 ;
  assign n2638 = ( n1553 & n1555 ) | ( n1553 & ~n2637 ) | ( n1555 & ~n2637 ) ;
  assign n2639 = n2444 ^ n1569 ^ 1'b0 ;
  assign n2640 = ( n1569 & n1571 ) | ( n1569 & ~n2639 ) | ( n1571 & ~n2639 ) ;
  assign n2641 = n2444 ^ n1560 ^ 1'b0 ;
  assign n2642 = ( n1558 & n1560 ) | ( n1558 & ~n2641 ) | ( n1560 & ~n2641 ) ;
  assign n2643 = n2444 ^ n1563 ^ 1'b0 ;
  assign n2644 = ( n1563 & n1565 ) | ( n1563 & ~n2643 ) | ( n1565 & ~n2643 ) ;
  assign n2645 = n2444 ^ n2307 ^ 1'b0 ;
  assign n2646 = ( n2307 & n2309 ) | ( n2307 & ~n2645 ) | ( n2309 & ~n2645 ) ;
  assign n2647 = n2444 ^ n2302 ^ 1'b0 ;
  assign n2648 = ( n2302 & n2304 ) | ( n2302 & ~n2647 ) | ( n2304 & ~n2647 ) ;
  assign n2649 = n2444 ^ n1549 ^ 1'b0 ;
  assign n2650 = ( n1547 & n1549 ) | ( n1547 & ~n2649 ) | ( n1549 & ~n2649 ) ;
  assign n2651 = n2444 ^ n1542 ^ 1'b0 ;
  assign n2652 = ( n1542 & n1544 ) | ( n1542 & ~n2651 ) | ( n1544 & ~n2651 ) ;
  assign n2653 = n2444 ^ n2343 ^ 1'b0 ;
  assign n2654 = ( n2341 & n2343 ) | ( n2341 & ~n2653 ) | ( n2343 & ~n2653 ) ;
  assign n2655 = n2444 ^ n2337 ^ 1'b0 ;
  assign n2656 = ( n2337 & n2339 ) | ( n2337 & ~n2655 ) | ( n2339 & ~n2655 ) ;
  assign n2657 = n2444 ^ n2330 ^ 1'b0 ;
  assign n2658 = ( n2328 & n2330 ) | ( n2328 & ~n2657 ) | ( n2330 & ~n2657 ) ;
  assign n2659 = n2444 ^ n2326 ^ 1'b0 ;
  assign n2660 = ( n2326 & n2333 ) | ( n2326 & ~n2659 ) | ( n2333 & ~n2659 ) ;
  assign n2661 = n2444 ^ n2363 ^ 1'b0 ;
  assign n2662 = ( n2363 & n2365 ) | ( n2363 & ~n2661 ) | ( n2365 & ~n2661 ) ;
  assign n2663 = n2444 ^ n2358 ^ 1'b0 ;
  assign n2664 = ( n2358 & n2360 ) | ( n2358 & ~n2663 ) | ( n2360 & ~n2663 ) ;
  assign n2665 = n2444 ^ n1538 ^ 1'b0 ;
  assign n2666 = ( n1536 & n1538 ) | ( n1536 & ~n2665 ) | ( n1538 & ~n2665 ) ;
  assign n2667 = n2444 ^ n1530 ^ 1'b0 ;
  assign n2668 = ( n1530 & n1532 ) | ( n1530 & ~n2667 ) | ( n1532 & ~n2667 ) ;
  assign n2669 = n2444 ^ n1511 ^ 1'b0 ;
  assign n2670 = ( n1509 & n1511 ) | ( n1509 & ~n2669 ) | ( n1511 & ~n2669 ) ;
  assign n2671 = n2444 ^ n1525 ^ 1'b0 ;
  assign n2672 = ( n1525 & n1527 ) | ( n1525 & ~n2671 ) | ( n1527 & ~n2671 ) ;
  assign n2673 = n2444 ^ n1516 ^ 1'b0 ;
  assign n2674 = ( n1514 & n1516 ) | ( n1514 & ~n2673 ) | ( n1516 & ~n2673 ) ;
  assign n2675 = n2444 ^ n1519 ^ 1'b0 ;
  assign n2676 = ( n1519 & n1521 ) | ( n1519 & ~n2675 ) | ( n1521 & ~n2675 ) ;
  assign n2677 = n2444 ^ n1500 ^ 1'b0 ;
  assign n2678 = ( n1500 & n1503 ) | ( n1500 & ~n2677 ) | ( n1503 & ~n2677 ) ;
  assign n2679 = n2444 ^ n1495 ^ 1'b0 ;
  assign n2680 = ( n1495 & n1497 ) | ( n1495 & ~n2679 ) | ( n1497 & ~n2679 ) ;
  assign n2681 = n2444 ^ n1491 ^ 1'b0 ;
  assign n2682 = ( n1489 & n1491 ) | ( n1489 & ~n2681 ) | ( n1491 & ~n2681 ) ;
  assign n2683 = n2444 ^ n1484 ^ 1'b0 ;
  assign n2684 = ( n1484 & n1486 ) | ( n1484 & ~n2683 ) | ( n1486 & ~n2683 ) ;
  assign n2685 = n2444 ^ n1480 ^ 1'b0 ;
  assign n2686 = ( n1478 & n1480 ) | ( n1478 & ~n2685 ) | ( n1480 & ~n2685 ) ;
  assign n2687 = n2444 ^ n1473 ^ 1'b0 ;
  assign n2688 = ( n1473 & n1475 ) | ( n1473 & ~n2687 ) | ( n1475 & ~n2687 ) ;
  assign n2689 = n2444 ^ n1468 ^ 1'b0 ;
  assign n2690 = ( n1466 & n1468 ) | ( n1466 & ~n2689 ) | ( n1468 & ~n2689 ) ;
  assign n2691 = n2444 ^ n1461 ^ 1'b0 ;
  assign n2692 = ( n1461 & n1463 ) | ( n1461 & ~n2691 ) | ( n1463 & ~n2691 ) ;
  assign n2693 = n2444 ^ n2431 ^ 1'b0 ;
  assign n2694 = ( n2431 & n2433 ) | ( n2431 & ~n2693 ) | ( n2433 & ~n2693 ) ;
  assign n2695 = n2444 ^ n2424 ^ 1'b0 ;
  assign n2696 = ( n2424 & n2426 ) | ( n2424 & ~n2695 ) | ( n2426 & ~n2695 ) ;
  assign n2697 = n2444 ^ n2418 ^ 1'b0 ;
  assign n2698 = ( n2418 & n2420 ) | ( n2418 & ~n2697 ) | ( n2420 & ~n2697 ) ;
  assign n2699 = n1456 | n2443 ;
  assign n2700 = n1458 & n2699 ;
  assign n2701 = n2444 ^ n979 ^ 1'b0 ;
  assign n2702 = ( n979 & n1452 ) | ( n979 & ~n2701 ) | ( n1452 & ~n2701 ) ;
  assign y0 = n2446 ;
  assign y1 = n2448 ;
  assign y2 = n2450 ;
  assign y3 = n2452 ;
  assign y4 = n2454 ;
  assign y5 = n2456 ;
  assign y6 = n2458 ;
  assign y7 = n2460 ;
  assign y8 = n2462 ;
  assign y9 = n2464 ;
  assign y10 = n2466 ;
  assign y11 = n2468 ;
  assign y12 = n2470 ;
  assign y13 = n2472 ;
  assign y14 = n2474 ;
  assign y15 = n2476 ;
  assign y16 = n2478 ;
  assign y17 = n2480 ;
  assign y18 = n2482 ;
  assign y19 = n2484 ;
  assign y20 = n2486 ;
  assign y21 = n2488 ;
  assign y22 = n2490 ;
  assign y23 = n2492 ;
  assign y24 = n2494 ;
  assign y25 = n2496 ;
  assign y26 = n2498 ;
  assign y27 = n2500 ;
  assign y28 = n2502 ;
  assign y29 = n2504 ;
  assign y30 = n2506 ;
  assign y31 = n2508 ;
  assign y32 = n2510 ;
  assign y33 = n2512 ;
  assign y34 = n2514 ;
  assign y35 = n2516 ;
  assign y36 = n2518 ;
  assign y37 = n2520 ;
  assign y38 = n2522 ;
  assign y39 = n2524 ;
  assign y40 = n2526 ;
  assign y41 = n2528 ;
  assign y42 = n2530 ;
  assign y43 = n2532 ;
  assign y44 = n2534 ;
  assign y45 = n2536 ;
  assign y46 = n2538 ;
  assign y47 = n2540 ;
  assign y48 = n2542 ;
  assign y49 = n2544 ;
  assign y50 = n2546 ;
  assign y51 = n2548 ;
  assign y52 = n2550 ;
  assign y53 = n2552 ;
  assign y54 = n2554 ;
  assign y55 = n2556 ;
  assign y56 = n2558 ;
  assign y57 = n2560 ;
  assign y58 = n2562 ;
  assign y59 = n2564 ;
  assign y60 = n2566 ;
  assign y61 = n2568 ;
  assign y62 = n2570 ;
  assign y63 = n2572 ;
  assign y64 = n2574 ;
  assign y65 = n2576 ;
  assign y66 = n2578 ;
  assign y67 = n2580 ;
  assign y68 = n2582 ;
  assign y69 = n2584 ;
  assign y70 = n2586 ;
  assign y71 = n2588 ;
  assign y72 = n2590 ;
  assign y73 = n2592 ;
  assign y74 = n2594 ;
  assign y75 = n2596 ;
  assign y76 = n2598 ;
  assign y77 = n2600 ;
  assign y78 = n2602 ;
  assign y79 = n2604 ;
  assign y80 = n2606 ;
  assign y81 = n2608 ;
  assign y82 = n2610 ;
  assign y83 = n2612 ;
  assign y84 = n2614 ;
  assign y85 = n2616 ;
  assign y86 = n2618 ;
  assign y87 = n2620 ;
  assign y88 = n2622 ;
  assign y89 = n2624 ;
  assign y90 = n2626 ;
  assign y91 = n2628 ;
  assign y92 = n2630 ;
  assign y93 = n2632 ;
  assign y94 = n2634 ;
  assign y95 = n2636 ;
  assign y96 = n2638 ;
  assign y97 = n2640 ;
  assign y98 = n2642 ;
  assign y99 = n2644 ;
  assign y100 = n2646 ;
  assign y101 = n2648 ;
  assign y102 = n2650 ;
  assign y103 = n2652 ;
  assign y104 = n2654 ;
  assign y105 = n2656 ;
  assign y106 = n2658 ;
  assign y107 = n2660 ;
  assign y108 = n2662 ;
  assign y109 = n2664 ;
  assign y110 = n2666 ;
  assign y111 = n2668 ;
  assign y112 = n2670 ;
  assign y113 = n2672 ;
  assign y114 = n2674 ;
  assign y115 = n2676 ;
  assign y116 = n2678 ;
  assign y117 = n2680 ;
  assign y118 = n2682 ;
  assign y119 = n2684 ;
  assign y120 = n2686 ;
  assign y121 = n2688 ;
  assign y122 = n2690 ;
  assign y123 = n2692 ;
  assign y124 = n2694 ;
  assign y125 = n2696 ;
  assign y126 = n2698 ;
  assign y127 = n2700 ;
  assign y128 = ~n2702 ;
  assign y129 = ~n2444 ;
endmodule
