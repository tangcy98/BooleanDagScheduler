module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , n77825 , n77826 , n77827 , n77828 , n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , n77835 , n77836 , n77837 , n77838 , n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , n77845 , n77846 , n77847 , n77848 , n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , n77855 , n77856 , n77857 , n77858 , n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , n77865 , n77866 , n77867 , n77868 , n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , n77875 , n77876 , n77877 , n77878 , n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , n77885 , n77886 , n77887 , n77888 , n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , n77895 , n77896 , n77897 , n77898 , n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , n77905 , n77906 , n77907 , n77908 , n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , n77915 , n77916 , n77917 , n77918 , n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , n77925 , n77926 , n77927 , n77928 , n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , n77935 , n77936 , n77937 , n77938 , n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , n77945 , n77946 , n77947 , n77948 , n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , n77955 , n77956 , n77957 , n77958 , n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , n77965 , n77966 , n77967 , n77968 , n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , n77975 , n77976 , n77977 , n77978 , n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , n77985 , n77986 , n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , n78005 , n78006 , n78007 , n78008 , n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , n78015 , n78016 , n78017 , n78018 , n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , n78025 , n78026 , n78027 , n78028 , n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , n78035 , n78036 , n78037 , n78038 , n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , n78045 , n78046 , n78047 , n78048 , n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , n78055 , n78056 , n78057 , n78058 , n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , n78065 , n78066 , n78067 , n78068 , n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , n78075 , n78076 , n78077 , n78078 , n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , n78085 , n78086 , n78087 , n78088 , n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , n78095 , n78096 , n78097 , n78098 , n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , n78105 , n78106 , n78107 , n78108 , n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , n78115 , n78116 , n78117 , n78118 , n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , n78125 , n78126 , n78127 , n78128 , n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , n78135 , n78136 , n78137 , n78138 , n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , n78145 , n78146 , n78147 , n78148 , n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , n78155 , n78156 , n78157 , n78158 , n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , n78165 , n78166 , n78167 , n78168 , n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , n78175 , n78176 , n78177 , n78178 , n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , n78185 , n78186 , n78187 , n78188 , n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , n78195 , n78196 , n78197 , n78198 , n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , n78205 , n78206 , n78207 , n78208 , n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , n78215 , n78216 , n78217 , n78218 , n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , n78225 , n78226 , n78227 , n78228 , n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , n78235 , n78236 , n78237 , n78238 , n78239 , n78240 , n78241 , n78242 , n78243 , n78244 , n78245 , n78246 , n78247 , n78248 , n78249 , n78250 , n78251 , n78252 , n78253 , n78254 , n78255 , n78256 , n78257 , n78258 , n78259 , n78260 , n78261 , n78262 , n78263 , n78264 , n78265 , n78266 , n78267 , n78268 , n78269 , n78270 , n78271 , n78272 , n78273 , n78274 , n78275 , n78276 , n78277 , n78278 , n78279 , n78280 , n78281 , n78282 , n78283 , n78284 , n78285 , n78286 , n78287 , n78288 , n78289 , n78290 , n78291 , n78292 , n78293 , n78294 , n78295 , n78296 , n78297 , n78298 , n78299 , n78300 , n78301 , n78302 , n78303 , n78304 , n78305 , n78306 , n78307 , n78308 , n78309 , n78310 , n78311 , n78312 , n78313 , n78314 , n78315 , n78316 , n78317 , n78318 , n78319 , n78320 , n78321 , n78322 , n78323 , n78324 , n78325 , n78326 , n78327 , n78328 , n78329 , n78330 , n78331 , n78332 , n78333 , n78334 , n78335 , n78336 , n78337 , n78338 , n78339 , n78340 , n78341 , n78342 , n78343 , n78344 , n78345 , n78346 , n78347 , n78348 , n78349 , n78350 , n78351 , n78352 , n78353 , n78354 , n78355 , n78356 , n78357 , n78358 , n78359 , n78360 , n78361 , n78362 , n78363 , n78364 , n78365 , n78366 , n78367 , n78368 , n78369 , n78370 , n78371 , n78372 , n78373 , n78374 , n78375 , n78376 , n78377 , n78378 , n78379 , n78380 , n78381 , n78382 , n78383 , n78384 , n78385 , n78386 , n78387 , n78388 , n78389 , n78390 , n78391 , n78392 , n78393 , n78394 , n78395 , n78396 , n78397 , n78398 , n78399 , n78400 , n78401 , n78402 , n78403 , n78404 , n78405 , n78406 , n78407 , n78408 , n78409 , n78410 , n78411 , n78412 , n78413 , n78414 , n78415 , n78416 , n78417 , n78418 , n78419 , n78420 , n78421 , n78422 , n78423 , n78424 , n78425 , n78426 , n78427 , n78428 , n78429 , n78430 , n78431 , n78432 , n78433 , n78434 , n78435 , n78436 , n78437 , n78438 , n78439 , n78440 , n78441 , n78442 , n78443 , n78444 , n78445 , n78446 , n78447 , n78448 , n78449 , n78450 , n78451 , n78452 , n78453 , n78454 , n78455 , n78456 , n78457 , n78458 , n78459 , n78460 , n78461 , n78462 , n78463 , n78464 , n78465 , n78466 , n78467 , n78468 , n78469 , n78470 , n78471 , n78472 , n78473 , n78474 , n78475 , n78476 , n78477 , n78478 , n78479 , n78480 , n78481 , n78482 , n78483 , n78484 , n78485 , n78486 , n78487 , n78488 , n78489 , n78490 , n78491 , n78492 , n78493 , n78494 , n78495 , n78496 , n78497 , n78498 , n78499 , n78500 , n78501 , n78502 , n78503 , n78504 , n78505 , n78506 , n78507 , n78508 , n78509 , n78510 , n78511 , n78512 , n78513 , n78514 , n78515 , n78516 , n78517 , n78518 , n78519 , n78520 , n78521 , n78522 , n78523 , n78524 , n78525 , n78526 , n78527 , n78528 , n78529 , n78530 , n78531 , n78532 , n78533 , n78534 , n78535 , n78536 , n78537 , n78538 , n78539 , n78540 , n78541 , n78542 , n78543 , n78544 , n78545 , n78546 , n78547 , n78548 , n78549 , n78550 , n78551 , n78552 , n78553 , n78554 , n78555 , n78556 , n78557 , n78558 , n78559 , n78560 , n78561 , n78562 , n78563 , n78564 , n78565 , n78566 , n78567 , n78568 , n78569 , n78570 , n78571 , n78572 , n78573 , n78574 , n78575 , n78576 , n78577 , n78578 , n78579 , n78580 , n78581 , n78582 , n78583 , n78584 , n78585 , n78586 , n78587 , n78588 , n78589 , n78590 , n78591 , n78592 , n78593 , n78594 , n78595 , n78596 , n78597 , n78598 , n78599 , n78600 , n78601 , n78602 , n78603 , n78604 , n78605 , n78606 , n78607 , n78608 , n78609 , n78610 , n78611 , n78612 , n78613 , n78614 , n78615 , n78616 , n78617 , n78618 , n78619 , n78620 , n78621 , n78622 , n78623 , n78624 , n78625 , n78626 , n78627 , n78628 , n78629 , n78630 , n78631 , n78632 , n78633 , n78634 , n78635 , n78636 , n78637 , n78638 , n78639 , n78640 , n78641 , n78642 , n78643 , n78644 , n78645 , n78646 , n78647 , n78648 , n78649 , n78650 , n78651 , n78652 , n78653 , n78654 , n78655 , n78656 , n78657 , n78658 , n78659 , n78660 , n78661 , n78662 , n78663 , n78664 , n78665 , n78666 , n78667 , n78668 , n78669 , n78670 , n78671 , n78672 , n78673 , n78674 , n78675 , n78676 , n78677 , n78678 , n78679 , n78680 , n78681 , n78682 , n78683 , n78684 , n78685 , n78686 , n78687 , n78688 , n78689 , n78690 , n78691 , n78692 , n78693 , n78694 , n78695 , n78696 , n78697 , n78698 , n78699 , n78700 , n78701 , n78702 , n78703 , n78704 , n78705 , n78706 , n78707 , n78708 , n78709 , n78710 , n78711 , n78712 , n78713 , n78714 , n78715 , n78716 , n78717 , n78718 , n78719 , n78720 , n78721 , n78722 , n78723 , n78724 , n78725 , n78726 , n78727 , n78728 , n78729 , n78730 , n78731 , n78732 , n78733 , n78734 , n78735 , n78736 , n78737 , n78738 , n78739 , n78740 , n78741 , n78742 , n78743 , n78744 , n78745 , n78746 , n78747 , n78748 , n78749 , n78750 , n78751 , n78752 , n78753 , n78754 , n78755 , n78756 , n78757 , n78758 , n78759 , n78760 , n78761 , n78762 , n78763 , n78764 , n78765 , n78766 , n78767 , n78768 , n78769 , n78770 , n78771 , n78772 , n78773 , n78774 , n78775 , n78776 , n78777 , n78778 , n78779 , n78780 , n78781 , n78782 , n78783 , n78784 , n78785 , n78786 , n78787 , n78788 , n78789 , n78790 , n78791 , n78792 , n78793 , n78794 , n78795 , n78796 , n78797 , n78798 , n78799 , n78800 , n78801 , n78802 , n78803 , n78804 , n78805 , n78806 , n78807 , n78808 , n78809 , n78810 , n78811 , n78812 , n78813 , n78814 , n78815 , n78816 , n78817 , n78818 , n78819 , n78820 , n78821 , n78822 , n78823 , n78824 , n78825 , n78826 , n78827 , n78828 , n78829 , n78830 , n78831 , n78832 , n78833 , n78834 , n78835 , n78836 , n78837 , n78838 , n78839 , n78840 , n78841 , n78842 , n78843 , n78844 , n78845 , n78846 , n78847 , n78848 , n78849 , n78850 , n78851 , n78852 , n78853 , n78854 , n78855 , n78856 , n78857 , n78858 , n78859 , n78860 , n78861 , n78862 , n78863 , n78864 , n78865 , n78866 , n78867 , n78868 , n78869 , n78870 , n78871 , n78872 , n78873 , n78874 , n78875 , n78876 , n78877 , n78878 , n78879 , n78880 , n78881 , n78882 , n78883 , n78884 , n78885 , n78886 , n78887 , n78888 , n78889 , n78890 , n78891 , n78892 , n78893 , n78894 , n78895 , n78896 , n78897 , n78898 , n78899 , n78900 , n78901 , n78902 , n78903 , n78904 , n78905 , n78906 , n78907 , n78908 , n78909 , n78910 , n78911 , n78912 , n78913 , n78914 , n78915 , n78916 , n78917 , n78918 , n78919 , n78920 , n78921 , n78922 , n78923 , n78924 , n78925 , n78926 , n78927 , n78928 , n78929 , n78930 , n78931 , n78932 , n78933 , n78934 , n78935 , n78936 , n78937 , n78938 , n78939 , n78940 , n78941 , n78942 , n78943 , n78944 , n78945 , n78946 , n78947 , n78948 , n78949 , n78950 , n78951 , n78952 , n78953 , n78954 , n78955 , n78956 , n78957 , n78958 , n78959 , n78960 , n78961 , n78962 , n78963 , n78964 , n78965 , n78966 , n78967 , n78968 , n78969 , n78970 , n78971 , n78972 , n78973 , n78974 , n78975 , n78976 , n78977 , n78978 , n78979 , n78980 , n78981 , n78982 , n78983 , n78984 , n78985 , n78986 , n78987 , n78988 , n78989 , n78990 , n78991 , n78992 , n78993 , n78994 , n78995 , n78996 , n78997 , n78998 , n78999 , n79000 , n79001 , n79002 , n79003 , n79004 , n79005 , n79006 , n79007 , n79008 , n79009 , n79010 , n79011 , n79012 , n79013 , n79014 , n79015 , n79016 , n79017 , n79018 , n79019 , n79020 , n79021 , n79022 , n79023 , n79024 , n79025 , n79026 , n79027 , n79028 , n79029 , n79030 , n79031 , n79032 , n79033 , n79034 , n79035 , n79036 , n79037 , n79038 , n79039 , n79040 , n79041 , n79042 , n79043 , n79044 , n79045 , n79046 , n79047 , n79048 , n79049 , n79050 , n79051 , n79052 , n79053 , n79054 , n79055 , n79056 , n79057 , n79058 , n79059 , n79060 , n79061 , n79062 , n79063 , n79064 , n79065 , n79066 , n79067 , n79068 , n79069 , n79070 , n79071 , n79072 , n79073 , n79074 , n79075 , n79076 , n79077 , n79078 , n79079 , n79080 , n79081 , n79082 , n79083 , n79084 , n79085 , n79086 , n79087 , n79088 , n79089 , n79090 , n79091 , n79092 , n79093 , n79094 , n79095 , n79096 , n79097 , n79098 , n79099 , n79100 , n79101 , n79102 , n79103 , n79104 , n79105 , n79106 , n79107 , n79108 , n79109 , n79110 , n79111 , n79112 , n79113 , n79114 , n79115 , n79116 , n79117 , n79118 , n79119 , n79120 , n79121 , n79122 , n79123 , n79124 , n79125 , n79126 , n79127 , n79128 , n79129 , n79130 , n79131 , n79132 , n79133 , n79134 , n79135 , n79136 , n79137 , n79138 , n79139 , n79140 , n79141 , n79142 , n79143 , n79144 , n79145 , n79146 , n79147 , n79148 , n79149 , n79150 , n79151 , n79152 , n79153 , n79154 , n79155 , n79156 , n79157 , n79158 , n79159 , n79160 , n79161 , n79162 , n79163 , n79164 , n79165 , n79166 , n79167 , n79168 , n79169 , n79170 , n79171 , n79172 , n79173 , n79174 , n79175 , n79176 , n79177 , n79178 , n79179 , n79180 , n79181 , n79182 , n79183 , n79184 , n79185 , n79186 , n79187 , n79188 , n79189 , n79190 , n79191 , n79192 , n79193 , n79194 , n79195 , n79196 , n79197 , n79198 , n79199 , n79200 , n79201 , n79202 , n79203 , n79204 , n79205 , n79206 , n79207 , n79208 , n79209 , n79210 , n79211 , n79212 , n79213 , n79214 , n79215 , n79216 , n79217 , n79218 , n79219 , n79220 , n79221 , n79222 , n79223 , n79224 , n79225 , n79226 , n79227 , n79228 , n79229 , n79230 , n79231 , n79232 , n79233 , n79234 , n79235 , n79236 , n79237 , n79238 , n79239 , n79240 , n79241 , n79242 , n79243 , n79244 , n79245 , n79246 , n79247 , n79248 , n79249 , n79250 , n79251 , n79252 , n79253 , n79254 , n79255 , n79256 , n79257 , n79258 , n79259 , n79260 , n79261 , n79262 , n79263 , n79264 , n79265 , n79266 , n79267 , n79268 , n79269 , n79270 , n79271 , n79272 , n79273 , n79274 , n79275 , n79276 , n79277 , n79278 , n79279 , n79280 , n79281 , n79282 , n79283 , n79284 , n79285 , n79286 , n79287 , n79288 , n79289 , n79290 , n79291 , n79292 , n79293 , n79294 , n79295 , n79296 , n79297 , n79298 , n79299 , n79300 , n79301 , n79302 , n79303 , n79304 , n79305 , n79306 , n79307 , n79308 , n79309 , n79310 , n79311 , n79312 , n79313 , n79314 , n79315 , n79316 , n79317 , n79318 , n79319 , n79320 , n79321 , n79322 , n79323 , n79324 , n79325 , n79326 , n79327 , n79328 , n79329 , n79330 , n79331 , n79332 , n79333 , n79334 , n79335 , n79336 , n79337 , n79338 , n79339 , n79340 , n79341 , n79342 , n79343 , n79344 , n79345 , n79346 , n79347 , n79348 , n79349 , n79350 , n79351 , n79352 , n79353 , n79354 , n79355 , n79356 , n79357 , n79358 , n79359 , n79360 , n79361 , n79362 , n79363 , n79364 , n79365 , n79366 , n79367 , n79368 , n79369 , n79370 , n79371 , n79372 , n79373 , n79374 , n79375 , n79376 , n79377 , n79378 , n79379 , n79380 , n79381 , n79382 , n79383 , n79384 , n79385 , n79386 , n79387 , n79388 , n79389 , n79390 , n79391 , n79392 , n79393 , n79394 , n79395 , n79396 , n79397 , n79398 , n79399 , n79400 , n79401 , n79402 , n79403 , n79404 , n79405 , n79406 , n79407 , n79408 , n79409 , n79410 , n79411 , n79412 , n79413 , n79414 , n79415 , n79416 , n79417 , n79418 , n79419 , n79420 , n79421 , n79422 , n79423 , n79424 , n79425 , n79426 , n79427 , n79428 , n79429 , n79430 , n79431 , n79432 , n79433 , n79434 , n79435 , n79436 , n79437 , n79438 , n79439 , n79440 , n79441 , n79442 , n79443 , n79444 , n79445 , n79446 , n79447 , n79448 , n79449 , n79450 , n79451 , n79452 , n79453 , n79454 , n79455 , n79456 , n79457 , n79458 , n79459 , n79460 , n79461 , n79462 , n79463 , n79464 , n79465 , n79466 , n79467 , n79468 , n79469 , n79470 , n79471 , n79472 , n79473 , n79474 , n79475 , n79476 , n79477 , n79478 , n79479 , n79480 , n79481 , n79482 , n79483 , n79484 , n79485 , n79486 , n79487 , n79488 , n79489 , n79490 , n79491 , n79492 , n79493 , n79494 , n79495 , n79496 , n79497 , n79498 , n79499 , n79500 , n79501 , n79502 , n79503 , n79504 , n79505 , n79506 , n79507 , n79508 , n79509 , n79510 , n79511 , n79512 , n79513 , n79514 , n79515 , n79516 , n79517 , n79518 , n79519 , n79520 , n79521 , n79522 , n79523 , n79524 , n79525 , n79526 , n79527 , n79528 , n79529 , n79530 , n79531 , n79532 , n79533 , n79534 , n79535 , n79536 , n79537 , n79538 , n79539 , n79540 , n79541 , n79542 , n79543 , n79544 , n79545 , n79546 , n79547 , n79548 , n79549 , n79550 , n79551 , n79552 , n79553 , n79554 , n79555 , n79556 , n79557 , n79558 , n79559 , n79560 , n79561 , n79562 , n79563 , n79564 , n79565 , n79566 , n79567 , n79568 , n79569 , n79570 , n79571 , n79572 , n79573 , n79574 , n79575 , n79576 , n79577 , n79578 , n79579 , n79580 , n79581 , n79582 , n79583 , n79584 , n79585 , n79586 , n79587 , n79588 , n79589 , n79590 , n79591 , n79592 , n79593 , n79594 , n79595 , n79596 , n79597 , n79598 , n79599 , n79600 , n79601 , n79602 , n79603 , n79604 , n79605 , n79606 , n79607 , n79608 , n79609 , n79610 , n79611 , n79612 , n79613 , n79614 , n79615 , n79616 , n79617 , n79618 , n79619 , n79620 , n79621 , n79622 , n79623 , n79624 , n79625 , n79626 , n79627 , n79628 , n79629 , n79630 , n79631 , n79632 , n79633 , n79634 , n79635 , n79636 , n79637 , n79638 , n79639 , n79640 , n79641 , n79642 , n79643 , n79644 , n79645 , n79646 , n79647 , n79648 , n79649 , n79650 , n79651 , n79652 , n79653 , n79654 , n79655 , n79656 , n79657 , n79658 , n79659 , n79660 , n79661 , n79662 , n79663 , n79664 , n79665 , n79666 , n79667 , n79668 , n79669 , n79670 , n79671 , n79672 , n79673 , n79674 , n79675 , n79676 , n79677 , n79678 , n79679 , n79680 , n79681 , n79682 , n79683 , n79684 , n79685 , n79686 , n79687 , n79688 , n79689 , n79690 , n79691 , n79692 , n79693 , n79694 , n79695 , n79696 , n79697 , n79698 , n79699 , n79700 , n79701 , n79702 , n79703 , n79704 , n79705 , n79706 , n79707 , n79708 , n79709 , n79710 , n79711 , n79712 , n79713 , n79714 , n79715 , n79716 , n79717 , n79718 , n79719 , n79720 , n79721 , n79722 , n79723 , n79724 , n79725 , n79726 , n79727 , n79728 , n79729 , n79730 , n79731 , n79732 , n79733 , n79734 , n79735 , n79736 , n79737 , n79738 , n79739 , n79740 , n79741 , n79742 , n79743 , n79744 , n79745 , n79746 , n79747 , n79748 , n79749 , n79750 , n79751 , n79752 , n79753 , n79754 , n79755 , n79756 , n79757 , n79758 , n79759 , n79760 , n79761 , n79762 , n79763 , n79764 , n79765 , n79766 , n79767 , n79768 , n79769 , n79770 , n79771 , n79772 , n79773 , n79774 , n79775 , n79776 , n79777 , n79778 , n79779 , n79780 , n79781 , n79782 , n79783 , n79784 , n79785 , n79786 , n79787 , n79788 , n79789 , n79790 , n79791 , n79792 , n79793 , n79794 , n79795 , n79796 , n79797 , n79798 , n79799 , n79800 , n79801 , n79802 , n79803 , n79804 , n79805 , n79806 , n79807 , n79808 , n79809 , n79810 , n79811 , n79812 , n79813 , n79814 , n79815 , n79816 , n79817 , n79818 , n79819 , n79820 , n79821 , n79822 , n79823 , n79824 , n79825 , n79826 , n79827 , n79828 , n79829 , n79830 , n79831 , n79832 , n79833 , n79834 , n79835 , n79836 , n79837 , n79838 , n79839 , n79840 , n79841 , n79842 , n79843 , n79844 , n79845 , n79846 , n79847 , n79848 , n79849 , n79850 , n79851 , n79852 , n79853 , n79854 , n79855 , n79856 , n79857 , n79858 , n79859 , n79860 , n79861 , n79862 , n79863 , n79864 , n79865 , n79866 , n79867 , n79868 , n79869 , n79870 , n79871 , n79872 , n79873 , n79874 , n79875 , n79876 , n79877 , n79878 , n79879 , n79880 , n79881 , n79882 , n79883 , n79884 , n79885 , n79886 , n79887 , n79888 , n79889 , n79890 , n79891 , n79892 , n79893 , n79894 , n79895 , n79896 , n79897 , n79898 , n79899 , n79900 , n79901 , n79902 , n79903 , n79904 , n79905 , n79906 , n79907 , n79908 , n79909 , n79910 , n79911 , n79912 , n79913 , n79914 , n79915 , n79916 , n79917 , n79918 , n79919 , n79920 , n79921 , n79922 , n79923 , n79924 , n79925 , n79926 , n79927 , n79928 , n79929 , n79930 , n79931 , n79932 , n79933 , n79934 , n79935 , n79936 , n79937 , n79938 , n79939 , n79940 , n79941 , n79942 , n79943 , n79944 , n79945 , n79946 , n79947 , n79948 , n79949 , n79950 , n79951 , n79952 , n79953 , n79954 , n79955 , n79956 , n79957 , n79958 , n79959 , n79960 , n79961 , n79962 , n79963 , n79964 , n79965 , n79966 , n79967 , n79968 , n79969 , n79970 , n79971 , n79972 , n79973 , n79974 , n79975 , n79976 , n79977 , n79978 , n79979 , n79980 , n79981 , n79982 , n79983 , n79984 , n79985 , n79986 , n79987 , n79988 , n79989 , n79990 , n79991 , n79992 , n79993 , n79994 , n79995 , n79996 , n79997 , n79998 , n79999 , n80000 , n80001 , n80002 , n80003 , n80004 , n80005 , n80006 , n80007 , n80008 , n80009 , n80010 , n80011 , n80012 , n80013 , n80014 , n80015 , n80016 , n80017 , n80018 , n80019 , n80020 , n80021 , n80022 , n80023 , n80024 , n80025 , n80026 , n80027 , n80028 , n80029 , n80030 , n80031 , n80032 , n80033 , n80034 , n80035 , n80036 , n80037 , n80038 , n80039 , n80040 , n80041 , n80042 , n80043 , n80044 , n80045 , n80046 , n80047 , n80048 , n80049 , n80050 , n80051 , n80052 , n80053 , n80054 , n80055 , n80056 , n80057 , n80058 , n80059 , n80060 , n80061 , n80062 , n80063 , n80064 , n80065 , n80066 , n80067 , n80068 , n80069 , n80070 , n80071 , n80072 , n80073 , n80074 , n80075 , n80076 , n80077 , n80078 , n80079 , n80080 , n80081 , n80082 , n80083 , n80084 , n80085 , n80086 , n80087 , n80088 , n80089 , n80090 , n80091 , n80092 , n80093 , n80094 , n80095 , n80096 , n80097 , n80098 , n80099 , n80100 , n80101 , n80102 , n80103 , n80104 , n80105 , n80106 , n80107 , n80108 , n80109 , n80110 , n80111 , n80112 , n80113 , n80114 , n80115 , n80116 , n80117 , n80118 , n80119 , n80120 , n80121 , n80122 , n80123 , n80124 , n80125 , n80126 , n80127 , n80128 , n80129 , n80130 , n80131 , n80132 , n80133 , n80134 , n80135 , n80136 , n80137 , n80138 , n80139 , n80140 , n80141 , n80142 , n80143 , n80144 , n80145 , n80146 , n80147 , n80148 , n80149 , n80150 , n80151 , n80152 , n80153 , n80154 , n80155 , n80156 , n80157 , n80158 , n80159 , n80160 , n80161 , n80162 , n80163 , n80164 , n80165 , n80166 , n80167 , n80168 , n80169 , n80170 , n80171 , n80172 , n80173 , n80174 , n80175 , n80176 , n80177 , n80178 , n80179 , n80180 , n80181 , n80182 , n80183 , n80184 , n80185 , n80186 , n80187 , n80188 , n80189 , n80190 , n80191 , n80192 , n80193 , n80194 , n80195 , n80196 , n80197 , n80198 , n80199 , n80200 , n80201 , n80202 , n80203 , n80204 , n80205 , n80206 , n80207 , n80208 , n80209 , n80210 , n80211 , n80212 , n80213 , n80214 , n80215 , n80216 , n80217 , n80218 , n80219 , n80220 , n80221 , n80222 , n80223 , n80224 , n80225 , n80226 , n80227 , n80228 , n80229 , n80230 , n80231 , n80232 , n80233 , n80234 , n80235 , n80236 , n80237 , n80238 , n80239 , n80240 , n80241 , n80242 , n80243 , n80244 , n80245 , n80246 , n80247 , n80248 , n80249 , n80250 , n80251 , n80252 , n80253 , n80254 , n80255 , n80256 , n80257 , n80258 , n80259 , n80260 , n80261 , n80262 , n80263 , n80264 , n80265 , n80266 , n80267 , n80268 , n80269 , n80270 , n80271 , n80272 , n80273 , n80274 , n80275 , n80276 , n80277 , n80278 , n80279 , n80280 , n80281 , n80282 , n80283 , n80284 , n80285 , n80286 , n80287 , n80288 , n80289 , n80290 , n80291 , n80292 , n80293 , n80294 , n80295 , n80296 , n80297 , n80298 , n80299 , n80300 , n80301 , n80302 , n80303 , n80304 , n80305 , n80306 , n80307 , n80308 , n80309 , n80310 , n80311 , n80312 , n80313 , n80314 , n80315 , n80316 , n80317 , n80318 , n80319 , n80320 , n80321 , n80322 , n80323 , n80324 , n80325 , n80326 , n80327 , n80328 , n80329 , n80330 , n80331 , n80332 , n80333 , n80334 , n80335 , n80336 , n80337 , n80338 , n80339 , n80340 , n80341 , n80342 , n80343 , n80344 , n80345 , n80346 , n80347 , n80348 , n80349 , n80350 , n80351 , n80352 , n80353 , n80354 , n80355 , n80356 , n80357 , n80358 , n80359 , n80360 , n80361 , n80362 , n80363 , n80364 , n80365 , n80366 , n80367 , n80368 , n80369 , n80370 , n80371 , n80372 , n80373 , n80374 , n80375 , n80376 , n80377 , n80378 , n80379 , n80380 , n80381 , n80382 , n80383 , n80384 , n80385 , n80386 , n80387 , n80388 , n80389 , n80390 , n80391 , n80392 , n80393 , n80394 , n80395 , n80396 , n80397 , n80398 , n80399 , n80400 , n80401 , n80402 , n80403 , n80404 , n80405 , n80406 , n80407 , n80408 , n80409 , n80410 , n80411 , n80412 , n80413 , n80414 , n80415 , n80416 , n80417 , n80418 , n80419 , n80420 , n80421 , n80422 , n80423 , n80424 , n80425 , n80426 , n80427 , n80428 , n80429 , n80430 , n80431 , n80432 , n80433 , n80434 , n80435 , n80436 , n80437 , n80438 , n80439 , n80440 , n80441 , n80442 , n80443 , n80444 , n80445 , n80446 , n80447 , n80448 , n80449 , n80450 , n80451 , n80452 , n80453 , n80454 , n80455 , n80456 , n80457 , n80458 , n80459 , n80460 , n80461 , n80462 , n80463 , n80464 , n80465 , n80466 , n80467 , n80468 , n80469 , n80470 , n80471 , n80472 , n80473 , n80474 , n80475 , n80476 , n80477 , n80478 , n80479 , n80480 , n80481 , n80482 , n80483 , n80484 , n80485 , n80486 , n80487 , n80488 , n80489 , n80490 , n80491 , n80492 , n80493 , n80494 , n80495 , n80496 , n80497 , n80498 , n80499 , n80500 , n80501 , n80502 , n80503 , n80504 , n80505 , n80506 , n80507 , n80508 , n80509 , n80510 , n80511 , n80512 , n80513 , n80514 , n80515 , n80516 , n80517 , n80518 , n80519 , n80520 , n80521 , n80522 , n80523 , n80524 , n80525 , n80526 , n80527 , n80528 , n80529 , n80530 , n80531 , n80532 , n80533 , n80534 , n80535 , n80536 , n80537 , n80538 , n80539 , n80540 , n80541 , n80542 , n80543 , n80544 , n80545 , n80546 , n80547 , n80548 , n80549 , n80550 , n80551 , n80552 , n80553 , n80554 , n80555 , n80556 , n80557 , n80558 , n80559 , n80560 , n80561 , n80562 , n80563 , n80564 , n80565 , n80566 , n80567 , n80568 , n80569 , n80570 , n80571 , n80572 , n80573 , n80574 , n80575 , n80576 , n80577 , n80578 , n80579 , n80580 , n80581 , n80582 , n80583 , n80584 , n80585 , n80586 , n80587 , n80588 , n80589 , n80590 , n80591 , n80592 , n80593 , n80594 , n80595 , n80596 , n80597 , n80598 , n80599 , n80600 , n80601 , n80602 , n80603 , n80604 , n80605 , n80606 , n80607 , n80608 , n80609 , n80610 , n80611 , n80612 , n80613 , n80614 , n80615 , n80616 , n80617 , n80618 , n80619 , n80620 , n80621 , n80622 , n80623 , n80624 , n80625 , n80626 , n80627 , n80628 , n80629 , n80630 , n80631 , n80632 , n80633 , n80634 , n80635 , n80636 , n80637 , n80638 , n80639 , n80640 , n80641 , n80642 , n80643 , n80644 , n80645 , n80646 , n80647 , n80648 , n80649 , n80650 , n80651 , n80652 , n80653 , n80654 , n80655 , n80656 , n80657 , n80658 , n80659 , n80660 , n80661 , n80662 , n80663 , n80664 , n80665 , n80666 , n80667 , n80668 , n80669 , n80670 , n80671 , n80672 , n80673 , n80674 , n80675 , n80676 , n80677 , n80678 , n80679 , n80680 , n80681 , n80682 , n80683 , n80684 , n80685 , n80686 , n80687 , n80688 , n80689 , n80690 , n80691 , n80692 , n80693 , n80694 , n80695 , n80696 , n80697 , n80698 , n80699 , n80700 , n80701 , n80702 , n80703 , n80704 , n80705 , n80706 , n80707 , n80708 , n80709 , n80710 , n80711 , n80712 , n80713 , n80714 , n80715 , n80716 , n80717 , n80718 , n80719 , n80720 , n80721 , n80722 , n80723 , n80724 , n80725 , n80726 , n80727 , n80728 , n80729 , n80730 , n80731 , n80732 , n80733 , n80734 , n80735 , n80736 , n80737 , n80738 , n80739 , n80740 , n80741 , n80742 , n80743 , n80744 , n80745 , n80746 , n80747 , n80748 , n80749 , n80750 , n80751 , n80752 , n80753 , n80754 , n80755 , n80756 , n80757 , n80758 , n80759 , n80760 , n80761 , n80762 , n80763 , n80764 , n80765 , n80766 , n80767 , n80768 , n80769 , n80770 , n80771 , n80772 , n80773 , n80774 , n80775 , n80776 , n80777 , n80778 , n80779 , n80780 , n80781 , n80782 , n80783 , n80784 , n80785 , n80786 , n80787 , n80788 , n80789 , n80790 , n80791 , n80792 , n80793 , n80794 , n80795 , n80796 , n80797 , n80798 , n80799 , n80800 , n80801 , n80802 , n80803 , n80804 , n80805 , n80806 , n80807 , n80808 , n80809 , n80810 , n80811 , n80812 , n80813 , n80814 , n80815 , n80816 , n80817 , n80818 , n80819 , n80820 , n80821 , n80822 , n80823 , n80824 , n80825 , n80826 , n80827 , n80828 , n80829 , n80830 , n80831 , n80832 , n80833 , n80834 , n80835 , n80836 , n80837 , n80838 , n80839 , n80840 , n80841 , n80842 , n80843 , n80844 , n80845 , n80846 , n80847 , n80848 , n80849 , n80850 , n80851 , n80852 , n80853 , n80854 , n80855 , n80856 , n80857 , n80858 , n80859 , n80860 , n80861 , n80862 , n80863 , n80864 , n80865 , n80866 , n80867 , n80868 , n80869 , n80870 , n80871 , n80872 , n80873 , n80874 , n80875 , n80876 , n80877 , n80878 , n80879 , n80880 , n80881 , n80882 , n80883 , n80884 , n80885 , n80886 , n80887 , n80888 , n80889 , n80890 , n80891 , n80892 , n80893 , n80894 , n80895 , n80896 , n80897 , n80898 , n80899 , n80900 , n80901 , n80902 , n80903 , n80904 , n80905 , n80906 , n80907 , n80908 , n80909 , n80910 , n80911 , n80912 , n80913 , n80914 , n80915 , n80916 , n80917 , n80918 , n80919 , n80920 , n80921 , n80922 , n80923 , n80924 , n80925 , n80926 , n80927 , n80928 , n80929 , n80930 , n80931 , n80932 , n80933 , n80934 , n80935 , n80936 , n80937 , n80938 , n80939 , n80940 , n80941 , n80942 , n80943 , n80944 , n80945 , n80946 , n80947 , n80948 , n80949 , n80950 , n80951 , n80952 , n80953 , n80954 , n80955 , n80956 , n80957 , n80958 , n80959 , n80960 , n80961 , n80962 , n80963 , n80964 , n80965 , n80966 , n80967 , n80968 , n80969 , n80970 , n80971 , n80972 , n80973 , n80974 , n80975 , n80976 , n80977 , n80978 , n80979 , n80980 , n80981 , n80982 , n80983 , n80984 , n80985 , n80986 , n80987 , n80988 , n80989 , n80990 , n80991 , n80992 , n80993 , n80994 , n80995 , n80996 , n80997 , n80998 , n80999 , n81000 , n81001 , n81002 , n81003 , n81004 , n81005 , n81006 , n81007 , n81008 , n81009 , n81010 , n81011 , n81012 , n81013 , n81014 , n81015 , n81016 , n81017 , n81018 , n81019 , n81020 , n81021 , n81022 , n81023 , n81024 , n81025 , n81026 , n81027 , n81028 , n81029 , n81030 , n81031 , n81032 , n81033 , n81034 , n81035 , n81036 , n81037 , n81038 , n81039 , n81040 , n81041 , n81042 , n81043 , n81044 , n81045 , n81046 , n81047 , n81048 , n81049 , n81050 , n81051 , n81052 , n81053 , n81054 , n81055 , n81056 , n81057 , n81058 , n81059 , n81060 , n81061 , n81062 , n81063 , n81064 , n81065 , n81066 , n81067 , n81068 , n81069 , n81070 , n81071 , n81072 , n81073 , n81074 , n81075 , n81076 , n81077 , n81078 , n81079 , n81080 , n81081 , n81082 , n81083 , n81084 , n81085 , n81086 , n81087 , n81088 , n81089 , n81090 , n81091 , n81092 , n81093 , n81094 , n81095 , n81096 , n81097 , n81098 , n81099 , n81100 , n81101 , n81102 , n81103 , n81104 , n81105 , n81106 , n81107 , n81108 , n81109 , n81110 , n81111 , n81112 , n81113 , n81114 , n81115 , n81116 , n81117 , n81118 , n81119 , n81120 , n81121 , n81122 , n81123 , n81124 , n81125 , n81126 , n81127 , n81128 , n81129 , n81130 , n81131 , n81132 , n81133 , n81134 , n81135 , n81136 , n81137 , n81138 , n81139 , n81140 , n81141 , n81142 , n81143 , n81144 , n81145 , n81146 , n81147 , n81148 , n81149 , n81150 , n81151 , n81152 , n81153 , n81154 , n81155 , n81156 , n81157 , n81158 , n81159 , n81160 , n81161 , n81162 , n81163 , n81164 , n81165 , n81166 , n81167 , n81168 , n81169 , n81170 , n81171 , n81172 , n81173 , n81174 , n81175 , n81176 , n81177 , n81178 , n81179 , n81180 , n81181 , n81182 , n81183 , n81184 , n81185 , n81186 , n81187 , n81188 , n81189 , n81190 , n81191 , n81192 , n81193 , n81194 , n81195 , n81196 , n81197 , n81198 , n81199 , n81200 , n81201 , n81202 , n81203 , n81204 , n81205 , n81206 , n81207 , n81208 , n81209 , n81210 , n81211 , n81212 , n81213 , n81214 , n81215 , n81216 , n81217 , n81218 , n81219 , n81220 , n81221 , n81222 , n81223 , n81224 , n81225 , n81226 , n81227 , n81228 , n81229 , n81230 , n81231 , n81232 , n81233 , n81234 , n81235 , n81236 , n81237 , n81238 , n81239 , n81240 , n81241 , n81242 , n81243 , n81244 , n81245 , n81246 , n81247 , n81248 , n81249 , n81250 , n81251 , n81252 , n81253 , n81254 , n81255 , n81256 , n81257 , n81258 , n81259 , n81260 , n81261 , n81262 , n81263 , n81264 , n81265 , n81266 , n81267 , n81268 , n81269 , n81270 , n81271 , n81272 , n81273 , n81274 , n81275 , n81276 , n81277 , n81278 , n81279 , n81280 , n81281 , n81282 , n81283 , n81284 , n81285 , n81286 , n81287 , n81288 , n81289 , n81290 , n81291 , n81292 , n81293 , n81294 , n81295 , n81296 , n81297 , n81298 , n81299 , n81300 , n81301 , n81302 , n81303 , n81304 , n81305 , n81306 , n81307 , n81308 , n81309 , n81310 , n81311 , n81312 , n81313 , n81314 , n81315 , n81316 , n81317 , n81318 , n81319 , n81320 , n81321 , n81322 , n81323 , n81324 , n81325 , n81326 , n81327 , n81328 , n81329 , n81330 , n81331 , n81332 , n81333 , n81334 , n81335 , n81336 , n81337 , n81338 , n81339 , n81340 , n81341 , n81342 , n81343 , n81344 , n81345 , n81346 , n81347 , n81348 , n81349 , n81350 , n81351 , n81352 , n81353 , n81354 , n81355 , n81356 , n81357 , n81358 , n81359 , n81360 , n81361 , n81362 , n81363 , n81364 , n81365 , n81366 , n81367 , n81368 , n81369 , n81370 , n81371 , n81372 , n81373 , n81374 , n81375 , n81376 , n81377 , n81378 , n81379 , n81380 , n81381 , n81382 , n81383 , n81384 , n81385 , n81386 , n81387 , n81388 , n81389 , n81390 , n81391 , n81392 , n81393 , n81394 , n81395 , n81396 , n81397 , n81398 , n81399 , n81400 , n81401 , n81402 , n81403 , n81404 , n81405 , n81406 , n81407 , n81408 , n81409 , n81410 , n81411 , n81412 , n81413 , n81414 , n81415 , n81416 , n81417 , n81418 , n81419 , n81420 , n81421 , n81422 , n81423 , n81424 , n81425 , n81426 , n81427 , n81428 , n81429 , n81430 , n81431 , n81432 , n81433 , n81434 , n81435 , n81436 , n81437 , n81438 , n81439 , n81440 , n81441 , n81442 , n81443 , n81444 , n81445 , n81446 , n81447 , n81448 , n81449 , n81450 , n81451 , n81452 , n81453 , n81454 , n81455 , n81456 , n81457 , n81458 , n81459 , n81460 , n81461 , n81462 , n81463 , n81464 , n81465 , n81466 , n81467 , n81468 , n81469 , n81470 , n81471 , n81472 , n81473 , n81474 , n81475 , n81476 , n81477 , n81478 , n81479 , n81480 , n81481 , n81482 , n81483 , n81484 , n81485 , n81486 , n81487 , n81488 , n81489 , n81490 , n81491 , n81492 , n81493 , n81494 , n81495 , n81496 , n81497 , n81498 , n81499 , n81500 , n81501 , n81502 , n81503 , n81504 , n81505 , n81506 , n81507 , n81508 , n81509 , n81510 , n81511 , n81512 , n81513 , n81514 , n81515 , n81516 , n81517 , n81518 , n81519 , n81520 , n81521 , n81522 , n81523 , n81524 , n81525 , n81526 , n81527 , n81528 , n81529 , n81530 , n81531 , n81532 , n81533 , n81534 , n81535 , n81536 , n81537 , n81538 , n81539 , n81540 , n81541 , n81542 , n81543 , n81544 , n81545 , n81546 , n81547 , n81548 , n81549 , n81550 , n81551 , n81552 , n81553 , n81554 , n81555 , n81556 , n81557 , n81558 , n81559 , n81560 , n81561 , n81562 , n81563 , n81564 , n81565 , n81566 , n81567 , n81568 , n81569 , n81570 , n81571 , n81572 , n81573 , n81574 , n81575 , n81576 , n81577 , n81578 , n81579 , n81580 , n81581 , n81582 , n81583 , n81584 , n81585 , n81586 , n81587 , n81588 , n81589 , n81590 , n81591 , n81592 , n81593 , n81594 , n81595 , n81596 , n81597 , n81598 , n81599 , n81600 , n81601 , n81602 , n81603 , n81604 , n81605 , n81606 , n81607 , n81608 , n81609 , n81610 , n81611 , n81612 , n81613 , n81614 , n81615 , n81616 , n81617 , n81618 , n81619 , n81620 , n81621 , n81622 , n81623 , n81624 , n81625 , n81626 , n81627 , n81628 , n81629 , n81630 , n81631 , n81632 , n81633 , n81634 , n81635 , n81636 , n81637 , n81638 , n81639 , n81640 , n81641 , n81642 , n81643 , n81644 , n81645 , n81646 , n81647 , n81648 , n81649 , n81650 , n81651 , n81652 , n81653 , n81654 , n81655 , n81656 , n81657 , n81658 , n81659 , n81660 , n81661 , n81662 , n81663 , n81664 , n81665 , n81666 , n81667 , n81668 , n81669 , n81670 , n81671 , n81672 , n81673 , n81674 , n81675 , n81676 , n81677 , n81678 , n81679 , n81680 , n81681 , n81682 , n81683 , n81684 , n81685 , n81686 , n81687 , n81688 , n81689 , n81690 , n81691 , n81692 , n81693 , n81694 , n81695 , n81696 , n81697 , n81698 , n81699 , n81700 , n81701 , n81702 , n81703 , n81704 , n81705 , n81706 , n81707 , n81708 , n81709 , n81710 , n81711 , n81712 , n81713 , n81714 , n81715 , n81716 , n81717 , n81718 , n81719 , n81720 , n81721 , n81722 , n81723 , n81724 , n81725 , n81726 , n81727 , n81728 , n81729 , n81730 , n81731 , n81732 , n81733 , n81734 , n81735 , n81736 , n81737 , n81738 , n81739 , n81740 , n81741 , n81742 , n81743 , n81744 , n81745 , n81746 , n81747 , n81748 , n81749 , n81750 , n81751 , n81752 , n81753 , n81754 , n81755 , n81756 , n81757 , n81758 , n81759 , n81760 , n81761 , n81762 , n81763 , n81764 , n81765 , n81766 , n81767 , n81768 , n81769 , n81770 , n81771 , n81772 , n81773 , n81774 , n81775 , n81776 , n81777 , n81778 , n81779 , n81780 , n81781 , n81782 , n81783 , n81784 , n81785 , n81786 , n81787 , n81788 , n81789 , n81790 , n81791 , n81792 , n81793 , n81794 , n81795 , n81796 , n81797 , n81798 , n81799 , n81800 , n81801 , n81802 , n81803 , n81804 , n81805 , n81806 , n81807 , n81808 , n81809 , n81810 , n81811 , n81812 , n81813 , n81814 , n81815 , n81816 , n81817 , n81818 , n81819 , n81820 , n81821 , n81822 , n81823 , n81824 , n81825 , n81826 , n81827 , n81828 , n81829 , n81830 , n81831 , n81832 , n81833 , n81834 , n81835 , n81836 , n81837 , n81838 , n81839 , n81840 , n81841 , n81842 , n81843 , n81844 , n81845 , n81846 , n81847 , n81848 , n81849 , n81850 , n81851 , n81852 , n81853 , n81854 , n81855 , n81856 , n81857 , n81858 , n81859 , n81860 , n81861 , n81862 , n81863 , n81864 , n81865 , n81866 , n81867 , n81868 , n81869 , n81870 , n81871 , n81872 , n81873 , n81874 , n81875 , n81876 , n81877 , n81878 , n81879 , n81880 , n81881 , n81882 , n81883 , n81884 , n81885 , n81886 , n81887 , n81888 , n81889 , n81890 , n81891 , n81892 , n81893 , n81894 , n81895 , n81896 , n81897 , n81898 , n81899 , n81900 , n81901 , n81902 , n81903 , n81904 , n81905 , n81906 , n81907 , n81908 , n81909 , n81910 , n81911 , n81912 , n81913 , n81914 , n81915 , n81916 , n81917 , n81918 , n81919 , n81920 , n81921 , n81922 , n81923 , n81924 , n81925 , n81926 , n81927 , n81928 , n81929 , n81930 , n81931 , n81932 , n81933 , n81934 , n81935 , n81936 , n81937 , n81938 , n81939 , n81940 , n81941 , n81942 , n81943 , n81944 , n81945 , n81946 , n81947 , n81948 , n81949 , n81950 , n81951 , n81952 , n81953 , n81954 , n81955 , n81956 , n81957 , n81958 , n81959 , n81960 , n81961 , n81962 , n81963 , n81964 , n81965 , n81966 , n81967 , n81968 , n81969 , n81970 , n81971 , n81972 , n81973 , n81974 , n81975 , n81976 , n81977 , n81978 , n81979 , n81980 , n81981 , n81982 , n81983 , n81984 , n81985 , n81986 , n81987 , n81988 , n81989 , n81990 , n81991 , n81992 , n81993 , n81994 , n81995 , n81996 , n81997 , n81998 , n81999 , n82000 , n82001 , n82002 , n82003 , n82004 , n82005 , n82006 , n82007 , n82008 , n82009 , n82010 , n82011 , n82012 , n82013 , n82014 , n82015 , n82016 , n82017 , n82018 , n82019 , n82020 , n82021 , n82022 , n82023 , n82024 , n82025 , n82026 , n82027 , n82028 , n82029 , n82030 , n82031 , n82032 , n82033 , n82034 , n82035 , n82036 , n82037 , n82038 , n82039 , n82040 , n82041 , n82042 , n82043 , n82044 , n82045 , n82046 , n82047 , n82048 , n82049 , n82050 , n82051 , n82052 , n82053 , n82054 , n82055 , n82056 , n82057 , n82058 , n82059 , n82060 , n82061 , n82062 , n82063 , n82064 , n82065 , n82066 , n82067 , n82068 , n82069 , n82070 , n82071 , n82072 , n82073 , n82074 , n82075 , n82076 , n82077 , n82078 , n82079 , n82080 , n82081 , n82082 , n82083 , n82084 , n82085 , n82086 , n82087 , n82088 , n82089 , n82090 , n82091 , n82092 , n82093 , n82094 , n82095 , n82096 , n82097 , n82098 , n82099 , n82100 , n82101 , n82102 , n82103 , n82104 , n82105 , n82106 , n82107 , n82108 , n82109 , n82110 , n82111 , n82112 , n82113 , n82114 , n82115 , n82116 , n82117 , n82118 , n82119 , n82120 , n82121 , n82122 , n82123 , n82124 , n82125 , n82126 , n82127 , n82128 , n82129 , n82130 , n82131 , n82132 , n82133 , n82134 , n82135 , n82136 , n82137 , n82138 , n82139 , n82140 , n82141 , n82142 , n82143 , n82144 , n82145 , n82146 , n82147 , n82148 , n82149 , n82150 , n82151 , n82152 , n82153 , n82154 , n82155 , n82156 , n82157 , n82158 , n82159 , n82160 , n82161 , n82162 , n82163 , n82164 , n82165 , n82166 , n82167 , n82168 , n82169 , n82170 , n82171 , n82172 , n82173 , n82174 , n82175 , n82176 , n82177 , n82178 , n82179 , n82180 , n82181 , n82182 , n82183 , n82184 , n82185 , n82186 , n82187 , n82188 , n82189 , n82190 , n82191 , n82192 , n82193 , n82194 , n82195 , n82196 , n82197 , n82198 , n82199 , n82200 , n82201 , n82202 , n82203 , n82204 , n82205 , n82206 , n82207 , n82208 , n82209 , n82210 , n82211 , n82212 , n82213 , n82214 , n82215 , n82216 , n82217 , n82218 , n82219 , n82220 , n82221 , n82222 , n82223 , n82224 , n82225 , n82226 , n82227 , n82228 , n82229 , n82230 , n82231 , n82232 , n82233 , n82234 , n82235 , n82236 , n82237 , n82238 , n82239 , n82240 , n82241 , n82242 , n82243 , n82244 , n82245 , n82246 , n82247 , n82248 , n82249 , n82250 , n82251 , n82252 , n82253 , n82254 , n82255 , n82256 , n82257 , n82258 , n82259 , n82260 , n82261 , n82262 , n82263 , n82264 , n82265 , n82266 , n82267 , n82268 , n82269 , n82270 , n82271 , n82272 , n82273 , n82274 , n82275 , n82276 , n82277 , n82278 , n82279 , n82280 , n82281 , n82282 , n82283 , n82284 , n82285 , n82286 , n82287 , n82288 , n82289 , n82290 , n82291 , n82292 , n82293 , n82294 , n82295 , n82296 , n82297 , n82298 , n82299 , n82300 , n82301 , n82302 , n82303 , n82304 , n82305 , n82306 , n82307 , n82308 , n82309 , n82310 , n82311 , n82312 , n82313 , n82314 , n82315 , n82316 , n82317 , n82318 , n82319 , n82320 , n82321 , n82322 , n82323 , n82324 , n82325 , n82326 , n82327 , n82328 , n82329 , n82330 , n82331 , n82332 , n82333 , n82334 , n82335 , n82336 , n82337 , n82338 , n82339 , n82340 , n82341 , n82342 , n82343 , n82344 , n82345 , n82346 , n82347 , n82348 , n82349 , n82350 , n82351 , n82352 , n82353 , n82354 , n82355 , n82356 , n82357 , n82358 , n82359 , n82360 , n82361 , n82362 , n82363 , n82364 , n82365 , n82366 , n82367 , n82368 , n82369 , n82370 , n82371 , n82372 , n82373 , n82374 , n82375 , n82376 , n82377 , n82378 , n82379 , n82380 , n82381 , n82382 , n82383 , n82384 , n82385 , n82386 , n82387 , n82388 , n82389 , n82390 , n82391 , n82392 , n82393 , n82394 , n82395 , n82396 , n82397 , n82398 , n82399 , n82400 , n82401 , n82402 , n82403 , n82404 , n82405 , n82406 , n82407 , n82408 , n82409 , n82410 , n82411 , n82412 , n82413 , n82414 , n82415 , n82416 , n82417 , n82418 , n82419 , n82420 , n82421 , n82422 , n82423 , n82424 , n82425 , n82426 , n82427 , n82428 , n82429 , n82430 , n82431 , n82432 , n82433 , n82434 , n82435 , n82436 , n82437 , n82438 , n82439 , n82440 , n82441 , n82442 , n82443 , n82444 , n82445 , n82446 , n82447 , n82448 , n82449 , n82450 , n82451 , n82452 , n82453 , n82454 , n82455 , n82456 , n82457 , n82458 , n82459 , n82460 , n82461 , n82462 , n82463 , n82464 , n82465 , n82466 , n82467 , n82468 , n82469 , n82470 , n82471 , n82472 , n82473 , n82474 , n82475 , n82476 , n82477 , n82478 , n82479 , n82480 , n82481 , n82482 , n82483 , n82484 , n82485 , n82486 , n82487 , n82488 , n82489 , n82490 , n82491 , n82492 , n82493 , n82494 , n82495 , n82496 , n82497 , n82498 , n82499 , n82500 , n82501 , n82502 , n82503 , n82504 , n82505 , n82506 , n82507 , n82508 , n82509 , n82510 , n82511 , n82512 , n82513 , n82514 , n82515 , n82516 , n82517 , n82518 , n82519 , n82520 , n82521 , n82522 , n82523 , n82524 , n82525 , n82526 , n82527 , n82528 , n82529 , n82530 , n82531 , n82532 , n82533 , n82534 , n82535 , n82536 , n82537 , n82538 , n82539 , n82540 , n82541 , n82542 , n82543 , n82544 , n82545 , n82546 , n82547 , n82548 , n82549 , n82550 , n82551 , n82552 , n82553 , n82554 , n82555 , n82556 , n82557 , n82558 , n82559 , n82560 , n82561 , n82562 , n82563 , n82564 , n82565 , n82566 , n82567 , n82568 , n82569 , n82570 , n82571 , n82572 , n82573 , n82574 , n82575 , n82576 , n82577 , n82578 , n82579 , n82580 , n82581 , n82582 , n82583 , n82584 , n82585 , n82586 , n82587 , n82588 , n82589 , n82590 , n82591 , n82592 , n82593 , n82594 , n82595 , n82596 , n82597 , n82598 , n82599 , n82600 , n82601 , n82602 , n82603 , n82604 , n82605 , n82606 , n82607 , n82608 , n82609 , n82610 , n82611 , n82612 , n82613 , n82614 , n82615 , n82616 , n82617 , n82618 , n82619 , n82620 , n82621 , n82622 , n82623 , n82624 , n82625 , n82626 , n82627 , n82628 , n82629 , n82630 , n82631 , n82632 , n82633 , n82634 , n82635 , n82636 , n82637 , n82638 , n82639 , n82640 , n82641 , n82642 , n82643 , n82644 , n82645 , n82646 , n82647 , n82648 , n82649 , n82650 , n82651 , n82652 , n82653 , n82654 , n82655 , n82656 , n82657 , n82658 , n82659 , n82660 , n82661 , n82662 , n82663 , n82664 , n82665 , n82666 , n82667 , n82668 , n82669 , n82670 , n82671 , n82672 , n82673 , n82674 , n82675 , n82676 , n82677 , n82678 , n82679 , n82680 , n82681 , n82682 , n82683 , n82684 , n82685 , n82686 , n82687 , n82688 , n82689 , n82690 , n82691 , n82692 , n82693 , n82694 , n82695 , n82696 , n82697 , n82698 , n82699 , n82700 , n82701 , n82702 , n82703 , n82704 , n82705 , n82706 , n82707 , n82708 , n82709 , n82710 , n82711 , n82712 , n82713 , n82714 , n82715 , n82716 , n82717 , n82718 , n82719 , n82720 , n82721 , n82722 , n82723 , n82724 , n82725 , n82726 , n82727 , n82728 , n82729 , n82730 , n82731 , n82732 , n82733 , n82734 , n82735 , n82736 , n82737 , n82738 , n82739 , n82740 , n82741 , n82742 , n82743 , n82744 , n82745 , n82746 , n82747 , n82748 , n82749 , n82750 , n82751 , n82752 , n82753 , n82754 , n82755 , n82756 , n82757 , n82758 , n82759 , n82760 , n82761 , n82762 , n82763 , n82764 , n82765 , n82766 , n82767 , n82768 , n82769 , n82770 , n82771 , n82772 , n82773 , n82774 , n82775 , n82776 , n82777 , n82778 , n82779 , n82780 , n82781 , n82782 , n82783 , n82784 , n82785 , n82786 , n82787 , n82788 , n82789 , n82790 , n82791 , n82792 , n82793 , n82794 , n82795 , n82796 , n82797 , n82798 , n82799 , n82800 , n82801 , n82802 , n82803 , n82804 , n82805 , n82806 , n82807 , n82808 , n82809 , n82810 , n82811 , n82812 , n82813 , n82814 , n82815 , n82816 , n82817 , n82818 , n82819 , n82820 , n82821 , n82822 , n82823 , n82824 , n82825 , n82826 , n82827 , n82828 , n82829 , n82830 , n82831 , n82832 , n82833 , n82834 , n82835 , n82836 , n82837 , n82838 , n82839 , n82840 , n82841 , n82842 , n82843 , n82844 , n82845 , n82846 , n82847 , n82848 , n82849 , n82850 , n82851 , n82852 , n82853 , n82854 , n82855 , n82856 , n82857 , n82858 , n82859 , n82860 , n82861 , n82862 , n82863 , n82864 , n82865 , n82866 , n82867 , n82868 , n82869 , n82870 , n82871 , n82872 , n82873 , n82874 , n82875 , n82876 , n82877 , n82878 , n82879 , n82880 , n82881 , n82882 , n82883 , n82884 , n82885 , n82886 , n82887 , n82888 , n82889 , n82890 , n82891 , n82892 , n82893 , n82894 , n82895 , n82896 , n82897 , n82898 , n82899 , n82900 , n82901 , n82902 , n82903 , n82904 , n82905 , n82906 , n82907 , n82908 , n82909 , n82910 , n82911 , n82912 , n82913 , n82914 , n82915 , n82916 , n82917 , n82918 , n82919 , n82920 , n82921 , n82922 , n82923 , n82924 , n82925 , n82926 , n82927 , n82928 , n82929 , n82930 , n82931 , n82932 , n82933 , n82934 , n82935 , n82936 , n82937 , n82938 , n82939 , n82940 , n82941 , n82942 , n82943 , n82944 , n82945 , n82946 , n82947 , n82948 , n82949 , n82950 , n82951 , n82952 , n82953 , n82954 , n82955 , n82956 , n82957 , n82958 , n82959 , n82960 , n82961 , n82962 , n82963 , n82964 , n82965 , n82966 , n82967 , n82968 , n82969 , n82970 , n82971 , n82972 , n82973 , n82974 , n82975 , n82976 , n82977 , n82978 , n82979 , n82980 , n82981 , n82982 , n82983 , n82984 , n82985 , n82986 , n82987 , n82988 , n82989 , n82990 , n82991 , n82992 , n82993 , n82994 , n82995 , n82996 , n82997 , n82998 , n82999 , n83000 , n83001 , n83002 , n83003 , n83004 , n83005 , n83006 , n83007 , n83008 , n83009 , n83010 , n83011 , n83012 , n83013 , n83014 , n83015 , n83016 , n83017 , n83018 , n83019 , n83020 , n83021 , n83022 , n83023 , n83024 , n83025 , n83026 , n83027 , n83028 , n83029 , n83030 , n83031 , n83032 , n83033 , n83034 , n83035 , n83036 , n83037 , n83038 , n83039 , n83040 , n83041 , n83042 , n83043 , n83044 , n83045 , n83046 , n83047 , n83048 , n83049 , n83050 , n83051 , n83052 , n83053 , n83054 , n83055 , n83056 , n83057 , n83058 , n83059 , n83060 , n83061 , n83062 , n83063 , n83064 , n83065 , n83066 , n83067 , n83068 , n83069 , n83070 , n83071 , n83072 , n83073 , n83074 , n83075 , n83076 , n83077 , n83078 , n83079 , n83080 , n83081 , n83082 , n83083 , n83084 , n83085 , n83086 , n83087 , n83088 , n83089 , n83090 , n83091 , n83092 , n83093 , n83094 , n83095 , n83096 , n83097 , n83098 , n83099 , n83100 , n83101 , n83102 , n83103 , n83104 , n83105 , n83106 , n83107 , n83108 , n83109 , n83110 , n83111 , n83112 , n83113 , n83114 , n83115 , n83116 , n83117 , n83118 , n83119 , n83120 , n83121 , n83122 , n83123 , n83124 , n83125 , n83126 , n83127 , n83128 , n83129 , n83130 , n83131 , n83132 , n83133 , n83134 , n83135 , n83136 , n83137 , n83138 , n83139 , n83140 , n83141 , n83142 , n83143 , n83144 , n83145 , n83146 , n83147 , n83148 , n83149 , n83150 , n83151 , n83152 , n83153 , n83154 , n83155 , n83156 , n83157 , n83158 , n83159 , n83160 , n83161 , n83162 , n83163 , n83164 , n83165 , n83166 , n83167 , n83168 , n83169 , n83170 , n83171 , n83172 , n83173 , n83174 , n83175 , n83176 , n83177 , n83178 , n83179 , n83180 , n83181 , n83182 , n83183 , n83184 , n83185 , n83186 , n83187 , n83188 , n83189 , n83190 , n83191 , n83192 , n83193 , n83194 , n83195 , n83196 , n83197 , n83198 , n83199 , n83200 , n83201 , n83202 , n83203 , n83204 , n83205 , n83206 , n83207 , n83208 , n83209 , n83210 , n83211 , n83212 , n83213 , n83214 , n83215 , n83216 , n83217 , n83218 , n83219 , n83220 , n83221 , n83222 , n83223 , n83224 , n83225 , n83226 , n83227 , n83228 , n83229 , n83230 , n83231 , n83232 , n83233 , n83234 , n83235 , n83236 , n83237 , n83238 , n83239 , n83240 , n83241 , n83242 , n83243 , n83244 , n83245 , n83246 , n83247 , n83248 , n83249 , n83250 , n83251 , n83252 , n83253 , n83254 , n83255 , n83256 , n83257 , n83258 , n83259 , n83260 , n83261 , n83262 , n83263 , n83264 , n83265 , n83266 , n83267 , n83268 , n83269 , n83270 , n83271 , n83272 , n83273 , n83274 , n83275 , n83276 , n83277 , n83278 , n83279 , n83280 , n83281 , n83282 , n83283 , n83284 , n83285 , n83286 , n83287 , n83288 , n83289 , n83290 , n83291 , n83292 , n83293 , n83294 , n83295 , n83296 , n83297 , n83298 , n83299 , n83300 , n83301 , n83302 , n83303 , n83304 , n83305 , n83306 , n83307 , n83308 , n83309 , n83310 , n83311 , n83312 , n83313 , n83314 , n83315 , n83316 , n83317 , n83318 , n83319 , n83320 , n83321 , n83322 , n83323 , n83324 , n83325 , n83326 , n83327 , n83328 , n83329 , n83330 , n83331 , n83332 , n83333 , n83334 , n83335 , n83336 , n83337 , n83338 , n83339 , n83340 , n83341 , n83342 , n83343 , n83344 , n83345 , n83346 , n83347 , n83348 , n83349 , n83350 , n83351 , n83352 , n83353 , n83354 , n83355 , n83356 , n83357 , n83358 , n83359 , n83360 , n83361 , n83362 , n83363 , n83364 , n83365 , n83366 , n83367 , n83368 , n83369 , n83370 , n83371 , n83372 , n83373 , n83374 , n83375 , n83376 , n83377 , n83378 , n83379 , n83380 , n83381 , n83382 , n83383 , n83384 , n83385 , n83386 , n83387 , n83388 , n83389 , n83390 , n83391 , n83392 , n83393 , n83394 , n83395 , n83396 , n83397 , n83398 , n83399 , n83400 , n83401 , n83402 , n83403 , n83404 , n83405 , n83406 , n83407 , n83408 , n83409 , n83410 , n83411 , n83412 , n83413 , n83414 , n83415 , n83416 , n83417 , n83418 , n83419 , n83420 , n83421 , n83422 , n83423 , n83424 , n83425 , n83426 , n83427 , n83428 , n83429 , n83430 , n83431 , n83432 , n83433 , n83434 , n83435 , n83436 , n83437 , n83438 , n83439 , n83440 , n83441 , n83442 , n83443 , n83444 , n83445 , n83446 , n83447 , n83448 , n83449 , n83450 , n83451 , n83452 , n83453 , n83454 , n83455 , n83456 , n83457 , n83458 , n83459 , n83460 , n83461 , n83462 , n83463 , n83464 , n83465 , n83466 , n83467 , n83468 , n83469 , n83470 , n83471 , n83472 , n83473 , n83474 , n83475 , n83476 , n83477 , n83478 , n83479 , n83480 , n83481 , n83482 , n83483 , n83484 , n83485 , n83486 , n83487 , n83488 , n83489 , n83490 , n83491 , n83492 , n83493 , n83494 , n83495 , n83496 , n83497 , n83498 , n83499 , n83500 , n83501 , n83502 , n83503 , n83504 , n83505 , n83506 , n83507 , n83508 , n83509 , n83510 , n83511 , n83512 , n83513 , n83514 , n83515 , n83516 , n83517 , n83518 , n83519 , n83520 , n83521 , n83522 , n83523 , n83524 , n83525 , n83526 , n83527 , n83528 , n83529 , n83530 , n83531 , n83532 , n83533 , n83534 , n83535 , n83536 , n83537 , n83538 , n83539 , n83540 , n83541 , n83542 , n83543 , n83544 , n83545 , n83546 , n83547 , n83548 , n83549 , n83550 , n83551 , n83552 , n83553 , n83554 , n83555 , n83556 , n83557 , n83558 , n83559 , n83560 , n83561 , n83562 , n83563 , n83564 , n83565 , n83566 , n83567 , n83568 , n83569 , n83570 , n83571 , n83572 , n83573 , n83574 , n83575 , n83576 , n83577 , n83578 , n83579 , n83580 , n83581 , n83582 , n83583 , n83584 , n83585 , n83586 , n83587 , n83588 , n83589 , n83590 , n83591 , n83592 , n83593 , n83594 , n83595 , n83596 , n83597 , n83598 , n83599 , n83600 , n83601 , n83602 , n83603 , n83604 , n83605 , n83606 , n83607 , n83608 , n83609 , n83610 , n83611 , n83612 , n83613 , n83614 , n83615 , n83616 , n83617 , n83618 , n83619 , n83620 , n83621 , n83622 , n83623 , n83624 , n83625 , n83626 , n83627 , n83628 , n83629 , n83630 , n83631 , n83632 , n83633 , n83634 , n83635 , n83636 , n83637 , n83638 , n83639 , n83640 , n83641 , n83642 , n83643 , n83644 , n83645 , n83646 , n83647 , n83648 , n83649 , n83650 , n83651 , n83652 , n83653 , n83654 , n83655 , n83656 , n83657 , n83658 , n83659 , n83660 , n83661 , n83662 , n83663 , n83664 , n83665 , n83666 , n83667 , n83668 , n83669 , n83670 , n83671 , n83672 , n83673 , n83674 , n83675 , n83676 , n83677 , n83678 , n83679 , n83680 , n83681 , n83682 , n83683 , n83684 , n83685 , n83686 , n83687 , n83688 , n83689 , n83690 , n83691 , n83692 , n83693 , n83694 , n83695 , n83696 , n83697 , n83698 , n83699 , n83700 , n83701 , n83702 , n83703 , n83704 , n83705 , n83706 , n83707 , n83708 , n83709 , n83710 , n83711 , n83712 , n83713 , n83714 , n83715 , n83716 , n83717 , n83718 , n83719 , n83720 , n83721 , n83722 , n83723 , n83724 , n83725 , n83726 , n83727 , n83728 , n83729 , n83730 , n83731 , n83732 , n83733 , n83734 , n83735 , n83736 , n83737 , n83738 , n83739 , n83740 , n83741 , n83742 , n83743 , n83744 , n83745 , n83746 , n83747 , n83748 , n83749 , n83750 , n83751 , n83752 , n83753 , n83754 , n83755 , n83756 , n83757 , n83758 , n83759 , n83760 , n83761 , n83762 , n83763 , n83764 , n83765 , n83766 , n83767 , n83768 , n83769 , n83770 , n83771 , n83772 , n83773 , n83774 , n83775 , n83776 , n83777 , n83778 , n83779 , n83780 , n83781 , n83782 , n83783 , n83784 , n83785 , n83786 , n83787 , n83788 , n83789 , n83790 , n83791 , n83792 , n83793 , n83794 , n83795 , n83796 , n83797 , n83798 , n83799 , n83800 , n83801 , n83802 , n83803 , n83804 , n83805 , n83806 , n83807 , n83808 , n83809 , n83810 , n83811 , n83812 , n83813 , n83814 , n83815 , n83816 , n83817 , n83818 , n83819 , n83820 , n83821 , n83822 , n83823 , n83824 , n83825 , n83826 , n83827 , n83828 , n83829 , n83830 , n83831 , n83832 , n83833 , n83834 , n83835 , n83836 , n83837 , n83838 , n83839 , n83840 , n83841 , n83842 , n83843 , n83844 , n83845 , n83846 , n83847 , n83848 , n83849 , n83850 , n83851 , n83852 , n83853 , n83854 , n83855 , n83856 , n83857 , n83858 , n83859 , n83860 , n83861 , n83862 , n83863 , n83864 , n83865 , n83866 , n83867 , n83868 , n83869 , n83870 , n83871 , n83872 , n83873 , n83874 , n83875 , n83876 , n83877 , n83878 , n83879 , n83880 , n83881 , n83882 , n83883 , n83884 , n83885 , n83886 , n83887 , n83888 , n83889 , n83890 , n83891 , n83892 , n83893 , n83894 , n83895 , n83896 , n83897 , n83898 , n83899 , n83900 , n83901 , n83902 , n83903 , n83904 , n83905 , n83906 , n83907 , n83908 , n83909 , n83910 , n83911 , n83912 , n83913 , n83914 , n83915 , n83916 , n83917 , n83918 , n83919 , n83920 , n83921 , n83922 , n83923 , n83924 , n83925 , n83926 , n83927 , n83928 , n83929 , n83930 , n83931 , n83932 , n83933 , n83934 , n83935 , n83936 , n83937 , n83938 , n83939 , n83940 , n83941 , n83942 , n83943 , n83944 , n83945 , n83946 , n83947 , n83948 , n83949 , n83950 , n83951 , n83952 , n83953 , n83954 , n83955 , n83956 , n83957 , n83958 , n83959 , n83960 , n83961 , n83962 , n83963 , n83964 , n83965 , n83966 , n83967 , n83968 , n83969 , n83970 , n83971 , n83972 , n83973 , n83974 , n83975 , n83976 , n83977 , n83978 , n83979 , n83980 , n83981 , n83982 , n83983 , n83984 , n83985 , n83986 , n83987 , n83988 , n83989 , n83990 , n83991 , n83992 , n83993 , n83994 , n83995 , n83996 , n83997 , n83998 , n83999 , n84000 , n84001 , n84002 , n84003 , n84004 , n84005 , n84006 , n84007 , n84008 , n84009 , n84010 , n84011 , n84012 , n84013 , n84014 , n84015 , n84016 , n84017 , n84018 , n84019 , n84020 , n84021 , n84022 , n84023 , n84024 , n84025 , n84026 , n84027 , n84028 , n84029 , n84030 , n84031 , n84032 , n84033 , n84034 , n84035 , n84036 , n84037 , n84038 , n84039 , n84040 , n84041 , n84042 , n84043 , n84044 , n84045 , n84046 , n84047 , n84048 , n84049 , n84050 , n84051 , n84052 , n84053 , n84054 , n84055 , n84056 , n84057 , n84058 , n84059 , n84060 , n84061 , n84062 , n84063 , n84064 , n84065 , n84066 , n84067 , n84068 , n84069 , n84070 , n84071 , n84072 , n84073 , n84074 , n84075 , n84076 , n84077 , n84078 , n84079 , n84080 , n84081 , n84082 , n84083 , n84084 , n84085 , n84086 , n84087 , n84088 , n84089 , n84090 , n84091 , n84092 , n84093 , n84094 , n84095 , n84096 , n84097 , n84098 , n84099 , n84100 , n84101 , n84102 , n84103 , n84104 , n84105 , n84106 , n84107 , n84108 , n84109 , n84110 , n84111 , n84112 , n84113 , n84114 , n84115 , n84116 , n84117 , n84118 , n84119 , n84120 , n84121 , n84122 , n84123 , n84124 , n84125 , n84126 , n84127 , n84128 , n84129 , n84130 , n84131 , n84132 , n84133 , n84134 , n84135 , n84136 , n84137 , n84138 , n84139 , n84140 , n84141 , n84142 , n84143 , n84144 , n84145 , n84146 , n84147 , n84148 , n84149 , n84150 , n84151 , n84152 , n84153 , n84154 , n84155 , n84156 , n84157 , n84158 , n84159 , n84160 , n84161 , n84162 , n84163 , n84164 , n84165 , n84166 , n84167 , n84168 , n84169 , n84170 , n84171 , n84172 , n84173 , n84174 , n84175 , n84176 , n84177 , n84178 , n84179 , n84180 , n84181 , n84182 , n84183 , n84184 , n84185 , n84186 , n84187 , n84188 , n84189 , n84190 , n84191 , n84192 , n84193 , n84194 , n84195 , n84196 , n84197 , n84198 , n84199 , n84200 , n84201 , n84202 , n84203 , n84204 , n84205 , n84206 , n84207 , n84208 , n84209 , n84210 , n84211 , n84212 , n84213 , n84214 , n84215 , n84216 , n84217 , n84218 , n84219 , n84220 , n84221 , n84222 , n84223 , n84224 , n84225 , n84226 , n84227 , n84228 , n84229 , n84230 , n84231 , n84232 , n84233 , n84234 , n84235 , n84236 , n84237 , n84238 , n84239 , n84240 , n84241 , n84242 , n84243 , n84244 , n84245 , n84246 , n84247 , n84248 , n84249 , n84250 , n84251 , n84252 , n84253 , n84254 , n84255 , n84256 , n84257 , n84258 , n84259 , n84260 , n84261 , n84262 , n84263 , n84264 , n84265 , n84266 , n84267 , n84268 , n84269 , n84270 , n84271 , n84272 , n84273 , n84274 , n84275 , n84276 , n84277 , n84278 , n84279 , n84280 , n84281 , n84282 , n84283 , n84284 , n84285 , n84286 , n84287 , n84288 , n84289 , n84290 , n84291 , n84292 , n84293 , n84294 , n84295 , n84296 , n84297 , n84298 , n84299 , n84300 , n84301 , n84302 , n84303 , n84304 , n84305 , n84306 , n84307 , n84308 , n84309 , n84310 , n84311 , n84312 , n84313 , n84314 , n84315 , n84316 , n84317 , n84318 , n84319 , n84320 , n84321 , n84322 , n84323 , n84324 , n84325 , n84326 , n84327 , n84328 , n84329 , n84330 , n84331 , n84332 , n84333 , n84334 , n84335 , n84336 , n84337 , n84338 , n84339 , n84340 , n84341 , n84342 , n84343 , n84344 , n84345 , n84346 , n84347 , n84348 , n84349 , n84350 , n84351 , n84352 , n84353 , n84354 , n84355 , n84356 , n84357 , n84358 , n84359 , n84360 , n84361 , n84362 , n84363 , n84364 , n84365 , n84366 , n84367 , n84368 , n84369 , n84370 , n84371 , n84372 , n84373 , n84374 , n84375 , n84376 , n84377 , n84378 , n84379 , n84380 , n84381 , n84382 , n84383 , n84384 , n84385 , n84386 , n84387 , n84388 , n84389 , n84390 , n84391 , n84392 , n84393 , n84394 , n84395 , n84396 , n84397 , n84398 , n84399 , n84400 , n84401 , n84402 , n84403 , n84404 , n84405 , n84406 , n84407 , n84408 , n84409 , n84410 , n84411 , n84412 , n84413 , n84414 , n84415 , n84416 , n84417 , n84418 , n84419 , n84420 , n84421 , n84422 , n84423 , n84424 , n84425 , n84426 , n84427 , n84428 , n84429 , n84430 , n84431 , n84432 , n84433 , n84434 , n84435 , n84436 , n84437 , n84438 , n84439 , n84440 , n84441 , n84442 , n84443 , n84444 , n84445 , n84446 , n84447 , n84448 , n84449 , n84450 , n84451 , n84452 , n84453 , n84454 , n84455 , n84456 , n84457 , n84458 , n84459 , n84460 , n84461 , n84462 , n84463 , n84464 , n84465 , n84466 , n84467 , n84468 , n84469 , n84470 , n84471 , n84472 , n84473 , n84474 , n84475 , n84476 , n84477 , n84478 , n84479 , n84480 , n84481 , n84482 , n84483 , n84484 , n84485 , n84486 , n84487 , n84488 , n84489 , n84490 , n84491 , n84492 , n84493 , n84494 , n84495 , n84496 , n84497 , n84498 , n84499 , n84500 , n84501 , n84502 , n84503 , n84504 , n84505 , n84506 , n84507 , n84508 , n84509 , n84510 , n84511 , n84512 , n84513 , n84514 , n84515 , n84516 , n84517 , n84518 , n84519 , n84520 , n84521 , n84522 , n84523 , n84524 , n84525 , n84526 , n84527 , n84528 , n84529 , n84530 , n84531 , n84532 , n84533 , n84534 , n84535 , n84536 , n84537 , n84538 , n84539 , n84540 , n84541 , n84542 , n84543 , n84544 , n84545 , n84546 , n84547 , n84548 , n84549 , n84550 , n84551 , n84552 , n84553 , n84554 , n84555 , n84556 , n84557 , n84558 , n84559 , n84560 , n84561 , n84562 , n84563 , n84564 , n84565 , n84566 , n84567 , n84568 , n84569 , n84570 , n84571 , n84572 , n84573 , n84574 , n84575 , n84576 , n84577 , n84578 , n84579 , n84580 , n84581 , n84582 , n84583 , n84584 , n84585 , n84586 , n84587 , n84588 , n84589 , n84590 , n84591 , n84592 , n84593 , n84594 , n84595 , n84596 , n84597 , n84598 , n84599 , n84600 , n84601 , n84602 , n84603 , n84604 , n84605 , n84606 , n84607 , n84608 , n84609 , n84610 , n84611 , n84612 , n84613 , n84614 , n84615 , n84616 , n84617 , n84618 , n84619 , n84620 , n84621 , n84622 , n84623 , n84624 , n84625 , n84626 , n84627 , n84628 , n84629 , n84630 , n84631 , n84632 , n84633 , n84634 , n84635 , n84636 , n84637 , n84638 , n84639 , n84640 , n84641 , n84642 , n84643 , n84644 , n84645 , n84646 , n84647 , n84648 , n84649 , n84650 , n84651 , n84652 , n84653 , n84654 , n84655 , n84656 , n84657 , n84658 , n84659 , n84660 , n84661 , n84662 , n84663 , n84664 , n84665 , n84666 , n84667 , n84668 , n84669 , n84670 , n84671 , n84672 , n84673 , n84674 , n84675 , n84676 , n84677 , n84678 , n84679 , n84680 , n84681 , n84682 , n84683 , n84684 , n84685 , n84686 , n84687 , n84688 , n84689 , n84690 , n84691 , n84692 , n84693 , n84694 , n84695 , n84696 , n84697 , n84698 , n84699 , n84700 , n84701 , n84702 , n84703 , n84704 , n84705 , n84706 , n84707 , n84708 , n84709 , n84710 , n84711 , n84712 , n84713 , n84714 , n84715 , n84716 , n84717 , n84718 , n84719 , n84720 , n84721 , n84722 , n84723 , n84724 , n84725 , n84726 , n84727 , n84728 , n84729 , n84730 , n84731 , n84732 , n84733 , n84734 , n84735 , n84736 , n84737 , n84738 , n84739 , n84740 , n84741 , n84742 , n84743 , n84744 , n84745 , n84746 , n84747 , n84748 , n84749 , n84750 , n84751 , n84752 , n84753 , n84754 , n84755 , n84756 , n84757 , n84758 , n84759 , n84760 , n84761 , n84762 , n84763 , n84764 , n84765 , n84766 , n84767 , n84768 , n84769 , n84770 , n84771 , n84772 , n84773 , n84774 , n84775 , n84776 , n84777 , n84778 , n84779 , n84780 , n84781 , n84782 , n84783 , n84784 , n84785 , n84786 , n84787 , n84788 , n84789 , n84790 , n84791 , n84792 , n84793 , n84794 , n84795 , n84796 , n84797 , n84798 , n84799 , n84800 , n84801 , n84802 , n84803 , n84804 , n84805 , n84806 , n84807 , n84808 , n84809 , n84810 , n84811 , n84812 , n84813 , n84814 , n84815 , n84816 , n84817 , n84818 , n84819 , n84820 , n84821 , n84822 , n84823 , n84824 , n84825 , n84826 , n84827 , n84828 , n84829 , n84830 , n84831 , n84832 , n84833 , n84834 , n84835 , n84836 , n84837 , n84838 , n84839 , n84840 , n84841 , n84842 , n84843 , n84844 , n84845 , n84846 , n84847 , n84848 , n84849 , n84850 , n84851 , n84852 , n84853 , n84854 , n84855 , n84856 , n84857 , n84858 , n84859 , n84860 , n84861 , n84862 , n84863 , n84864 , n84865 , n84866 , n84867 , n84868 , n84869 , n84870 , n84871 , n84872 , n84873 , n84874 , n84875 , n84876 , n84877 , n84878 , n84879 , n84880 , n84881 , n84882 , n84883 , n84884 , n84885 , n84886 , n84887 , n84888 , n84889 , n84890 , n84891 , n84892 , n84893 , n84894 , n84895 , n84896 , n84897 , n84898 , n84899 , n84900 , n84901 , n84902 , n84903 , n84904 , n84905 , n84906 , n84907 , n84908 , n84909 , n84910 , n84911 , n84912 , n84913 , n84914 , n84915 , n84916 , n84917 , n84918 , n84919 , n84920 , n84921 , n84922 , n84923 , n84924 , n84925 , n84926 , n84927 , n84928 , n84929 , n84930 , n84931 , n84932 , n84933 , n84934 , n84935 , n84936 , n84937 , n84938 , n84939 , n84940 , n84941 , n84942 , n84943 , n84944 , n84945 , n84946 , n84947 , n84948 , n84949 , n84950 , n84951 , n84952 , n84953 , n84954 , n84955 , n84956 , n84957 , n84958 , n84959 , n84960 , n84961 , n84962 , n84963 , n84964 , n84965 , n84966 , n84967 , n84968 , n84969 , n84970 , n84971 , n84972 , n84973 , n84974 , n84975 , n84976 , n84977 , n84978 , n84979 , n84980 , n84981 , n84982 , n84983 , n84984 , n84985 , n84986 , n84987 , n84988 , n84989 , n84990 , n84991 , n84992 , n84993 , n84994 , n84995 , n84996 , n84997 , n84998 , n84999 , n85000 , n85001 , n85002 , n85003 , n85004 , n85005 , n85006 , n85007 , n85008 , n85009 , n85010 , n85011 , n85012 , n85013 , n85014 , n85015 , n85016 , n85017 , n85018 , n85019 , n85020 , n85021 , n85022 , n85023 , n85024 , n85025 , n85026 , n85027 , n85028 , n85029 , n85030 , n85031 , n85032 , n85033 , n85034 , n85035 , n85036 , n85037 , n85038 , n85039 , n85040 , n85041 , n85042 , n85043 , n85044 , n85045 , n85046 , n85047 , n85048 , n85049 , n85050 , n85051 , n85052 , n85053 , n85054 , n85055 , n85056 , n85057 , n85058 , n85059 , n85060 , n85061 , n85062 , n85063 , n85064 , n85065 , n85066 , n85067 , n85068 , n85069 , n85070 , n85071 , n85072 , n85073 , n85074 , n85075 , n85076 , n85077 , n85078 , n85079 , n85080 , n85081 , n85082 , n85083 , n85084 , n85085 , n85086 , n85087 , n85088 , n85089 , n85090 , n85091 , n85092 , n85093 , n85094 , n85095 , n85096 , n85097 , n85098 , n85099 , n85100 , n85101 , n85102 , n85103 , n85104 , n85105 , n85106 , n85107 , n85108 , n85109 , n85110 , n85111 , n85112 , n85113 , n85114 , n85115 , n85116 , n85117 , n85118 , n85119 , n85120 , n85121 , n85122 , n85123 , n85124 , n85125 , n85126 , n85127 , n85128 , n85129 , n85130 , n85131 , n85132 , n85133 , n85134 , n85135 , n85136 , n85137 , n85138 , n85139 , n85140 , n85141 , n85142 , n85143 , n85144 , n85145 , n85146 , n85147 , n85148 , n85149 , n85150 , n85151 , n85152 , n85153 , n85154 , n85155 , n85156 , n85157 , n85158 , n85159 , n85160 , n85161 , n85162 , n85163 , n85164 , n85165 , n85166 , n85167 , n85168 , n85169 , n85170 , n85171 , n85172 , n85173 , n85174 , n85175 , n85176 , n85177 , n85178 , n85179 , n85180 , n85181 , n85182 , n85183 , n85184 , n85185 , n85186 , n85187 , n85188 , n85189 , n85190 , n85191 , n85192 , n85193 , n85194 , n85195 , n85196 , n85197 , n85198 , n85199 , n85200 , n85201 , n85202 , n85203 , n85204 , n85205 , n85206 , n85207 , n85208 , n85209 , n85210 , n85211 , n85212 , n85213 , n85214 , n85215 , n85216 , n85217 , n85218 , n85219 , n85220 , n85221 , n85222 , n85223 , n85224 , n85225 , n85226 , n85227 , n85228 , n85229 , n85230 , n85231 , n85232 , n85233 , n85234 , n85235 , n85236 , n85237 , n85238 , n85239 , n85240 , n85241 , n85242 , n85243 , n85244 , n85245 , n85246 , n85247 , n85248 , n85249 , n85250 , n85251 , n85252 , n85253 , n85254 , n85255 , n85256 , n85257 , n85258 , n85259 , n85260 , n85261 , n85262 , n85263 , n85264 , n85265 , n85266 , n85267 , n85268 , n85269 , n85270 , n85271 , n85272 , n85273 , n85274 , n85275 , n85276 , n85277 , n85278 , n85279 , n85280 , n85281 , n85282 , n85283 , n85284 , n85285 , n85286 , n85287 , n85288 , n85289 , n85290 , n85291 , n85292 , n85293 , n85294 , n85295 , n85296 , n85297 , n85298 , n85299 , n85300 , n85301 , n85302 , n85303 , n85304 , n85305 , n85306 , n85307 , n85308 , n85309 , n85310 , n85311 , n85312 , n85313 , n85314 , n85315 , n85316 , n85317 , n85318 , n85319 , n85320 , n85321 , n85322 , n85323 , n85324 , n85325 , n85326 , n85327 , n85328 , n85329 , n85330 , n85331 , n85332 , n85333 , n85334 , n85335 , n85336 , n85337 , n85338 , n85339 , n85340 , n85341 , n85342 , n85343 , n85344 , n85345 , n85346 , n85347 , n85348 , n85349 , n85350 , n85351 , n85352 , n85353 , n85354 , n85355 , n85356 , n85357 , n85358 , n85359 , n85360 , n85361 , n85362 , n85363 , n85364 , n85365 , n85366 , n85367 , n85368 , n85369 , n85370 , n85371 , n85372 , n85373 , n85374 , n85375 , n85376 , n85377 , n85378 , n85379 , n85380 , n85381 , n85382 , n85383 , n85384 , n85385 , n85386 , n85387 , n85388 , n85389 , n85390 , n85391 , n85392 , n85393 , n85394 , n85395 , n85396 , n85397 , n85398 , n85399 , n85400 , n85401 , n85402 , n85403 , n85404 , n85405 , n85406 , n85407 , n85408 , n85409 , n85410 , n85411 , n85412 , n85413 , n85414 , n85415 , n85416 , n85417 , n85418 , n85419 , n85420 , n85421 , n85422 , n85423 , n85424 , n85425 , n85426 , n85427 , n85428 , n85429 , n85430 , n85431 , n85432 , n85433 , n85434 , n85435 , n85436 , n85437 , n85438 , n85439 , n85440 , n85441 , n85442 , n85443 , n85444 , n85445 , n85446 , n85447 , n85448 , n85449 , n85450 , n85451 , n85452 , n85453 , n85454 , n85455 , n85456 , n85457 , n85458 , n85459 , n85460 , n85461 , n85462 , n85463 , n85464 , n85465 , n85466 , n85467 , n85468 , n85469 , n85470 , n85471 , n85472 , n85473 , n85474 , n85475 , n85476 , n85477 , n85478 , n85479 , n85480 , n85481 , n85482 , n85483 , n85484 , n85485 , n85486 , n85487 , n85488 , n85489 , n85490 , n85491 , n85492 , n85493 , n85494 , n85495 , n85496 , n85497 , n85498 , n85499 , n85500 , n85501 , n85502 , n85503 , n85504 , n85505 , n85506 , n85507 , n85508 , n85509 , n85510 , n85511 , n85512 , n85513 , n85514 , n85515 , n85516 , n85517 , n85518 , n85519 , n85520 , n85521 , n85522 , n85523 , n85524 , n85525 , n85526 , n85527 , n85528 , n85529 , n85530 , n85531 , n85532 , n85533 , n85534 , n85535 , n85536 , n85537 , n85538 , n85539 , n85540 , n85541 , n85542 , n85543 , n85544 , n85545 , n85546 , n85547 , n85548 , n85549 , n85550 , n85551 , n85552 , n85553 , n85554 , n85555 , n85556 , n85557 , n85558 , n85559 , n85560 , n85561 , n85562 , n85563 , n85564 , n85565 , n85566 , n85567 , n85568 , n85569 , n85570 , n85571 , n85572 , n85573 , n85574 , n85575 , n85576 , n85577 , n85578 , n85579 , n85580 , n85581 , n85582 , n85583 , n85584 , n85585 , n85586 , n85587 , n85588 , n85589 , n85590 , n85591 , n85592 , n85593 , n85594 , n85595 , n85596 , n85597 , n85598 , n85599 , n85600 , n85601 , n85602 , n85603 , n85604 , n85605 , n85606 , n85607 , n85608 , n85609 , n85610 , n85611 , n85612 , n85613 , n85614 , n85615 , n85616 , n85617 , n85618 , n85619 , n85620 , n85621 , n85622 , n85623 , n85624 , n85625 , n85626 , n85627 , n85628 , n85629 , n85630 , n85631 , n85632 , n85633 , n85634 , n85635 , n85636 , n85637 , n85638 , n85639 , n85640 , n85641 , n85642 , n85643 , n85644 , n85645 , n85646 , n85647 , n85648 , n85649 , n85650 , n85651 , n85652 , n85653 , n85654 , n85655 , n85656 , n85657 , n85658 , n85659 , n85660 , n85661 , n85662 , n85663 , n85664 , n85665 , n85666 , n85667 , n85668 , n85669 , n85670 , n85671 , n85672 , n85673 , n85674 , n85675 , n85676 , n85677 , n85678 , n85679 , n85680 , n85681 , n85682 , n85683 , n85684 , n85685 , n85686 , n85687 , n85688 , n85689 , n85690 , n85691 , n85692 , n85693 , n85694 , n85695 , n85696 , n85697 , n85698 , n85699 , n85700 , n85701 , n85702 , n85703 , n85704 , n85705 , n85706 , n85707 , n85708 , n85709 , n85710 , n85711 , n85712 , n85713 , n85714 , n85715 , n85716 , n85717 , n85718 , n85719 , n85720 , n85721 , n85722 , n85723 , n85724 , n85725 , n85726 , n85727 , n85728 , n85729 , n85730 , n85731 , n85732 , n85733 , n85734 , n85735 , n85736 , n85737 , n85738 , n85739 , n85740 , n85741 , n85742 , n85743 , n85744 , n85745 , n85746 , n85747 , n85748 , n85749 , n85750 , n85751 , n85752 , n85753 , n85754 , n85755 , n85756 , n85757 , n85758 , n85759 , n85760 , n85761 , n85762 , n85763 , n85764 , n85765 , n85766 , n85767 , n85768 , n85769 , n85770 , n85771 , n85772 , n85773 , n85774 , n85775 , n85776 , n85777 , n85778 , n85779 , n85780 , n85781 , n85782 , n85783 , n85784 , n85785 , n85786 , n85787 , n85788 , n85789 , n85790 , n85791 , n85792 , n85793 , n85794 , n85795 , n85796 , n85797 , n85798 , n85799 , n85800 , n85801 , n85802 , n85803 , n85804 , n85805 , n85806 , n85807 , n85808 , n85809 , n85810 , n85811 , n85812 , n85813 , n85814 , n85815 , n85816 , n85817 , n85818 , n85819 , n85820 , n85821 , n85822 , n85823 , n85824 , n85825 , n85826 , n85827 , n85828 , n85829 , n85830 , n85831 , n85832 , n85833 , n85834 , n85835 , n85836 , n85837 , n85838 , n85839 , n85840 , n85841 , n85842 , n85843 , n85844 , n85845 , n85846 , n85847 , n85848 , n85849 , n85850 , n85851 , n85852 , n85853 , n85854 , n85855 , n85856 , n85857 , n85858 , n85859 , n85860 , n85861 , n85862 , n85863 , n85864 , n85865 , n85866 , n85867 , n85868 , n85869 , n85870 , n85871 , n85872 , n85873 , n85874 , n85875 , n85876 , n85877 , n85878 , n85879 , n85880 , n85881 , n85882 , n85883 , n85884 , n85885 , n85886 , n85887 , n85888 , n85889 , n85890 , n85891 , n85892 , n85893 , n85894 , n85895 , n85896 , n85897 , n85898 , n85899 , n85900 , n85901 , n85902 , n85903 , n85904 , n85905 , n85906 , n85907 , n85908 , n85909 , n85910 , n85911 , n85912 , n85913 , n85914 , n85915 , n85916 , n85917 , n85918 , n85919 , n85920 , n85921 , n85922 , n85923 , n85924 , n85925 , n85926 , n85927 , n85928 , n85929 , n85930 , n85931 , n85932 , n85933 , n85934 , n85935 , n85936 , n85937 , n85938 , n85939 , n85940 , n85941 , n85942 , n85943 , n85944 , n85945 , n85946 , n85947 , n85948 , n85949 , n85950 , n85951 , n85952 , n85953 , n85954 , n85955 , n85956 , n85957 , n85958 , n85959 , n85960 , n85961 , n85962 , n85963 , n85964 , n85965 , n85966 , n85967 , n85968 , n85969 , n85970 , n85971 , n85972 , n85973 , n85974 , n85975 , n85976 , n85977 , n85978 , n85979 , n85980 , n85981 , n85982 , n85983 , n85984 , n85985 , n85986 , n85987 , n85988 , n85989 , n85990 , n85991 , n85992 , n85993 , n85994 , n85995 , n85996 , n85997 , n85998 , n85999 , n86000 , n86001 , n86002 , n86003 , n86004 , n86005 , n86006 , n86007 , n86008 , n86009 , n86010 , n86011 , n86012 , n86013 , n86014 , n86015 , n86016 , n86017 , n86018 , n86019 , n86020 , n86021 , n86022 , n86023 , n86024 , n86025 , n86026 , n86027 , n86028 , n86029 , n86030 , n86031 , n86032 , n86033 , n86034 , n86035 , n86036 , n86037 , n86038 , n86039 , n86040 , n86041 , n86042 , n86043 , n86044 , n86045 , n86046 , n86047 , n86048 , n86049 , n86050 , n86051 , n86052 , n86053 , n86054 , n86055 , n86056 , n86057 , n86058 , n86059 , n86060 , n86061 , n86062 , n86063 , n86064 , n86065 , n86066 , n86067 , n86068 , n86069 , n86070 , n86071 , n86072 , n86073 , n86074 , n86075 , n86076 , n86077 , n86078 , n86079 , n86080 , n86081 , n86082 , n86083 , n86084 , n86085 , n86086 , n86087 , n86088 , n86089 , n86090 , n86091 , n86092 , n86093 , n86094 , n86095 , n86096 , n86097 , n86098 , n86099 , n86100 , n86101 , n86102 , n86103 , n86104 , n86105 , n86106 , n86107 , n86108 , n86109 , n86110 , n86111 , n86112 , n86113 , n86114 , n86115 , n86116 , n86117 , n86118 , n86119 , n86120 , n86121 , n86122 , n86123 , n86124 , n86125 , n86126 , n86127 , n86128 , n86129 , n86130 , n86131 , n86132 , n86133 , n86134 , n86135 , n86136 , n86137 , n86138 , n86139 , n86140 , n86141 , n86142 , n86143 , n86144 , n86145 , n86146 , n86147 , n86148 , n86149 , n86150 , n86151 , n86152 , n86153 , n86154 , n86155 , n86156 , n86157 , n86158 , n86159 , n86160 , n86161 , n86162 , n86163 , n86164 , n86165 , n86166 , n86167 , n86168 , n86169 , n86170 , n86171 , n86172 , n86173 , n86174 , n86175 , n86176 , n86177 , n86178 , n86179 , n86180 , n86181 , n86182 , n86183 , n86184 , n86185 , n86186 , n86187 , n86188 , n86189 , n86190 , n86191 , n86192 , n86193 , n86194 , n86195 , n86196 , n86197 , n86198 , n86199 , n86200 , n86201 , n86202 , n86203 , n86204 , n86205 , n86206 , n86207 , n86208 , n86209 , n86210 , n86211 , n86212 , n86213 , n86214 , n86215 , n86216 , n86217 , n86218 , n86219 , n86220 , n86221 , n86222 , n86223 , n86224 , n86225 , n86226 , n86227 , n86228 , n86229 , n86230 , n86231 , n86232 , n86233 , n86234 , n86235 , n86236 , n86237 , n86238 , n86239 , n86240 , n86241 , n86242 , n86243 , n86244 , n86245 , n86246 , n86247 , n86248 , n86249 , n86250 , n86251 , n86252 , n86253 , n86254 , n86255 , n86256 , n86257 , n86258 , n86259 , n86260 , n86261 , n86262 , n86263 , n86264 , n86265 , n86266 , n86267 , n86268 , n86269 , n86270 , n86271 , n86272 , n86273 , n86274 , n86275 , n86276 , n86277 , n86278 , n86279 , n86280 , n86281 , n86282 , n86283 , n86284 , n86285 , n86286 , n86287 , n86288 , n86289 , n86290 , n86291 , n86292 , n86293 , n86294 , n86295 , n86296 , n86297 , n86298 , n86299 , n86300 , n86301 , n86302 , n86303 , n86304 , n86305 , n86306 , n86307 , n86308 , n86309 , n86310 , n86311 , n86312 , n86313 , n86314 , n86315 , n86316 , n86317 , n86318 , n86319 , n86320 , n86321 , n86322 , n86323 , n86324 , n86325 , n86326 , n86327 , n86328 , n86329 , n86330 , n86331 , n86332 , n86333 , n86334 , n86335 , n86336 , n86337 , n86338 , n86339 , n86340 , n86341 , n86342 , n86343 , n86344 , n86345 , n86346 , n86347 , n86348 , n86349 , n86350 , n86351 , n86352 , n86353 , n86354 , n86355 , n86356 , n86357 , n86358 , n86359 , n86360 , n86361 , n86362 , n86363 , n86364 , n86365 , n86366 , n86367 , n86368 , n86369 , n86370 , n86371 , n86372 , n86373 , n86374 , n86375 , n86376 , n86377 , n86378 , n86379 , n86380 , n86381 , n86382 , n86383 , n86384 , n86385 , n86386 , n86387 , n86388 , n86389 , n86390 , n86391 , n86392 , n86393 , n86394 , n86395 , n86396 , n86397 , n86398 , n86399 , n86400 , n86401 , n86402 , n86403 , n86404 , n86405 , n86406 , n86407 , n86408 , n86409 , n86410 , n86411 , n86412 , n86413 , n86414 , n86415 , n86416 , n86417 , n86418 , n86419 , n86420 , n86421 , n86422 , n86423 , n86424 , n86425 , n86426 , n86427 , n86428 , n86429 , n86430 , n86431 , n86432 , n86433 , n86434 , n86435 , n86436 , n86437 , n86438 , n86439 , n86440 , n86441 , n86442 , n86443 , n86444 , n86445 , n86446 , n86447 , n86448 , n86449 , n86450 , n86451 , n86452 , n86453 , n86454 , n86455 , n86456 , n86457 , n86458 , n86459 , n86460 , n86461 , n86462 , n86463 , n86464 , n86465 , n86466 , n86467 , n86468 , n86469 , n86470 , n86471 , n86472 , n86473 , n86474 , n86475 , n86476 , n86477 , n86478 , n86479 , n86480 , n86481 , n86482 , n86483 , n86484 , n86485 , n86486 , n86487 , n86488 ;
  assign n65362 = x126 | x127 ;
  assign n65354 = x124 | x125 ;
  assign n65369 = n65354 | n65362 ;
  assign n65384 = x122 | x123 ;
  assign n27311 = n65369 | n65384 ;
  assign n65377 = x120 | x121 ;
  assign n65392 = n65377 | n65384 ;
  assign n66655 = n65369 | n65392 ;
  assign n65399 = x116 | x117 ;
  assign n65407 = x118 | x119 ;
  assign n65414 = n65399 | n65407 ;
  assign n65422 = n65392 | n65414 ;
  assign n65429 = n65369 | n65422 ;
  assign n65497 = x114 | x115 ;
  assign n20357 = n65414 | n65497 ;
  assign n20358 = n66655 | n20357 ;
  assign n65489 = x112 | x113 ;
  assign n65504 = n65489 | n65497 ;
  assign n65519 = x110 | x111 ;
  assign n17323 = n65504 | n65519 ;
  assign n17324 = n65429 | n17323 ;
  assign n65512 = x108 | x109 ;
  assign n65527 = n65512 | n65519 ;
  assign n65534 = n65504 | n65527 ;
  assign n15856 = n65429 | n65534 ;
  assign n65437 = x104 | x105 ;
  assign n65444 = x106 | x107 ;
  assign n65452 = n65437 | n65444 ;
  assign n65467 = x102 | x103 ;
  assign n11927 = n65452 | n65467 ;
  assign n11928 = n65534 | n11927 ;
  assign n11929 = n65429 | n11928 ;
  assign n273 = x125 | x126 ;
  assign n274 = x127 | n273 ;
  assign n266 = x117 | x118 ;
  assign n267 = x119 | x120 ;
  assign n268 = n266 | n267 ;
  assign n275 = x121 | x122 ;
  assign n276 = x123 | x124 ;
  assign n277 = n275 | n276 ;
  assign n464 = n268 | n277 ;
  assign n465 = n274 | n464 ;
  assign n280 = x101 | x102 ;
  assign n281 = x103 | x104 ;
  assign n282 = n280 | n281 ;
  assign n290 = x105 | x106 ;
  assign n291 = x107 | x108 ;
  assign n292 = n290 | n291 ;
  assign n466 = n282 | n292 ;
  assign n269 = x113 | x114 ;
  assign n270 = x115 | x116 ;
  assign n271 = n269 | n270 ;
  assign n287 = x109 | x110 ;
  assign n288 = x111 | x112 ;
  assign n289 = n287 | n288 ;
  assign n467 = n271 | n289 ;
  assign n468 = n466 | n467 ;
  assign n469 = n465 | n468 ;
  assign n66559 = n65414 | n65504 ;
  assign n66858 = n66559 | n66655 ;
  assign n65459 = x100 | x101 ;
  assign n65474 = n65459 | n65467 ;
  assign n65602 = x96 | x97 ;
  assign n65609 = x98 | x99 ;
  assign n65617 = n65602 | n65609 ;
  assign n66865 = n65474 | n65617 ;
  assign n67093 = n65452 | n65527 ;
  assign n67215 = n66865 | n67093 ;
  assign n303 = n66858 | n67215 ;
  assign n65557 = x90 | x91 ;
  assign n65624 = x92 | x93 ;
  assign n65632 = x94 | x95 ;
  assign n65639 = n65624 | n65632 ;
  assign n5741 = n65557 | n65639 ;
  assign n5742 = n67215 | n5741 ;
  assign n5743 = n66858 | n5742 ;
  assign n65482 = n65452 | n65474 ;
  assign n65542 = n65482 | n65534 ;
  assign n65549 = x88 | x89 ;
  assign n65564 = n65549 | n65557 ;
  assign n65572 = x84 | x85 ;
  assign n65579 = x86 | x87 ;
  assign n65587 = n65572 | n65579 ;
  assign n65594 = n65564 | n65587 ;
  assign n65647 = n65617 | n65639 ;
  assign n65654 = n65594 | n65647 ;
  assign n65662 = n65542 | n65654 ;
  assign n65666 = n65429 | n65662 ;
  assign n380 = n65429 | n65542 ;
  assign n65287 = x80 | x81 ;
  assign n65294 = x82 | x83 ;
  assign n65302 = n65287 | n65294 ;
  assign n65317 = x78 | x79 ;
  assign n1837 = n65302 | n65317 ;
  assign n1838 = n65654 | n1837 ;
  assign n1839 = n380 | n1838 ;
  assign n65235 = x72 | x73 ;
  assign n65243 = x74 | x75 ;
  assign n65249 = n65235 | n65243 ;
  assign n65309 = x76 | x77 ;
  assign n65324 = n65309 | n65317 ;
  assign n66296 = n65249 | n65324 ;
  assign n67221 = n65302 | n65587 ;
  assign n67349 = n65564 | n65639 ;
  assign n67612 = n67221 | n67349 ;
  assign n767 = n66296 | n67612 ;
  assign n768 = n303 | n767 ;
  assign n65667 = ~x62 ;
  assign n65702 = n65667 & x64 ;
  assign n65790 = x65 & n65702 ;
  assign n65668 = ~n65790 ;
  assign n65821 = x63 & n65668 ;
  assign n65669 = ~x63 ;
  assign n65199 = n65669 & x64 ;
  assign n65670 = ~x65 ;
  assign n65206 = x64 & n65670 ;
  assign n65214 = x66 | x67 ;
  assign n65671 = ~n65214 ;
  assign n65221 = n65206 & n65671 ;
  assign n65672 = ~n65199 ;
  assign n65229 = n65672 & n65221 ;
  assign n65257 = x68 | x69 ;
  assign n65264 = x70 | x71 ;
  assign n65272 = n65257 | n65264 ;
  assign n65279 = n65249 | n65272 ;
  assign n65332 = n65302 | n65324 ;
  assign n65339 = n65279 | n65332 ;
  assign n65673 = ~n65339 ;
  assign n65347 = n65229 & n65673 ;
  assign n65674 = ~n65666 ;
  assign n65900 = n65347 & n65674 ;
  assign n65675 = ~n65900 ;
  assign n65906 = n65821 & n65675 ;
  assign n66008 = x65 | n65702 ;
  assign n65676 = ~n65906 ;
  assign n66070 = n65676 & n66008 ;
  assign n66146 = x63 & n65675 ;
  assign n66080 = n65668 & n66008 ;
  assign n66289 = n65214 | n65272 ;
  assign n66453 = n66289 | n66296 ;
  assign n65677 = ~n66453 ;
  assign n66549 = n66080 & n65677 ;
  assign n67619 = n67215 | n67612 ;
  assign n67897 = n66858 | n67619 ;
  assign n65678 = ~n67897 ;
  assign n68051 = n66549 & n65678 ;
  assign n65679 = ~n66146 ;
  assign n68057 = n65679 & n68051 ;
  assign n65680 = ~n66070 ;
  assign n68215 = n65680 & n68057 ;
  assign n68535 = n66296 | n67221 ;
  assign n68542 = n66289 | n68535 ;
  assign n65681 = ~n66655 ;
  assign n68886 = n66080 & n65681 ;
  assign n69068 = n66559 | n67093 ;
  assign n69074 = n66865 | n67349 ;
  assign n69262 = n69068 | n69074 ;
  assign n65682 = ~n69262 ;
  assign n69646 = n68886 & n65682 ;
  assign n65683 = ~n68542 ;
  assign n69653 = n65683 & n69646 ;
  assign n70051 = n65680 & n69653 ;
  assign n65684 = ~n70051 ;
  assign n70265 = n66146 & n65684 ;
  assign n70273 = n68215 | n70265 ;
  assign n65685 = ~x61 ;
  assign n70710 = n65685 & x64 ;
  assign n307 = x65 | n70710 ;
  assign n71396 = x65 & n70710 ;
  assign n71403 = x85 | x86 ;
  assign n71642 = x87 | x88 ;
  assign n72130 = n71403 | n71642 ;
  assign n72138 = x81 | x82 ;
  assign n72392 = x83 | x84 ;
  assign n72910 = n72138 | n72392 ;
  assign n72917 = n72130 | n72910 ;
  assign n73185 = x93 | x94 ;
  assign n73737 = x95 | x96 ;
  assign n73745 = n73185 | n73737 ;
  assign n74028 = x89 | x90 ;
  assign n74608 = x91 | x92 ;
  assign n74615 = n74028 | n74608 ;
  assign n74914 = n73745 | n74615 ;
  assign n75217 = n72917 | n74914 ;
  assign n75525 = x69 | x70 ;
  assign n75838 = x71 | x72 ;
  assign n86484 = n75525 | n75838 ;
  assign n65686 = ~x66 ;
  assign n86485 = x64 & n65686 ;
  assign n86486 = x67 | x68 ;
  assign n65687 = ~n86486 ;
  assign n86487 = n86485 & n65687 ;
  assign n65688 = ~n86484 ;
  assign n86488 = n65688 & n86487 ;
  assign n257 = x77 | x78 ;
  assign n258 = x79 | x80 ;
  assign n259 = n257 | n258 ;
  assign n260 = x73 | x74 ;
  assign n261 = x75 | x76 ;
  assign n262 = n260 | n261 ;
  assign n263 = n259 | n262 ;
  assign n65689 = ~n263 ;
  assign n264 = n86488 & n65689 ;
  assign n65690 = ~n75217 ;
  assign n265 = n65690 & n264 ;
  assign n272 = n268 | n271 ;
  assign n278 = n274 | n277 ;
  assign n279 = n272 | n278 ;
  assign n283 = x97 | x98 ;
  assign n284 = x99 | x100 ;
  assign n285 = n283 | n284 ;
  assign n286 = n282 | n285 ;
  assign n293 = n289 | n292 ;
  assign n294 = n286 | n293 ;
  assign n295 = n279 | n294 ;
  assign n65691 = ~n295 ;
  assign n296 = n265 & n65691 ;
  assign n297 = n65680 & n296 ;
  assign n65692 = ~n297 ;
  assign n298 = x62 & n65692 ;
  assign n299 = n65671 & n65702 ;
  assign n65693 = ~n65272 ;
  assign n300 = n65693 & n299 ;
  assign n65694 = ~n66296 ;
  assign n301 = n65694 & n300 ;
  assign n65695 = ~n67612 ;
  assign n302 = n65695 & n301 ;
  assign n65696 = ~n303 ;
  assign n304 = n302 & n65696 ;
  assign n305 = n65680 & n304 ;
  assign n306 = n298 | n305 ;
  assign n65697 = ~n71396 ;
  assign n308 = n65697 & n306 ;
  assign n65698 = ~n308 ;
  assign n309 = n307 & n65698 ;
  assign n70702 = n65686 & n70273 ;
  assign n65699 = ~n68215 ;
  assign n310 = x66 & n65699 ;
  assign n65700 = ~n70265 ;
  assign n311 = n65700 & n310 ;
  assign n313 = n70702 | n311 ;
  assign n314 = n309 & n313 ;
  assign n315 = x66 | n314 ;
  assign n312 = n309 | n311 ;
  assign n65701 = ~n70702 ;
  assign n316 = n65701 & n312 ;
  assign n317 = n86484 | n86486 ;
  assign n318 = n263 | n317 ;
  assign n319 = n75217 | n318 ;
  assign n320 = n295 | n319 ;
  assign n321 = n316 | n320 ;
  assign n190 = ~n321 ;
  assign n322 = n315 & n190 ;
  assign n65703 = ~n322 ;
  assign n323 = n70273 & n65703 ;
  assign n65704 = ~n320 ;
  assign n324 = n312 & n65704 ;
  assign n65705 = ~n314 ;
  assign n325 = n65705 & n324 ;
  assign n65706 = ~n316 ;
  assign n326 = n65706 & n325 ;
  assign n65707 = ~n326 ;
  assign n327 = x67 & n65707 ;
  assign n65708 = ~n323 ;
  assign n328 = n65708 & n327 ;
  assign n329 = n72917 | n263 ;
  assign n330 = n317 | n329 ;
  assign n331 = n65697 & n307 ;
  assign n65709 = ~n278 ;
  assign n332 = n65709 & n331 ;
  assign n333 = n272 | n293 ;
  assign n334 = n74914 | n286 ;
  assign n335 = n333 | n334 ;
  assign n65710 = ~n335 ;
  assign n336 = n332 & n65710 ;
  assign n65711 = ~n330 ;
  assign n337 = n65711 & n336 ;
  assign n338 = n65706 & n337 ;
  assign n65712 = ~n338 ;
  assign n339 = n306 & n65712 ;
  assign n70934 = n65670 & n70710 ;
  assign n65713 = ~n70710 ;
  assign n340 = x65 & n65713 ;
  assign n341 = n70934 | n340 ;
  assign n65714 = ~n318 ;
  assign n342 = n65714 & n341 ;
  assign n343 = n75217 | n294 ;
  assign n344 = n279 | n343 ;
  assign n65715 = ~n344 ;
  assign n345 = n342 & n65715 ;
  assign n65716 = ~n305 ;
  assign n346 = n65716 & n345 ;
  assign n65717 = ~n298 ;
  assign n347 = n65717 & n346 ;
  assign n348 = n65706 & n347 ;
  assign n349 = n339 | n348 ;
  assign n350 = n65686 & n349 ;
  assign n65718 = ~n348 ;
  assign n351 = x66 & n65718 ;
  assign n65719 = ~n339 ;
  assign n352 = n65719 & n351 ;
  assign n65720 = ~x60 ;
  assign n366 = n65720 & x64 ;
  assign n368 = x65 & n366 ;
  assign n65721 = ~x67 ;
  assign n353 = x64 & n65721 ;
  assign n354 = n65693 & n353 ;
  assign n355 = n65694 & n354 ;
  assign n356 = n65695 & n355 ;
  assign n357 = n65696 & n356 ;
  assign n358 = n65706 & n357 ;
  assign n65722 = ~n358 ;
  assign n359 = x61 & n65722 ;
  assign n360 = n70710 & n65687 ;
  assign n361 = n65688 & n360 ;
  assign n362 = n65689 & n361 ;
  assign n363 = n65690 & n362 ;
  assign n364 = n65691 & n363 ;
  assign n365 = n65706 & n364 ;
  assign n369 = n359 | n365 ;
  assign n65723 = ~n368 ;
  assign n370 = n65723 & n369 ;
  assign n371 = x65 | n366 ;
  assign n65724 = ~n370 ;
  assign n372 = n65724 & n371 ;
  assign n373 = n352 | n372 ;
  assign n65725 = ~n350 ;
  assign n374 = n65725 & n373 ;
  assign n375 = n328 | n374 ;
  assign n376 = n323 | n326 ;
  assign n377 = n65721 & n376 ;
  assign n65726 = ~n377 ;
  assign n378 = n375 & n65726 ;
  assign n383 = n350 | n352 ;
  assign n384 = n372 & n383 ;
  assign n379 = n65339 | n65654 ;
  assign n381 = n379 | n380 ;
  assign n65727 = ~n381 ;
  assign n386 = n373 & n65727 ;
  assign n65728 = ~n384 ;
  assign n387 = n65728 & n386 ;
  assign n65729 = ~n378 ;
  assign n388 = n65729 & n387 ;
  assign n385 = x66 | n384 ;
  assign n389 = n65727 & n385 ;
  assign n390 = n65729 & n389 ;
  assign n65730 = ~n390 ;
  assign n391 = n349 & n65730 ;
  assign n392 = n388 | n391 ;
  assign n393 = n328 | n377 ;
  assign n394 = n374 | n393 ;
  assign n395 = n374 & n393 ;
  assign n396 = n381 | n395 ;
  assign n65731 = ~n396 ;
  assign n397 = n394 & n65731 ;
  assign n398 = n65729 & n397 ;
  assign n382 = n378 | n381 ;
  assign n399 = n376 & n382 ;
  assign n65732 = ~n399 ;
  assign n400 = x68 & n65732 ;
  assign n65733 = ~n398 ;
  assign n401 = n65733 & n400 ;
  assign n402 = n65721 & n392 ;
  assign n65734 = ~n388 ;
  assign n403 = x67 & n65734 ;
  assign n65735 = ~n391 ;
  assign n404 = n65735 & n403 ;
  assign n405 = n65332 | n65594 ;
  assign n406 = n65279 | n405 ;
  assign n407 = n65369 | n368 ;
  assign n65736 = ~n407 ;
  assign n408 = n371 & n65736 ;
  assign n409 = n65422 | n65534 ;
  assign n410 = n65482 | n65647 ;
  assign n411 = n409 | n410 ;
  assign n65737 = ~n411 ;
  assign n412 = n408 & n65737 ;
  assign n65738 = ~n406 ;
  assign n413 = n65738 & n412 ;
  assign n414 = n65729 & n413 ;
  assign n65739 = ~n414 ;
  assign n415 = n369 & n65739 ;
  assign n367 = n65670 & n366 ;
  assign n65740 = ~n366 ;
  assign n416 = x65 & n65740 ;
  assign n417 = n367 | n416 ;
  assign n418 = n65673 & n417 ;
  assign n419 = n65674 & n418 ;
  assign n65741 = ~n365 ;
  assign n420 = n65741 & n419 ;
  assign n65742 = ~n359 ;
  assign n421 = n65742 & n420 ;
  assign n422 = n65729 & n421 ;
  assign n423 = n415 | n422 ;
  assign n424 = n65686 & n423 ;
  assign n65743 = ~n422 ;
  assign n425 = x66 & n65743 ;
  assign n65744 = ~n415 ;
  assign n426 = n65744 & n425 ;
  assign n65745 = ~x59 ;
  assign n427 = n65745 & x64 ;
  assign n429 = x65 & n427 ;
  assign n436 = n65693 & n366 ;
  assign n437 = n65694 & n436 ;
  assign n438 = n65695 & n437 ;
  assign n439 = n65696 & n438 ;
  assign n440 = n65729 & n439 ;
  assign n65746 = ~x68 ;
  assign n430 = x64 & n65746 ;
  assign n431 = n65688 & n430 ;
  assign n432 = n65689 & n431 ;
  assign n433 = n65690 & n432 ;
  assign n434 = n65691 & n433 ;
  assign n435 = n65729 & n434 ;
  assign n65747 = ~n435 ;
  assign n441 = x60 & n65747 ;
  assign n442 = n440 | n441 ;
  assign n65748 = ~n429 ;
  assign n443 = n65748 & n442 ;
  assign n444 = x65 | n427 ;
  assign n65749 = ~n443 ;
  assign n445 = n65749 & n444 ;
  assign n446 = n426 | n445 ;
  assign n65750 = ~n424 ;
  assign n447 = n65750 & n446 ;
  assign n448 = n404 | n447 ;
  assign n65751 = ~n402 ;
  assign n449 = n65751 & n448 ;
  assign n451 = n401 | n449 ;
  assign n450 = n398 | n399 ;
  assign n452 = n65746 & n450 ;
  assign n65752 = ~n452 ;
  assign n453 = n451 & n65752 ;
  assign n457 = n72130 | n74615 ;
  assign n458 = n73745 | n285 ;
  assign n459 = n457 | n458 ;
  assign n460 = n86484 | n262 ;
  assign n461 = n72910 | n259 ;
  assign n462 = n460 | n461 ;
  assign n463 = n459 | n462 ;
  assign n470 = n463 | n469 ;
  assign n454 = n402 | n404 ;
  assign n455 = n65750 & n454 ;
  assign n456 = n446 & n455 ;
  assign n472 = x67 | n456 ;
  assign n65753 = ~n470 ;
  assign n473 = n65753 & n472 ;
  assign n65754 = ~n453 ;
  assign n474 = n65754 & n473 ;
  assign n65755 = ~n474 ;
  assign n475 = n392 & n65755 ;
  assign n476 = n456 | n470 ;
  assign n65756 = ~n476 ;
  assign n477 = n448 & n65756 ;
  assign n478 = n65754 & n477 ;
  assign n479 = n475 | n478 ;
  assign n481 = x68 & n479 ;
  assign n480 = x68 | n478 ;
  assign n482 = n475 | n480 ;
  assign n65757 = ~n481 ;
  assign n483 = n65757 & n482 ;
  assign n484 = n424 | n426 ;
  assign n485 = n445 & n484 ;
  assign n487 = n446 & n65753 ;
  assign n65758 = ~n485 ;
  assign n488 = n65758 & n487 ;
  assign n489 = n65754 & n488 ;
  assign n486 = x66 | n485 ;
  assign n490 = n65753 & n486 ;
  assign n491 = n65754 & n490 ;
  assign n65759 = ~n491 ;
  assign n492 = n423 & n65759 ;
  assign n493 = n489 | n492 ;
  assign n494 = x67 & n493 ;
  assign n495 = x67 | n489 ;
  assign n496 = n492 | n495 ;
  assign n65760 = ~n494 ;
  assign n497 = n65760 & n496 ;
  assign n498 = n457 | n461 ;
  assign n499 = n460 | n498 ;
  assign n500 = n274 | n429 ;
  assign n65761 = ~n500 ;
  assign n501 = n444 & n65761 ;
  assign n502 = n464 | n467 ;
  assign n503 = n458 | n466 ;
  assign n504 = n502 | n503 ;
  assign n65762 = ~n504 ;
  assign n505 = n501 & n65762 ;
  assign n65763 = ~n499 ;
  assign n506 = n65763 & n505 ;
  assign n507 = n65754 & n506 ;
  assign n65764 = ~n507 ;
  assign n508 = n442 & n65764 ;
  assign n428 = n65670 & n427 ;
  assign n65765 = ~n427 ;
  assign n509 = x65 & n65765 ;
  assign n510 = n428 | n509 ;
  assign n65766 = ~n462 ;
  assign n511 = n65766 & n510 ;
  assign n512 = n459 | n468 ;
  assign n513 = n465 | n512 ;
  assign n65767 = ~n513 ;
  assign n514 = n511 & n65767 ;
  assign n65768 = ~n440 ;
  assign n515 = n65768 & n514 ;
  assign n65769 = ~n441 ;
  assign n516 = n65769 & n515 ;
  assign n517 = n65754 & n516 ;
  assign n518 = n508 | n517 ;
  assign n519 = n65686 & n518 ;
  assign n65770 = ~n517 ;
  assign n541 = x66 & n65770 ;
  assign n65771 = ~n508 ;
  assign n542 = n65771 & n541 ;
  assign n543 = n519 | n542 ;
  assign n65772 = ~x69 ;
  assign n520 = x64 & n65772 ;
  assign n65773 = ~n65264 ;
  assign n521 = n65773 & n520 ;
  assign n65774 = ~n65249 ;
  assign n522 = n65774 & n521 ;
  assign n65775 = ~n65332 ;
  assign n523 = n65775 & n522 ;
  assign n65776 = ~n65654 ;
  assign n524 = n65776 & n523 ;
  assign n65777 = ~n380 ;
  assign n525 = n65777 & n524 ;
  assign n526 = n65754 & n525 ;
  assign n65778 = ~n526 ;
  assign n527 = x59 & n65778 ;
  assign n528 = n65688 & n427 ;
  assign n529 = n65689 & n528 ;
  assign n530 = n65690 & n529 ;
  assign n531 = n65691 & n530 ;
  assign n532 = n65754 & n531 ;
  assign n533 = n527 | n532 ;
  assign n534 = x65 & n533 ;
  assign n535 = x65 | n532 ;
  assign n536 = n527 | n535 ;
  assign n65779 = ~n534 ;
  assign n537 = n65779 & n536 ;
  assign n65780 = ~x58 ;
  assign n538 = n65780 & x64 ;
  assign n539 = n537 | n538 ;
  assign n540 = n65670 & n533 ;
  assign n65781 = ~n540 ;
  assign n544 = n539 & n65781 ;
  assign n545 = n543 | n544 ;
  assign n65782 = ~n519 ;
  assign n546 = n65782 & n545 ;
  assign n547 = n497 | n546 ;
  assign n548 = n65721 & n493 ;
  assign n65783 = ~n548 ;
  assign n549 = n547 & n65783 ;
  assign n550 = n483 | n549 ;
  assign n551 = n65746 & n479 ;
  assign n65784 = ~n551 ;
  assign n552 = n550 & n65784 ;
  assign n567 = n65249 | n65264 ;
  assign n568 = n65332 | n567 ;
  assign n569 = n65654 | n568 ;
  assign n570 = n380 | n569 ;
  assign n553 = n401 | n452 ;
  assign n554 = n65751 & n553 ;
  assign n555 = n448 & n554 ;
  assign n556 = n470 | n555 ;
  assign n65785 = ~n556 ;
  assign n557 = n451 & n65785 ;
  assign n558 = n65754 & n557 ;
  assign n559 = x68 | n555 ;
  assign n560 = n65753 & n559 ;
  assign n561 = n65754 & n560 ;
  assign n65786 = ~n561 ;
  assign n562 = n450 & n65786 ;
  assign n563 = n558 | n562 ;
  assign n564 = x69 & n563 ;
  assign n565 = x69 | n558 ;
  assign n566 = n562 | n565 ;
  assign n65787 = ~n564 ;
  assign n571 = n65787 & n566 ;
  assign n572 = n570 | n571 ;
  assign n573 = n552 | n572 ;
  assign n574 = n65753 & n563 ;
  assign n65788 = ~n574 ;
  assign n575 = n573 & n65788 ;
  assign n579 = n552 | n571 ;
  assign n578 = n65784 & n571 ;
  assign n580 = n550 & n578 ;
  assign n65789 = ~n580 ;
  assign n581 = n579 & n65789 ;
  assign n187 = ~n575 ;
  assign n582 = n187 & n581 ;
  assign n583 = n470 & n563 ;
  assign n584 = n573 & n583 ;
  assign n585 = n582 | n584 ;
  assign n65791 = ~x70 ;
  assign n586 = n65791 & n585 ;
  assign n587 = n483 & n65783 ;
  assign n588 = n547 & n587 ;
  assign n65792 = ~n588 ;
  assign n589 = n550 & n65792 ;
  assign n590 = n187 & n589 ;
  assign n591 = n479 & n65788 ;
  assign n592 = n573 & n591 ;
  assign n593 = n590 | n592 ;
  assign n594 = n65772 & n593 ;
  assign n595 = n497 & n65782 ;
  assign n596 = n545 & n595 ;
  assign n65793 = ~n596 ;
  assign n597 = n547 & n65793 ;
  assign n598 = n187 & n597 ;
  assign n599 = n493 & n65788 ;
  assign n600 = n573 & n599 ;
  assign n601 = n598 | n600 ;
  assign n602 = n65746 & n601 ;
  assign n65794 = ~n544 ;
  assign n603 = n543 & n65794 ;
  assign n577 = n540 | n543 ;
  assign n65795 = ~n577 ;
  assign n604 = n539 & n65795 ;
  assign n605 = n603 | n604 ;
  assign n606 = n187 & n605 ;
  assign n607 = n518 & n65788 ;
  assign n608 = n573 & n607 ;
  assign n609 = n606 | n608 ;
  assign n610 = n65721 & n609 ;
  assign n611 = n536 & n538 ;
  assign n612 = n65779 & n611 ;
  assign n65796 = ~n612 ;
  assign n613 = n539 & n65796 ;
  assign n614 = n187 & n613 ;
  assign n615 = n533 & n65788 ;
  assign n616 = n573 & n615 ;
  assign n617 = n614 | n616 ;
  assign n618 = n65686 & n617 ;
  assign n576 = n538 & n187 ;
  assign n619 = x64 & n187 ;
  assign n65797 = ~n619 ;
  assign n620 = x58 & n65797 ;
  assign n621 = n576 | n620 ;
  assign n627 = n65670 & n621 ;
  assign n622 = x65 & n621 ;
  assign n623 = x65 | n576 ;
  assign n624 = n620 | n623 ;
  assign n65798 = ~n622 ;
  assign n625 = n65798 & n624 ;
  assign n65799 = ~x57 ;
  assign n626 = n65799 & x64 ;
  assign n628 = n625 | n626 ;
  assign n65800 = ~n627 ;
  assign n629 = n65800 & n628 ;
  assign n65801 = ~n616 ;
  assign n630 = x66 & n65801 ;
  assign n65802 = ~n614 ;
  assign n631 = n65802 & n630 ;
  assign n632 = n618 | n631 ;
  assign n633 = n629 | n632 ;
  assign n65803 = ~n618 ;
  assign n634 = n65803 & n633 ;
  assign n65804 = ~n608 ;
  assign n635 = x67 & n65804 ;
  assign n65805 = ~n606 ;
  assign n636 = n65805 & n635 ;
  assign n637 = n610 | n636 ;
  assign n638 = n634 | n637 ;
  assign n65806 = ~n610 ;
  assign n639 = n65806 & n638 ;
  assign n65807 = ~n600 ;
  assign n640 = x68 & n65807 ;
  assign n65808 = ~n598 ;
  assign n641 = n65808 & n640 ;
  assign n642 = n602 | n641 ;
  assign n643 = n639 | n642 ;
  assign n65809 = ~n602 ;
  assign n644 = n65809 & n643 ;
  assign n65810 = ~n592 ;
  assign n645 = x69 & n65810 ;
  assign n65811 = ~n590 ;
  assign n646 = n65811 & n645 ;
  assign n647 = n594 | n646 ;
  assign n648 = n644 | n647 ;
  assign n65812 = ~n594 ;
  assign n649 = n65812 & n648 ;
  assign n65813 = ~n584 ;
  assign n650 = x70 & n65813 ;
  assign n65814 = ~n582 ;
  assign n651 = n65814 & n650 ;
  assign n652 = n586 | n651 ;
  assign n654 = n649 | n652 ;
  assign n65815 = ~n586 ;
  assign n655 = n65815 & n654 ;
  assign n656 = n75838 | n262 ;
  assign n657 = n461 | n656 ;
  assign n658 = n459 | n657 ;
  assign n659 = n469 | n658 ;
  assign n660 = n655 | n659 ;
  assign n65816 = ~n649 ;
  assign n653 = n65816 & n652 ;
  assign n664 = n594 | n652 ;
  assign n65817 = ~n664 ;
  assign n665 = n648 & n65817 ;
  assign n666 = n653 | n665 ;
  assign n667 = n660 | n666 ;
  assign n65818 = ~n585 ;
  assign n668 = n65818 & n660 ;
  assign n65819 = ~n668 ;
  assign n669 = n667 & n65819 ;
  assign n65820 = ~x71 ;
  assign n670 = n65820 & n669 ;
  assign n186 = ~n660 ;
  assign n759 = n186 & n666 ;
  assign n760 = n585 & n660 ;
  assign n65822 = ~n760 ;
  assign n761 = x71 & n65822 ;
  assign n65823 = ~n759 ;
  assign n762 = n65823 & n761 ;
  assign n763 = n670 | n762 ;
  assign n671 = n593 & n660 ;
  assign n65824 = ~n644 ;
  assign n663 = n65824 & n647 ;
  assign n672 = n602 | n647 ;
  assign n65825 = ~n672 ;
  assign n673 = n643 & n65825 ;
  assign n674 = n663 | n673 ;
  assign n65826 = ~n659 ;
  assign n675 = n65826 & n674 ;
  assign n65827 = ~n655 ;
  assign n676 = n65827 & n675 ;
  assign n677 = n671 | n676 ;
  assign n678 = n65791 & n677 ;
  assign n679 = n601 & n660 ;
  assign n65828 = ~n639 ;
  assign n662 = n65828 & n642 ;
  assign n680 = n610 | n642 ;
  assign n65829 = ~n680 ;
  assign n681 = n638 & n65829 ;
  assign n682 = n662 | n681 ;
  assign n683 = n65826 & n682 ;
  assign n684 = n65827 & n683 ;
  assign n685 = n679 | n684 ;
  assign n686 = n65772 & n685 ;
  assign n65830 = ~n684 ;
  assign n748 = x69 & n65830 ;
  assign n65831 = ~n679 ;
  assign n749 = n65831 & n748 ;
  assign n750 = n686 | n749 ;
  assign n687 = n609 & n660 ;
  assign n65832 = ~n634 ;
  assign n661 = n65832 & n637 ;
  assign n688 = n618 | n637 ;
  assign n65833 = ~n688 ;
  assign n689 = n633 & n65833 ;
  assign n690 = n661 | n689 ;
  assign n691 = n65826 & n690 ;
  assign n692 = n65827 & n691 ;
  assign n693 = n687 | n692 ;
  assign n694 = n65746 & n693 ;
  assign n695 = n617 & n660 ;
  assign n696 = n627 | n632 ;
  assign n65834 = ~n696 ;
  assign n697 = n628 & n65834 ;
  assign n65835 = ~n629 ;
  assign n698 = n65835 & n632 ;
  assign n699 = n697 | n698 ;
  assign n700 = n65826 & n699 ;
  assign n701 = n65827 & n700 ;
  assign n702 = n695 | n701 ;
  assign n703 = n65721 & n702 ;
  assign n65836 = ~n701 ;
  assign n738 = x67 & n65836 ;
  assign n65837 = ~n695 ;
  assign n739 = n65837 & n738 ;
  assign n740 = n703 | n739 ;
  assign n704 = n621 & n660 ;
  assign n705 = n624 & n626 ;
  assign n706 = n65798 & n705 ;
  assign n707 = n659 | n706 ;
  assign n65838 = ~n707 ;
  assign n708 = n628 & n65838 ;
  assign n709 = n65827 & n708 ;
  assign n710 = n704 | n709 ;
  assign n711 = n65686 & n710 ;
  assign n65839 = ~x56 ;
  assign n729 = n65839 & x64 ;
  assign n712 = x64 & n65820 ;
  assign n713 = n65774 & n712 ;
  assign n714 = n65775 & n713 ;
  assign n715 = n65776 & n714 ;
  assign n716 = n65777 & n715 ;
  assign n717 = n65827 & n716 ;
  assign n65840 = ~n717 ;
  assign n718 = x57 & n65840 ;
  assign n65841 = ~n75838 ;
  assign n719 = n65841 & n626 ;
  assign n65842 = ~n262 ;
  assign n720 = n65842 & n719 ;
  assign n65843 = ~n461 ;
  assign n721 = n65843 & n720 ;
  assign n65844 = ~n459 ;
  assign n722 = n65844 & n721 ;
  assign n65845 = ~n469 ;
  assign n723 = n65845 & n722 ;
  assign n724 = n65827 & n723 ;
  assign n725 = n718 | n724 ;
  assign n726 = x65 & n725 ;
  assign n727 = x65 | n724 ;
  assign n728 = n718 | n727 ;
  assign n65846 = ~n726 ;
  assign n730 = n65846 & n728 ;
  assign n731 = n729 | n730 ;
  assign n732 = n65670 & n725 ;
  assign n65847 = ~n732 ;
  assign n733 = n731 & n65847 ;
  assign n65848 = ~n709 ;
  assign n734 = x66 & n65848 ;
  assign n65849 = ~n704 ;
  assign n735 = n65849 & n734 ;
  assign n736 = n711 | n735 ;
  assign n737 = n733 | n736 ;
  assign n65850 = ~n711 ;
  assign n741 = n65850 & n737 ;
  assign n742 = n740 | n741 ;
  assign n65851 = ~n703 ;
  assign n743 = n65851 & n742 ;
  assign n65852 = ~n692 ;
  assign n744 = x68 & n65852 ;
  assign n65853 = ~n687 ;
  assign n745 = n65853 & n744 ;
  assign n746 = n694 | n745 ;
  assign n747 = n743 | n746 ;
  assign n65854 = ~n694 ;
  assign n751 = n65854 & n747 ;
  assign n752 = n750 | n751 ;
  assign n65855 = ~n686 ;
  assign n753 = n65855 & n752 ;
  assign n65856 = ~n676 ;
  assign n754 = x70 & n65856 ;
  assign n65857 = ~n671 ;
  assign n755 = n65857 & n754 ;
  assign n756 = n678 | n755 ;
  assign n758 = n753 | n756 ;
  assign n65858 = ~n678 ;
  assign n764 = n65858 & n758 ;
  assign n765 = n763 | n764 ;
  assign n65859 = ~n670 ;
  assign n766 = n65859 & n765 ;
  assign n769 = n766 | n768 ;
  assign n65860 = ~n669 ;
  assign n798 = n65860 & n769 ;
  assign n65861 = ~n764 ;
  assign n874 = n763 & n65861 ;
  assign n875 = n678 | n763 ;
  assign n65862 = ~n875 ;
  assign n876 = n758 & n65862 ;
  assign n877 = n874 | n876 ;
  assign n878 = n769 | n877 ;
  assign n65863 = ~n798 ;
  assign n879 = n65863 & n878 ;
  assign n65864 = ~n768 ;
  assign n889 = n65864 & n879 ;
  assign n770 = n677 & n769 ;
  assign n757 = n686 | n756 ;
  assign n65865 = ~n757 ;
  assign n771 = n752 & n65865 ;
  assign n65866 = ~n753 ;
  assign n772 = n65866 & n756 ;
  assign n773 = n771 | n772 ;
  assign n774 = n65864 & n773 ;
  assign n65867 = ~n766 ;
  assign n775 = n65867 & n774 ;
  assign n776 = n770 | n775 ;
  assign n777 = n65820 & n776 ;
  assign n778 = n685 & n769 ;
  assign n779 = n694 | n750 ;
  assign n65868 = ~n779 ;
  assign n780 = n747 & n65868 ;
  assign n65869 = ~n751 ;
  assign n782 = n750 & n65869 ;
  assign n783 = n780 | n782 ;
  assign n784 = n65864 & n783 ;
  assign n785 = n65867 & n784 ;
  assign n786 = n778 | n785 ;
  assign n787 = n65791 & n786 ;
  assign n788 = n693 & n769 ;
  assign n789 = n703 | n746 ;
  assign n65870 = ~n789 ;
  assign n790 = n742 & n65870 ;
  assign n65871 = ~n743 ;
  assign n791 = n65871 & n746 ;
  assign n792 = n790 | n791 ;
  assign n793 = n65864 & n792 ;
  assign n794 = n65867 & n793 ;
  assign n795 = n788 | n794 ;
  assign n796 = n65772 & n795 ;
  assign n799 = n702 & n769 ;
  assign n800 = n711 | n740 ;
  assign n65872 = ~n800 ;
  assign n801 = n737 & n65872 ;
  assign n65873 = ~n741 ;
  assign n802 = n740 & n65873 ;
  assign n803 = n801 | n802 ;
  assign n804 = n65864 & n803 ;
  assign n805 = n65867 & n804 ;
  assign n806 = n799 | n805 ;
  assign n807 = n65746 & n806 ;
  assign n808 = n710 & n769 ;
  assign n65874 = ~n733 ;
  assign n809 = n65874 & n736 ;
  assign n810 = n732 | n736 ;
  assign n65875 = ~n810 ;
  assign n811 = n731 & n65875 ;
  assign n812 = n809 | n811 ;
  assign n813 = n65864 & n812 ;
  assign n814 = n65867 & n813 ;
  assign n815 = n808 | n814 ;
  assign n816 = n65721 & n815 ;
  assign n797 = n725 & n769 ;
  assign n781 = n728 & n729 ;
  assign n817 = n65846 & n781 ;
  assign n818 = n768 | n817 ;
  assign n65876 = ~n818 ;
  assign n819 = n731 & n65876 ;
  assign n820 = n65867 & n819 ;
  assign n821 = n797 | n820 ;
  assign n822 = n65686 & n821 ;
  assign n65877 = ~x72 ;
  assign n823 = x64 & n65877 ;
  assign n824 = n65842 & n823 ;
  assign n825 = n65843 & n824 ;
  assign n826 = n65844 & n825 ;
  assign n827 = n65845 & n826 ;
  assign n828 = n65867 & n827 ;
  assign n65878 = ~n828 ;
  assign n829 = x56 & n65878 ;
  assign n830 = n65774 & n729 ;
  assign n831 = n65775 & n830 ;
  assign n832 = n65776 & n831 ;
  assign n833 = n65777 & n832 ;
  assign n834 = n65867 & n833 ;
  assign n835 = n829 | n834 ;
  assign n837 = x65 & n835 ;
  assign n836 = x65 | n834 ;
  assign n838 = n829 | n836 ;
  assign n65879 = ~n837 ;
  assign n839 = n65879 & n838 ;
  assign n65880 = ~x55 ;
  assign n840 = n65880 & x64 ;
  assign n841 = n839 | n840 ;
  assign n842 = n65670 & n835 ;
  assign n65881 = ~n842 ;
  assign n843 = n841 & n65881 ;
  assign n65882 = ~n820 ;
  assign n844 = x66 & n65882 ;
  assign n65883 = ~n797 ;
  assign n845 = n65883 & n844 ;
  assign n846 = n822 | n845 ;
  assign n847 = n843 | n846 ;
  assign n65884 = ~n822 ;
  assign n848 = n65884 & n847 ;
  assign n65885 = ~n814 ;
  assign n849 = x67 & n65885 ;
  assign n65886 = ~n808 ;
  assign n850 = n65886 & n849 ;
  assign n851 = n848 | n850 ;
  assign n65887 = ~n816 ;
  assign n852 = n65887 & n851 ;
  assign n65888 = ~n805 ;
  assign n853 = x68 & n65888 ;
  assign n65889 = ~n799 ;
  assign n854 = n65889 & n853 ;
  assign n855 = n807 | n854 ;
  assign n856 = n852 | n855 ;
  assign n65890 = ~n807 ;
  assign n857 = n65890 & n856 ;
  assign n65891 = ~n794 ;
  assign n858 = x69 & n65891 ;
  assign n65892 = ~n788 ;
  assign n859 = n65892 & n858 ;
  assign n860 = n796 | n859 ;
  assign n861 = n857 | n860 ;
  assign n65893 = ~n796 ;
  assign n862 = n65893 & n861 ;
  assign n65894 = ~n785 ;
  assign n863 = x70 & n65894 ;
  assign n65895 = ~n778 ;
  assign n864 = n65895 & n863 ;
  assign n865 = n787 | n864 ;
  assign n866 = n862 | n865 ;
  assign n65896 = ~n787 ;
  assign n867 = n65896 & n866 ;
  assign n65897 = ~n775 ;
  assign n868 = x71 & n65897 ;
  assign n65898 = ~n770 ;
  assign n869 = n65898 & n868 ;
  assign n870 = n777 | n869 ;
  assign n872 = n867 | n870 ;
  assign n65899 = ~n777 ;
  assign n873 = n65899 & n872 ;
  assign n880 = n65877 & n879 ;
  assign n185 = ~n769 ;
  assign n881 = n185 & n877 ;
  assign n882 = n669 & n769 ;
  assign n65901 = ~n882 ;
  assign n883 = x72 & n65901 ;
  assign n65902 = ~n881 ;
  assign n884 = n65902 & n883 ;
  assign n885 = n75217 | n263 ;
  assign n886 = n295 | n885 ;
  assign n887 = n884 | n886 ;
  assign n888 = n880 | n887 ;
  assign n890 = n873 | n888 ;
  assign n65903 = ~n889 ;
  assign n891 = n65903 & n890 ;
  assign n65904 = ~n867 ;
  assign n871 = n65904 & n870 ;
  assign n895 = n843 | n845 ;
  assign n896 = n65884 & n895 ;
  assign n897 = n816 | n850 ;
  assign n899 = n896 | n897 ;
  assign n900 = n65887 & n899 ;
  assign n902 = n855 | n900 ;
  assign n903 = n65890 & n902 ;
  assign n905 = n860 | n903 ;
  assign n906 = n65893 & n905 ;
  assign n907 = n865 | n906 ;
  assign n924 = n787 | n870 ;
  assign n65905 = ~n924 ;
  assign n925 = n907 & n65905 ;
  assign n926 = n871 | n925 ;
  assign n184 = ~n891 ;
  assign n927 = n184 & n926 ;
  assign n909 = n65896 & n907 ;
  assign n910 = n870 | n909 ;
  assign n911 = n65899 & n910 ;
  assign n912 = n888 | n911 ;
  assign n928 = n776 & n65903 ;
  assign n929 = n912 & n928 ;
  assign n930 = n927 | n929 ;
  assign n913 = n777 | n884 ;
  assign n914 = n880 | n913 ;
  assign n65907 = ~n914 ;
  assign n915 = n872 & n65907 ;
  assign n916 = n880 | n884 ;
  assign n65908 = ~n911 ;
  assign n917 = n65908 & n916 ;
  assign n918 = n915 | n917 ;
  assign n919 = n184 & n918 ;
  assign n920 = n768 & n879 ;
  assign n921 = n912 & n920 ;
  assign n922 = n919 | n921 ;
  assign n65909 = ~x73 ;
  assign n923 = n65909 & n922 ;
  assign n65910 = ~n921 ;
  assign n1033 = x73 & n65910 ;
  assign n65911 = ~n919 ;
  assign n1034 = n65911 & n1033 ;
  assign n1035 = n923 | n1034 ;
  assign n931 = n65877 & n930 ;
  assign n65912 = ~n906 ;
  assign n908 = n865 & n65912 ;
  assign n932 = n796 | n865 ;
  assign n65913 = ~n932 ;
  assign n933 = n861 & n65913 ;
  assign n934 = n908 | n933 ;
  assign n935 = n184 & n934 ;
  assign n936 = n786 & n65903 ;
  assign n937 = n912 & n936 ;
  assign n938 = n935 | n937 ;
  assign n939 = n65820 & n938 ;
  assign n65914 = ~n937 ;
  assign n1021 = x71 & n65914 ;
  assign n65915 = ~n935 ;
  assign n1022 = n65915 & n1021 ;
  assign n1023 = n939 | n1022 ;
  assign n65916 = ~n857 ;
  assign n904 = n65916 & n860 ;
  assign n940 = n807 | n860 ;
  assign n65917 = ~n940 ;
  assign n941 = n902 & n65917 ;
  assign n942 = n904 | n941 ;
  assign n943 = n184 & n942 ;
  assign n944 = n795 & n65903 ;
  assign n945 = n912 & n944 ;
  assign n946 = n943 | n945 ;
  assign n947 = n65791 & n946 ;
  assign n65918 = ~n900 ;
  assign n901 = n855 & n65918 ;
  assign n948 = n848 | n897 ;
  assign n949 = n816 | n855 ;
  assign n65919 = ~n949 ;
  assign n950 = n948 & n65919 ;
  assign n951 = n901 | n950 ;
  assign n952 = n184 & n951 ;
  assign n953 = n806 & n65903 ;
  assign n954 = n912 & n953 ;
  assign n955 = n952 | n954 ;
  assign n956 = n65772 & n955 ;
  assign n65920 = ~n954 ;
  assign n1010 = x69 & n65920 ;
  assign n65921 = ~n952 ;
  assign n1011 = n65921 & n1010 ;
  assign n1012 = n956 | n1011 ;
  assign n65922 = ~n848 ;
  assign n898 = n65922 & n897 ;
  assign n957 = n822 | n897 ;
  assign n65923 = ~n957 ;
  assign n958 = n847 & n65923 ;
  assign n959 = n898 | n958 ;
  assign n960 = n184 & n959 ;
  assign n961 = n815 & n65903 ;
  assign n962 = n912 & n961 ;
  assign n963 = n960 | n962 ;
  assign n964 = n65746 & n963 ;
  assign n65924 = ~n843 ;
  assign n894 = n65924 & n846 ;
  assign n965 = n842 | n846 ;
  assign n65925 = ~n965 ;
  assign n966 = n841 & n65925 ;
  assign n967 = n894 | n966 ;
  assign n968 = n184 & n967 ;
  assign n969 = n821 & n65903 ;
  assign n970 = n912 & n969 ;
  assign n971 = n968 | n970 ;
  assign n972 = n65721 & n971 ;
  assign n65926 = ~n970 ;
  assign n1000 = x67 & n65926 ;
  assign n65927 = ~n968 ;
  assign n1001 = n65927 & n1000 ;
  assign n1002 = n972 | n1001 ;
  assign n973 = n838 & n840 ;
  assign n974 = n65879 & n973 ;
  assign n65928 = ~n974 ;
  assign n975 = n841 & n65928 ;
  assign n976 = n184 & n975 ;
  assign n977 = n835 & n65903 ;
  assign n978 = n912 & n977 ;
  assign n979 = n976 | n978 ;
  assign n980 = n65686 & n979 ;
  assign n65929 = ~x54 ;
  assign n990 = n65929 & x64 ;
  assign n892 = n840 & n184 ;
  assign n981 = n65903 & n912 ;
  assign n65930 = ~n981 ;
  assign n982 = x64 & n65930 ;
  assign n65931 = ~n982 ;
  assign n983 = x55 & n65931 ;
  assign n984 = n892 | n983 ;
  assign n985 = x65 & n984 ;
  assign n893 = x64 & n184 ;
  assign n65932 = ~n893 ;
  assign n986 = x55 & n65932 ;
  assign n987 = n840 & n65930 ;
  assign n988 = x65 | n987 ;
  assign n989 = n986 | n988 ;
  assign n65933 = ~n985 ;
  assign n991 = n65933 & n989 ;
  assign n992 = n990 | n991 ;
  assign n993 = n892 | n986 ;
  assign n994 = n65670 & n993 ;
  assign n65934 = ~n994 ;
  assign n995 = n992 & n65934 ;
  assign n65935 = ~n978 ;
  assign n996 = x66 & n65935 ;
  assign n65936 = ~n976 ;
  assign n997 = n65936 & n996 ;
  assign n998 = n980 | n997 ;
  assign n999 = n995 | n998 ;
  assign n65937 = ~n980 ;
  assign n1003 = n65937 & n999 ;
  assign n1004 = n1002 | n1003 ;
  assign n65938 = ~n972 ;
  assign n1005 = n65938 & n1004 ;
  assign n65939 = ~n962 ;
  assign n1006 = x68 & n65939 ;
  assign n65940 = ~n960 ;
  assign n1007 = n65940 & n1006 ;
  assign n1008 = n964 | n1007 ;
  assign n1009 = n1005 | n1008 ;
  assign n65941 = ~n964 ;
  assign n1013 = n65941 & n1009 ;
  assign n1014 = n1012 | n1013 ;
  assign n65942 = ~n956 ;
  assign n1015 = n65942 & n1014 ;
  assign n65943 = ~n945 ;
  assign n1016 = x70 & n65943 ;
  assign n65944 = ~n943 ;
  assign n1017 = n65944 & n1016 ;
  assign n1018 = n947 | n1017 ;
  assign n1020 = n1015 | n1018 ;
  assign n65945 = ~n947 ;
  assign n1025 = n65945 & n1020 ;
  assign n1026 = n1023 | n1025 ;
  assign n65946 = ~n939 ;
  assign n1027 = n65946 & n1026 ;
  assign n65947 = ~n929 ;
  assign n1028 = x72 & n65947 ;
  assign n65948 = ~n927 ;
  assign n1029 = n65948 & n1028 ;
  assign n1030 = n931 | n1029 ;
  assign n1032 = n1027 | n1030 ;
  assign n65949 = ~n931 ;
  assign n1036 = n65949 & n1032 ;
  assign n1037 = n1035 | n1036 ;
  assign n65950 = ~n923 ;
  assign n1038 = n65950 & n1037 ;
  assign n1039 = n65243 | n65324 ;
  assign n1040 = n67612 | n1039 ;
  assign n1041 = n303 | n1040 ;
  assign n1042 = n1038 | n1041 ;
  assign n1073 = n930 & n1042 ;
  assign n1031 = n939 | n1030 ;
  assign n1046 = x65 & n993 ;
  assign n65951 = ~n1046 ;
  assign n1047 = n989 & n65951 ;
  assign n1049 = n990 | n1047 ;
  assign n1051 = n65934 & n1049 ;
  assign n1052 = n998 | n1051 ;
  assign n1053 = n65937 & n1052 ;
  assign n1054 = n1002 | n1053 ;
  assign n1055 = n65938 & n1054 ;
  assign n1056 = n1008 | n1055 ;
  assign n1057 = n65941 & n1056 ;
  assign n1058 = n1012 | n1057 ;
  assign n1059 = n65942 & n1058 ;
  assign n1060 = n1018 | n1059 ;
  assign n1061 = n65945 & n1060 ;
  assign n1062 = n1023 | n1061 ;
  assign n65952 = ~n1031 ;
  assign n1074 = n65952 & n1062 ;
  assign n65953 = ~n1027 ;
  assign n1075 = n65953 & n1030 ;
  assign n1076 = n1074 | n1075 ;
  assign n65954 = ~n1041 ;
  assign n1077 = n65954 & n1076 ;
  assign n65955 = ~n1038 ;
  assign n1078 = n65955 & n1077 ;
  assign n1079 = n1073 | n1078 ;
  assign n65956 = ~n922 ;
  assign n1043 = n65956 & n1042 ;
  assign n65957 = ~n1036 ;
  assign n1066 = n1035 & n65957 ;
  assign n1063 = n65946 & n1062 ;
  assign n1064 = n1030 | n1063 ;
  assign n1067 = n931 | n1035 ;
  assign n65958 = ~n1067 ;
  assign n1068 = n1064 & n65958 ;
  assign n1069 = n1066 | n1068 ;
  assign n1070 = n1042 | n1069 ;
  assign n65959 = ~n1043 ;
  assign n1071 = n65959 & n1070 ;
  assign n65960 = ~x74 ;
  assign n1072 = n65960 & n1071 ;
  assign n1080 = n65909 & n1079 ;
  assign n1081 = n938 & n1042 ;
  assign n1024 = n947 | n1023 ;
  assign n65961 = ~n1024 ;
  assign n1082 = n1020 & n65961 ;
  assign n65962 = ~n1061 ;
  assign n1083 = n1023 & n65962 ;
  assign n1084 = n1082 | n1083 ;
  assign n1085 = n65954 & n1084 ;
  assign n1086 = n65955 & n1085 ;
  assign n1087 = n1081 | n1086 ;
  assign n1088 = n65877 & n1087 ;
  assign n1089 = n946 & n1042 ;
  assign n1019 = n956 | n1018 ;
  assign n65963 = ~n1019 ;
  assign n1090 = n65963 & n1058 ;
  assign n65964 = ~n1015 ;
  assign n1091 = n65964 & n1018 ;
  assign n1092 = n1090 | n1091 ;
  assign n1093 = n65954 & n1092 ;
  assign n1094 = n65955 & n1093 ;
  assign n1095 = n1089 | n1094 ;
  assign n1096 = n65820 & n1095 ;
  assign n1097 = n955 & n1042 ;
  assign n1045 = n964 | n1012 ;
  assign n65965 = ~n1045 ;
  assign n1098 = n1009 & n65965 ;
  assign n65966 = ~n1057 ;
  assign n1099 = n1012 & n65966 ;
  assign n1100 = n1098 | n1099 ;
  assign n1101 = n65954 & n1100 ;
  assign n1102 = n65955 & n1101 ;
  assign n1103 = n1097 | n1102 ;
  assign n1104 = n65791 & n1103 ;
  assign n1105 = n963 & n1042 ;
  assign n1106 = n972 | n1008 ;
  assign n65967 = ~n1106 ;
  assign n1107 = n1054 & n65967 ;
  assign n65968 = ~n1005 ;
  assign n1108 = n65968 & n1008 ;
  assign n1109 = n1107 | n1108 ;
  assign n1110 = n65954 & n1109 ;
  assign n1111 = n65955 & n1110 ;
  assign n1112 = n1105 | n1111 ;
  assign n1113 = n65772 & n1112 ;
  assign n1114 = n971 & n1042 ;
  assign n1115 = n980 | n1002 ;
  assign n65969 = ~n1115 ;
  assign n1116 = n1052 & n65969 ;
  assign n65970 = ~n1053 ;
  assign n1117 = n1002 & n65970 ;
  assign n1118 = n1116 | n1117 ;
  assign n1119 = n65954 & n1118 ;
  assign n1120 = n65955 & n1119 ;
  assign n1121 = n1114 | n1120 ;
  assign n1122 = n65746 & n1121 ;
  assign n1123 = n979 & n1042 ;
  assign n1050 = n994 | n998 ;
  assign n65971 = ~n1050 ;
  assign n1124 = n992 & n65971 ;
  assign n65972 = ~n995 ;
  assign n1125 = n65972 & n998 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = n65954 & n1126 ;
  assign n1128 = n65955 & n1127 ;
  assign n1129 = n1123 | n1128 ;
  assign n1130 = n65721 & n1129 ;
  assign n1044 = n993 & n1042 ;
  assign n1048 = n989 & n990 ;
  assign n1131 = n65933 & n1048 ;
  assign n1132 = n1041 | n1131 ;
  assign n65973 = ~n1132 ;
  assign n1133 = n992 & n65973 ;
  assign n1134 = n65955 & n1133 ;
  assign n1135 = n1044 | n1134 ;
  assign n1136 = n65686 & n1135 ;
  assign n65974 = ~n65243 ;
  assign n1143 = n65974 & n990 ;
  assign n65975 = ~n65324 ;
  assign n1144 = n65975 & n1143 ;
  assign n1145 = n65695 & n1144 ;
  assign n1146 = n65696 & n1145 ;
  assign n1147 = n65955 & n1146 ;
  assign n1137 = x64 & n65960 ;
  assign n65976 = ~n261 ;
  assign n1138 = n65976 & n1137 ;
  assign n65977 = ~n259 ;
  assign n1139 = n65977 & n1138 ;
  assign n1140 = n65690 & n1139 ;
  assign n1141 = n65691 & n1140 ;
  assign n1142 = n65955 & n1141 ;
  assign n65978 = ~n1142 ;
  assign n1148 = x54 & n65978 ;
  assign n1149 = n1147 | n1148 ;
  assign n1150 = n65670 & n1149 ;
  assign n1065 = n65949 & n1064 ;
  assign n1152 = n1035 | n1065 ;
  assign n1153 = n65950 & n1152 ;
  assign n65979 = ~n1153 ;
  assign n1154 = n1141 & n65979 ;
  assign n65980 = ~n1154 ;
  assign n1155 = x54 & n65980 ;
  assign n1156 = n1147 | n1155 ;
  assign n1158 = x65 & n1156 ;
  assign n1157 = x65 | n1147 ;
  assign n1159 = n1148 | n1157 ;
  assign n65981 = ~n1158 ;
  assign n1160 = n65981 & n1159 ;
  assign n65982 = ~x53 ;
  assign n1161 = n65982 & x64 ;
  assign n1162 = n1160 | n1161 ;
  assign n65983 = ~n1150 ;
  assign n1163 = n65983 & n1162 ;
  assign n65984 = ~n1134 ;
  assign n1164 = x66 & n65984 ;
  assign n65985 = ~n1044 ;
  assign n1165 = n65985 & n1164 ;
  assign n1166 = n1136 | n1165 ;
  assign n1167 = n1163 | n1166 ;
  assign n65986 = ~n1136 ;
  assign n1168 = n65986 & n1167 ;
  assign n65987 = ~n1128 ;
  assign n1169 = x67 & n65987 ;
  assign n65988 = ~n1123 ;
  assign n1170 = n65988 & n1169 ;
  assign n1171 = n1168 | n1170 ;
  assign n65989 = ~n1130 ;
  assign n1172 = n65989 & n1171 ;
  assign n65990 = ~n1120 ;
  assign n1173 = x68 & n65990 ;
  assign n65991 = ~n1114 ;
  assign n1174 = n65991 & n1173 ;
  assign n1175 = n1122 | n1174 ;
  assign n1176 = n1172 | n1175 ;
  assign n65992 = ~n1122 ;
  assign n1177 = n65992 & n1176 ;
  assign n65993 = ~n1111 ;
  assign n1178 = x69 & n65993 ;
  assign n65994 = ~n1105 ;
  assign n1179 = n65994 & n1178 ;
  assign n1180 = n1113 | n1179 ;
  assign n1181 = n1177 | n1180 ;
  assign n65995 = ~n1113 ;
  assign n1182 = n65995 & n1181 ;
  assign n65996 = ~n1102 ;
  assign n1183 = x70 & n65996 ;
  assign n65997 = ~n1097 ;
  assign n1184 = n65997 & n1183 ;
  assign n1185 = n1104 | n1184 ;
  assign n1186 = n1182 | n1185 ;
  assign n65998 = ~n1104 ;
  assign n1187 = n65998 & n1186 ;
  assign n65999 = ~n1094 ;
  assign n1188 = x71 & n65999 ;
  assign n66000 = ~n1089 ;
  assign n1189 = n66000 & n1188 ;
  assign n1190 = n1096 | n1189 ;
  assign n1192 = n1187 | n1190 ;
  assign n66001 = ~n1096 ;
  assign n1193 = n66001 & n1192 ;
  assign n66002 = ~n1086 ;
  assign n1194 = x72 & n66002 ;
  assign n66003 = ~n1081 ;
  assign n1195 = n66003 & n1194 ;
  assign n1196 = n1088 | n1195 ;
  assign n1197 = n1193 | n1196 ;
  assign n66004 = ~n1088 ;
  assign n1198 = n66004 & n1197 ;
  assign n66005 = ~n1078 ;
  assign n1199 = x73 & n66005 ;
  assign n66006 = ~n1073 ;
  assign n1200 = n66006 & n1199 ;
  assign n1201 = n1080 | n1200 ;
  assign n1203 = n1198 | n1201 ;
  assign n66007 = ~n1080 ;
  assign n1204 = n66007 & n1203 ;
  assign n183 = ~n1042 ;
  assign n1205 = n183 & n1069 ;
  assign n1206 = n922 & n1042 ;
  assign n66009 = ~n1206 ;
  assign n1207 = x74 & n66009 ;
  assign n66010 = ~n1205 ;
  assign n1208 = n66010 & n1207 ;
  assign n1209 = n1072 | n1208 ;
  assign n1210 = n1204 | n1209 ;
  assign n66011 = ~n1072 ;
  assign n1211 = n66011 & n1210 ;
  assign n1212 = n259 | n261 ;
  assign n1213 = n75217 | n1212 ;
  assign n1214 = n295 | n1213 ;
  assign n1215 = n1211 | n1214 ;
  assign n1217 = n1079 & n1215 ;
  assign n66012 = ~n1198 ;
  assign n1202 = n66012 & n1201 ;
  assign n1219 = n65670 & n1156 ;
  assign n1151 = x65 & n1149 ;
  assign n66013 = ~n1151 ;
  assign n1218 = n66013 & n1159 ;
  assign n1220 = n1161 | n1218 ;
  assign n66014 = ~n1219 ;
  assign n1221 = n66014 & n1220 ;
  assign n1222 = n1166 | n1221 ;
  assign n1223 = n65986 & n1222 ;
  assign n1224 = n1130 | n1170 ;
  assign n1226 = n1223 | n1224 ;
  assign n1227 = n65989 & n1226 ;
  assign n1229 = n1175 | n1227 ;
  assign n1230 = n65992 & n1229 ;
  assign n1232 = n1180 | n1230 ;
  assign n1233 = n65995 & n1232 ;
  assign n1234 = n1185 | n1233 ;
  assign n1236 = n65998 & n1234 ;
  assign n1237 = n1190 | n1236 ;
  assign n1238 = n66001 & n1237 ;
  assign n1240 = n1196 | n1238 ;
  assign n1241 = n1088 | n1201 ;
  assign n66015 = ~n1241 ;
  assign n1242 = n1240 & n66015 ;
  assign n1243 = n1202 | n1242 ;
  assign n66016 = ~n1214 ;
  assign n1244 = n66016 & n1243 ;
  assign n66017 = ~n1211 ;
  assign n1245 = n66017 & n1244 ;
  assign n1246 = n1217 | n1245 ;
  assign n1247 = n65960 & n1246 ;
  assign n66018 = ~n1245 ;
  assign n1387 = x74 & n66018 ;
  assign n66019 = ~n1217 ;
  assign n1388 = n66019 & n1387 ;
  assign n1389 = n1247 | n1388 ;
  assign n1248 = n1087 & n1215 ;
  assign n66020 = ~n1238 ;
  assign n1239 = n1196 & n66020 ;
  assign n1249 = n1096 | n1196 ;
  assign n66021 = ~n1249 ;
  assign n1250 = n1192 & n66021 ;
  assign n1251 = n1239 | n1250 ;
  assign n1252 = n66016 & n1251 ;
  assign n1253 = n66017 & n1252 ;
  assign n1254 = n1248 | n1253 ;
  assign n1255 = n65909 & n1254 ;
  assign n1256 = n1095 & n1215 ;
  assign n66022 = ~n1187 ;
  assign n1191 = n66022 & n1190 ;
  assign n1257 = n1104 | n1190 ;
  assign n66023 = ~n1257 ;
  assign n1258 = n1234 & n66023 ;
  assign n1259 = n1191 | n1258 ;
  assign n1260 = n66016 & n1259 ;
  assign n1261 = n66017 & n1260 ;
  assign n1262 = n1256 | n1261 ;
  assign n1263 = n65877 & n1262 ;
  assign n66024 = ~n1261 ;
  assign n1375 = x72 & n66024 ;
  assign n66025 = ~n1256 ;
  assign n1376 = n66025 & n1375 ;
  assign n1377 = n1263 | n1376 ;
  assign n1264 = n1103 & n1215 ;
  assign n66026 = ~n1233 ;
  assign n1235 = n1185 & n66026 ;
  assign n1265 = n1113 | n1185 ;
  assign n66027 = ~n1265 ;
  assign n1266 = n1181 & n66027 ;
  assign n1267 = n1235 | n1266 ;
  assign n1268 = n66016 & n1267 ;
  assign n1269 = n66017 & n1268 ;
  assign n1270 = n1264 | n1269 ;
  assign n1271 = n65820 & n1270 ;
  assign n1272 = n1112 & n1215 ;
  assign n66028 = ~n1177 ;
  assign n1231 = n66028 & n1180 ;
  assign n1273 = n1122 | n1180 ;
  assign n66029 = ~n1273 ;
  assign n1274 = n1176 & n66029 ;
  assign n1275 = n1231 | n1274 ;
  assign n1276 = n66016 & n1275 ;
  assign n1277 = n66017 & n1276 ;
  assign n1278 = n1272 | n1277 ;
  assign n1279 = n65791 & n1278 ;
  assign n66030 = ~n1277 ;
  assign n1364 = x70 & n66030 ;
  assign n66031 = ~n1272 ;
  assign n1365 = n66031 & n1364 ;
  assign n1366 = n1279 | n1365 ;
  assign n1280 = n1121 & n1215 ;
  assign n66032 = ~n1227 ;
  assign n1228 = n1175 & n66032 ;
  assign n1281 = n1168 | n1224 ;
  assign n1282 = n1130 | n1175 ;
  assign n66033 = ~n1282 ;
  assign n1283 = n1281 & n66033 ;
  assign n1284 = n1228 | n1283 ;
  assign n1285 = n66016 & n1284 ;
  assign n1286 = n66017 & n1285 ;
  assign n1287 = n1280 | n1286 ;
  assign n1288 = n65772 & n1287 ;
  assign n1289 = n1129 & n1215 ;
  assign n66034 = ~n1168 ;
  assign n1225 = n66034 & n1224 ;
  assign n1290 = n1136 | n1224 ;
  assign n66035 = ~n1290 ;
  assign n1291 = n1167 & n66035 ;
  assign n1292 = n1225 | n1291 ;
  assign n1293 = n66016 & n1292 ;
  assign n1294 = n66017 & n1293 ;
  assign n1295 = n1289 | n1294 ;
  assign n1296 = n65746 & n1295 ;
  assign n66036 = ~n1294 ;
  assign n1354 = x68 & n66036 ;
  assign n66037 = ~n1289 ;
  assign n1355 = n66037 & n1354 ;
  assign n1356 = n1296 | n1355 ;
  assign n1297 = n1135 & n1215 ;
  assign n1298 = n1166 | n1219 ;
  assign n66038 = ~n1298 ;
  assign n1299 = n1162 & n66038 ;
  assign n66039 = ~n1221 ;
  assign n1300 = n1166 & n66039 ;
  assign n1301 = n1299 | n1300 ;
  assign n1302 = n66016 & n1301 ;
  assign n1303 = n66017 & n1302 ;
  assign n1304 = n1297 | n1303 ;
  assign n1305 = n65721 & n1304 ;
  assign n1306 = n1156 & n1215 ;
  assign n1307 = n1159 & n1161 ;
  assign n1308 = n65981 & n1307 ;
  assign n1309 = n1214 | n1308 ;
  assign n66040 = ~n1309 ;
  assign n1310 = n1162 & n66040 ;
  assign n1311 = n66017 & n1310 ;
  assign n1312 = n1306 | n1311 ;
  assign n1313 = n65686 & n1312 ;
  assign n1327 = n66004 & n1240 ;
  assign n1328 = n1201 | n1327 ;
  assign n1329 = n66007 & n1328 ;
  assign n1330 = n1209 | n1329 ;
  assign n1332 = n66011 & n1330 ;
  assign n1340 = n1214 | n1332 ;
  assign n1341 = n1149 & n1340 ;
  assign n1342 = n1311 | n1341 ;
  assign n1343 = n65686 & n1342 ;
  assign n66041 = ~n1311 ;
  assign n1344 = x66 & n66041 ;
  assign n66042 = ~n1341 ;
  assign n1345 = n66042 & n1344 ;
  assign n1346 = n1343 | n1345 ;
  assign n66043 = ~x75 ;
  assign n1314 = x64 & n66043 ;
  assign n1315 = n65975 & n1314 ;
  assign n1316 = n65695 & n1315 ;
  assign n1317 = n65696 & n1316 ;
  assign n1318 = n66017 & n1317 ;
  assign n66044 = ~n1318 ;
  assign n1319 = x53 & n66044 ;
  assign n1320 = n65976 & n1161 ;
  assign n1321 = n65977 & n1320 ;
  assign n1322 = n65690 & n1321 ;
  assign n1323 = n65691 & n1322 ;
  assign n1324 = n66017 & n1323 ;
  assign n1325 = n1319 | n1324 ;
  assign n1326 = x65 & n1325 ;
  assign n66045 = ~n1332 ;
  assign n1333 = n1323 & n66045 ;
  assign n1334 = x65 | n1333 ;
  assign n1335 = n1319 | n1334 ;
  assign n66046 = ~n1326 ;
  assign n1336 = n66046 & n1335 ;
  assign n66047 = ~x52 ;
  assign n1337 = n66047 & x64 ;
  assign n1338 = n1336 | n1337 ;
  assign n1339 = n65670 & n1325 ;
  assign n66048 = ~n1339 ;
  assign n1347 = n1338 & n66048 ;
  assign n1348 = n1346 | n1347 ;
  assign n66049 = ~n1313 ;
  assign n1349 = n66049 & n1348 ;
  assign n66050 = ~n1303 ;
  assign n1350 = x67 & n66050 ;
  assign n66051 = ~n1297 ;
  assign n1351 = n66051 & n1350 ;
  assign n1352 = n1305 | n1351 ;
  assign n1353 = n1349 | n1352 ;
  assign n66052 = ~n1305 ;
  assign n1357 = n66052 & n1353 ;
  assign n1358 = n1356 | n1357 ;
  assign n66053 = ~n1296 ;
  assign n1359 = n66053 & n1358 ;
  assign n66054 = ~n1286 ;
  assign n1360 = x69 & n66054 ;
  assign n66055 = ~n1280 ;
  assign n1361 = n66055 & n1360 ;
  assign n1362 = n1288 | n1361 ;
  assign n1363 = n1359 | n1362 ;
  assign n66056 = ~n1288 ;
  assign n1367 = n66056 & n1363 ;
  assign n1368 = n1366 | n1367 ;
  assign n66057 = ~n1279 ;
  assign n1369 = n66057 & n1368 ;
  assign n66058 = ~n1269 ;
  assign n1370 = x71 & n66058 ;
  assign n66059 = ~n1264 ;
  assign n1371 = n66059 & n1370 ;
  assign n1372 = n1271 | n1371 ;
  assign n1374 = n1369 | n1372 ;
  assign n66060 = ~n1271 ;
  assign n1379 = n66060 & n1374 ;
  assign n1380 = n1377 | n1379 ;
  assign n66061 = ~n1263 ;
  assign n1381 = n66061 & n1380 ;
  assign n66062 = ~n1253 ;
  assign n1382 = x73 & n66062 ;
  assign n66063 = ~n1248 ;
  assign n1383 = n66063 & n1382 ;
  assign n1384 = n1255 | n1383 ;
  assign n1386 = n1381 | n1384 ;
  assign n66064 = ~n1255 ;
  assign n1391 = n66064 & n1386 ;
  assign n1392 = n1389 | n1391 ;
  assign n66065 = ~n1247 ;
  assign n1393 = n66065 & n1392 ;
  assign n66066 = ~n1071 ;
  assign n1216 = n66066 & n1215 ;
  assign n66067 = ~n1329 ;
  assign n1331 = n1209 & n66067 ;
  assign n1394 = n1080 | n1209 ;
  assign n66068 = ~n1394 ;
  assign n1395 = n1203 & n66068 ;
  assign n1396 = n1331 | n1395 ;
  assign n1397 = n1215 | n1396 ;
  assign n66069 = ~n1216 ;
  assign n1398 = n66069 & n1397 ;
  assign n1399 = n66043 & n1398 ;
  assign n182 = ~n1215 ;
  assign n1400 = n182 & n1396 ;
  assign n1401 = n1071 & n1215 ;
  assign n66071 = ~n1401 ;
  assign n1402 = x75 & n66071 ;
  assign n66072 = ~n1400 ;
  assign n1403 = n66072 & n1402 ;
  assign n1404 = n65332 | n65654 ;
  assign n1405 = n380 | n1404 ;
  assign n1406 = n1403 | n1405 ;
  assign n1407 = n1399 | n1406 ;
  assign n1408 = n1393 | n1407 ;
  assign n1409 = n66016 & n1398 ;
  assign n66073 = ~n1409 ;
  assign n1410 = n1408 & n66073 ;
  assign n1412 = n1247 | n1403 ;
  assign n1413 = n1399 | n1412 ;
  assign n66074 = ~n1413 ;
  assign n1414 = n1392 & n66074 ;
  assign n1416 = n1317 & n66045 ;
  assign n66075 = ~n1416 ;
  assign n1417 = x53 & n66075 ;
  assign n1418 = n1324 | n1417 ;
  assign n1419 = x65 & n1418 ;
  assign n66076 = ~n1419 ;
  assign n1420 = n1335 & n66076 ;
  assign n1421 = n1337 | n1420 ;
  assign n1422 = n66048 & n1421 ;
  assign n66077 = ~n1306 ;
  assign n1423 = n66077 & n1344 ;
  assign n1424 = n1313 | n1423 ;
  assign n1425 = n1422 | n1424 ;
  assign n66078 = ~n1343 ;
  assign n1426 = n66078 & n1425 ;
  assign n1427 = n1352 | n1426 ;
  assign n1428 = n66052 & n1427 ;
  assign n1429 = n1356 | n1428 ;
  assign n1430 = n66053 & n1429 ;
  assign n1431 = n1362 | n1430 ;
  assign n1432 = n66056 & n1431 ;
  assign n1433 = n1366 | n1432 ;
  assign n1434 = n66057 & n1433 ;
  assign n1435 = n1372 | n1434 ;
  assign n1436 = n66060 & n1435 ;
  assign n1437 = n1377 | n1436 ;
  assign n1438 = n66061 & n1437 ;
  assign n1439 = n1384 | n1438 ;
  assign n1440 = n66064 & n1439 ;
  assign n1441 = n1389 | n1440 ;
  assign n1442 = n66065 & n1441 ;
  assign n1443 = n1399 | n1403 ;
  assign n66079 = ~n1442 ;
  assign n1444 = n66079 & n1443 ;
  assign n1445 = n1414 | n1444 ;
  assign n181 = ~n1410 ;
  assign n1446 = n181 & n1445 ;
  assign n1447 = n1214 & n1398 ;
  assign n1448 = n1408 & n1447 ;
  assign n1449 = n1446 | n1448 ;
  assign n66081 = ~x76 ;
  assign n1450 = n66081 & n1449 ;
  assign n66082 = ~n1391 ;
  assign n1451 = n1389 & n66082 ;
  assign n1390 = n1255 | n1389 ;
  assign n66083 = ~n1390 ;
  assign n1452 = n1386 & n66083 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = n181 & n1453 ;
  assign n1455 = n1246 & n66073 ;
  assign n1456 = n1408 & n1455 ;
  assign n1457 = n1454 | n1456 ;
  assign n1458 = n66043 & n1457 ;
  assign n66084 = ~n1438 ;
  assign n1459 = n1384 & n66084 ;
  assign n1385 = n1263 | n1384 ;
  assign n66085 = ~n1385 ;
  assign n1460 = n66085 & n1437 ;
  assign n1461 = n1459 | n1460 ;
  assign n1462 = n181 & n1461 ;
  assign n1463 = n1254 & n66073 ;
  assign n1464 = n1408 & n1463 ;
  assign n1465 = n1462 | n1464 ;
  assign n1466 = n65960 & n1465 ;
  assign n66086 = ~n1379 ;
  assign n1467 = n1377 & n66086 ;
  assign n1378 = n1271 | n1377 ;
  assign n66087 = ~n1378 ;
  assign n1468 = n1374 & n66087 ;
  assign n1469 = n1467 | n1468 ;
  assign n1470 = n181 & n1469 ;
  assign n1471 = n1262 & n66073 ;
  assign n1472 = n1408 & n1471 ;
  assign n1473 = n1470 | n1472 ;
  assign n1474 = n65909 & n1473 ;
  assign n66088 = ~n1434 ;
  assign n1475 = n1372 & n66088 ;
  assign n1373 = n1279 | n1372 ;
  assign n66089 = ~n1373 ;
  assign n1476 = n66089 & n1433 ;
  assign n1477 = n1475 | n1476 ;
  assign n1478 = n181 & n1477 ;
  assign n1479 = n1270 & n66073 ;
  assign n1480 = n1408 & n1479 ;
  assign n1481 = n1478 | n1480 ;
  assign n1482 = n65877 & n1481 ;
  assign n66090 = ~n1367 ;
  assign n1483 = n1366 & n66090 ;
  assign n1415 = n1288 | n1366 ;
  assign n66091 = ~n1415 ;
  assign n1484 = n1363 & n66091 ;
  assign n1485 = n1483 | n1484 ;
  assign n1486 = n181 & n1485 ;
  assign n1487 = n1278 & n66073 ;
  assign n1488 = n1408 & n1487 ;
  assign n1489 = n1486 | n1488 ;
  assign n1490 = n65820 & n1489 ;
  assign n66092 = ~n1430 ;
  assign n1492 = n1362 & n66092 ;
  assign n1491 = n1296 | n1362 ;
  assign n66093 = ~n1491 ;
  assign n1493 = n1429 & n66093 ;
  assign n1494 = n1492 | n1493 ;
  assign n1495 = n181 & n1494 ;
  assign n1496 = n1287 & n66073 ;
  assign n1497 = n1408 & n1496 ;
  assign n1498 = n1495 | n1497 ;
  assign n1499 = n65791 & n1498 ;
  assign n66094 = ~n1357 ;
  assign n1501 = n1356 & n66094 ;
  assign n1500 = n1305 | n1356 ;
  assign n66095 = ~n1500 ;
  assign n1502 = n1353 & n66095 ;
  assign n1503 = n1501 | n1502 ;
  assign n1504 = n181 & n1503 ;
  assign n1505 = n1295 & n66073 ;
  assign n1506 = n1408 & n1505 ;
  assign n1507 = n1504 | n1506 ;
  assign n1508 = n65772 & n1507 ;
  assign n1509 = n66049 & n1425 ;
  assign n66096 = ~n1509 ;
  assign n1511 = n1352 & n66096 ;
  assign n1510 = n1313 | n1352 ;
  assign n66097 = ~n1510 ;
  assign n1512 = n1425 & n66097 ;
  assign n1513 = n1511 | n1512 ;
  assign n1514 = n181 & n1513 ;
  assign n1515 = n1304 & n66073 ;
  assign n1516 = n1408 & n1515 ;
  assign n1517 = n1514 | n1516 ;
  assign n1518 = n65746 & n1517 ;
  assign n66098 = ~n1347 ;
  assign n1520 = n1346 & n66098 ;
  assign n1519 = n1339 | n1424 ;
  assign n66099 = ~n1519 ;
  assign n1521 = n1338 & n66099 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = n181 & n1522 ;
  assign n1524 = n1312 & n66073 ;
  assign n1525 = n1408 & n1524 ;
  assign n1526 = n1523 | n1525 ;
  assign n1527 = n65721 & n1526 ;
  assign n1528 = n1335 & n1337 ;
  assign n1529 = n66046 & n1528 ;
  assign n66100 = ~n1529 ;
  assign n1530 = n1338 & n66100 ;
  assign n1531 = n181 & n1530 ;
  assign n1532 = n1325 & n66073 ;
  assign n1533 = n1408 & n1532 ;
  assign n1534 = n1531 | n1533 ;
  assign n1535 = n65686 & n1534 ;
  assign n1411 = n1337 & n181 ;
  assign n1540 = x64 & n181 ;
  assign n66101 = ~n1540 ;
  assign n1541 = x52 & n66101 ;
  assign n1542 = n1411 | n1541 ;
  assign n1544 = x65 & n1542 ;
  assign n1536 = n1407 | n1442 ;
  assign n1537 = n66073 & n1536 ;
  assign n66102 = ~n1537 ;
  assign n1538 = x64 & n66102 ;
  assign n66103 = ~n1538 ;
  assign n1539 = x52 & n66103 ;
  assign n1543 = x65 | n1411 ;
  assign n1545 = n1539 | n1543 ;
  assign n66104 = ~n1544 ;
  assign n1546 = n66104 & n1545 ;
  assign n66105 = ~x51 ;
  assign n1547 = n66105 & x64 ;
  assign n1548 = n1546 | n1547 ;
  assign n1549 = n65670 & n1542 ;
  assign n66106 = ~n1549 ;
  assign n1550 = n1548 & n66106 ;
  assign n66107 = ~n1533 ;
  assign n1551 = x66 & n66107 ;
  assign n66108 = ~n1531 ;
  assign n1552 = n66108 & n1551 ;
  assign n1553 = n1535 | n1552 ;
  assign n1554 = n1550 | n1553 ;
  assign n66109 = ~n1535 ;
  assign n1555 = n66109 & n1554 ;
  assign n66110 = ~n1525 ;
  assign n1556 = x67 & n66110 ;
  assign n66111 = ~n1523 ;
  assign n1557 = n66111 & n1556 ;
  assign n1558 = n1527 | n1557 ;
  assign n1559 = n1555 | n1558 ;
  assign n66112 = ~n1527 ;
  assign n1560 = n66112 & n1559 ;
  assign n66113 = ~n1516 ;
  assign n1561 = x68 & n66113 ;
  assign n66114 = ~n1514 ;
  assign n1562 = n66114 & n1561 ;
  assign n1563 = n1518 | n1562 ;
  assign n1564 = n1560 | n1563 ;
  assign n66115 = ~n1518 ;
  assign n1565 = n66115 & n1564 ;
  assign n66116 = ~n1506 ;
  assign n1566 = x69 & n66116 ;
  assign n66117 = ~n1504 ;
  assign n1567 = n66117 & n1566 ;
  assign n1568 = n1508 | n1567 ;
  assign n1570 = n1565 | n1568 ;
  assign n66118 = ~n1508 ;
  assign n1571 = n66118 & n1570 ;
  assign n66119 = ~n1497 ;
  assign n1572 = x70 & n66119 ;
  assign n66120 = ~n1495 ;
  assign n1573 = n66120 & n1572 ;
  assign n1574 = n1499 | n1573 ;
  assign n1575 = n1571 | n1574 ;
  assign n66121 = ~n1499 ;
  assign n1576 = n66121 & n1575 ;
  assign n66122 = ~n1488 ;
  assign n1577 = x71 & n66122 ;
  assign n66123 = ~n1486 ;
  assign n1578 = n66123 & n1577 ;
  assign n1579 = n1490 | n1578 ;
  assign n1581 = n1576 | n1579 ;
  assign n66124 = ~n1490 ;
  assign n1582 = n66124 & n1581 ;
  assign n66125 = ~n1480 ;
  assign n1583 = x72 & n66125 ;
  assign n66126 = ~n1478 ;
  assign n1584 = n66126 & n1583 ;
  assign n1585 = n1482 | n1584 ;
  assign n1586 = n1582 | n1585 ;
  assign n66127 = ~n1482 ;
  assign n1587 = n66127 & n1586 ;
  assign n66128 = ~n1472 ;
  assign n1588 = x73 & n66128 ;
  assign n66129 = ~n1470 ;
  assign n1589 = n66129 & n1588 ;
  assign n1590 = n1474 | n1589 ;
  assign n1592 = n1587 | n1590 ;
  assign n66130 = ~n1474 ;
  assign n1593 = n66130 & n1592 ;
  assign n66131 = ~n1464 ;
  assign n1594 = x74 & n66131 ;
  assign n66132 = ~n1462 ;
  assign n1595 = n66132 & n1594 ;
  assign n1596 = n1466 | n1595 ;
  assign n1597 = n1593 | n1596 ;
  assign n66133 = ~n1466 ;
  assign n1598 = n66133 & n1597 ;
  assign n66134 = ~n1456 ;
  assign n1599 = x75 & n66134 ;
  assign n66135 = ~n1454 ;
  assign n1600 = n66135 & n1599 ;
  assign n1601 = n1458 | n1600 ;
  assign n1603 = n1598 | n1601 ;
  assign n66136 = ~n1458 ;
  assign n1604 = n66136 & n1603 ;
  assign n66137 = ~n1448 ;
  assign n1605 = x76 & n66137 ;
  assign n66138 = ~n1446 ;
  assign n1606 = n66138 & n1605 ;
  assign n1607 = n1450 | n1606 ;
  assign n1608 = n1604 | n1607 ;
  assign n66139 = ~n1450 ;
  assign n1609 = n66139 & n1608 ;
  assign n1610 = n459 | n461 ;
  assign n1611 = n469 | n1610 ;
  assign n1612 = n1609 | n1611 ;
  assign n1613 = n1411 | n1539 ;
  assign n1614 = x65 & n1613 ;
  assign n66140 = ~n1614 ;
  assign n1615 = n1545 & n66140 ;
  assign n1616 = n1547 | n1615 ;
  assign n1617 = n66106 & n1616 ;
  assign n1618 = n1553 | n1617 ;
  assign n1619 = n66109 & n1618 ;
  assign n1621 = n1558 | n1619 ;
  assign n1622 = n66112 & n1621 ;
  assign n1624 = n1563 | n1622 ;
  assign n1625 = n66115 & n1624 ;
  assign n1626 = n1568 | n1625 ;
  assign n1627 = n66118 & n1626 ;
  assign n1628 = n1574 | n1627 ;
  assign n1630 = n66121 & n1628 ;
  assign n1631 = n1579 | n1630 ;
  assign n1632 = n66124 & n1631 ;
  assign n1633 = n1585 | n1632 ;
  assign n1635 = n66127 & n1633 ;
  assign n1636 = n1590 | n1635 ;
  assign n1637 = n66130 & n1636 ;
  assign n1638 = n1596 | n1637 ;
  assign n1640 = n66133 & n1638 ;
  assign n1641 = n1601 | n1640 ;
  assign n1642 = n66136 & n1641 ;
  assign n66141 = ~n1642 ;
  assign n1643 = n1607 & n66141 ;
  assign n1645 = n1458 | n1607 ;
  assign n66142 = ~n1645 ;
  assign n1646 = n1603 & n66142 ;
  assign n1647 = n1643 | n1646 ;
  assign n1648 = n1612 | n1647 ;
  assign n66143 = ~n1449 ;
  assign n1649 = n66143 & n1612 ;
  assign n66144 = ~n1649 ;
  assign n1650 = n1648 & n66144 ;
  assign n66145 = ~x77 ;
  assign n1651 = n66145 & n1650 ;
  assign n180 = ~n1612 ;
  assign n1829 = n180 & n1647 ;
  assign n1830 = n1449 & n1612 ;
  assign n66147 = ~n1830 ;
  assign n1831 = x77 & n66147 ;
  assign n66148 = ~n1829 ;
  assign n1832 = n66148 & n1831 ;
  assign n1833 = n1651 | n1832 ;
  assign n1652 = n1457 & n1612 ;
  assign n66149 = ~n1598 ;
  assign n1602 = n66149 & n1601 ;
  assign n1653 = n1466 | n1601 ;
  assign n66150 = ~n1653 ;
  assign n1654 = n1638 & n66150 ;
  assign n1655 = n1602 | n1654 ;
  assign n66151 = ~n1611 ;
  assign n1656 = n66151 & n1655 ;
  assign n66152 = ~n1609 ;
  assign n1657 = n66152 & n1656 ;
  assign n1658 = n1652 | n1657 ;
  assign n1659 = n66081 & n1658 ;
  assign n1660 = n1465 & n1612 ;
  assign n66153 = ~n1637 ;
  assign n1639 = n1596 & n66153 ;
  assign n1661 = n1474 | n1596 ;
  assign n66154 = ~n1661 ;
  assign n1662 = n1592 & n66154 ;
  assign n1663 = n1639 | n1662 ;
  assign n1664 = n66151 & n1663 ;
  assign n1665 = n66152 & n1664 ;
  assign n1666 = n1660 | n1665 ;
  assign n1667 = n66043 & n1666 ;
  assign n66155 = ~n1665 ;
  assign n1817 = x75 & n66155 ;
  assign n66156 = ~n1660 ;
  assign n1818 = n66156 & n1817 ;
  assign n1819 = n1667 | n1818 ;
  assign n1668 = n1473 & n1612 ;
  assign n66157 = ~n1587 ;
  assign n1591 = n66157 & n1590 ;
  assign n1669 = n1482 | n1590 ;
  assign n66158 = ~n1669 ;
  assign n1670 = n1633 & n66158 ;
  assign n1671 = n1591 | n1670 ;
  assign n1672 = n66151 & n1671 ;
  assign n1673 = n66152 & n1672 ;
  assign n1674 = n1668 | n1673 ;
  assign n1675 = n65960 & n1674 ;
  assign n1676 = n1481 & n1612 ;
  assign n66159 = ~n1632 ;
  assign n1634 = n1585 & n66159 ;
  assign n1677 = n1490 | n1585 ;
  assign n66160 = ~n1677 ;
  assign n1678 = n1581 & n66160 ;
  assign n1679 = n1634 | n1678 ;
  assign n1680 = n66151 & n1679 ;
  assign n1681 = n66152 & n1680 ;
  assign n1682 = n1676 | n1681 ;
  assign n1683 = n65909 & n1682 ;
  assign n66161 = ~n1681 ;
  assign n1805 = x73 & n66161 ;
  assign n66162 = ~n1676 ;
  assign n1806 = n66162 & n1805 ;
  assign n1807 = n1683 | n1806 ;
  assign n1684 = n1489 & n1612 ;
  assign n66163 = ~n1576 ;
  assign n1580 = n66163 & n1579 ;
  assign n1685 = n1499 | n1579 ;
  assign n66164 = ~n1685 ;
  assign n1686 = n1628 & n66164 ;
  assign n1687 = n1580 | n1686 ;
  assign n1688 = n66151 & n1687 ;
  assign n1689 = n66152 & n1688 ;
  assign n1690 = n1684 | n1689 ;
  assign n1691 = n65877 & n1690 ;
  assign n1692 = n1498 & n1612 ;
  assign n66165 = ~n1627 ;
  assign n1629 = n1574 & n66165 ;
  assign n1693 = n1508 | n1574 ;
  assign n66166 = ~n1693 ;
  assign n1694 = n1570 & n66166 ;
  assign n1695 = n1629 | n1694 ;
  assign n1696 = n66151 & n1695 ;
  assign n1697 = n66152 & n1696 ;
  assign n1698 = n1692 | n1697 ;
  assign n1699 = n65820 & n1698 ;
  assign n66167 = ~n1697 ;
  assign n1793 = x71 & n66167 ;
  assign n66168 = ~n1692 ;
  assign n1794 = n66168 & n1793 ;
  assign n1795 = n1699 | n1794 ;
  assign n1700 = n1507 & n1612 ;
  assign n66169 = ~n1565 ;
  assign n1569 = n66169 & n1568 ;
  assign n1701 = n1518 | n1568 ;
  assign n66170 = ~n1701 ;
  assign n1702 = n1624 & n66170 ;
  assign n1703 = n1569 | n1702 ;
  assign n1704 = n66151 & n1703 ;
  assign n1705 = n66152 & n1704 ;
  assign n1706 = n1700 | n1705 ;
  assign n1707 = n65791 & n1706 ;
  assign n1708 = n1517 & n1612 ;
  assign n66171 = ~n1622 ;
  assign n1623 = n1563 & n66171 ;
  assign n1709 = n1527 | n1563 ;
  assign n66172 = ~n1709 ;
  assign n1710 = n1559 & n66172 ;
  assign n1711 = n1623 | n1710 ;
  assign n1712 = n66151 & n1711 ;
  assign n1713 = n66152 & n1712 ;
  assign n1714 = n1708 | n1713 ;
  assign n1715 = n65772 & n1714 ;
  assign n66173 = ~n1713 ;
  assign n1782 = x69 & n66173 ;
  assign n66174 = ~n1708 ;
  assign n1783 = n66174 & n1782 ;
  assign n1784 = n1715 | n1783 ;
  assign n1716 = n1526 & n1612 ;
  assign n66175 = ~n1555 ;
  assign n1620 = n66175 & n1558 ;
  assign n1717 = n1535 | n1558 ;
  assign n66176 = ~n1717 ;
  assign n1718 = n1554 & n66176 ;
  assign n1719 = n1620 | n1718 ;
  assign n1720 = n66151 & n1719 ;
  assign n1721 = n66152 & n1720 ;
  assign n1722 = n1716 | n1721 ;
  assign n1723 = n65746 & n1722 ;
  assign n1724 = n1534 & n1612 ;
  assign n1725 = n1549 | n1553 ;
  assign n66177 = ~n1725 ;
  assign n1726 = n1548 & n66177 ;
  assign n66178 = ~n1617 ;
  assign n1727 = n1553 & n66178 ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = n66151 & n1728 ;
  assign n1730 = n66152 & n1729 ;
  assign n1731 = n1724 | n1730 ;
  assign n1732 = n65721 & n1731 ;
  assign n66179 = ~n1730 ;
  assign n1772 = x67 & n66179 ;
  assign n66180 = ~n1724 ;
  assign n1773 = n66180 & n1772 ;
  assign n1774 = n1732 | n1773 ;
  assign n1644 = n1607 | n1642 ;
  assign n1733 = n66139 & n1644 ;
  assign n1734 = n1611 | n1733 ;
  assign n1735 = n1613 & n1734 ;
  assign n1736 = n1545 & n1547 ;
  assign n1737 = n66104 & n1736 ;
  assign n1738 = n1611 | n1737 ;
  assign n66181 = ~n1738 ;
  assign n1739 = n1548 & n66181 ;
  assign n1740 = n66152 & n1739 ;
  assign n1741 = n1735 | n1740 ;
  assign n1742 = n65686 & n1741 ;
  assign n66182 = ~x50 ;
  assign n1761 = n66182 & x64 ;
  assign n1743 = x64 & n66145 ;
  assign n66183 = ~n65317 ;
  assign n1744 = n66183 & n1743 ;
  assign n66184 = ~n65302 ;
  assign n1745 = n66184 & n1744 ;
  assign n1746 = n65776 & n1745 ;
  assign n1747 = n65777 & n1746 ;
  assign n66185 = ~n1733 ;
  assign n1749 = n66185 & n1747 ;
  assign n66186 = ~n1749 ;
  assign n1750 = x51 & n66186 ;
  assign n1751 = n65977 & n1547 ;
  assign n1752 = n65690 & n1751 ;
  assign n1753 = n65691 & n1752 ;
  assign n1754 = n66152 & n1753 ;
  assign n1755 = n1750 | n1754 ;
  assign n1756 = x65 & n1755 ;
  assign n1748 = n66152 & n1747 ;
  assign n66187 = ~n1748 ;
  assign n1757 = x51 & n66187 ;
  assign n1758 = n66185 & n1753 ;
  assign n1759 = x65 | n1758 ;
  assign n1760 = n1757 | n1759 ;
  assign n66188 = ~n1756 ;
  assign n1762 = n66188 & n1760 ;
  assign n1763 = n1761 | n1762 ;
  assign n1764 = n1754 | n1757 ;
  assign n1765 = n65670 & n1764 ;
  assign n66189 = ~n1765 ;
  assign n1766 = n1763 & n66189 ;
  assign n1767 = n66185 & n1739 ;
  assign n66190 = ~n1767 ;
  assign n1768 = x66 & n66190 ;
  assign n66191 = ~n1735 ;
  assign n1769 = n66191 & n1768 ;
  assign n1770 = n1742 | n1769 ;
  assign n1771 = n1766 | n1770 ;
  assign n66192 = ~n1742 ;
  assign n1775 = n66192 & n1771 ;
  assign n1776 = n1774 | n1775 ;
  assign n66193 = ~n1732 ;
  assign n1777 = n66193 & n1776 ;
  assign n66194 = ~n1721 ;
  assign n1778 = x68 & n66194 ;
  assign n66195 = ~n1716 ;
  assign n1779 = n66195 & n1778 ;
  assign n1780 = n1723 | n1779 ;
  assign n1781 = n1777 | n1780 ;
  assign n66196 = ~n1723 ;
  assign n1785 = n66196 & n1781 ;
  assign n1786 = n1784 | n1785 ;
  assign n66197 = ~n1715 ;
  assign n1787 = n66197 & n1786 ;
  assign n66198 = ~n1705 ;
  assign n1788 = x70 & n66198 ;
  assign n66199 = ~n1700 ;
  assign n1789 = n66199 & n1788 ;
  assign n1790 = n1707 | n1789 ;
  assign n1792 = n1787 | n1790 ;
  assign n66200 = ~n1707 ;
  assign n1797 = n66200 & n1792 ;
  assign n1798 = n1795 | n1797 ;
  assign n66201 = ~n1699 ;
  assign n1799 = n66201 & n1798 ;
  assign n66202 = ~n1689 ;
  assign n1800 = x72 & n66202 ;
  assign n66203 = ~n1684 ;
  assign n1801 = n66203 & n1800 ;
  assign n1802 = n1691 | n1801 ;
  assign n1804 = n1799 | n1802 ;
  assign n66204 = ~n1691 ;
  assign n1809 = n66204 & n1804 ;
  assign n1810 = n1807 | n1809 ;
  assign n66205 = ~n1683 ;
  assign n1811 = n66205 & n1810 ;
  assign n66206 = ~n1673 ;
  assign n1812 = x74 & n66206 ;
  assign n66207 = ~n1668 ;
  assign n1813 = n66207 & n1812 ;
  assign n1814 = n1675 | n1813 ;
  assign n1816 = n1811 | n1814 ;
  assign n66208 = ~n1675 ;
  assign n1821 = n66208 & n1816 ;
  assign n1822 = n1819 | n1821 ;
  assign n66209 = ~n1667 ;
  assign n1823 = n66209 & n1822 ;
  assign n66210 = ~n1657 ;
  assign n1824 = x76 & n66210 ;
  assign n66211 = ~n1652 ;
  assign n1825 = n66211 & n1824 ;
  assign n1826 = n1659 | n1825 ;
  assign n1828 = n1823 | n1826 ;
  assign n66212 = ~n1659 ;
  assign n1834 = n66212 & n1828 ;
  assign n1835 = n1833 | n1834 ;
  assign n66213 = ~n1651 ;
  assign n1836 = n66213 & n1835 ;
  assign n1840 = n1836 | n1839 ;
  assign n66214 = ~n1650 ;
  assign n1842 = n66214 & n1840 ;
  assign n66215 = ~n1834 ;
  assign n2056 = n1833 & n66215 ;
  assign n1844 = x65 & n1764 ;
  assign n66216 = ~n1844 ;
  assign n1845 = n1760 & n66216 ;
  assign n1847 = n1761 | n1845 ;
  assign n1848 = n66189 & n1847 ;
  assign n1849 = n1770 | n1848 ;
  assign n1850 = n66192 & n1849 ;
  assign n1851 = n1774 | n1850 ;
  assign n1852 = n66193 & n1851 ;
  assign n1853 = n1780 | n1852 ;
  assign n1854 = n66196 & n1853 ;
  assign n1855 = n1784 | n1854 ;
  assign n1856 = n66197 & n1855 ;
  assign n1857 = n1790 | n1856 ;
  assign n1858 = n66200 & n1857 ;
  assign n1859 = n1795 | n1858 ;
  assign n1860 = n66201 & n1859 ;
  assign n1861 = n1802 | n1860 ;
  assign n1862 = n66204 & n1861 ;
  assign n1863 = n1807 | n1862 ;
  assign n1864 = n66205 & n1863 ;
  assign n1865 = n1814 | n1864 ;
  assign n1866 = n66208 & n1865 ;
  assign n1867 = n1819 | n1866 ;
  assign n1972 = n66209 & n1867 ;
  assign n1973 = n1826 | n1972 ;
  assign n2057 = n1659 | n1833 ;
  assign n66217 = ~n2057 ;
  assign n2058 = n1973 & n66217 ;
  assign n2059 = n2056 | n2058 ;
  assign n2060 = n1840 | n2059 ;
  assign n66218 = ~n1842 ;
  assign n2061 = n66218 & n2060 ;
  assign n66219 = ~n1839 ;
  assign n2072 = n66219 & n2061 ;
  assign n1843 = n1658 & n1840 ;
  assign n1827 = n1667 | n1826 ;
  assign n66220 = ~n1827 ;
  assign n1868 = n66220 & n1867 ;
  assign n66221 = ~n1823 ;
  assign n1869 = n66221 & n1826 ;
  assign n1870 = n1868 | n1869 ;
  assign n1871 = n66219 & n1870 ;
  assign n66222 = ~n1836 ;
  assign n1872 = n66222 & n1871 ;
  assign n1873 = n1843 | n1872 ;
  assign n1874 = n66145 & n1873 ;
  assign n1875 = n1666 & n1840 ;
  assign n1820 = n1675 | n1819 ;
  assign n66223 = ~n1820 ;
  assign n1876 = n1816 & n66223 ;
  assign n66224 = ~n1866 ;
  assign n1877 = n1819 & n66224 ;
  assign n1878 = n1876 | n1877 ;
  assign n1879 = n66219 & n1878 ;
  assign n1880 = n66222 & n1879 ;
  assign n1881 = n1875 | n1880 ;
  assign n1882 = n66081 & n1881 ;
  assign n1883 = n1674 & n1840 ;
  assign n1815 = n1683 | n1814 ;
  assign n66225 = ~n1815 ;
  assign n1884 = n66225 & n1863 ;
  assign n66226 = ~n1811 ;
  assign n1885 = n66226 & n1814 ;
  assign n1886 = n1884 | n1885 ;
  assign n1887 = n66219 & n1886 ;
  assign n1888 = n66222 & n1887 ;
  assign n1889 = n1883 | n1888 ;
  assign n1890 = n66043 & n1889 ;
  assign n1891 = n1682 & n1840 ;
  assign n1808 = n1691 | n1807 ;
  assign n66227 = ~n1808 ;
  assign n1892 = n1804 & n66227 ;
  assign n66228 = ~n1862 ;
  assign n1893 = n1807 & n66228 ;
  assign n1894 = n1892 | n1893 ;
  assign n1895 = n66219 & n1894 ;
  assign n1896 = n66222 & n1895 ;
  assign n1897 = n1891 | n1896 ;
  assign n1898 = n65960 & n1897 ;
  assign n1899 = n1690 & n1840 ;
  assign n1803 = n1699 | n1802 ;
  assign n66229 = ~n1803 ;
  assign n1900 = n66229 & n1859 ;
  assign n66230 = ~n1799 ;
  assign n1901 = n66230 & n1802 ;
  assign n1902 = n1900 | n1901 ;
  assign n1903 = n66219 & n1902 ;
  assign n1904 = n66222 & n1903 ;
  assign n1905 = n1899 | n1904 ;
  assign n1906 = n65909 & n1905 ;
  assign n1907 = n1698 & n1840 ;
  assign n1796 = n1707 | n1795 ;
  assign n66231 = ~n1796 ;
  assign n1908 = n1792 & n66231 ;
  assign n66232 = ~n1858 ;
  assign n1909 = n1795 & n66232 ;
  assign n1910 = n1908 | n1909 ;
  assign n1911 = n66219 & n1910 ;
  assign n1912 = n66222 & n1911 ;
  assign n1913 = n1907 | n1912 ;
  assign n1914 = n65877 & n1913 ;
  assign n1915 = n1706 & n1840 ;
  assign n1791 = n1715 | n1790 ;
  assign n66233 = ~n1791 ;
  assign n1916 = n1786 & n66233 ;
  assign n66234 = ~n1787 ;
  assign n1917 = n66234 & n1790 ;
  assign n1918 = n1916 | n1917 ;
  assign n1919 = n66219 & n1918 ;
  assign n1920 = n66222 & n1919 ;
  assign n1921 = n1915 | n1920 ;
  assign n1922 = n65820 & n1921 ;
  assign n1923 = n1714 & n1840 ;
  assign n1924 = n1723 | n1784 ;
  assign n66235 = ~n1924 ;
  assign n1925 = n1781 & n66235 ;
  assign n66236 = ~n1854 ;
  assign n1926 = n1784 & n66236 ;
  assign n1927 = n1925 | n1926 ;
  assign n1928 = n66219 & n1927 ;
  assign n1929 = n66222 & n1928 ;
  assign n1930 = n1923 | n1929 ;
  assign n1931 = n65791 & n1930 ;
  assign n1932 = n1722 & n1840 ;
  assign n1933 = n1732 | n1780 ;
  assign n66237 = ~n1933 ;
  assign n1934 = n1776 & n66237 ;
  assign n66238 = ~n1777 ;
  assign n1935 = n66238 & n1780 ;
  assign n1936 = n1934 | n1935 ;
  assign n1937 = n66219 & n1936 ;
  assign n1938 = n66222 & n1937 ;
  assign n1939 = n1932 | n1938 ;
  assign n1940 = n65772 & n1939 ;
  assign n1941 = n1731 & n1840 ;
  assign n1942 = n1742 | n1774 ;
  assign n66239 = ~n1942 ;
  assign n1943 = n1771 & n66239 ;
  assign n66240 = ~n1850 ;
  assign n1944 = n1774 & n66240 ;
  assign n1945 = n1943 | n1944 ;
  assign n1946 = n66219 & n1945 ;
  assign n1947 = n66222 & n1946 ;
  assign n1948 = n1941 | n1947 ;
  assign n1949 = n65746 & n1948 ;
  assign n1950 = n1741 & n1840 ;
  assign n66241 = ~n1766 ;
  assign n1951 = n66241 & n1770 ;
  assign n1952 = n1765 | n1770 ;
  assign n66242 = ~n1952 ;
  assign n1953 = n1763 & n66242 ;
  assign n1954 = n1951 | n1953 ;
  assign n1955 = n66219 & n1954 ;
  assign n1956 = n66222 & n1955 ;
  assign n1957 = n1950 | n1956 ;
  assign n1958 = n65721 & n1957 ;
  assign n1841 = n1764 & n1840 ;
  assign n1846 = n1760 & n1761 ;
  assign n1959 = n66188 & n1846 ;
  assign n1960 = n1839 | n1959 ;
  assign n66243 = ~n1960 ;
  assign n1961 = n1763 & n66243 ;
  assign n1962 = n66222 & n1961 ;
  assign n1963 = n1841 | n1962 ;
  assign n1964 = n65686 & n1963 ;
  assign n66244 = ~x78 ;
  assign n1965 = x64 & n66244 ;
  assign n66245 = ~n258 ;
  assign n1966 = n66245 & n1965 ;
  assign n66246 = ~n72910 ;
  assign n1967 = n66246 & n1966 ;
  assign n1968 = n65844 & n1967 ;
  assign n1969 = n65845 & n1968 ;
  assign n1974 = n66212 & n1973 ;
  assign n1975 = n1833 | n1974 ;
  assign n1976 = n66213 & n1975 ;
  assign n66247 = ~n1976 ;
  assign n1977 = n1969 & n66247 ;
  assign n66248 = ~n1977 ;
  assign n1978 = x50 & n66248 ;
  assign n1979 = n66183 & n1761 ;
  assign n1980 = n66184 & n1979 ;
  assign n1981 = n65776 & n1980 ;
  assign n1982 = n65777 & n1981 ;
  assign n1983 = n66222 & n1982 ;
  assign n1984 = n1978 | n1983 ;
  assign n1986 = x65 & n1984 ;
  assign n1970 = n66222 & n1969 ;
  assign n66249 = ~n1970 ;
  assign n1971 = x50 & n66249 ;
  assign n1985 = x65 | n1983 ;
  assign n1987 = n1971 | n1985 ;
  assign n66250 = ~n1986 ;
  assign n1988 = n66250 & n1987 ;
  assign n66251 = ~x49 ;
  assign n1989 = n66251 & x64 ;
  assign n1990 = n1988 | n1989 ;
  assign n1991 = n65670 & n1984 ;
  assign n66252 = ~n1991 ;
  assign n1992 = n1990 & n66252 ;
  assign n66253 = ~n1962 ;
  assign n1993 = x66 & n66253 ;
  assign n66254 = ~n1841 ;
  assign n1994 = n66254 & n1993 ;
  assign n1995 = n1964 | n1994 ;
  assign n1996 = n1992 | n1995 ;
  assign n66255 = ~n1964 ;
  assign n1997 = n66255 & n1996 ;
  assign n66256 = ~n1956 ;
  assign n1998 = x67 & n66256 ;
  assign n66257 = ~n1950 ;
  assign n1999 = n66257 & n1998 ;
  assign n2000 = n1997 | n1999 ;
  assign n66258 = ~n1958 ;
  assign n2001 = n66258 & n2000 ;
  assign n66259 = ~n1947 ;
  assign n2002 = x68 & n66259 ;
  assign n66260 = ~n1941 ;
  assign n2003 = n66260 & n2002 ;
  assign n2004 = n1949 | n2003 ;
  assign n2005 = n2001 | n2004 ;
  assign n66261 = ~n1949 ;
  assign n2006 = n66261 & n2005 ;
  assign n66262 = ~n1938 ;
  assign n2007 = x69 & n66262 ;
  assign n66263 = ~n1932 ;
  assign n2008 = n66263 & n2007 ;
  assign n2009 = n1940 | n2008 ;
  assign n2010 = n2006 | n2009 ;
  assign n66264 = ~n1940 ;
  assign n2011 = n66264 & n2010 ;
  assign n66265 = ~n1929 ;
  assign n2012 = x70 & n66265 ;
  assign n66266 = ~n1923 ;
  assign n2013 = n66266 & n2012 ;
  assign n2014 = n1931 | n2013 ;
  assign n2015 = n2011 | n2014 ;
  assign n66267 = ~n1931 ;
  assign n2016 = n66267 & n2015 ;
  assign n66268 = ~n1920 ;
  assign n2017 = x71 & n66268 ;
  assign n66269 = ~n1915 ;
  assign n2018 = n66269 & n2017 ;
  assign n2019 = n1922 | n2018 ;
  assign n2021 = n2016 | n2019 ;
  assign n66270 = ~n1922 ;
  assign n2022 = n66270 & n2021 ;
  assign n66271 = ~n1912 ;
  assign n2023 = x72 & n66271 ;
  assign n66272 = ~n1907 ;
  assign n2024 = n66272 & n2023 ;
  assign n2025 = n1914 | n2024 ;
  assign n2026 = n2022 | n2025 ;
  assign n66273 = ~n1914 ;
  assign n2027 = n66273 & n2026 ;
  assign n66274 = ~n1904 ;
  assign n2028 = x73 & n66274 ;
  assign n66275 = ~n1899 ;
  assign n2029 = n66275 & n2028 ;
  assign n2030 = n1906 | n2029 ;
  assign n2032 = n2027 | n2030 ;
  assign n66276 = ~n1906 ;
  assign n2033 = n66276 & n2032 ;
  assign n66277 = ~n1896 ;
  assign n2034 = x74 & n66277 ;
  assign n66278 = ~n1891 ;
  assign n2035 = n66278 & n2034 ;
  assign n2036 = n1898 | n2035 ;
  assign n2037 = n2033 | n2036 ;
  assign n66279 = ~n1898 ;
  assign n2038 = n66279 & n2037 ;
  assign n66280 = ~n1888 ;
  assign n2039 = x75 & n66280 ;
  assign n66281 = ~n1883 ;
  assign n2040 = n66281 & n2039 ;
  assign n2041 = n1890 | n2040 ;
  assign n2043 = n2038 | n2041 ;
  assign n66282 = ~n1890 ;
  assign n2044 = n66282 & n2043 ;
  assign n66283 = ~n1880 ;
  assign n2045 = x76 & n66283 ;
  assign n66284 = ~n1875 ;
  assign n2046 = n66284 & n2045 ;
  assign n2047 = n1882 | n2046 ;
  assign n2048 = n2044 | n2047 ;
  assign n66285 = ~n1882 ;
  assign n2049 = n66285 & n2048 ;
  assign n66286 = ~n1872 ;
  assign n2050 = x77 & n66286 ;
  assign n66287 = ~n1843 ;
  assign n2051 = n66287 & n2050 ;
  assign n2052 = n1874 | n2051 ;
  assign n2054 = n2049 | n2052 ;
  assign n66288 = ~n1874 ;
  assign n2055 = n66288 & n2054 ;
  assign n2062 = n66244 & n2061 ;
  assign n179 = ~n1840 ;
  assign n2063 = n179 & n2059 ;
  assign n2064 = n1650 & n1840 ;
  assign n66290 = ~n2064 ;
  assign n2065 = x78 & n66290 ;
  assign n66291 = ~n2063 ;
  assign n2066 = n66291 & n2065 ;
  assign n2067 = n72910 | n258 ;
  assign n2068 = n459 | n2067 ;
  assign n2069 = n469 | n2068 ;
  assign n2070 = n2066 | n2069 ;
  assign n2071 = n2062 | n2070 ;
  assign n2073 = n2055 | n2071 ;
  assign n66292 = ~n2072 ;
  assign n2074 = n66292 & n2073 ;
  assign n66293 = ~n2049 ;
  assign n2053 = n66293 & n2052 ;
  assign n2077 = n1971 | n1983 ;
  assign n2078 = x65 & n2077 ;
  assign n66294 = ~n2078 ;
  assign n2079 = n1987 & n66294 ;
  assign n2080 = n1989 | n2079 ;
  assign n2081 = n66252 & n2080 ;
  assign n2083 = n1994 | n2081 ;
  assign n2084 = n66255 & n2083 ;
  assign n2085 = n1958 | n1999 ;
  assign n2087 = n2084 | n2085 ;
  assign n2088 = n66258 & n2087 ;
  assign n2090 = n2004 | n2088 ;
  assign n2091 = n66261 & n2090 ;
  assign n2093 = n2009 | n2091 ;
  assign n2094 = n66264 & n2093 ;
  assign n2095 = n2014 | n2094 ;
  assign n2097 = n66267 & n2095 ;
  assign n2098 = n2019 | n2097 ;
  assign n2099 = n66270 & n2098 ;
  assign n2100 = n2025 | n2099 ;
  assign n2102 = n66273 & n2100 ;
  assign n2103 = n2030 | n2102 ;
  assign n2104 = n66276 & n2103 ;
  assign n2105 = n2036 | n2104 ;
  assign n2107 = n66279 & n2105 ;
  assign n2108 = n2041 | n2107 ;
  assign n2109 = n66282 & n2108 ;
  assign n2110 = n2047 | n2109 ;
  assign n2127 = n1882 | n2052 ;
  assign n66295 = ~n2127 ;
  assign n2128 = n2110 & n66295 ;
  assign n2129 = n2053 | n2128 ;
  assign n178 = ~n2074 ;
  assign n2130 = n178 & n2129 ;
  assign n2112 = n66285 & n2110 ;
  assign n2113 = n2052 | n2112 ;
  assign n2114 = n66288 & n2113 ;
  assign n2115 = n2071 | n2114 ;
  assign n2131 = n1873 & n66292 ;
  assign n2132 = n2115 & n2131 ;
  assign n2133 = n2130 | n2132 ;
  assign n2116 = n1874 | n2066 ;
  assign n2117 = n2062 | n2116 ;
  assign n66297 = ~n2117 ;
  assign n2118 = n2054 & n66297 ;
  assign n2119 = n2062 | n2066 ;
  assign n66298 = ~n2114 ;
  assign n2120 = n66298 & n2119 ;
  assign n2121 = n2118 | n2120 ;
  assign n2122 = n178 & n2121 ;
  assign n2123 = n1839 & n2061 ;
  assign n2124 = n2115 & n2123 ;
  assign n2125 = n2122 | n2124 ;
  assign n66299 = ~x79 ;
  assign n2126 = n66299 & n2125 ;
  assign n66300 = ~n2124 ;
  assign n2320 = x79 & n66300 ;
  assign n66301 = ~n2122 ;
  assign n2321 = n66301 & n2320 ;
  assign n2322 = n2126 | n2321 ;
  assign n2134 = n66244 & n2133 ;
  assign n66302 = ~n2109 ;
  assign n2111 = n2047 & n66302 ;
  assign n2135 = n1890 | n2047 ;
  assign n66303 = ~n2135 ;
  assign n2136 = n2043 & n66303 ;
  assign n2137 = n2111 | n2136 ;
  assign n2138 = n178 & n2137 ;
  assign n2139 = n1881 & n66292 ;
  assign n2140 = n2115 & n2139 ;
  assign n2141 = n2138 | n2140 ;
  assign n2142 = n66145 & n2141 ;
  assign n66304 = ~n2140 ;
  assign n2308 = x77 & n66304 ;
  assign n66305 = ~n2138 ;
  assign n2309 = n66305 & n2308 ;
  assign n2310 = n2142 | n2309 ;
  assign n66306 = ~n2038 ;
  assign n2042 = n66306 & n2041 ;
  assign n2143 = n1898 | n2041 ;
  assign n66307 = ~n2143 ;
  assign n2144 = n2105 & n66307 ;
  assign n2145 = n2042 | n2144 ;
  assign n2146 = n178 & n2145 ;
  assign n2147 = n1889 & n66292 ;
  assign n2148 = n2115 & n2147 ;
  assign n2149 = n2146 | n2148 ;
  assign n2150 = n66081 & n2149 ;
  assign n66308 = ~n2104 ;
  assign n2106 = n2036 & n66308 ;
  assign n2151 = n1906 | n2036 ;
  assign n66309 = ~n2151 ;
  assign n2152 = n2032 & n66309 ;
  assign n2153 = n2106 | n2152 ;
  assign n2154 = n178 & n2153 ;
  assign n2155 = n1897 & n66292 ;
  assign n2156 = n2115 & n2155 ;
  assign n2157 = n2154 | n2156 ;
  assign n2158 = n66043 & n2157 ;
  assign n66310 = ~n2156 ;
  assign n2296 = x75 & n66310 ;
  assign n66311 = ~n2154 ;
  assign n2297 = n66311 & n2296 ;
  assign n2298 = n2158 | n2297 ;
  assign n66312 = ~n2027 ;
  assign n2031 = n66312 & n2030 ;
  assign n2159 = n1914 | n2030 ;
  assign n66313 = ~n2159 ;
  assign n2160 = n2100 & n66313 ;
  assign n2161 = n2031 | n2160 ;
  assign n2162 = n178 & n2161 ;
  assign n2163 = n1905 & n66292 ;
  assign n2164 = n2115 & n2163 ;
  assign n2165 = n2162 | n2164 ;
  assign n2166 = n65960 & n2165 ;
  assign n66314 = ~n2099 ;
  assign n2101 = n2025 & n66314 ;
  assign n2167 = n1922 | n2025 ;
  assign n66315 = ~n2167 ;
  assign n2168 = n2021 & n66315 ;
  assign n2169 = n2101 | n2168 ;
  assign n2170 = n178 & n2169 ;
  assign n2171 = n1913 & n66292 ;
  assign n2172 = n2115 & n2171 ;
  assign n2173 = n2170 | n2172 ;
  assign n2174 = n65909 & n2173 ;
  assign n66316 = ~n2172 ;
  assign n2284 = x73 & n66316 ;
  assign n66317 = ~n2170 ;
  assign n2285 = n66317 & n2284 ;
  assign n2286 = n2174 | n2285 ;
  assign n66318 = ~n2016 ;
  assign n2020 = n66318 & n2019 ;
  assign n2175 = n1931 | n2019 ;
  assign n66319 = ~n2175 ;
  assign n2176 = n2095 & n66319 ;
  assign n2177 = n2020 | n2176 ;
  assign n2178 = n178 & n2177 ;
  assign n2179 = n1921 & n66292 ;
  assign n2180 = n2115 & n2179 ;
  assign n2181 = n2178 | n2180 ;
  assign n2182 = n65877 & n2181 ;
  assign n66320 = ~n2094 ;
  assign n2096 = n2014 & n66320 ;
  assign n2183 = n1940 | n2014 ;
  assign n66321 = ~n2183 ;
  assign n2184 = n2010 & n66321 ;
  assign n2185 = n2096 | n2184 ;
  assign n2186 = n178 & n2185 ;
  assign n2187 = n1930 & n66292 ;
  assign n2188 = n2115 & n2187 ;
  assign n2189 = n2186 | n2188 ;
  assign n2190 = n65820 & n2189 ;
  assign n66322 = ~n2188 ;
  assign n2272 = x71 & n66322 ;
  assign n66323 = ~n2186 ;
  assign n2273 = n66323 & n2272 ;
  assign n2274 = n2190 | n2273 ;
  assign n66324 = ~n2006 ;
  assign n2092 = n66324 & n2009 ;
  assign n2191 = n1949 | n2009 ;
  assign n66325 = ~n2191 ;
  assign n2192 = n2090 & n66325 ;
  assign n2193 = n2092 | n2192 ;
  assign n2194 = n178 & n2193 ;
  assign n2195 = n1939 & n66292 ;
  assign n2196 = n2115 & n2195 ;
  assign n2197 = n2194 | n2196 ;
  assign n2198 = n65791 & n2197 ;
  assign n66326 = ~n2088 ;
  assign n2089 = n2004 & n66326 ;
  assign n2199 = n1997 | n2085 ;
  assign n2200 = n1958 | n2004 ;
  assign n66327 = ~n2200 ;
  assign n2201 = n2199 & n66327 ;
  assign n2202 = n2089 | n2201 ;
  assign n2203 = n178 & n2202 ;
  assign n2204 = n1948 & n66292 ;
  assign n2205 = n2115 & n2204 ;
  assign n2206 = n2203 | n2205 ;
  assign n2207 = n65772 & n2206 ;
  assign n66328 = ~n2205 ;
  assign n2261 = x69 & n66328 ;
  assign n66329 = ~n2203 ;
  assign n2262 = n66329 & n2261 ;
  assign n2263 = n2207 | n2262 ;
  assign n66330 = ~n1997 ;
  assign n2086 = n66330 & n2085 ;
  assign n2208 = n1964 | n2085 ;
  assign n66331 = ~n2208 ;
  assign n2209 = n1996 & n66331 ;
  assign n2210 = n2086 | n2209 ;
  assign n2211 = n178 & n2210 ;
  assign n2212 = n1957 & n66292 ;
  assign n2213 = n2115 & n2212 ;
  assign n2214 = n2211 | n2213 ;
  assign n2215 = n65746 & n2214 ;
  assign n66332 = ~n2081 ;
  assign n2082 = n1995 & n66332 ;
  assign n2216 = n1991 | n1995 ;
  assign n66333 = ~n2216 ;
  assign n2217 = n1990 & n66333 ;
  assign n2218 = n2082 | n2217 ;
  assign n2219 = n178 & n2218 ;
  assign n2220 = n1963 & n66292 ;
  assign n2221 = n2115 & n2220 ;
  assign n2222 = n2219 | n2221 ;
  assign n2223 = n65721 & n2222 ;
  assign n66334 = ~n2221 ;
  assign n2251 = x67 & n66334 ;
  assign n66335 = ~n2219 ;
  assign n2252 = n66335 & n2251 ;
  assign n2253 = n2223 | n2252 ;
  assign n2224 = n1987 & n1989 ;
  assign n2225 = n66250 & n2224 ;
  assign n66336 = ~n2225 ;
  assign n2226 = n2080 & n66336 ;
  assign n2227 = n178 & n2226 ;
  assign n2228 = n1984 & n66292 ;
  assign n2229 = n2115 & n2228 ;
  assign n2230 = n2227 | n2229 ;
  assign n2231 = n65686 & n2230 ;
  assign n66337 = ~x48 ;
  assign n2241 = n66337 & x64 ;
  assign n2075 = n1989 & n178 ;
  assign n2232 = n66292 & n2115 ;
  assign n66338 = ~n2232 ;
  assign n2233 = x64 & n66338 ;
  assign n66339 = ~n2233 ;
  assign n2234 = x49 & n66339 ;
  assign n2235 = n2075 | n2234 ;
  assign n2236 = x65 & n2235 ;
  assign n2076 = x64 & n178 ;
  assign n66340 = ~n2076 ;
  assign n2237 = x49 & n66340 ;
  assign n2238 = n1989 & n66338 ;
  assign n2239 = x65 | n2238 ;
  assign n2240 = n2237 | n2239 ;
  assign n66341 = ~n2236 ;
  assign n2242 = n66341 & n2240 ;
  assign n2243 = n2241 | n2242 ;
  assign n2244 = n2075 | n2237 ;
  assign n2245 = n65670 & n2244 ;
  assign n66342 = ~n2245 ;
  assign n2246 = n2243 & n66342 ;
  assign n66343 = ~n2229 ;
  assign n2247 = x66 & n66343 ;
  assign n66344 = ~n2227 ;
  assign n2248 = n66344 & n2247 ;
  assign n2249 = n2231 | n2248 ;
  assign n2250 = n2246 | n2249 ;
  assign n66345 = ~n2231 ;
  assign n2254 = n66345 & n2250 ;
  assign n2255 = n2253 | n2254 ;
  assign n66346 = ~n2223 ;
  assign n2256 = n66346 & n2255 ;
  assign n66347 = ~n2213 ;
  assign n2257 = x68 & n66347 ;
  assign n66348 = ~n2211 ;
  assign n2258 = n66348 & n2257 ;
  assign n2259 = n2215 | n2258 ;
  assign n2260 = n2256 | n2259 ;
  assign n66349 = ~n2215 ;
  assign n2264 = n66349 & n2260 ;
  assign n2265 = n2263 | n2264 ;
  assign n66350 = ~n2207 ;
  assign n2266 = n66350 & n2265 ;
  assign n66351 = ~n2196 ;
  assign n2267 = x70 & n66351 ;
  assign n66352 = ~n2194 ;
  assign n2268 = n66352 & n2267 ;
  assign n2269 = n2198 | n2268 ;
  assign n2271 = n2266 | n2269 ;
  assign n66353 = ~n2198 ;
  assign n2276 = n66353 & n2271 ;
  assign n2277 = n2274 | n2276 ;
  assign n66354 = ~n2190 ;
  assign n2278 = n66354 & n2277 ;
  assign n66355 = ~n2180 ;
  assign n2279 = x72 & n66355 ;
  assign n66356 = ~n2178 ;
  assign n2280 = n66356 & n2279 ;
  assign n2281 = n2182 | n2280 ;
  assign n2283 = n2278 | n2281 ;
  assign n66357 = ~n2182 ;
  assign n2288 = n66357 & n2283 ;
  assign n2289 = n2286 | n2288 ;
  assign n66358 = ~n2174 ;
  assign n2290 = n66358 & n2289 ;
  assign n66359 = ~n2164 ;
  assign n2291 = x74 & n66359 ;
  assign n66360 = ~n2162 ;
  assign n2292 = n66360 & n2291 ;
  assign n2293 = n2166 | n2292 ;
  assign n2295 = n2290 | n2293 ;
  assign n66361 = ~n2166 ;
  assign n2300 = n66361 & n2295 ;
  assign n2301 = n2298 | n2300 ;
  assign n66362 = ~n2158 ;
  assign n2302 = n66362 & n2301 ;
  assign n66363 = ~n2148 ;
  assign n2303 = x76 & n66363 ;
  assign n66364 = ~n2146 ;
  assign n2304 = n66364 & n2303 ;
  assign n2305 = n2150 | n2304 ;
  assign n2307 = n2302 | n2305 ;
  assign n66365 = ~n2150 ;
  assign n2312 = n66365 & n2307 ;
  assign n2313 = n2310 | n2312 ;
  assign n66366 = ~n2142 ;
  assign n2314 = n66366 & n2313 ;
  assign n66367 = ~n2132 ;
  assign n2315 = x78 & n66367 ;
  assign n66368 = ~n2130 ;
  assign n2316 = n66368 & n2315 ;
  assign n2317 = n2134 | n2316 ;
  assign n2319 = n2314 | n2317 ;
  assign n66369 = ~n2134 ;
  assign n2323 = n66369 & n2319 ;
  assign n2324 = n2322 | n2323 ;
  assign n66370 = ~n2126 ;
  assign n2325 = n66370 & n2324 ;
  assign n2326 = n67897 | n2325 ;
  assign n2369 = n2133 & n2326 ;
  assign n2318 = n2142 | n2317 ;
  assign n2330 = x65 & n2244 ;
  assign n66371 = ~n2330 ;
  assign n2331 = n2240 & n66371 ;
  assign n2333 = n2241 | n2331 ;
  assign n2335 = n66342 & n2333 ;
  assign n2336 = n2249 | n2335 ;
  assign n2337 = n66345 & n2336 ;
  assign n2338 = n2253 | n2337 ;
  assign n2339 = n66346 & n2338 ;
  assign n2340 = n2259 | n2339 ;
  assign n2341 = n66349 & n2340 ;
  assign n2342 = n2263 | n2341 ;
  assign n2343 = n66350 & n2342 ;
  assign n2344 = n2269 | n2343 ;
  assign n2345 = n66353 & n2344 ;
  assign n2346 = n2274 | n2345 ;
  assign n2347 = n66354 & n2346 ;
  assign n2348 = n2281 | n2347 ;
  assign n2349 = n66357 & n2348 ;
  assign n2350 = n2286 | n2349 ;
  assign n2351 = n66358 & n2350 ;
  assign n2352 = n2293 | n2351 ;
  assign n2353 = n66361 & n2352 ;
  assign n2354 = n2298 | n2353 ;
  assign n2355 = n66362 & n2354 ;
  assign n2356 = n2305 | n2355 ;
  assign n2357 = n66365 & n2356 ;
  assign n2358 = n2310 | n2357 ;
  assign n66372 = ~n2318 ;
  assign n2370 = n66372 & n2358 ;
  assign n66373 = ~n2314 ;
  assign n2371 = n66373 & n2317 ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = n65678 & n2372 ;
  assign n66374 = ~n2325 ;
  assign n2374 = n66374 & n2373 ;
  assign n2375 = n2369 | n2374 ;
  assign n66375 = ~n2125 ;
  assign n2327 = n66375 & n2326 ;
  assign n66376 = ~n2323 ;
  assign n2362 = n2322 & n66376 ;
  assign n2359 = n66366 & n2358 ;
  assign n2360 = n2317 | n2359 ;
  assign n2363 = n2134 | n2322 ;
  assign n66377 = ~n2363 ;
  assign n2364 = n2360 & n66377 ;
  assign n2365 = n2362 | n2364 ;
  assign n2366 = n2326 | n2365 ;
  assign n66378 = ~n2327 ;
  assign n2367 = n66378 & n2366 ;
  assign n66379 = ~x80 ;
  assign n2368 = n66379 & n2367 ;
  assign n2376 = n66299 & n2375 ;
  assign n2377 = n2141 & n2326 ;
  assign n2311 = n2150 | n2310 ;
  assign n66380 = ~n2311 ;
  assign n2378 = n2307 & n66380 ;
  assign n66381 = ~n2357 ;
  assign n2379 = n2310 & n66381 ;
  assign n2380 = n2378 | n2379 ;
  assign n2381 = n65678 & n2380 ;
  assign n2382 = n66374 & n2381 ;
  assign n2383 = n2377 | n2382 ;
  assign n2384 = n66244 & n2383 ;
  assign n2385 = n2149 & n2326 ;
  assign n2306 = n2158 | n2305 ;
  assign n66382 = ~n2306 ;
  assign n2386 = n66382 & n2354 ;
  assign n66383 = ~n2302 ;
  assign n2387 = n66383 & n2305 ;
  assign n2388 = n2386 | n2387 ;
  assign n2389 = n65678 & n2388 ;
  assign n2390 = n66374 & n2389 ;
  assign n2391 = n2385 | n2390 ;
  assign n2392 = n66145 & n2391 ;
  assign n2393 = n2157 & n2326 ;
  assign n2299 = n2166 | n2298 ;
  assign n66384 = ~n2299 ;
  assign n2394 = n2295 & n66384 ;
  assign n66385 = ~n2353 ;
  assign n2395 = n2298 & n66385 ;
  assign n2396 = n2394 | n2395 ;
  assign n2397 = n65678 & n2396 ;
  assign n2398 = n66374 & n2397 ;
  assign n2399 = n2393 | n2398 ;
  assign n2400 = n66081 & n2399 ;
  assign n2401 = n2165 & n2326 ;
  assign n2294 = n2174 | n2293 ;
  assign n66386 = ~n2294 ;
  assign n2402 = n66386 & n2350 ;
  assign n66387 = ~n2290 ;
  assign n2403 = n66387 & n2293 ;
  assign n2404 = n2402 | n2403 ;
  assign n2405 = n65678 & n2404 ;
  assign n2406 = n66374 & n2405 ;
  assign n2407 = n2401 | n2406 ;
  assign n2408 = n66043 & n2407 ;
  assign n2409 = n2173 & n2326 ;
  assign n2287 = n2182 | n2286 ;
  assign n66388 = ~n2287 ;
  assign n2410 = n2283 & n66388 ;
  assign n66389 = ~n2349 ;
  assign n2411 = n2286 & n66389 ;
  assign n2412 = n2410 | n2411 ;
  assign n2413 = n65678 & n2412 ;
  assign n2414 = n66374 & n2413 ;
  assign n2415 = n2409 | n2414 ;
  assign n2416 = n65960 & n2415 ;
  assign n2417 = n2181 & n2326 ;
  assign n2282 = n2190 | n2281 ;
  assign n66390 = ~n2282 ;
  assign n2418 = n66390 & n2346 ;
  assign n66391 = ~n2278 ;
  assign n2419 = n66391 & n2281 ;
  assign n2420 = n2418 | n2419 ;
  assign n2421 = n65678 & n2420 ;
  assign n2422 = n66374 & n2421 ;
  assign n2423 = n2417 | n2422 ;
  assign n2424 = n65909 & n2423 ;
  assign n2425 = n2189 & n2326 ;
  assign n2275 = n2198 | n2274 ;
  assign n66392 = ~n2275 ;
  assign n2426 = n2271 & n66392 ;
  assign n66393 = ~n2345 ;
  assign n2427 = n2274 & n66393 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n65678 & n2428 ;
  assign n2430 = n66374 & n2429 ;
  assign n2431 = n2425 | n2430 ;
  assign n2432 = n65877 & n2431 ;
  assign n2433 = n2197 & n2326 ;
  assign n2270 = n2207 | n2269 ;
  assign n66394 = ~n2270 ;
  assign n2434 = n66394 & n2342 ;
  assign n66395 = ~n2266 ;
  assign n2435 = n66395 & n2269 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n65678 & n2436 ;
  assign n2438 = n66374 & n2437 ;
  assign n2439 = n2433 | n2438 ;
  assign n2440 = n65820 & n2439 ;
  assign n2441 = n2206 & n2326 ;
  assign n2329 = n2215 | n2263 ;
  assign n66396 = ~n2329 ;
  assign n2442 = n2260 & n66396 ;
  assign n66397 = ~n2341 ;
  assign n2443 = n2263 & n66397 ;
  assign n2444 = n2442 | n2443 ;
  assign n2445 = n65678 & n2444 ;
  assign n2446 = n66374 & n2445 ;
  assign n2447 = n2441 | n2446 ;
  assign n2448 = n65791 & n2447 ;
  assign n2449 = n2214 & n2326 ;
  assign n2450 = n2223 | n2259 ;
  assign n66398 = ~n2450 ;
  assign n2451 = n2338 & n66398 ;
  assign n66399 = ~n2256 ;
  assign n2452 = n66399 & n2259 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = n65678 & n2453 ;
  assign n2455 = n66374 & n2454 ;
  assign n2456 = n2449 | n2455 ;
  assign n2457 = n65772 & n2456 ;
  assign n2458 = n2222 & n2326 ;
  assign n2459 = n2231 | n2253 ;
  assign n66400 = ~n2459 ;
  assign n2460 = n2336 & n66400 ;
  assign n66401 = ~n2337 ;
  assign n2461 = n2253 & n66401 ;
  assign n2462 = n2460 | n2461 ;
  assign n2463 = n65678 & n2462 ;
  assign n2464 = n66374 & n2463 ;
  assign n2465 = n2458 | n2464 ;
  assign n2466 = n65746 & n2465 ;
  assign n2467 = n2230 & n2326 ;
  assign n2334 = n2245 | n2249 ;
  assign n66402 = ~n2334 ;
  assign n2468 = n2243 & n66402 ;
  assign n66403 = ~n2246 ;
  assign n2469 = n66403 & n2249 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = n65678 & n2470 ;
  assign n2472 = n66374 & n2471 ;
  assign n2473 = n2467 | n2472 ;
  assign n2474 = n65721 & n2473 ;
  assign n2328 = n2244 & n2326 ;
  assign n2332 = n2240 & n2241 ;
  assign n2475 = n66341 & n2332 ;
  assign n2476 = n67897 | n2475 ;
  assign n66404 = ~n2476 ;
  assign n2477 = n2243 & n66404 ;
  assign n2478 = n66374 & n2477 ;
  assign n2479 = n2328 | n2478 ;
  assign n2480 = n65686 & n2479 ;
  assign n2487 = n66184 & n2241 ;
  assign n2488 = n65776 & n2487 ;
  assign n2489 = n65777 & n2488 ;
  assign n2490 = n66374 & n2489 ;
  assign n2481 = x64 & n66379 ;
  assign n2482 = n66246 & n2481 ;
  assign n2483 = n65844 & n2482 ;
  assign n2484 = n65845 & n2483 ;
  assign n2361 = n66369 & n2360 ;
  assign n2498 = n2322 | n2361 ;
  assign n2499 = n66370 & n2498 ;
  assign n66405 = ~n2499 ;
  assign n2500 = n2484 & n66405 ;
  assign n66406 = ~n2500 ;
  assign n2501 = x48 & n66406 ;
  assign n2502 = n2490 | n2501 ;
  assign n2503 = n65670 & n2502 ;
  assign n2485 = n66374 & n2484 ;
  assign n66407 = ~n2485 ;
  assign n2486 = x48 & n66407 ;
  assign n2491 = n2486 | n2490 ;
  assign n2492 = x65 & n2491 ;
  assign n2494 = x65 | n2490 ;
  assign n2495 = n2486 | n2494 ;
  assign n66408 = ~n2492 ;
  assign n2496 = n66408 & n2495 ;
  assign n66409 = ~x47 ;
  assign n2497 = n66409 & x64 ;
  assign n2504 = n2496 | n2497 ;
  assign n66410 = ~n2503 ;
  assign n2505 = n66410 & n2504 ;
  assign n66411 = ~n2478 ;
  assign n2506 = x66 & n66411 ;
  assign n66412 = ~n2328 ;
  assign n2507 = n66412 & n2506 ;
  assign n2508 = n2480 | n2507 ;
  assign n2509 = n2505 | n2508 ;
  assign n66413 = ~n2480 ;
  assign n2510 = n66413 & n2509 ;
  assign n66414 = ~n2472 ;
  assign n2511 = x67 & n66414 ;
  assign n66415 = ~n2467 ;
  assign n2512 = n66415 & n2511 ;
  assign n2513 = n2474 | n2512 ;
  assign n2514 = n2510 | n2513 ;
  assign n66416 = ~n2474 ;
  assign n2515 = n66416 & n2514 ;
  assign n66417 = ~n2464 ;
  assign n2516 = x68 & n66417 ;
  assign n66418 = ~n2458 ;
  assign n2517 = n66418 & n2516 ;
  assign n2518 = n2466 | n2517 ;
  assign n2519 = n2515 | n2518 ;
  assign n66419 = ~n2466 ;
  assign n2520 = n66419 & n2519 ;
  assign n66420 = ~n2455 ;
  assign n2521 = x69 & n66420 ;
  assign n66421 = ~n2449 ;
  assign n2522 = n66421 & n2521 ;
  assign n2523 = n2457 | n2522 ;
  assign n2524 = n2520 | n2523 ;
  assign n66422 = ~n2457 ;
  assign n2525 = n66422 & n2524 ;
  assign n66423 = ~n2446 ;
  assign n2526 = x70 & n66423 ;
  assign n66424 = ~n2441 ;
  assign n2527 = n66424 & n2526 ;
  assign n2528 = n2448 | n2527 ;
  assign n2530 = n2525 | n2528 ;
  assign n66425 = ~n2448 ;
  assign n2531 = n66425 & n2530 ;
  assign n66426 = ~n2438 ;
  assign n2532 = x71 & n66426 ;
  assign n66427 = ~n2433 ;
  assign n2533 = n66427 & n2532 ;
  assign n2534 = n2440 | n2533 ;
  assign n2535 = n2531 | n2534 ;
  assign n66428 = ~n2440 ;
  assign n2536 = n66428 & n2535 ;
  assign n66429 = ~n2430 ;
  assign n2537 = x72 & n66429 ;
  assign n66430 = ~n2425 ;
  assign n2538 = n66430 & n2537 ;
  assign n2539 = n2432 | n2538 ;
  assign n2541 = n2536 | n2539 ;
  assign n66431 = ~n2432 ;
  assign n2542 = n66431 & n2541 ;
  assign n66432 = ~n2422 ;
  assign n2543 = x73 & n66432 ;
  assign n66433 = ~n2417 ;
  assign n2544 = n66433 & n2543 ;
  assign n2545 = n2424 | n2544 ;
  assign n2546 = n2542 | n2545 ;
  assign n66434 = ~n2424 ;
  assign n2547 = n66434 & n2546 ;
  assign n66435 = ~n2414 ;
  assign n2548 = x74 & n66435 ;
  assign n66436 = ~n2409 ;
  assign n2549 = n66436 & n2548 ;
  assign n2550 = n2416 | n2549 ;
  assign n2552 = n2547 | n2550 ;
  assign n66437 = ~n2416 ;
  assign n2553 = n66437 & n2552 ;
  assign n66438 = ~n2406 ;
  assign n2554 = x75 & n66438 ;
  assign n66439 = ~n2401 ;
  assign n2555 = n66439 & n2554 ;
  assign n2556 = n2408 | n2555 ;
  assign n2557 = n2553 | n2556 ;
  assign n66440 = ~n2408 ;
  assign n2558 = n66440 & n2557 ;
  assign n66441 = ~n2398 ;
  assign n2559 = x76 & n66441 ;
  assign n66442 = ~n2393 ;
  assign n2560 = n66442 & n2559 ;
  assign n2561 = n2400 | n2560 ;
  assign n2563 = n2558 | n2561 ;
  assign n66443 = ~n2400 ;
  assign n2564 = n66443 & n2563 ;
  assign n66444 = ~n2390 ;
  assign n2565 = x77 & n66444 ;
  assign n66445 = ~n2385 ;
  assign n2566 = n66445 & n2565 ;
  assign n2567 = n2392 | n2566 ;
  assign n2568 = n2564 | n2567 ;
  assign n66446 = ~n2392 ;
  assign n2569 = n66446 & n2568 ;
  assign n66447 = ~n2382 ;
  assign n2570 = x78 & n66447 ;
  assign n66448 = ~n2377 ;
  assign n2571 = n66448 & n2570 ;
  assign n2572 = n2384 | n2571 ;
  assign n2574 = n2569 | n2572 ;
  assign n66449 = ~n2384 ;
  assign n2575 = n66449 & n2574 ;
  assign n66450 = ~n2374 ;
  assign n2576 = x79 & n66450 ;
  assign n66451 = ~n2369 ;
  assign n2577 = n66451 & n2576 ;
  assign n2578 = n2376 | n2577 ;
  assign n2579 = n2575 | n2578 ;
  assign n66452 = ~n2376 ;
  assign n2580 = n66452 & n2579 ;
  assign n177 = ~n2326 ;
  assign n2581 = n177 & n2365 ;
  assign n2582 = n2125 & n2326 ;
  assign n66454 = ~n2582 ;
  assign n2583 = x80 & n66454 ;
  assign n66455 = ~n2581 ;
  assign n2584 = n66455 & n2583 ;
  assign n2585 = n2368 | n2584 ;
  assign n2587 = n2580 | n2585 ;
  assign n66456 = ~n2368 ;
  assign n2588 = n66456 & n2587 ;
  assign n2589 = n344 | n2588 ;
  assign n2591 = n2375 & n2589 ;
  assign n2493 = n65670 & n2491 ;
  assign n2592 = x65 & n2502 ;
  assign n66457 = ~n2592 ;
  assign n2593 = n2495 & n66457 ;
  assign n2594 = n2497 | n2593 ;
  assign n66458 = ~n2493 ;
  assign n2595 = n66458 & n2594 ;
  assign n2596 = n2508 | n2595 ;
  assign n2597 = n66413 & n2596 ;
  assign n2598 = n2512 | n2597 ;
  assign n2600 = n66416 & n2598 ;
  assign n2602 = n2518 | n2600 ;
  assign n2603 = n66419 & n2602 ;
  assign n2605 = n2523 | n2603 ;
  assign n2606 = n66422 & n2605 ;
  assign n2607 = n2528 | n2606 ;
  assign n2608 = n66425 & n2607 ;
  assign n2609 = n2534 | n2608 ;
  assign n2611 = n66428 & n2609 ;
  assign n2612 = n2539 | n2611 ;
  assign n2613 = n66431 & n2612 ;
  assign n2614 = n2545 | n2613 ;
  assign n2616 = n66434 & n2614 ;
  assign n2617 = n2550 | n2616 ;
  assign n2618 = n66437 & n2617 ;
  assign n2619 = n2556 | n2618 ;
  assign n2621 = n66440 & n2619 ;
  assign n2622 = n2561 | n2621 ;
  assign n2623 = n66443 & n2622 ;
  assign n2624 = n2567 | n2623 ;
  assign n2626 = n66446 & n2624 ;
  assign n2627 = n2572 | n2626 ;
  assign n2628 = n66449 & n2627 ;
  assign n66459 = ~n2628 ;
  assign n2629 = n2578 & n66459 ;
  assign n2631 = n2384 | n2578 ;
  assign n66460 = ~n2631 ;
  assign n2632 = n2574 & n66460 ;
  assign n2633 = n2629 | n2632 ;
  assign n2634 = n65715 & n2633 ;
  assign n66461 = ~n2588 ;
  assign n2635 = n66461 & n2634 ;
  assign n2636 = n2591 | n2635 ;
  assign n2637 = n66379 & n2636 ;
  assign n66462 = ~n2635 ;
  assign n2855 = x80 & n66462 ;
  assign n66463 = ~n2591 ;
  assign n2856 = n66463 & n2855 ;
  assign n2857 = n2637 | n2856 ;
  assign n2638 = n2383 & n2589 ;
  assign n66464 = ~n2569 ;
  assign n2573 = n66464 & n2572 ;
  assign n2639 = n2392 | n2572 ;
  assign n66465 = ~n2639 ;
  assign n2640 = n2624 & n66465 ;
  assign n2641 = n2573 | n2640 ;
  assign n2642 = n65715 & n2641 ;
  assign n2643 = n66461 & n2642 ;
  assign n2644 = n2638 | n2643 ;
  assign n2645 = n66299 & n2644 ;
  assign n2646 = n2391 & n2589 ;
  assign n66466 = ~n2623 ;
  assign n2625 = n2567 & n66466 ;
  assign n2647 = n2400 | n2567 ;
  assign n66467 = ~n2647 ;
  assign n2648 = n2563 & n66467 ;
  assign n2649 = n2625 | n2648 ;
  assign n2650 = n65715 & n2649 ;
  assign n2651 = n66461 & n2650 ;
  assign n2652 = n2646 | n2651 ;
  assign n2653 = n66244 & n2652 ;
  assign n66468 = ~n2651 ;
  assign n2844 = x78 & n66468 ;
  assign n66469 = ~n2646 ;
  assign n2845 = n66469 & n2844 ;
  assign n2846 = n2653 | n2845 ;
  assign n2654 = n2399 & n2589 ;
  assign n66470 = ~n2558 ;
  assign n2562 = n66470 & n2561 ;
  assign n2655 = n2408 | n2561 ;
  assign n66471 = ~n2655 ;
  assign n2656 = n2619 & n66471 ;
  assign n2657 = n2562 | n2656 ;
  assign n2658 = n65715 & n2657 ;
  assign n2659 = n66461 & n2658 ;
  assign n2660 = n2654 | n2659 ;
  assign n2661 = n66145 & n2660 ;
  assign n2662 = n2407 & n2589 ;
  assign n66472 = ~n2618 ;
  assign n2620 = n2556 & n66472 ;
  assign n2663 = n2416 | n2556 ;
  assign n66473 = ~n2663 ;
  assign n2664 = n2552 & n66473 ;
  assign n2665 = n2620 | n2664 ;
  assign n2666 = n65715 & n2665 ;
  assign n2667 = n66461 & n2666 ;
  assign n2668 = n2662 | n2667 ;
  assign n2669 = n66081 & n2668 ;
  assign n66474 = ~n2667 ;
  assign n2833 = x76 & n66474 ;
  assign n66475 = ~n2662 ;
  assign n2834 = n66475 & n2833 ;
  assign n2835 = n2669 | n2834 ;
  assign n2670 = n2415 & n2589 ;
  assign n66476 = ~n2547 ;
  assign n2551 = n66476 & n2550 ;
  assign n2671 = n2424 | n2550 ;
  assign n66477 = ~n2671 ;
  assign n2672 = n2614 & n66477 ;
  assign n2673 = n2551 | n2672 ;
  assign n2674 = n65715 & n2673 ;
  assign n2675 = n66461 & n2674 ;
  assign n2676 = n2670 | n2675 ;
  assign n2677 = n66043 & n2676 ;
  assign n2678 = n2423 & n2589 ;
  assign n66478 = ~n2613 ;
  assign n2615 = n2545 & n66478 ;
  assign n2679 = n2432 | n2545 ;
  assign n66479 = ~n2679 ;
  assign n2680 = n2541 & n66479 ;
  assign n2681 = n2615 | n2680 ;
  assign n2682 = n65715 & n2681 ;
  assign n2683 = n66461 & n2682 ;
  assign n2684 = n2678 | n2683 ;
  assign n2685 = n65960 & n2684 ;
  assign n66480 = ~n2683 ;
  assign n2821 = x74 & n66480 ;
  assign n66481 = ~n2678 ;
  assign n2822 = n66481 & n2821 ;
  assign n2823 = n2685 | n2822 ;
  assign n2686 = n2431 & n2589 ;
  assign n66482 = ~n2536 ;
  assign n2540 = n66482 & n2539 ;
  assign n2687 = n2440 | n2539 ;
  assign n66483 = ~n2687 ;
  assign n2688 = n2609 & n66483 ;
  assign n2689 = n2540 | n2688 ;
  assign n2690 = n65715 & n2689 ;
  assign n2691 = n66461 & n2690 ;
  assign n2692 = n2686 | n2691 ;
  assign n2693 = n65909 & n2692 ;
  assign n2694 = n2439 & n2589 ;
  assign n66484 = ~n2608 ;
  assign n2610 = n2534 & n66484 ;
  assign n2695 = n2448 | n2534 ;
  assign n66485 = ~n2695 ;
  assign n2696 = n2530 & n66485 ;
  assign n2697 = n2610 | n2696 ;
  assign n2698 = n65715 & n2697 ;
  assign n2699 = n66461 & n2698 ;
  assign n2700 = n2694 | n2699 ;
  assign n2701 = n65877 & n2700 ;
  assign n66486 = ~n2699 ;
  assign n2810 = x72 & n66486 ;
  assign n66487 = ~n2694 ;
  assign n2811 = n66487 & n2810 ;
  assign n2812 = n2701 | n2811 ;
  assign n2702 = n2447 & n2589 ;
  assign n66488 = ~n2525 ;
  assign n2529 = n66488 & n2528 ;
  assign n2703 = n2457 | n2528 ;
  assign n66489 = ~n2703 ;
  assign n2704 = n2605 & n66489 ;
  assign n2705 = n2529 | n2704 ;
  assign n2706 = n65715 & n2705 ;
  assign n2707 = n66461 & n2706 ;
  assign n2708 = n2702 | n2707 ;
  assign n2709 = n65820 & n2708 ;
  assign n2710 = n2456 & n2589 ;
  assign n66490 = ~n2603 ;
  assign n2604 = n2523 & n66490 ;
  assign n2711 = n2466 | n2523 ;
  assign n66491 = ~n2711 ;
  assign n2712 = n2602 & n66491 ;
  assign n2713 = n2604 | n2712 ;
  assign n2714 = n65715 & n2713 ;
  assign n2715 = n66461 & n2714 ;
  assign n2716 = n2710 | n2715 ;
  assign n2717 = n65791 & n2716 ;
  assign n66492 = ~n2715 ;
  assign n2799 = x70 & n66492 ;
  assign n66493 = ~n2710 ;
  assign n2800 = n66493 & n2799 ;
  assign n2801 = n2717 | n2800 ;
  assign n2718 = n2465 & n2589 ;
  assign n66494 = ~n2515 ;
  assign n2601 = n66494 & n2518 ;
  assign n2719 = n2513 | n2597 ;
  assign n2720 = n2474 | n2518 ;
  assign n66495 = ~n2720 ;
  assign n2721 = n2719 & n66495 ;
  assign n2722 = n2601 | n2721 ;
  assign n2723 = n65715 & n2722 ;
  assign n2724 = n66461 & n2723 ;
  assign n2725 = n2718 | n2724 ;
  assign n2726 = n65772 & n2725 ;
  assign n2727 = n2473 & n2589 ;
  assign n66496 = ~n2597 ;
  assign n2599 = n2513 & n66496 ;
  assign n2728 = n2480 | n2513 ;
  assign n66497 = ~n2728 ;
  assign n2729 = n2596 & n66497 ;
  assign n2730 = n2599 | n2729 ;
  assign n2731 = n65715 & n2730 ;
  assign n2732 = n66461 & n2731 ;
  assign n2733 = n2727 | n2732 ;
  assign n2734 = n65746 & n2733 ;
  assign n66498 = ~n2732 ;
  assign n2789 = x68 & n66498 ;
  assign n66499 = ~n2727 ;
  assign n2790 = n66499 & n2789 ;
  assign n2791 = n2734 | n2790 ;
  assign n2735 = n2479 & n2589 ;
  assign n2736 = n2503 | n2508 ;
  assign n66500 = ~n2736 ;
  assign n2737 = n2594 & n66500 ;
  assign n66501 = ~n2505 ;
  assign n2738 = n66501 & n2508 ;
  assign n2739 = n2737 | n2738 ;
  assign n2740 = n65715 & n2739 ;
  assign n2741 = n66461 & n2740 ;
  assign n2742 = n2735 | n2741 ;
  assign n2743 = n65721 & n2742 ;
  assign n2630 = n2578 | n2628 ;
  assign n2744 = n66452 & n2630 ;
  assign n2745 = n2585 | n2744 ;
  assign n2746 = n66456 & n2745 ;
  assign n2747 = n344 | n2746 ;
  assign n2748 = n2502 & n2747 ;
  assign n2749 = n2495 & n2497 ;
  assign n2750 = n66457 & n2749 ;
  assign n2751 = n344 | n2750 ;
  assign n66502 = ~n2751 ;
  assign n2752 = n2594 & n66502 ;
  assign n2753 = n66461 & n2752 ;
  assign n2754 = n2748 | n2753 ;
  assign n2755 = n65686 & n2754 ;
  assign n2776 = n2491 & n2589 ;
  assign n2777 = n2753 | n2776 ;
  assign n2778 = n65686 & n2777 ;
  assign n66503 = ~n2753 ;
  assign n2779 = x66 & n66503 ;
  assign n66504 = ~n2776 ;
  assign n2780 = n66504 & n2779 ;
  assign n2781 = n2778 | n2780 ;
  assign n66505 = ~x81 ;
  assign n2756 = x64 & n66505 ;
  assign n66506 = ~n65294 ;
  assign n2757 = n66506 & n2756 ;
  assign n66507 = ~n65587 ;
  assign n2758 = n66507 & n2757 ;
  assign n66508 = ~n67349 ;
  assign n2759 = n66508 & n2758 ;
  assign n66509 = ~n67215 ;
  assign n2760 = n66509 & n2759 ;
  assign n66510 = ~n66858 ;
  assign n2761 = n66510 & n2760 ;
  assign n66511 = ~n2746 ;
  assign n2762 = n66511 & n2761 ;
  assign n66512 = ~n2762 ;
  assign n2763 = x47 & n66512 ;
  assign n2764 = n66246 & n2497 ;
  assign n2765 = n65844 & n2764 ;
  assign n2766 = n65845 & n2765 ;
  assign n2767 = n66461 & n2766 ;
  assign n2768 = n2763 | n2767 ;
  assign n2769 = x65 & n2768 ;
  assign n2770 = x65 | n2767 ;
  assign n2771 = n2763 | n2770 ;
  assign n66513 = ~n2769 ;
  assign n2772 = n66513 & n2771 ;
  assign n66514 = ~x46 ;
  assign n2773 = n66514 & x64 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = n65670 & n2768 ;
  assign n66515 = ~n2775 ;
  assign n2782 = n2774 & n66515 ;
  assign n2783 = n2781 | n2782 ;
  assign n66516 = ~n2755 ;
  assign n2784 = n66516 & n2783 ;
  assign n66517 = ~n2741 ;
  assign n2785 = x67 & n66517 ;
  assign n66518 = ~n2735 ;
  assign n2786 = n66518 & n2785 ;
  assign n2787 = n2743 | n2786 ;
  assign n2788 = n2784 | n2787 ;
  assign n66519 = ~n2743 ;
  assign n2792 = n66519 & n2788 ;
  assign n2793 = n2791 | n2792 ;
  assign n66520 = ~n2734 ;
  assign n2794 = n66520 & n2793 ;
  assign n66521 = ~n2724 ;
  assign n2795 = x69 & n66521 ;
  assign n66522 = ~n2718 ;
  assign n2796 = n66522 & n2795 ;
  assign n2797 = n2726 | n2796 ;
  assign n2798 = n2794 | n2797 ;
  assign n66523 = ~n2726 ;
  assign n2802 = n66523 & n2798 ;
  assign n2803 = n2801 | n2802 ;
  assign n66524 = ~n2717 ;
  assign n2804 = n66524 & n2803 ;
  assign n66525 = ~n2707 ;
  assign n2805 = x71 & n66525 ;
  assign n66526 = ~n2702 ;
  assign n2806 = n66526 & n2805 ;
  assign n2807 = n2709 | n2806 ;
  assign n2809 = n2804 | n2807 ;
  assign n66527 = ~n2709 ;
  assign n2814 = n66527 & n2809 ;
  assign n2815 = n2812 | n2814 ;
  assign n66528 = ~n2701 ;
  assign n2816 = n66528 & n2815 ;
  assign n66529 = ~n2691 ;
  assign n2817 = x73 & n66529 ;
  assign n66530 = ~n2686 ;
  assign n2818 = n66530 & n2817 ;
  assign n2819 = n2693 | n2818 ;
  assign n2820 = n2816 | n2819 ;
  assign n66531 = ~n2693 ;
  assign n2825 = n66531 & n2820 ;
  assign n2826 = n2823 | n2825 ;
  assign n66532 = ~n2685 ;
  assign n2827 = n66532 & n2826 ;
  assign n66533 = ~n2675 ;
  assign n2828 = x75 & n66533 ;
  assign n66534 = ~n2670 ;
  assign n2829 = n66534 & n2828 ;
  assign n2830 = n2677 | n2829 ;
  assign n2832 = n2827 | n2830 ;
  assign n66535 = ~n2677 ;
  assign n2837 = n66535 & n2832 ;
  assign n2838 = n2835 | n2837 ;
  assign n66536 = ~n2669 ;
  assign n2839 = n66536 & n2838 ;
  assign n66537 = ~n2659 ;
  assign n2840 = x77 & n66537 ;
  assign n66538 = ~n2654 ;
  assign n2841 = n66538 & n2840 ;
  assign n2842 = n2661 | n2841 ;
  assign n2843 = n2839 | n2842 ;
  assign n66539 = ~n2661 ;
  assign n2848 = n66539 & n2843 ;
  assign n2849 = n2846 | n2848 ;
  assign n66540 = ~n2653 ;
  assign n2850 = n66540 & n2849 ;
  assign n66541 = ~n2643 ;
  assign n2851 = x79 & n66541 ;
  assign n66542 = ~n2638 ;
  assign n2852 = n66542 & n2851 ;
  assign n2853 = n2645 | n2852 ;
  assign n2854 = n2850 | n2853 ;
  assign n66543 = ~n2645 ;
  assign n2859 = n66543 & n2854 ;
  assign n2860 = n2857 | n2859 ;
  assign n66544 = ~n2637 ;
  assign n2861 = n66544 & n2860 ;
  assign n66545 = ~n2367 ;
  assign n2590 = n66545 & n2589 ;
  assign n66546 = ~n2580 ;
  assign n2586 = n66546 & n2585 ;
  assign n2862 = n2376 | n2585 ;
  assign n66547 = ~n2862 ;
  assign n2863 = n2630 & n66547 ;
  assign n2864 = n2586 | n2863 ;
  assign n2865 = n2589 | n2864 ;
  assign n66548 = ~n2590 ;
  assign n2866 = n66548 & n2865 ;
  assign n2867 = n66505 & n2866 ;
  assign n176 = ~n2589 ;
  assign n2868 = n176 & n2864 ;
  assign n2869 = n2367 & n2589 ;
  assign n66550 = ~n2869 ;
  assign n2870 = x81 & n66550 ;
  assign n66551 = ~n2868 ;
  assign n2871 = n66551 & n2870 ;
  assign n2872 = n65294 | n65587 ;
  assign n2873 = n67349 | n2872 ;
  assign n2874 = n67215 | n2873 ;
  assign n2875 = n66858 | n2874 ;
  assign n2876 = n2871 | n2875 ;
  assign n2877 = n2867 | n2876 ;
  assign n2878 = n2861 | n2877 ;
  assign n2879 = n65715 & n2866 ;
  assign n66552 = ~n2879 ;
  assign n2880 = n2878 & n66552 ;
  assign n2882 = n2637 | n2871 ;
  assign n2883 = n2867 | n2882 ;
  assign n66553 = ~n2883 ;
  assign n2884 = n2860 & n66553 ;
  assign n2885 = n66461 & n2761 ;
  assign n66554 = ~n2885 ;
  assign n2886 = x47 & n66554 ;
  assign n2887 = n2767 | n2886 ;
  assign n2888 = x65 & n2887 ;
  assign n66555 = ~n2888 ;
  assign n2889 = n2771 & n66555 ;
  assign n2890 = n2773 | n2889 ;
  assign n2891 = n66515 & n2890 ;
  assign n66556 = ~n2748 ;
  assign n2892 = n66556 & n2779 ;
  assign n2893 = n2755 | n2892 ;
  assign n2894 = n2891 | n2893 ;
  assign n66557 = ~n2778 ;
  assign n2895 = n66557 & n2894 ;
  assign n2896 = n2787 | n2895 ;
  assign n2897 = n66519 & n2896 ;
  assign n2898 = n2791 | n2897 ;
  assign n2899 = n66520 & n2898 ;
  assign n2900 = n2797 | n2899 ;
  assign n2901 = n66523 & n2900 ;
  assign n2902 = n2801 | n2901 ;
  assign n2903 = n66524 & n2902 ;
  assign n2904 = n2807 | n2903 ;
  assign n2905 = n66527 & n2904 ;
  assign n2906 = n2812 | n2905 ;
  assign n2907 = n66528 & n2906 ;
  assign n2908 = n2819 | n2907 ;
  assign n2909 = n66531 & n2908 ;
  assign n2910 = n2823 | n2909 ;
  assign n2911 = n66532 & n2910 ;
  assign n2912 = n2830 | n2911 ;
  assign n2913 = n66535 & n2912 ;
  assign n2914 = n2835 | n2913 ;
  assign n2915 = n66536 & n2914 ;
  assign n2916 = n2842 | n2915 ;
  assign n2917 = n66539 & n2916 ;
  assign n2918 = n2846 | n2917 ;
  assign n2919 = n66540 & n2918 ;
  assign n2920 = n2853 | n2919 ;
  assign n2921 = n66543 & n2920 ;
  assign n2922 = n2857 | n2921 ;
  assign n2923 = n66544 & n2922 ;
  assign n2924 = n2867 | n2871 ;
  assign n66558 = ~n2923 ;
  assign n2925 = n66558 & n2924 ;
  assign n2926 = n2884 | n2925 ;
  assign n175 = ~n2880 ;
  assign n2927 = n175 & n2926 ;
  assign n2928 = n344 & n2367 ;
  assign n2929 = n2878 & n2928 ;
  assign n2930 = n2927 | n2929 ;
  assign n66560 = ~x82 ;
  assign n2931 = n66560 & n2930 ;
  assign n66561 = ~n2859 ;
  assign n2932 = n2857 & n66561 ;
  assign n2858 = n2645 | n2857 ;
  assign n66562 = ~n2858 ;
  assign n2933 = n2854 & n66562 ;
  assign n2934 = n2932 | n2933 ;
  assign n2935 = n175 & n2934 ;
  assign n2936 = n2636 & n66552 ;
  assign n2937 = n2878 & n2936 ;
  assign n2938 = n2935 | n2937 ;
  assign n2939 = n66505 & n2938 ;
  assign n66563 = ~n2919 ;
  assign n2940 = n2853 & n66563 ;
  assign n2941 = n2653 | n2853 ;
  assign n66564 = ~n2941 ;
  assign n2942 = n2849 & n66564 ;
  assign n2943 = n2940 | n2942 ;
  assign n2944 = n175 & n2943 ;
  assign n2945 = n2644 & n66552 ;
  assign n2946 = n2878 & n2945 ;
  assign n2947 = n2944 | n2946 ;
  assign n2948 = n66379 & n2947 ;
  assign n66565 = ~n2848 ;
  assign n2949 = n2846 & n66565 ;
  assign n2847 = n2661 | n2846 ;
  assign n66566 = ~n2847 ;
  assign n2950 = n2843 & n66566 ;
  assign n2951 = n2949 | n2950 ;
  assign n2952 = n175 & n2951 ;
  assign n2953 = n2652 & n66552 ;
  assign n2954 = n2878 & n2953 ;
  assign n2955 = n2952 | n2954 ;
  assign n2956 = n66299 & n2955 ;
  assign n66567 = ~n2915 ;
  assign n2957 = n2842 & n66567 ;
  assign n2958 = n2669 | n2842 ;
  assign n66568 = ~n2958 ;
  assign n2959 = n2838 & n66568 ;
  assign n2960 = n2957 | n2959 ;
  assign n2961 = n175 & n2960 ;
  assign n2962 = n2660 & n66552 ;
  assign n2963 = n2878 & n2962 ;
  assign n2964 = n2961 | n2963 ;
  assign n2965 = n66244 & n2964 ;
  assign n66569 = ~n2837 ;
  assign n2966 = n2835 & n66569 ;
  assign n2836 = n2677 | n2835 ;
  assign n66570 = ~n2836 ;
  assign n2967 = n2832 & n66570 ;
  assign n2968 = n2966 | n2967 ;
  assign n2969 = n175 & n2968 ;
  assign n2970 = n2668 & n66552 ;
  assign n2971 = n2878 & n2970 ;
  assign n2972 = n2969 | n2971 ;
  assign n2973 = n66145 & n2972 ;
  assign n66571 = ~n2911 ;
  assign n2974 = n2830 & n66571 ;
  assign n2831 = n2685 | n2830 ;
  assign n66572 = ~n2831 ;
  assign n2975 = n66572 & n2910 ;
  assign n2976 = n2974 | n2975 ;
  assign n2977 = n175 & n2976 ;
  assign n2978 = n2676 & n66552 ;
  assign n2979 = n2878 & n2978 ;
  assign n2980 = n2977 | n2979 ;
  assign n2981 = n66081 & n2980 ;
  assign n66573 = ~n2825 ;
  assign n2982 = n2823 & n66573 ;
  assign n2824 = n2693 | n2823 ;
  assign n66574 = ~n2824 ;
  assign n2983 = n2820 & n66574 ;
  assign n2984 = n2982 | n2983 ;
  assign n2985 = n175 & n2984 ;
  assign n2986 = n2684 & n66552 ;
  assign n2987 = n2878 & n2986 ;
  assign n2988 = n2985 | n2987 ;
  assign n2989 = n66043 & n2988 ;
  assign n66575 = ~n2907 ;
  assign n2990 = n2819 & n66575 ;
  assign n2991 = n2701 | n2819 ;
  assign n66576 = ~n2991 ;
  assign n2992 = n2815 & n66576 ;
  assign n2993 = n2990 | n2992 ;
  assign n2994 = n175 & n2993 ;
  assign n2995 = n2692 & n66552 ;
  assign n2996 = n2878 & n2995 ;
  assign n2997 = n2994 | n2996 ;
  assign n2998 = n65960 & n2997 ;
  assign n66577 = ~n2814 ;
  assign n2999 = n2812 & n66577 ;
  assign n2813 = n2709 | n2812 ;
  assign n66578 = ~n2813 ;
  assign n3000 = n2809 & n66578 ;
  assign n3001 = n2999 | n3000 ;
  assign n3002 = n175 & n3001 ;
  assign n3003 = n2700 & n66552 ;
  assign n3004 = n2878 & n3003 ;
  assign n3005 = n3002 | n3004 ;
  assign n3006 = n65909 & n3005 ;
  assign n66579 = ~n2903 ;
  assign n3007 = n2807 & n66579 ;
  assign n2808 = n2717 | n2807 ;
  assign n66580 = ~n2808 ;
  assign n3008 = n66580 & n2902 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = n175 & n3009 ;
  assign n3011 = n2708 & n66552 ;
  assign n3012 = n2878 & n3011 ;
  assign n3013 = n3010 | n3012 ;
  assign n3014 = n65877 & n3013 ;
  assign n66581 = ~n2802 ;
  assign n3015 = n2801 & n66581 ;
  assign n3016 = n2726 | n2801 ;
  assign n66582 = ~n3016 ;
  assign n3017 = n2900 & n66582 ;
  assign n3018 = n3015 | n3017 ;
  assign n3019 = n175 & n3018 ;
  assign n3020 = n2716 & n66552 ;
  assign n3021 = n2878 & n3020 ;
  assign n3022 = n3019 | n3021 ;
  assign n3023 = n65820 & n3022 ;
  assign n66583 = ~n2899 ;
  assign n3025 = n2797 & n66583 ;
  assign n3024 = n2734 | n2797 ;
  assign n66584 = ~n3024 ;
  assign n3026 = n2898 & n66584 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = n175 & n3027 ;
  assign n3029 = n2725 & n66552 ;
  assign n3030 = n2878 & n3029 ;
  assign n3031 = n3028 | n3030 ;
  assign n3032 = n65791 & n3031 ;
  assign n66585 = ~n2792 ;
  assign n3034 = n2791 & n66585 ;
  assign n3033 = n2743 | n2791 ;
  assign n66586 = ~n3033 ;
  assign n3035 = n2788 & n66586 ;
  assign n3036 = n3034 | n3035 ;
  assign n3037 = n175 & n3036 ;
  assign n3038 = n2733 & n66552 ;
  assign n3039 = n2878 & n3038 ;
  assign n3040 = n3037 | n3039 ;
  assign n3041 = n65772 & n3040 ;
  assign n3042 = n66516 & n2894 ;
  assign n66587 = ~n3042 ;
  assign n3044 = n2787 & n66587 ;
  assign n3043 = n2755 | n2787 ;
  assign n66588 = ~n3043 ;
  assign n3045 = n2894 & n66588 ;
  assign n3046 = n3044 | n3045 ;
  assign n3047 = n175 & n3046 ;
  assign n3048 = n2742 & n66552 ;
  assign n3049 = n2878 & n3048 ;
  assign n3050 = n3047 | n3049 ;
  assign n3051 = n65746 & n3050 ;
  assign n66589 = ~n2782 ;
  assign n3052 = n66589 & n2893 ;
  assign n3053 = n2775 | n2893 ;
  assign n66590 = ~n3053 ;
  assign n3054 = n2890 & n66590 ;
  assign n3055 = n3052 | n3054 ;
  assign n3056 = n175 & n3055 ;
  assign n3057 = n2754 & n66552 ;
  assign n3058 = n2878 & n3057 ;
  assign n3059 = n3056 | n3058 ;
  assign n3060 = n65721 & n3059 ;
  assign n3061 = n2771 & n2773 ;
  assign n3062 = n66513 & n3061 ;
  assign n66591 = ~n3062 ;
  assign n3063 = n2774 & n66591 ;
  assign n3064 = n175 & n3063 ;
  assign n3065 = n2768 & n66552 ;
  assign n3066 = n2878 & n3065 ;
  assign n3067 = n3064 | n3066 ;
  assign n3068 = n65686 & n3067 ;
  assign n2881 = n2773 & n175 ;
  assign n3069 = x64 & n175 ;
  assign n66592 = ~n3069 ;
  assign n3070 = x46 & n66592 ;
  assign n3071 = n2881 | n3070 ;
  assign n3082 = n65670 & n3071 ;
  assign n3072 = n2877 | n2923 ;
  assign n3073 = n66552 & n3072 ;
  assign n66593 = ~n3073 ;
  assign n3074 = x64 & n66593 ;
  assign n66594 = ~n3074 ;
  assign n3075 = x46 & n66594 ;
  assign n3076 = n2881 | n3075 ;
  assign n3077 = x65 & n3076 ;
  assign n3078 = x65 | n2881 ;
  assign n3079 = n3075 | n3078 ;
  assign n66595 = ~n3077 ;
  assign n3080 = n66595 & n3079 ;
  assign n66596 = ~x45 ;
  assign n3081 = n66596 & x64 ;
  assign n3083 = n3080 | n3081 ;
  assign n66597 = ~n3082 ;
  assign n3084 = n66597 & n3083 ;
  assign n66598 = ~n3066 ;
  assign n3085 = x66 & n66598 ;
  assign n66599 = ~n3064 ;
  assign n3086 = n66599 & n3085 ;
  assign n3087 = n3068 | n3086 ;
  assign n3088 = n3084 | n3087 ;
  assign n66600 = ~n3068 ;
  assign n3089 = n66600 & n3088 ;
  assign n66601 = ~n3058 ;
  assign n3090 = x67 & n66601 ;
  assign n66602 = ~n3056 ;
  assign n3091 = n66602 & n3090 ;
  assign n3092 = n3060 | n3091 ;
  assign n3093 = n3089 | n3092 ;
  assign n66603 = ~n3060 ;
  assign n3094 = n66603 & n3093 ;
  assign n66604 = ~n3049 ;
  assign n3095 = x68 & n66604 ;
  assign n66605 = ~n3047 ;
  assign n3096 = n66605 & n3095 ;
  assign n3097 = n3051 | n3096 ;
  assign n3098 = n3094 | n3097 ;
  assign n66606 = ~n3051 ;
  assign n3099 = n66606 & n3098 ;
  assign n66607 = ~n3039 ;
  assign n3100 = x69 & n66607 ;
  assign n66608 = ~n3037 ;
  assign n3101 = n66608 & n3100 ;
  assign n3102 = n3041 | n3101 ;
  assign n3103 = n3099 | n3102 ;
  assign n66609 = ~n3041 ;
  assign n3104 = n66609 & n3103 ;
  assign n66610 = ~n3030 ;
  assign n3105 = x70 & n66610 ;
  assign n66611 = ~n3028 ;
  assign n3106 = n66611 & n3105 ;
  assign n3107 = n3032 | n3106 ;
  assign n3109 = n3104 | n3107 ;
  assign n66612 = ~n3032 ;
  assign n3110 = n66612 & n3109 ;
  assign n66613 = ~n3021 ;
  assign n3111 = x71 & n66613 ;
  assign n66614 = ~n3019 ;
  assign n3112 = n66614 & n3111 ;
  assign n3113 = n3023 | n3112 ;
  assign n3114 = n3110 | n3113 ;
  assign n66615 = ~n3023 ;
  assign n3115 = n66615 & n3114 ;
  assign n66616 = ~n3012 ;
  assign n3116 = x72 & n66616 ;
  assign n66617 = ~n3010 ;
  assign n3117 = n66617 & n3116 ;
  assign n3118 = n3014 | n3117 ;
  assign n3120 = n3115 | n3118 ;
  assign n66618 = ~n3014 ;
  assign n3121 = n66618 & n3120 ;
  assign n66619 = ~n3004 ;
  assign n3122 = x73 & n66619 ;
  assign n66620 = ~n3002 ;
  assign n3123 = n66620 & n3122 ;
  assign n3124 = n3006 | n3123 ;
  assign n3125 = n3121 | n3124 ;
  assign n66621 = ~n3006 ;
  assign n3126 = n66621 & n3125 ;
  assign n66622 = ~n2996 ;
  assign n3127 = x74 & n66622 ;
  assign n66623 = ~n2994 ;
  assign n3128 = n66623 & n3127 ;
  assign n3129 = n2998 | n3128 ;
  assign n3131 = n3126 | n3129 ;
  assign n66624 = ~n2998 ;
  assign n3132 = n66624 & n3131 ;
  assign n66625 = ~n2987 ;
  assign n3133 = x75 & n66625 ;
  assign n66626 = ~n2985 ;
  assign n3134 = n66626 & n3133 ;
  assign n3135 = n2989 | n3134 ;
  assign n3136 = n3132 | n3135 ;
  assign n66627 = ~n2989 ;
  assign n3137 = n66627 & n3136 ;
  assign n66628 = ~n2979 ;
  assign n3138 = x76 & n66628 ;
  assign n66629 = ~n2977 ;
  assign n3139 = n66629 & n3138 ;
  assign n3140 = n2981 | n3139 ;
  assign n3142 = n3137 | n3140 ;
  assign n66630 = ~n2981 ;
  assign n3143 = n66630 & n3142 ;
  assign n66631 = ~n2971 ;
  assign n3144 = x77 & n66631 ;
  assign n66632 = ~n2969 ;
  assign n3145 = n66632 & n3144 ;
  assign n3146 = n2973 | n3145 ;
  assign n3147 = n3143 | n3146 ;
  assign n66633 = ~n2973 ;
  assign n3148 = n66633 & n3147 ;
  assign n66634 = ~n2963 ;
  assign n3149 = x78 & n66634 ;
  assign n66635 = ~n2961 ;
  assign n3150 = n66635 & n3149 ;
  assign n3151 = n2965 | n3150 ;
  assign n3153 = n3148 | n3151 ;
  assign n66636 = ~n2965 ;
  assign n3154 = n66636 & n3153 ;
  assign n66637 = ~n2954 ;
  assign n3155 = x79 & n66637 ;
  assign n66638 = ~n2952 ;
  assign n3156 = n66638 & n3155 ;
  assign n3157 = n2956 | n3156 ;
  assign n3158 = n3154 | n3157 ;
  assign n66639 = ~n2956 ;
  assign n3159 = n66639 & n3158 ;
  assign n66640 = ~n2946 ;
  assign n3160 = x80 & n66640 ;
  assign n66641 = ~n2944 ;
  assign n3161 = n66641 & n3160 ;
  assign n3162 = n2948 | n3161 ;
  assign n3164 = n3159 | n3162 ;
  assign n66642 = ~n2948 ;
  assign n3165 = n66642 & n3164 ;
  assign n66643 = ~n2937 ;
  assign n3166 = x81 & n66643 ;
  assign n66644 = ~n2935 ;
  assign n3167 = n66644 & n3166 ;
  assign n3168 = n2939 | n3167 ;
  assign n3169 = n3165 | n3168 ;
  assign n66645 = ~n2939 ;
  assign n3170 = n66645 & n3169 ;
  assign n66646 = ~n2929 ;
  assign n3171 = x82 & n66646 ;
  assign n66647 = ~n2927 ;
  assign n3172 = n66647 & n3171 ;
  assign n3173 = n2931 | n3172 ;
  assign n3175 = n3170 | n3173 ;
  assign n66648 = ~n2931 ;
  assign n3176 = n66648 & n3175 ;
  assign n3177 = n72130 | n72392 ;
  assign n3178 = n74914 | n3177 ;
  assign n3179 = n294 | n3178 ;
  assign n3180 = n279 | n3179 ;
  assign n3181 = n3176 | n3180 ;
  assign n66649 = ~n2930 ;
  assign n3182 = n66649 & n3181 ;
  assign n66650 = ~n3170 ;
  assign n3174 = n66650 & n3173 ;
  assign n3185 = x65 & n3071 ;
  assign n66651 = ~n3185 ;
  assign n3186 = n3079 & n66651 ;
  assign n3187 = n3081 | n3186 ;
  assign n3188 = n66597 & n3187 ;
  assign n3189 = n3087 | n3188 ;
  assign n3190 = n66600 & n3189 ;
  assign n3191 = n3091 | n3190 ;
  assign n3193 = n66603 & n3191 ;
  assign n3195 = n3097 | n3193 ;
  assign n3196 = n66606 & n3195 ;
  assign n3197 = n3102 | n3196 ;
  assign n3199 = n66609 & n3197 ;
  assign n3200 = n3107 | n3199 ;
  assign n3201 = n66612 & n3200 ;
  assign n3202 = n3113 | n3201 ;
  assign n3204 = n66615 & n3202 ;
  assign n3205 = n3118 | n3204 ;
  assign n3206 = n66618 & n3205 ;
  assign n3207 = n3124 | n3206 ;
  assign n3209 = n66621 & n3207 ;
  assign n3210 = n3129 | n3209 ;
  assign n3211 = n66624 & n3210 ;
  assign n3212 = n3135 | n3211 ;
  assign n3214 = n66627 & n3212 ;
  assign n3215 = n3140 | n3214 ;
  assign n3216 = n66630 & n3215 ;
  assign n3217 = n3146 | n3216 ;
  assign n3219 = n66633 & n3217 ;
  assign n3220 = n3151 | n3219 ;
  assign n3221 = n66636 & n3220 ;
  assign n3222 = n3157 | n3221 ;
  assign n3224 = n66639 & n3222 ;
  assign n3225 = n3162 | n3224 ;
  assign n3226 = n66642 & n3225 ;
  assign n3228 = n3168 | n3226 ;
  assign n3229 = n2939 | n3173 ;
  assign n66652 = ~n3229 ;
  assign n3230 = n3228 & n66652 ;
  assign n3231 = n3174 | n3230 ;
  assign n3232 = n3181 | n3231 ;
  assign n66653 = ~n3182 ;
  assign n3233 = n66653 & n3232 ;
  assign n66654 = ~x83 ;
  assign n3234 = n66654 & n3233 ;
  assign n174 = ~n3181 ;
  assign n3496 = n174 & n3231 ;
  assign n3497 = n2930 & n3181 ;
  assign n66656 = ~n3497 ;
  assign n3498 = x83 & n66656 ;
  assign n66657 = ~n3496 ;
  assign n3499 = n66657 & n3498 ;
  assign n3500 = n3234 | n3499 ;
  assign n3235 = n2938 & n3181 ;
  assign n66658 = ~n3226 ;
  assign n3227 = n3168 & n66658 ;
  assign n3236 = n2948 | n3168 ;
  assign n66659 = ~n3236 ;
  assign n3237 = n3164 & n66659 ;
  assign n3238 = n3227 | n3237 ;
  assign n66660 = ~n3180 ;
  assign n3239 = n66660 & n3238 ;
  assign n66661 = ~n3176 ;
  assign n3240 = n66661 & n3239 ;
  assign n3241 = n3235 | n3240 ;
  assign n3242 = n66560 & n3241 ;
  assign n3243 = n2947 & n3181 ;
  assign n66662 = ~n3159 ;
  assign n3163 = n66662 & n3162 ;
  assign n3244 = n2956 | n3162 ;
  assign n66663 = ~n3244 ;
  assign n3245 = n3222 & n66663 ;
  assign n3246 = n3163 | n3245 ;
  assign n3247 = n66660 & n3246 ;
  assign n3248 = n66661 & n3247 ;
  assign n3249 = n3243 | n3248 ;
  assign n3250 = n66505 & n3249 ;
  assign n66664 = ~n3248 ;
  assign n3484 = x81 & n66664 ;
  assign n66665 = ~n3243 ;
  assign n3485 = n66665 & n3484 ;
  assign n3486 = n3250 | n3485 ;
  assign n3251 = n2955 & n3181 ;
  assign n66666 = ~n3221 ;
  assign n3223 = n3157 & n66666 ;
  assign n3252 = n2965 | n3157 ;
  assign n66667 = ~n3252 ;
  assign n3253 = n3153 & n66667 ;
  assign n3254 = n3223 | n3253 ;
  assign n3255 = n66660 & n3254 ;
  assign n3256 = n66661 & n3255 ;
  assign n3257 = n3251 | n3256 ;
  assign n3258 = n66379 & n3257 ;
  assign n3259 = n2964 & n3181 ;
  assign n66668 = ~n3148 ;
  assign n3152 = n66668 & n3151 ;
  assign n3260 = n2973 | n3151 ;
  assign n66669 = ~n3260 ;
  assign n3261 = n3217 & n66669 ;
  assign n3262 = n3152 | n3261 ;
  assign n3263 = n66660 & n3262 ;
  assign n3264 = n66661 & n3263 ;
  assign n3265 = n3259 | n3264 ;
  assign n3266 = n66299 & n3265 ;
  assign n66670 = ~n3264 ;
  assign n3472 = x79 & n66670 ;
  assign n66671 = ~n3259 ;
  assign n3473 = n66671 & n3472 ;
  assign n3474 = n3266 | n3473 ;
  assign n3267 = n2972 & n3181 ;
  assign n66672 = ~n3216 ;
  assign n3218 = n3146 & n66672 ;
  assign n3268 = n2981 | n3146 ;
  assign n66673 = ~n3268 ;
  assign n3269 = n3142 & n66673 ;
  assign n3270 = n3218 | n3269 ;
  assign n3271 = n66660 & n3270 ;
  assign n3272 = n66661 & n3271 ;
  assign n3273 = n3267 | n3272 ;
  assign n3274 = n66244 & n3273 ;
  assign n3275 = n2980 & n3181 ;
  assign n66674 = ~n3137 ;
  assign n3141 = n66674 & n3140 ;
  assign n3276 = n2989 | n3140 ;
  assign n66675 = ~n3276 ;
  assign n3277 = n3212 & n66675 ;
  assign n3278 = n3141 | n3277 ;
  assign n3279 = n66660 & n3278 ;
  assign n3280 = n66661 & n3279 ;
  assign n3281 = n3275 | n3280 ;
  assign n3282 = n66145 & n3281 ;
  assign n66676 = ~n3280 ;
  assign n3460 = x77 & n66676 ;
  assign n66677 = ~n3275 ;
  assign n3461 = n66677 & n3460 ;
  assign n3462 = n3282 | n3461 ;
  assign n3283 = n2988 & n3181 ;
  assign n66678 = ~n3211 ;
  assign n3213 = n3135 & n66678 ;
  assign n3284 = n2998 | n3135 ;
  assign n66679 = ~n3284 ;
  assign n3285 = n3131 & n66679 ;
  assign n3286 = n3213 | n3285 ;
  assign n3287 = n66660 & n3286 ;
  assign n3288 = n66661 & n3287 ;
  assign n3289 = n3283 | n3288 ;
  assign n3290 = n66081 & n3289 ;
  assign n3291 = n2997 & n3181 ;
  assign n66680 = ~n3126 ;
  assign n3130 = n66680 & n3129 ;
  assign n3292 = n3006 | n3129 ;
  assign n66681 = ~n3292 ;
  assign n3293 = n3207 & n66681 ;
  assign n3294 = n3130 | n3293 ;
  assign n3295 = n66660 & n3294 ;
  assign n3296 = n66661 & n3295 ;
  assign n3297 = n3291 | n3296 ;
  assign n3298 = n66043 & n3297 ;
  assign n66682 = ~n3296 ;
  assign n3448 = x75 & n66682 ;
  assign n66683 = ~n3291 ;
  assign n3449 = n66683 & n3448 ;
  assign n3450 = n3298 | n3449 ;
  assign n3299 = n3005 & n3181 ;
  assign n66684 = ~n3206 ;
  assign n3208 = n3124 & n66684 ;
  assign n3300 = n3014 | n3124 ;
  assign n66685 = ~n3300 ;
  assign n3301 = n3120 & n66685 ;
  assign n3302 = n3208 | n3301 ;
  assign n3303 = n66660 & n3302 ;
  assign n3304 = n66661 & n3303 ;
  assign n3305 = n3299 | n3304 ;
  assign n3306 = n65960 & n3305 ;
  assign n3307 = n3013 & n3181 ;
  assign n66686 = ~n3115 ;
  assign n3119 = n66686 & n3118 ;
  assign n3308 = n3023 | n3118 ;
  assign n66687 = ~n3308 ;
  assign n3309 = n3202 & n66687 ;
  assign n3310 = n3119 | n3309 ;
  assign n3311 = n66660 & n3310 ;
  assign n3312 = n66661 & n3311 ;
  assign n3313 = n3307 | n3312 ;
  assign n3314 = n65909 & n3313 ;
  assign n66688 = ~n3312 ;
  assign n3436 = x73 & n66688 ;
  assign n66689 = ~n3307 ;
  assign n3437 = n66689 & n3436 ;
  assign n3438 = n3314 | n3437 ;
  assign n3315 = n3022 & n3181 ;
  assign n66690 = ~n3201 ;
  assign n3203 = n3113 & n66690 ;
  assign n3316 = n3032 | n3113 ;
  assign n66691 = ~n3316 ;
  assign n3317 = n3109 & n66691 ;
  assign n3318 = n3203 | n3317 ;
  assign n3319 = n66660 & n3318 ;
  assign n3320 = n66661 & n3319 ;
  assign n3321 = n3315 | n3320 ;
  assign n3322 = n65877 & n3321 ;
  assign n3323 = n3031 & n3181 ;
  assign n66692 = ~n3104 ;
  assign n3108 = n66692 & n3107 ;
  assign n3324 = n3041 | n3107 ;
  assign n66693 = ~n3324 ;
  assign n3325 = n3197 & n66693 ;
  assign n3326 = n3108 | n3325 ;
  assign n3327 = n66660 & n3326 ;
  assign n3328 = n66661 & n3327 ;
  assign n3329 = n3323 | n3328 ;
  assign n3330 = n65820 & n3329 ;
  assign n66694 = ~n3328 ;
  assign n3424 = x71 & n66694 ;
  assign n66695 = ~n3323 ;
  assign n3425 = n66695 & n3424 ;
  assign n3426 = n3330 | n3425 ;
  assign n3331 = n3040 & n3181 ;
  assign n66696 = ~n3196 ;
  assign n3198 = n3102 & n66696 ;
  assign n3332 = n3051 | n3102 ;
  assign n66697 = ~n3332 ;
  assign n3333 = n3098 & n66697 ;
  assign n3334 = n3198 | n3333 ;
  assign n3335 = n66660 & n3334 ;
  assign n3336 = n66661 & n3335 ;
  assign n3337 = n3331 | n3336 ;
  assign n3338 = n65791 & n3337 ;
  assign n3339 = n3050 & n3181 ;
  assign n66698 = ~n3094 ;
  assign n3194 = n66698 & n3097 ;
  assign n3340 = n3092 | n3190 ;
  assign n3341 = n3060 | n3097 ;
  assign n66699 = ~n3341 ;
  assign n3342 = n3340 & n66699 ;
  assign n3343 = n3194 | n3342 ;
  assign n3344 = n66660 & n3343 ;
  assign n3345 = n66661 & n3344 ;
  assign n3346 = n3339 | n3345 ;
  assign n3347 = n65772 & n3346 ;
  assign n66700 = ~n3345 ;
  assign n3413 = x69 & n66700 ;
  assign n66701 = ~n3339 ;
  assign n3414 = n66701 & n3413 ;
  assign n3415 = n3347 | n3414 ;
  assign n3183 = n3059 & n3181 ;
  assign n66702 = ~n3190 ;
  assign n3192 = n3092 & n66702 ;
  assign n3348 = n3068 | n3092 ;
  assign n66703 = ~n3348 ;
  assign n3349 = n3189 & n66703 ;
  assign n3350 = n3192 | n3349 ;
  assign n3351 = n66660 & n3350 ;
  assign n3352 = n66661 & n3351 ;
  assign n3353 = n3183 | n3352 ;
  assign n3354 = n65746 & n3353 ;
  assign n3184 = n3067 & n3181 ;
  assign n3355 = n3082 | n3087 ;
  assign n66704 = ~n3355 ;
  assign n3356 = n3187 & n66704 ;
  assign n66705 = ~n3084 ;
  assign n3357 = n66705 & n3087 ;
  assign n3358 = n3356 | n3357 ;
  assign n3359 = n66660 & n3358 ;
  assign n3360 = n66661 & n3359 ;
  assign n3361 = n3184 | n3360 ;
  assign n3362 = n65721 & n3361 ;
  assign n66706 = ~n3360 ;
  assign n3403 = x67 & n66706 ;
  assign n66707 = ~n3184 ;
  assign n3404 = n66707 & n3403 ;
  assign n3405 = n3362 | n3404 ;
  assign n3363 = n3076 & n3181 ;
  assign n3364 = n3079 & n3081 ;
  assign n3365 = n66651 & n3364 ;
  assign n3366 = n3180 | n3365 ;
  assign n66708 = ~n3366 ;
  assign n3367 = n3187 & n66708 ;
  assign n3368 = n66661 & n3367 ;
  assign n3369 = n3363 | n3368 ;
  assign n3370 = n65686 & n3369 ;
  assign n66709 = ~x44 ;
  assign n3393 = n66709 & x64 ;
  assign n3371 = x64 & n66654 ;
  assign n3372 = n66507 & n3371 ;
  assign n3373 = n66508 & n3372 ;
  assign n3374 = n66509 & n3373 ;
  assign n3375 = n66510 & n3374 ;
  assign n3376 = n66661 & n3375 ;
  assign n66710 = ~n3376 ;
  assign n3377 = x45 & n66710 ;
  assign n66711 = ~n72392 ;
  assign n3378 = n66711 & n3081 ;
  assign n66712 = ~n72130 ;
  assign n3379 = n66712 & n3378 ;
  assign n66713 = ~n74914 ;
  assign n3380 = n66713 & n3379 ;
  assign n66714 = ~n294 ;
  assign n3381 = n66714 & n3380 ;
  assign n66715 = ~n279 ;
  assign n3382 = n66715 & n3381 ;
  assign n3383 = n66661 & n3382 ;
  assign n3384 = n3377 | n3383 ;
  assign n3385 = x65 & n3384 ;
  assign n3386 = n66645 & n3228 ;
  assign n3387 = n3173 | n3386 ;
  assign n3388 = n66648 & n3387 ;
  assign n66716 = ~n3388 ;
  assign n3389 = n3375 & n66716 ;
  assign n66717 = ~n3389 ;
  assign n3390 = x45 & n66717 ;
  assign n3391 = x65 | n3383 ;
  assign n3392 = n3390 | n3391 ;
  assign n66718 = ~n3385 ;
  assign n3394 = n66718 & n3392 ;
  assign n3395 = n3393 | n3394 ;
  assign n3396 = n3383 | n3390 ;
  assign n3397 = n65670 & n3396 ;
  assign n66719 = ~n3397 ;
  assign n3398 = n3395 & n66719 ;
  assign n66720 = ~n3368 ;
  assign n3399 = x66 & n66720 ;
  assign n66721 = ~n3363 ;
  assign n3400 = n66721 & n3399 ;
  assign n3401 = n3370 | n3400 ;
  assign n3402 = n3398 | n3401 ;
  assign n66722 = ~n3370 ;
  assign n3406 = n66722 & n3402 ;
  assign n3407 = n3405 | n3406 ;
  assign n66723 = ~n3362 ;
  assign n3408 = n66723 & n3407 ;
  assign n66724 = ~n3352 ;
  assign n3409 = x68 & n66724 ;
  assign n66725 = ~n3183 ;
  assign n3410 = n66725 & n3409 ;
  assign n3411 = n3354 | n3410 ;
  assign n3412 = n3408 | n3411 ;
  assign n66726 = ~n3354 ;
  assign n3416 = n66726 & n3412 ;
  assign n3417 = n3415 | n3416 ;
  assign n66727 = ~n3347 ;
  assign n3418 = n66727 & n3417 ;
  assign n66728 = ~n3336 ;
  assign n3419 = x70 & n66728 ;
  assign n66729 = ~n3331 ;
  assign n3420 = n66729 & n3419 ;
  assign n3421 = n3338 | n3420 ;
  assign n3423 = n3418 | n3421 ;
  assign n66730 = ~n3338 ;
  assign n3428 = n66730 & n3423 ;
  assign n3429 = n3426 | n3428 ;
  assign n66731 = ~n3330 ;
  assign n3430 = n66731 & n3429 ;
  assign n66732 = ~n3320 ;
  assign n3431 = x72 & n66732 ;
  assign n66733 = ~n3315 ;
  assign n3432 = n66733 & n3431 ;
  assign n3433 = n3322 | n3432 ;
  assign n3435 = n3430 | n3433 ;
  assign n66734 = ~n3322 ;
  assign n3440 = n66734 & n3435 ;
  assign n3441 = n3438 | n3440 ;
  assign n66735 = ~n3314 ;
  assign n3442 = n66735 & n3441 ;
  assign n66736 = ~n3304 ;
  assign n3443 = x74 & n66736 ;
  assign n66737 = ~n3299 ;
  assign n3444 = n66737 & n3443 ;
  assign n3445 = n3306 | n3444 ;
  assign n3447 = n3442 | n3445 ;
  assign n66738 = ~n3306 ;
  assign n3452 = n66738 & n3447 ;
  assign n3453 = n3450 | n3452 ;
  assign n66739 = ~n3298 ;
  assign n3454 = n66739 & n3453 ;
  assign n66740 = ~n3288 ;
  assign n3455 = x76 & n66740 ;
  assign n66741 = ~n3283 ;
  assign n3456 = n66741 & n3455 ;
  assign n3457 = n3290 | n3456 ;
  assign n3459 = n3454 | n3457 ;
  assign n66742 = ~n3290 ;
  assign n3464 = n66742 & n3459 ;
  assign n3465 = n3462 | n3464 ;
  assign n66743 = ~n3282 ;
  assign n3466 = n66743 & n3465 ;
  assign n66744 = ~n3272 ;
  assign n3467 = x78 & n66744 ;
  assign n66745 = ~n3267 ;
  assign n3468 = n66745 & n3467 ;
  assign n3469 = n3274 | n3468 ;
  assign n3471 = n3466 | n3469 ;
  assign n66746 = ~n3274 ;
  assign n3476 = n66746 & n3471 ;
  assign n3477 = n3474 | n3476 ;
  assign n66747 = ~n3266 ;
  assign n3478 = n66747 & n3477 ;
  assign n66748 = ~n3256 ;
  assign n3479 = x80 & n66748 ;
  assign n66749 = ~n3251 ;
  assign n3480 = n66749 & n3479 ;
  assign n3481 = n3258 | n3480 ;
  assign n3483 = n3478 | n3481 ;
  assign n66750 = ~n3258 ;
  assign n3488 = n66750 & n3483 ;
  assign n3489 = n3486 | n3488 ;
  assign n66751 = ~n3250 ;
  assign n3490 = n66751 & n3489 ;
  assign n66752 = ~n3240 ;
  assign n3491 = x82 & n66752 ;
  assign n66753 = ~n3235 ;
  assign n3492 = n66753 & n3491 ;
  assign n3493 = n3242 | n3492 ;
  assign n3495 = n3490 | n3493 ;
  assign n66754 = ~n3242 ;
  assign n3501 = n66754 & n3495 ;
  assign n3502 = n3500 | n3501 ;
  assign n66755 = ~n3234 ;
  assign n3503 = n66755 & n3502 ;
  assign n3504 = n65666 | n3503 ;
  assign n66756 = ~n3233 ;
  assign n3506 = n66756 & n3504 ;
  assign n66757 = ~n3501 ;
  assign n3813 = n3500 & n66757 ;
  assign n3508 = x65 & n3396 ;
  assign n66758 = ~n3508 ;
  assign n3509 = n3392 & n66758 ;
  assign n3511 = n3393 | n3509 ;
  assign n3512 = n66719 & n3511 ;
  assign n3513 = n3401 | n3512 ;
  assign n3514 = n66722 & n3513 ;
  assign n3515 = n3405 | n3514 ;
  assign n3516 = n66723 & n3515 ;
  assign n3517 = n3411 | n3516 ;
  assign n3518 = n66726 & n3517 ;
  assign n3519 = n3415 | n3518 ;
  assign n3520 = n66727 & n3519 ;
  assign n3521 = n3421 | n3520 ;
  assign n3522 = n66730 & n3521 ;
  assign n3523 = n3426 | n3522 ;
  assign n3524 = n66731 & n3523 ;
  assign n3525 = n3433 | n3524 ;
  assign n3526 = n66734 & n3525 ;
  assign n3527 = n3438 | n3526 ;
  assign n3528 = n66735 & n3527 ;
  assign n3529 = n3445 | n3528 ;
  assign n3530 = n66738 & n3529 ;
  assign n3531 = n3450 | n3530 ;
  assign n3532 = n66739 & n3531 ;
  assign n3533 = n3457 | n3532 ;
  assign n3534 = n66742 & n3533 ;
  assign n3535 = n3462 | n3534 ;
  assign n3536 = n66743 & n3535 ;
  assign n3537 = n3469 | n3536 ;
  assign n3538 = n66746 & n3537 ;
  assign n3539 = n3474 | n3538 ;
  assign n3540 = n66747 & n3539 ;
  assign n3541 = n3481 | n3540 ;
  assign n3542 = n66750 & n3541 ;
  assign n3543 = n3486 | n3542 ;
  assign n3545 = n66751 & n3543 ;
  assign n3697 = n3493 | n3545 ;
  assign n3814 = n3242 | n3500 ;
  assign n66759 = ~n3814 ;
  assign n3815 = n3697 & n66759 ;
  assign n3816 = n3813 | n3815 ;
  assign n3817 = n3504 | n3816 ;
  assign n66760 = ~n3506 ;
  assign n3818 = n66760 & n3817 ;
  assign n3826 = n65674 & n3818 ;
  assign n3507 = n3241 & n3504 ;
  assign n3494 = n3250 | n3493 ;
  assign n66761 = ~n3494 ;
  assign n3544 = n66761 & n3543 ;
  assign n66762 = ~n3545 ;
  assign n3546 = n3493 & n66762 ;
  assign n3547 = n3544 | n3546 ;
  assign n3548 = n65674 & n3547 ;
  assign n66763 = ~n3503 ;
  assign n3549 = n66763 & n3548 ;
  assign n3550 = n3507 | n3549 ;
  assign n3551 = n66654 & n3550 ;
  assign n3552 = n3249 & n3504 ;
  assign n3487 = n3258 | n3486 ;
  assign n66764 = ~n3487 ;
  assign n3553 = n3483 & n66764 ;
  assign n66765 = ~n3488 ;
  assign n3554 = n3486 & n66765 ;
  assign n3555 = n3553 | n3554 ;
  assign n3556 = n65674 & n3555 ;
  assign n3557 = n66763 & n3556 ;
  assign n3558 = n3552 | n3557 ;
  assign n3559 = n66560 & n3558 ;
  assign n3560 = n3257 & n3504 ;
  assign n3482 = n3266 | n3481 ;
  assign n66766 = ~n3482 ;
  assign n3561 = n66766 & n3539 ;
  assign n66767 = ~n3540 ;
  assign n3562 = n3481 & n66767 ;
  assign n3563 = n3561 | n3562 ;
  assign n3564 = n65674 & n3563 ;
  assign n3565 = n66763 & n3564 ;
  assign n3566 = n3560 | n3565 ;
  assign n3567 = n66505 & n3566 ;
  assign n3568 = n3265 & n3504 ;
  assign n3475 = n3274 | n3474 ;
  assign n66768 = ~n3475 ;
  assign n3569 = n3471 & n66768 ;
  assign n66769 = ~n3476 ;
  assign n3570 = n3474 & n66769 ;
  assign n3571 = n3569 | n3570 ;
  assign n3572 = n65674 & n3571 ;
  assign n3573 = n66763 & n3572 ;
  assign n3574 = n3568 | n3573 ;
  assign n3575 = n66379 & n3574 ;
  assign n3576 = n3273 & n3504 ;
  assign n3470 = n3282 | n3469 ;
  assign n66770 = ~n3470 ;
  assign n3577 = n66770 & n3535 ;
  assign n66771 = ~n3536 ;
  assign n3578 = n3469 & n66771 ;
  assign n3579 = n3577 | n3578 ;
  assign n3580 = n65674 & n3579 ;
  assign n3581 = n66763 & n3580 ;
  assign n3582 = n3576 | n3581 ;
  assign n3583 = n66299 & n3582 ;
  assign n3584 = n3281 & n3504 ;
  assign n3463 = n3290 | n3462 ;
  assign n66772 = ~n3463 ;
  assign n3585 = n3459 & n66772 ;
  assign n66773 = ~n3464 ;
  assign n3586 = n3462 & n66773 ;
  assign n3587 = n3585 | n3586 ;
  assign n3588 = n65674 & n3587 ;
  assign n3589 = n66763 & n3588 ;
  assign n3590 = n3584 | n3589 ;
  assign n3591 = n66244 & n3590 ;
  assign n3592 = n3289 & n3504 ;
  assign n3458 = n3298 | n3457 ;
  assign n66774 = ~n3458 ;
  assign n3593 = n66774 & n3531 ;
  assign n66775 = ~n3532 ;
  assign n3594 = n3457 & n66775 ;
  assign n3595 = n3593 | n3594 ;
  assign n3596 = n65674 & n3595 ;
  assign n3597 = n66763 & n3596 ;
  assign n3598 = n3592 | n3597 ;
  assign n3599 = n66145 & n3598 ;
  assign n3600 = n3297 & n3504 ;
  assign n3451 = n3306 | n3450 ;
  assign n66776 = ~n3451 ;
  assign n3601 = n3447 & n66776 ;
  assign n66777 = ~n3452 ;
  assign n3602 = n3450 & n66777 ;
  assign n3603 = n3601 | n3602 ;
  assign n3604 = n65674 & n3603 ;
  assign n3605 = n66763 & n3604 ;
  assign n3606 = n3600 | n3605 ;
  assign n3607 = n66081 & n3606 ;
  assign n3608 = n3305 & n3504 ;
  assign n3446 = n3314 | n3445 ;
  assign n66778 = ~n3446 ;
  assign n3609 = n66778 & n3527 ;
  assign n66779 = ~n3528 ;
  assign n3610 = n3445 & n66779 ;
  assign n3611 = n3609 | n3610 ;
  assign n3612 = n65674 & n3611 ;
  assign n3613 = n66763 & n3612 ;
  assign n3614 = n3608 | n3613 ;
  assign n3615 = n66043 & n3614 ;
  assign n3616 = n3313 & n3504 ;
  assign n3439 = n3322 | n3438 ;
  assign n66780 = ~n3439 ;
  assign n3617 = n3435 & n66780 ;
  assign n66781 = ~n3440 ;
  assign n3618 = n3438 & n66781 ;
  assign n3619 = n3617 | n3618 ;
  assign n3620 = n65674 & n3619 ;
  assign n3621 = n66763 & n3620 ;
  assign n3622 = n3616 | n3621 ;
  assign n3623 = n65960 & n3622 ;
  assign n3624 = n3321 & n3504 ;
  assign n3434 = n3330 | n3433 ;
  assign n66782 = ~n3434 ;
  assign n3625 = n66782 & n3523 ;
  assign n66783 = ~n3524 ;
  assign n3626 = n3433 & n66783 ;
  assign n3627 = n3625 | n3626 ;
  assign n3628 = n65674 & n3627 ;
  assign n3629 = n66763 & n3628 ;
  assign n3630 = n3624 | n3629 ;
  assign n3631 = n65909 & n3630 ;
  assign n3632 = n3329 & n3504 ;
  assign n3427 = n3338 | n3426 ;
  assign n66784 = ~n3427 ;
  assign n3633 = n3423 & n66784 ;
  assign n66785 = ~n3428 ;
  assign n3634 = n3426 & n66785 ;
  assign n3635 = n3633 | n3634 ;
  assign n3636 = n65674 & n3635 ;
  assign n3637 = n66763 & n3636 ;
  assign n3638 = n3632 | n3637 ;
  assign n3639 = n65877 & n3638 ;
  assign n3640 = n3337 & n3504 ;
  assign n3422 = n3347 | n3421 ;
  assign n66786 = ~n3422 ;
  assign n3641 = n66786 & n3519 ;
  assign n66787 = ~n3520 ;
  assign n3642 = n3421 & n66787 ;
  assign n3643 = n3641 | n3642 ;
  assign n3644 = n65674 & n3643 ;
  assign n3645 = n66763 & n3644 ;
  assign n3646 = n3640 | n3645 ;
  assign n3647 = n65820 & n3646 ;
  assign n3648 = n3346 & n3504 ;
  assign n3649 = n3354 | n3415 ;
  assign n66788 = ~n3649 ;
  assign n3650 = n3412 & n66788 ;
  assign n66789 = ~n3416 ;
  assign n3651 = n3415 & n66789 ;
  assign n3652 = n3650 | n3651 ;
  assign n3653 = n65674 & n3652 ;
  assign n3654 = n66763 & n3653 ;
  assign n3655 = n3648 | n3654 ;
  assign n3656 = n65791 & n3655 ;
  assign n3657 = n3353 & n3504 ;
  assign n3658 = n3362 | n3411 ;
  assign n66790 = ~n3658 ;
  assign n3659 = n3407 & n66790 ;
  assign n66791 = ~n3516 ;
  assign n3660 = n3411 & n66791 ;
  assign n3661 = n3659 | n3660 ;
  assign n3662 = n65674 & n3661 ;
  assign n3663 = n66763 & n3662 ;
  assign n3664 = n3657 | n3663 ;
  assign n3665 = n65772 & n3664 ;
  assign n3666 = n3361 & n3504 ;
  assign n3667 = n3370 | n3405 ;
  assign n66792 = ~n3667 ;
  assign n3668 = n3402 & n66792 ;
  assign n66793 = ~n3406 ;
  assign n3669 = n3405 & n66793 ;
  assign n3670 = n3668 | n3669 ;
  assign n3671 = n65674 & n3670 ;
  assign n3672 = n66763 & n3671 ;
  assign n3673 = n3666 | n3672 ;
  assign n3674 = n65746 & n3673 ;
  assign n3675 = n3369 & n3504 ;
  assign n66794 = ~n3398 ;
  assign n3676 = n66794 & n3401 ;
  assign n3677 = n3397 | n3401 ;
  assign n66795 = ~n3677 ;
  assign n3678 = n3395 & n66795 ;
  assign n3679 = n3676 | n3678 ;
  assign n3680 = n65674 & n3679 ;
  assign n3681 = n66763 & n3680 ;
  assign n3682 = n3675 | n3681 ;
  assign n3683 = n65721 & n3682 ;
  assign n3505 = n3396 & n3504 ;
  assign n3510 = n3392 & n3393 ;
  assign n3684 = n66718 & n3510 ;
  assign n3685 = n65666 | n3684 ;
  assign n66796 = ~n3685 ;
  assign n3686 = n3395 & n66796 ;
  assign n3687 = n66763 & n3686 ;
  assign n3688 = n3505 | n3687 ;
  assign n3689 = n65686 & n3688 ;
  assign n66797 = ~x84 ;
  assign n3690 = x64 & n66797 ;
  assign n3691 = n66712 & n3690 ;
  assign n3692 = n66713 & n3691 ;
  assign n3693 = n66714 & n3692 ;
  assign n3694 = n66715 & n3693 ;
  assign n3698 = n66754 & n3697 ;
  assign n3699 = n3500 | n3698 ;
  assign n3700 = n66755 & n3699 ;
  assign n66798 = ~n3700 ;
  assign n3701 = n3694 & n66798 ;
  assign n66799 = ~n3701 ;
  assign n3702 = x44 & n66799 ;
  assign n3703 = n66507 & n3393 ;
  assign n3704 = n66508 & n3703 ;
  assign n3705 = n66509 & n3704 ;
  assign n3706 = n66510 & n3705 ;
  assign n3707 = n66763 & n3706 ;
  assign n3708 = n3702 | n3707 ;
  assign n3710 = x65 & n3708 ;
  assign n3695 = n66763 & n3694 ;
  assign n66800 = ~n3695 ;
  assign n3696 = x44 & n66800 ;
  assign n3709 = x65 | n3707 ;
  assign n3711 = n3696 | n3709 ;
  assign n66801 = ~n3710 ;
  assign n3712 = n66801 & n3711 ;
  assign n66802 = ~x43 ;
  assign n3713 = n66802 & x64 ;
  assign n3714 = n3712 | n3713 ;
  assign n3715 = n65670 & n3708 ;
  assign n66803 = ~n3715 ;
  assign n3716 = n3714 & n66803 ;
  assign n66804 = ~n3687 ;
  assign n3717 = x66 & n66804 ;
  assign n66805 = ~n3505 ;
  assign n3718 = n66805 & n3717 ;
  assign n3719 = n3689 | n3718 ;
  assign n3720 = n3716 | n3719 ;
  assign n66806 = ~n3689 ;
  assign n3721 = n66806 & n3720 ;
  assign n66807 = ~n3681 ;
  assign n3722 = x67 & n66807 ;
  assign n66808 = ~n3675 ;
  assign n3723 = n66808 & n3722 ;
  assign n3724 = n3721 | n3723 ;
  assign n66809 = ~n3683 ;
  assign n3725 = n66809 & n3724 ;
  assign n66810 = ~n3672 ;
  assign n3726 = x68 & n66810 ;
  assign n66811 = ~n3666 ;
  assign n3727 = n66811 & n3726 ;
  assign n3728 = n3674 | n3727 ;
  assign n3729 = n3725 | n3728 ;
  assign n66812 = ~n3674 ;
  assign n3730 = n66812 & n3729 ;
  assign n66813 = ~n3663 ;
  assign n3731 = x69 & n66813 ;
  assign n66814 = ~n3657 ;
  assign n3732 = n66814 & n3731 ;
  assign n3733 = n3665 | n3732 ;
  assign n3734 = n3730 | n3733 ;
  assign n66815 = ~n3665 ;
  assign n3735 = n66815 & n3734 ;
  assign n66816 = ~n3654 ;
  assign n3736 = x70 & n66816 ;
  assign n66817 = ~n3648 ;
  assign n3737 = n66817 & n3736 ;
  assign n3738 = n3656 | n3737 ;
  assign n3739 = n3735 | n3738 ;
  assign n66818 = ~n3656 ;
  assign n3740 = n66818 & n3739 ;
  assign n66819 = ~n3645 ;
  assign n3741 = x71 & n66819 ;
  assign n66820 = ~n3640 ;
  assign n3742 = n66820 & n3741 ;
  assign n3743 = n3647 | n3742 ;
  assign n3745 = n3740 | n3743 ;
  assign n66821 = ~n3647 ;
  assign n3746 = n66821 & n3745 ;
  assign n66822 = ~n3637 ;
  assign n3747 = x72 & n66822 ;
  assign n66823 = ~n3632 ;
  assign n3748 = n66823 & n3747 ;
  assign n3749 = n3639 | n3748 ;
  assign n3750 = n3746 | n3749 ;
  assign n66824 = ~n3639 ;
  assign n3751 = n66824 & n3750 ;
  assign n66825 = ~n3629 ;
  assign n3752 = x73 & n66825 ;
  assign n66826 = ~n3624 ;
  assign n3753 = n66826 & n3752 ;
  assign n3754 = n3631 | n3753 ;
  assign n3756 = n3751 | n3754 ;
  assign n66827 = ~n3631 ;
  assign n3757 = n66827 & n3756 ;
  assign n66828 = ~n3621 ;
  assign n3758 = x74 & n66828 ;
  assign n66829 = ~n3616 ;
  assign n3759 = n66829 & n3758 ;
  assign n3760 = n3623 | n3759 ;
  assign n3761 = n3757 | n3760 ;
  assign n66830 = ~n3623 ;
  assign n3762 = n66830 & n3761 ;
  assign n66831 = ~n3613 ;
  assign n3763 = x75 & n66831 ;
  assign n66832 = ~n3608 ;
  assign n3764 = n66832 & n3763 ;
  assign n3765 = n3615 | n3764 ;
  assign n3767 = n3762 | n3765 ;
  assign n66833 = ~n3615 ;
  assign n3768 = n66833 & n3767 ;
  assign n66834 = ~n3605 ;
  assign n3769 = x76 & n66834 ;
  assign n66835 = ~n3600 ;
  assign n3770 = n66835 & n3769 ;
  assign n3771 = n3607 | n3770 ;
  assign n3772 = n3768 | n3771 ;
  assign n66836 = ~n3607 ;
  assign n3773 = n66836 & n3772 ;
  assign n66837 = ~n3597 ;
  assign n3774 = x77 & n66837 ;
  assign n66838 = ~n3592 ;
  assign n3775 = n66838 & n3774 ;
  assign n3776 = n3599 | n3775 ;
  assign n3778 = n3773 | n3776 ;
  assign n66839 = ~n3599 ;
  assign n3779 = n66839 & n3778 ;
  assign n66840 = ~n3589 ;
  assign n3780 = x78 & n66840 ;
  assign n66841 = ~n3584 ;
  assign n3781 = n66841 & n3780 ;
  assign n3782 = n3591 | n3781 ;
  assign n3783 = n3779 | n3782 ;
  assign n66842 = ~n3591 ;
  assign n3784 = n66842 & n3783 ;
  assign n66843 = ~n3581 ;
  assign n3785 = x79 & n66843 ;
  assign n66844 = ~n3576 ;
  assign n3786 = n66844 & n3785 ;
  assign n3787 = n3583 | n3786 ;
  assign n3789 = n3784 | n3787 ;
  assign n66845 = ~n3583 ;
  assign n3790 = n66845 & n3789 ;
  assign n66846 = ~n3573 ;
  assign n3791 = x80 & n66846 ;
  assign n66847 = ~n3568 ;
  assign n3792 = n66847 & n3791 ;
  assign n3793 = n3575 | n3792 ;
  assign n3794 = n3790 | n3793 ;
  assign n66848 = ~n3575 ;
  assign n3795 = n66848 & n3794 ;
  assign n66849 = ~n3565 ;
  assign n3796 = x81 & n66849 ;
  assign n66850 = ~n3560 ;
  assign n3797 = n66850 & n3796 ;
  assign n3798 = n3567 | n3797 ;
  assign n3800 = n3795 | n3798 ;
  assign n66851 = ~n3567 ;
  assign n3801 = n66851 & n3800 ;
  assign n66852 = ~n3557 ;
  assign n3802 = x82 & n66852 ;
  assign n66853 = ~n3552 ;
  assign n3803 = n66853 & n3802 ;
  assign n3804 = n3559 | n3803 ;
  assign n3805 = n3801 | n3804 ;
  assign n66854 = ~n3559 ;
  assign n3806 = n66854 & n3805 ;
  assign n66855 = ~n3549 ;
  assign n3807 = x83 & n66855 ;
  assign n66856 = ~n3507 ;
  assign n3808 = n66856 & n3807 ;
  assign n3809 = n3551 | n3808 ;
  assign n3811 = n3806 | n3809 ;
  assign n66857 = ~n3551 ;
  assign n3812 = n66857 & n3811 ;
  assign n3819 = n66797 & n3818 ;
  assign n173 = ~n3504 ;
  assign n3820 = n173 & n3816 ;
  assign n3821 = n3233 & n3504 ;
  assign n66859 = ~n3821 ;
  assign n3822 = x84 & n66859 ;
  assign n66860 = ~n3820 ;
  assign n3823 = n66860 & n3822 ;
  assign n3824 = n513 | n3823 ;
  assign n3825 = n3819 | n3824 ;
  assign n3827 = n3812 | n3825 ;
  assign n66861 = ~n3826 ;
  assign n3828 = n66861 & n3827 ;
  assign n66862 = ~n3806 ;
  assign n3810 = n66862 & n3809 ;
  assign n3831 = n3696 | n3707 ;
  assign n3832 = x65 & n3831 ;
  assign n66863 = ~n3832 ;
  assign n3833 = n3711 & n66863 ;
  assign n3834 = n3713 | n3833 ;
  assign n3835 = n66803 & n3834 ;
  assign n3837 = n3718 | n3835 ;
  assign n3838 = n66806 & n3837 ;
  assign n3839 = n3683 | n3723 ;
  assign n3841 = n3838 | n3839 ;
  assign n3842 = n66809 & n3841 ;
  assign n3844 = n3728 | n3842 ;
  assign n3845 = n66812 & n3844 ;
  assign n3847 = n3733 | n3845 ;
  assign n3848 = n66815 & n3847 ;
  assign n3849 = n3738 | n3848 ;
  assign n3851 = n66818 & n3849 ;
  assign n3852 = n3743 | n3851 ;
  assign n3853 = n66821 & n3852 ;
  assign n3854 = n3749 | n3853 ;
  assign n3856 = n66824 & n3854 ;
  assign n3857 = n3754 | n3856 ;
  assign n3858 = n66827 & n3857 ;
  assign n3859 = n3760 | n3858 ;
  assign n3861 = n66830 & n3859 ;
  assign n3862 = n3765 | n3861 ;
  assign n3863 = n66833 & n3862 ;
  assign n3864 = n3771 | n3863 ;
  assign n3866 = n66836 & n3864 ;
  assign n3867 = n3776 | n3866 ;
  assign n3868 = n66839 & n3867 ;
  assign n3869 = n3782 | n3868 ;
  assign n3871 = n66842 & n3869 ;
  assign n3872 = n3787 | n3871 ;
  assign n3873 = n66845 & n3872 ;
  assign n3874 = n3793 | n3873 ;
  assign n3876 = n66848 & n3874 ;
  assign n3877 = n3798 | n3876 ;
  assign n3878 = n66851 & n3877 ;
  assign n3879 = n3804 | n3878 ;
  assign n3896 = n3559 | n3809 ;
  assign n66864 = ~n3896 ;
  assign n3897 = n3879 & n66864 ;
  assign n3898 = n3810 | n3897 ;
  assign n172 = ~n3828 ;
  assign n3899 = n172 & n3898 ;
  assign n3881 = n66854 & n3879 ;
  assign n3882 = n3809 | n3881 ;
  assign n3883 = n66857 & n3882 ;
  assign n3884 = n3825 | n3883 ;
  assign n3900 = n3550 & n66861 ;
  assign n3901 = n3884 & n3900 ;
  assign n3902 = n3899 | n3901 ;
  assign n3885 = n3551 | n3823 ;
  assign n3886 = n3819 | n3885 ;
  assign n66866 = ~n3886 ;
  assign n3887 = n3811 & n66866 ;
  assign n3888 = n3819 | n3823 ;
  assign n66867 = ~n3883 ;
  assign n3889 = n66867 & n3888 ;
  assign n3890 = n3887 | n3889 ;
  assign n3891 = n172 & n3890 ;
  assign n3892 = n65666 & n3233 ;
  assign n3893 = n3884 & n3892 ;
  assign n3894 = n3891 | n3893 ;
  assign n66868 = ~x85 ;
  assign n3895 = n66868 & n3894 ;
  assign n66869 = ~n3893 ;
  assign n4173 = x85 & n66869 ;
  assign n66870 = ~n3891 ;
  assign n4174 = n66870 & n4173 ;
  assign n4175 = n3895 | n4174 ;
  assign n3903 = n66797 & n3902 ;
  assign n66871 = ~n3878 ;
  assign n3880 = n3804 & n66871 ;
  assign n3904 = n3567 | n3804 ;
  assign n66872 = ~n3904 ;
  assign n3905 = n3800 & n66872 ;
  assign n3906 = n3880 | n3905 ;
  assign n3907 = n172 & n3906 ;
  assign n3908 = n3558 & n66861 ;
  assign n3909 = n3884 & n3908 ;
  assign n3910 = n3907 | n3909 ;
  assign n3911 = n66654 & n3910 ;
  assign n66873 = ~n3909 ;
  assign n4161 = x83 & n66873 ;
  assign n66874 = ~n3907 ;
  assign n4162 = n66874 & n4161 ;
  assign n4163 = n3911 | n4162 ;
  assign n66875 = ~n3795 ;
  assign n3799 = n66875 & n3798 ;
  assign n3912 = n3575 | n3798 ;
  assign n66876 = ~n3912 ;
  assign n3913 = n3874 & n66876 ;
  assign n3914 = n3799 | n3913 ;
  assign n3915 = n172 & n3914 ;
  assign n3916 = n3566 & n66861 ;
  assign n3917 = n3884 & n3916 ;
  assign n3918 = n3915 | n3917 ;
  assign n3919 = n66560 & n3918 ;
  assign n66877 = ~n3873 ;
  assign n3875 = n3793 & n66877 ;
  assign n3920 = n3583 | n3793 ;
  assign n66878 = ~n3920 ;
  assign n3921 = n3789 & n66878 ;
  assign n3922 = n3875 | n3921 ;
  assign n3923 = n172 & n3922 ;
  assign n3924 = n3574 & n66861 ;
  assign n3925 = n3884 & n3924 ;
  assign n3926 = n3923 | n3925 ;
  assign n3927 = n66505 & n3926 ;
  assign n66879 = ~n3925 ;
  assign n4149 = x81 & n66879 ;
  assign n66880 = ~n3923 ;
  assign n4150 = n66880 & n4149 ;
  assign n4151 = n3927 | n4150 ;
  assign n66881 = ~n3784 ;
  assign n3788 = n66881 & n3787 ;
  assign n3928 = n3591 | n3787 ;
  assign n66882 = ~n3928 ;
  assign n3929 = n3869 & n66882 ;
  assign n3930 = n3788 | n3929 ;
  assign n3931 = n172 & n3930 ;
  assign n3932 = n3582 & n66861 ;
  assign n3933 = n3884 & n3932 ;
  assign n3934 = n3931 | n3933 ;
  assign n3935 = n66379 & n3934 ;
  assign n66883 = ~n3868 ;
  assign n3870 = n3782 & n66883 ;
  assign n3936 = n3599 | n3782 ;
  assign n66884 = ~n3936 ;
  assign n3937 = n3778 & n66884 ;
  assign n3938 = n3870 | n3937 ;
  assign n3939 = n172 & n3938 ;
  assign n3940 = n3590 & n66861 ;
  assign n3941 = n3884 & n3940 ;
  assign n3942 = n3939 | n3941 ;
  assign n3943 = n66299 & n3942 ;
  assign n66885 = ~n3941 ;
  assign n4137 = x79 & n66885 ;
  assign n66886 = ~n3939 ;
  assign n4138 = n66886 & n4137 ;
  assign n4139 = n3943 | n4138 ;
  assign n66887 = ~n3773 ;
  assign n3777 = n66887 & n3776 ;
  assign n3944 = n3607 | n3776 ;
  assign n66888 = ~n3944 ;
  assign n3945 = n3864 & n66888 ;
  assign n3946 = n3777 | n3945 ;
  assign n3947 = n172 & n3946 ;
  assign n3948 = n3598 & n66861 ;
  assign n3949 = n3884 & n3948 ;
  assign n3950 = n3947 | n3949 ;
  assign n3951 = n66244 & n3950 ;
  assign n66889 = ~n3863 ;
  assign n3865 = n3771 & n66889 ;
  assign n3952 = n3615 | n3771 ;
  assign n66890 = ~n3952 ;
  assign n3953 = n3767 & n66890 ;
  assign n3954 = n3865 | n3953 ;
  assign n3955 = n172 & n3954 ;
  assign n3956 = n3606 & n66861 ;
  assign n3957 = n3884 & n3956 ;
  assign n3958 = n3955 | n3957 ;
  assign n3959 = n66145 & n3958 ;
  assign n66891 = ~n3957 ;
  assign n4125 = x77 & n66891 ;
  assign n66892 = ~n3955 ;
  assign n4126 = n66892 & n4125 ;
  assign n4127 = n3959 | n4126 ;
  assign n66893 = ~n3762 ;
  assign n3766 = n66893 & n3765 ;
  assign n3960 = n3623 | n3765 ;
  assign n66894 = ~n3960 ;
  assign n3961 = n3859 & n66894 ;
  assign n3962 = n3766 | n3961 ;
  assign n3963 = n172 & n3962 ;
  assign n3964 = n3614 & n66861 ;
  assign n3965 = n3884 & n3964 ;
  assign n3966 = n3963 | n3965 ;
  assign n3967 = n66081 & n3966 ;
  assign n66895 = ~n3858 ;
  assign n3860 = n3760 & n66895 ;
  assign n3968 = n3631 | n3760 ;
  assign n66896 = ~n3968 ;
  assign n3969 = n3756 & n66896 ;
  assign n3970 = n3860 | n3969 ;
  assign n3971 = n172 & n3970 ;
  assign n3972 = n3622 & n66861 ;
  assign n3973 = n3884 & n3972 ;
  assign n3974 = n3971 | n3973 ;
  assign n3975 = n66043 & n3974 ;
  assign n66897 = ~n3973 ;
  assign n4113 = x75 & n66897 ;
  assign n66898 = ~n3971 ;
  assign n4114 = n66898 & n4113 ;
  assign n4115 = n3975 | n4114 ;
  assign n66899 = ~n3751 ;
  assign n3755 = n66899 & n3754 ;
  assign n3976 = n3639 | n3754 ;
  assign n66900 = ~n3976 ;
  assign n3977 = n3854 & n66900 ;
  assign n3978 = n3755 | n3977 ;
  assign n3979 = n172 & n3978 ;
  assign n3980 = n3630 & n66861 ;
  assign n3981 = n3884 & n3980 ;
  assign n3982 = n3979 | n3981 ;
  assign n3983 = n65960 & n3982 ;
  assign n66901 = ~n3853 ;
  assign n3855 = n3749 & n66901 ;
  assign n3984 = n3647 | n3749 ;
  assign n66902 = ~n3984 ;
  assign n3985 = n3745 & n66902 ;
  assign n3986 = n3855 | n3985 ;
  assign n3987 = n172 & n3986 ;
  assign n3988 = n3638 & n66861 ;
  assign n3989 = n3884 & n3988 ;
  assign n3990 = n3987 | n3989 ;
  assign n3991 = n65909 & n3990 ;
  assign n66903 = ~n3989 ;
  assign n4101 = x73 & n66903 ;
  assign n66904 = ~n3987 ;
  assign n4102 = n66904 & n4101 ;
  assign n4103 = n3991 | n4102 ;
  assign n66905 = ~n3740 ;
  assign n3744 = n66905 & n3743 ;
  assign n3992 = n3656 | n3743 ;
  assign n66906 = ~n3992 ;
  assign n3993 = n3849 & n66906 ;
  assign n3994 = n3744 | n3993 ;
  assign n3995 = n172 & n3994 ;
  assign n3996 = n3646 & n66861 ;
  assign n3997 = n3884 & n3996 ;
  assign n3998 = n3995 | n3997 ;
  assign n3999 = n65877 & n3998 ;
  assign n66907 = ~n3848 ;
  assign n3850 = n3738 & n66907 ;
  assign n4000 = n3665 | n3738 ;
  assign n66908 = ~n4000 ;
  assign n4001 = n3734 & n66908 ;
  assign n4002 = n3850 | n4001 ;
  assign n4003 = n172 & n4002 ;
  assign n4004 = n3655 & n66861 ;
  assign n4005 = n3884 & n4004 ;
  assign n4006 = n4003 | n4005 ;
  assign n4007 = n65820 & n4006 ;
  assign n66909 = ~n4005 ;
  assign n4089 = x71 & n66909 ;
  assign n66910 = ~n4003 ;
  assign n4090 = n66910 & n4089 ;
  assign n4091 = n4007 | n4090 ;
  assign n66911 = ~n3730 ;
  assign n3846 = n66911 & n3733 ;
  assign n4008 = n3674 | n3733 ;
  assign n66912 = ~n4008 ;
  assign n4009 = n3844 & n66912 ;
  assign n4010 = n3846 | n4009 ;
  assign n4011 = n172 & n4010 ;
  assign n4012 = n3664 & n66861 ;
  assign n4013 = n3884 & n4012 ;
  assign n4014 = n4011 | n4013 ;
  assign n4015 = n65791 & n4014 ;
  assign n66913 = ~n3842 ;
  assign n3843 = n3728 & n66913 ;
  assign n4016 = n3721 | n3839 ;
  assign n4017 = n3683 | n3728 ;
  assign n66914 = ~n4017 ;
  assign n4018 = n4016 & n66914 ;
  assign n4019 = n3843 | n4018 ;
  assign n4020 = n172 & n4019 ;
  assign n4021 = n3673 & n66861 ;
  assign n4022 = n3884 & n4021 ;
  assign n4023 = n4020 | n4022 ;
  assign n4024 = n65772 & n4023 ;
  assign n66915 = ~n4022 ;
  assign n4078 = x69 & n66915 ;
  assign n66916 = ~n4020 ;
  assign n4079 = n66916 & n4078 ;
  assign n4080 = n4024 | n4079 ;
  assign n66917 = ~n3721 ;
  assign n3840 = n66917 & n3839 ;
  assign n4025 = n3689 | n3839 ;
  assign n66918 = ~n4025 ;
  assign n4026 = n3720 & n66918 ;
  assign n4027 = n3840 | n4026 ;
  assign n4028 = n172 & n4027 ;
  assign n4029 = n3682 & n66861 ;
  assign n4030 = n3884 & n4029 ;
  assign n4031 = n4028 | n4030 ;
  assign n4032 = n65746 & n4031 ;
  assign n66919 = ~n3835 ;
  assign n3836 = n3719 & n66919 ;
  assign n4033 = n3715 | n3719 ;
  assign n66920 = ~n4033 ;
  assign n4034 = n3714 & n66920 ;
  assign n4035 = n3836 | n4034 ;
  assign n4036 = n172 & n4035 ;
  assign n4037 = n3688 & n66861 ;
  assign n4038 = n3884 & n4037 ;
  assign n4039 = n4036 | n4038 ;
  assign n4040 = n65721 & n4039 ;
  assign n66921 = ~n4038 ;
  assign n4068 = x67 & n66921 ;
  assign n66922 = ~n4036 ;
  assign n4069 = n66922 & n4068 ;
  assign n4070 = n4040 | n4069 ;
  assign n4041 = n3711 & n3713 ;
  assign n4042 = n66801 & n4041 ;
  assign n66923 = ~n4042 ;
  assign n4043 = n3834 & n66923 ;
  assign n4044 = n172 & n4043 ;
  assign n4045 = n3708 & n66861 ;
  assign n4046 = n3884 & n4045 ;
  assign n4047 = n4044 | n4046 ;
  assign n4048 = n65686 & n4047 ;
  assign n66924 = ~x42 ;
  assign n4058 = n66924 & x64 ;
  assign n3829 = n3713 & n172 ;
  assign n4049 = n66861 & n3884 ;
  assign n66925 = ~n4049 ;
  assign n4050 = x64 & n66925 ;
  assign n66926 = ~n4050 ;
  assign n4051 = x43 & n66926 ;
  assign n4052 = n3829 | n4051 ;
  assign n4053 = x65 & n4052 ;
  assign n3830 = x64 & n172 ;
  assign n66927 = ~n3830 ;
  assign n4054 = x43 & n66927 ;
  assign n4055 = n3713 & n66925 ;
  assign n4056 = x65 | n4055 ;
  assign n4057 = n4054 | n4056 ;
  assign n66928 = ~n4053 ;
  assign n4059 = n66928 & n4057 ;
  assign n4060 = n4058 | n4059 ;
  assign n4061 = n3829 | n4054 ;
  assign n4062 = n65670 & n4061 ;
  assign n66929 = ~n4062 ;
  assign n4063 = n4060 & n66929 ;
  assign n66930 = ~n4046 ;
  assign n4064 = x66 & n66930 ;
  assign n66931 = ~n4044 ;
  assign n4065 = n66931 & n4064 ;
  assign n4066 = n4048 | n4065 ;
  assign n4067 = n4063 | n4066 ;
  assign n66932 = ~n4048 ;
  assign n4071 = n66932 & n4067 ;
  assign n4072 = n4070 | n4071 ;
  assign n66933 = ~n4040 ;
  assign n4073 = n66933 & n4072 ;
  assign n66934 = ~n4030 ;
  assign n4074 = x68 & n66934 ;
  assign n66935 = ~n4028 ;
  assign n4075 = n66935 & n4074 ;
  assign n4076 = n4032 | n4075 ;
  assign n4077 = n4073 | n4076 ;
  assign n66936 = ~n4032 ;
  assign n4081 = n66936 & n4077 ;
  assign n4082 = n4080 | n4081 ;
  assign n66937 = ~n4024 ;
  assign n4083 = n66937 & n4082 ;
  assign n66938 = ~n4013 ;
  assign n4084 = x70 & n66938 ;
  assign n66939 = ~n4011 ;
  assign n4085 = n66939 & n4084 ;
  assign n4086 = n4015 | n4085 ;
  assign n4088 = n4083 | n4086 ;
  assign n66940 = ~n4015 ;
  assign n4093 = n66940 & n4088 ;
  assign n4094 = n4091 | n4093 ;
  assign n66941 = ~n4007 ;
  assign n4095 = n66941 & n4094 ;
  assign n66942 = ~n3997 ;
  assign n4096 = x72 & n66942 ;
  assign n66943 = ~n3995 ;
  assign n4097 = n66943 & n4096 ;
  assign n4098 = n3999 | n4097 ;
  assign n4100 = n4095 | n4098 ;
  assign n66944 = ~n3999 ;
  assign n4105 = n66944 & n4100 ;
  assign n4106 = n4103 | n4105 ;
  assign n66945 = ~n3991 ;
  assign n4107 = n66945 & n4106 ;
  assign n66946 = ~n3981 ;
  assign n4108 = x74 & n66946 ;
  assign n66947 = ~n3979 ;
  assign n4109 = n66947 & n4108 ;
  assign n4110 = n3983 | n4109 ;
  assign n4112 = n4107 | n4110 ;
  assign n66948 = ~n3983 ;
  assign n4117 = n66948 & n4112 ;
  assign n4118 = n4115 | n4117 ;
  assign n66949 = ~n3975 ;
  assign n4119 = n66949 & n4118 ;
  assign n66950 = ~n3965 ;
  assign n4120 = x76 & n66950 ;
  assign n66951 = ~n3963 ;
  assign n4121 = n66951 & n4120 ;
  assign n4122 = n3967 | n4121 ;
  assign n4124 = n4119 | n4122 ;
  assign n66952 = ~n3967 ;
  assign n4129 = n66952 & n4124 ;
  assign n4130 = n4127 | n4129 ;
  assign n66953 = ~n3959 ;
  assign n4131 = n66953 & n4130 ;
  assign n66954 = ~n3949 ;
  assign n4132 = x78 & n66954 ;
  assign n66955 = ~n3947 ;
  assign n4133 = n66955 & n4132 ;
  assign n4134 = n3951 | n4133 ;
  assign n4136 = n4131 | n4134 ;
  assign n66956 = ~n3951 ;
  assign n4141 = n66956 & n4136 ;
  assign n4142 = n4139 | n4141 ;
  assign n66957 = ~n3943 ;
  assign n4143 = n66957 & n4142 ;
  assign n66958 = ~n3933 ;
  assign n4144 = x80 & n66958 ;
  assign n66959 = ~n3931 ;
  assign n4145 = n66959 & n4144 ;
  assign n4146 = n3935 | n4145 ;
  assign n4148 = n4143 | n4146 ;
  assign n66960 = ~n3935 ;
  assign n4153 = n66960 & n4148 ;
  assign n4154 = n4151 | n4153 ;
  assign n66961 = ~n3927 ;
  assign n4155 = n66961 & n4154 ;
  assign n66962 = ~n3917 ;
  assign n4156 = x82 & n66962 ;
  assign n66963 = ~n3915 ;
  assign n4157 = n66963 & n4156 ;
  assign n4158 = n3919 | n4157 ;
  assign n4160 = n4155 | n4158 ;
  assign n66964 = ~n3919 ;
  assign n4165 = n66964 & n4160 ;
  assign n4166 = n4163 | n4165 ;
  assign n66965 = ~n3911 ;
  assign n4167 = n66965 & n4166 ;
  assign n66966 = ~n3901 ;
  assign n4168 = x84 & n66966 ;
  assign n66967 = ~n3899 ;
  assign n4169 = n66967 & n4168 ;
  assign n4170 = n3903 | n4169 ;
  assign n4172 = n4167 | n4170 ;
  assign n66968 = ~n3903 ;
  assign n4176 = n66968 & n4172 ;
  assign n4177 = n4175 | n4176 ;
  assign n66969 = ~n3895 ;
  assign n4178 = n66969 & n4177 ;
  assign n4179 = n65564 | n65579 ;
  assign n4180 = n65647 | n4179 ;
  assign n4181 = n65542 | n4180 ;
  assign n4182 = n65429 | n4181 ;
  assign n4183 = n4178 | n4182 ;
  assign n4238 = n3902 & n4183 ;
  assign n4171 = n3911 | n4170 ;
  assign n4187 = x65 & n4061 ;
  assign n66970 = ~n4187 ;
  assign n4188 = n4057 & n66970 ;
  assign n4190 = n4058 | n4188 ;
  assign n4192 = n66929 & n4190 ;
  assign n4193 = n4066 | n4192 ;
  assign n4194 = n66932 & n4193 ;
  assign n4195 = n4070 | n4194 ;
  assign n4196 = n66933 & n4195 ;
  assign n4197 = n4076 | n4196 ;
  assign n4198 = n66936 & n4197 ;
  assign n4199 = n4080 | n4198 ;
  assign n4200 = n66937 & n4199 ;
  assign n4201 = n4086 | n4200 ;
  assign n4202 = n66940 & n4201 ;
  assign n4203 = n4091 | n4202 ;
  assign n4204 = n66941 & n4203 ;
  assign n4205 = n4098 | n4204 ;
  assign n4206 = n66944 & n4205 ;
  assign n4207 = n4103 | n4206 ;
  assign n4208 = n66945 & n4207 ;
  assign n4209 = n4110 | n4208 ;
  assign n4210 = n66948 & n4209 ;
  assign n4211 = n4115 | n4210 ;
  assign n4212 = n66949 & n4211 ;
  assign n4213 = n4122 | n4212 ;
  assign n4214 = n66952 & n4213 ;
  assign n4215 = n4127 | n4214 ;
  assign n4216 = n66953 & n4215 ;
  assign n4217 = n4134 | n4216 ;
  assign n4218 = n66956 & n4217 ;
  assign n4219 = n4139 | n4218 ;
  assign n4220 = n66957 & n4219 ;
  assign n4221 = n4146 | n4220 ;
  assign n4222 = n66960 & n4221 ;
  assign n4223 = n4151 | n4222 ;
  assign n4224 = n66961 & n4223 ;
  assign n4225 = n4158 | n4224 ;
  assign n4226 = n66964 & n4225 ;
  assign n4227 = n4163 | n4226 ;
  assign n66971 = ~n4171 ;
  assign n4239 = n66971 & n4227 ;
  assign n4228 = n66965 & n4227 ;
  assign n66972 = ~n4228 ;
  assign n4240 = n4170 & n66972 ;
  assign n4241 = n4239 | n4240 ;
  assign n66973 = ~n4182 ;
  assign n4242 = n66973 & n4241 ;
  assign n66974 = ~n4178 ;
  assign n4243 = n66974 & n4242 ;
  assign n4244 = n4238 | n4243 ;
  assign n66975 = ~n3894 ;
  assign n4184 = n66975 & n4183 ;
  assign n66976 = ~n4176 ;
  assign n4231 = n4175 & n66976 ;
  assign n4229 = n4170 | n4228 ;
  assign n4232 = n3903 | n4175 ;
  assign n66977 = ~n4232 ;
  assign n4233 = n4229 & n66977 ;
  assign n4234 = n4231 | n4233 ;
  assign n4235 = n4183 | n4234 ;
  assign n66978 = ~n4184 ;
  assign n4236 = n66978 & n4235 ;
  assign n66979 = ~x86 ;
  assign n4237 = n66979 & n4236 ;
  assign n4245 = n66868 & n4244 ;
  assign n4246 = n3910 & n4183 ;
  assign n4164 = n3919 | n4163 ;
  assign n66980 = ~n4164 ;
  assign n4247 = n4160 & n66980 ;
  assign n66981 = ~n4165 ;
  assign n4248 = n4163 & n66981 ;
  assign n4249 = n4247 | n4248 ;
  assign n4250 = n66973 & n4249 ;
  assign n4251 = n66974 & n4250 ;
  assign n4252 = n4246 | n4251 ;
  assign n4253 = n66797 & n4252 ;
  assign n4254 = n3918 & n4183 ;
  assign n4159 = n3927 | n4158 ;
  assign n66982 = ~n4159 ;
  assign n4255 = n66982 & n4223 ;
  assign n66983 = ~n4224 ;
  assign n4256 = n4158 & n66983 ;
  assign n4257 = n4255 | n4256 ;
  assign n4258 = n66973 & n4257 ;
  assign n4259 = n66974 & n4258 ;
  assign n4260 = n4254 | n4259 ;
  assign n4261 = n66654 & n4260 ;
  assign n4262 = n3926 & n4183 ;
  assign n4152 = n3935 | n4151 ;
  assign n66984 = ~n4152 ;
  assign n4263 = n4148 & n66984 ;
  assign n66985 = ~n4153 ;
  assign n4264 = n4151 & n66985 ;
  assign n4265 = n4263 | n4264 ;
  assign n4266 = n66973 & n4265 ;
  assign n4267 = n66974 & n4266 ;
  assign n4268 = n4262 | n4267 ;
  assign n4269 = n66560 & n4268 ;
  assign n4270 = n3934 & n4183 ;
  assign n4147 = n3943 | n4146 ;
  assign n66986 = ~n4147 ;
  assign n4271 = n66986 & n4219 ;
  assign n66987 = ~n4220 ;
  assign n4272 = n4146 & n66987 ;
  assign n4273 = n4271 | n4272 ;
  assign n4274 = n66973 & n4273 ;
  assign n4275 = n66974 & n4274 ;
  assign n4276 = n4270 | n4275 ;
  assign n4277 = n66505 & n4276 ;
  assign n4278 = n3942 & n4183 ;
  assign n4140 = n3951 | n4139 ;
  assign n66988 = ~n4140 ;
  assign n4279 = n4136 & n66988 ;
  assign n66989 = ~n4141 ;
  assign n4280 = n4139 & n66989 ;
  assign n4281 = n4279 | n4280 ;
  assign n4282 = n66973 & n4281 ;
  assign n4283 = n66974 & n4282 ;
  assign n4284 = n4278 | n4283 ;
  assign n4285 = n66379 & n4284 ;
  assign n4286 = n3950 & n4183 ;
  assign n4135 = n3959 | n4134 ;
  assign n66990 = ~n4135 ;
  assign n4287 = n66990 & n4215 ;
  assign n66991 = ~n4216 ;
  assign n4288 = n4134 & n66991 ;
  assign n4289 = n4287 | n4288 ;
  assign n4290 = n66973 & n4289 ;
  assign n4291 = n66974 & n4290 ;
  assign n4292 = n4286 | n4291 ;
  assign n4293 = n66299 & n4292 ;
  assign n4294 = n3958 & n4183 ;
  assign n4128 = n3967 | n4127 ;
  assign n66992 = ~n4128 ;
  assign n4295 = n4124 & n66992 ;
  assign n66993 = ~n4129 ;
  assign n4296 = n4127 & n66993 ;
  assign n4297 = n4295 | n4296 ;
  assign n4298 = n66973 & n4297 ;
  assign n4299 = n66974 & n4298 ;
  assign n4300 = n4294 | n4299 ;
  assign n4301 = n66244 & n4300 ;
  assign n4302 = n3966 & n4183 ;
  assign n4123 = n3975 | n4122 ;
  assign n66994 = ~n4123 ;
  assign n4303 = n66994 & n4211 ;
  assign n66995 = ~n4212 ;
  assign n4304 = n4122 & n66995 ;
  assign n4305 = n4303 | n4304 ;
  assign n4306 = n66973 & n4305 ;
  assign n4307 = n66974 & n4306 ;
  assign n4308 = n4302 | n4307 ;
  assign n4309 = n66145 & n4308 ;
  assign n4310 = n3974 & n4183 ;
  assign n4116 = n3983 | n4115 ;
  assign n66996 = ~n4116 ;
  assign n4311 = n4112 & n66996 ;
  assign n66997 = ~n4117 ;
  assign n4312 = n4115 & n66997 ;
  assign n4313 = n4311 | n4312 ;
  assign n4314 = n66973 & n4313 ;
  assign n4315 = n66974 & n4314 ;
  assign n4316 = n4310 | n4315 ;
  assign n4317 = n66081 & n4316 ;
  assign n4318 = n3982 & n4183 ;
  assign n4111 = n3991 | n4110 ;
  assign n66998 = ~n4111 ;
  assign n4319 = n66998 & n4207 ;
  assign n66999 = ~n4208 ;
  assign n4320 = n4110 & n66999 ;
  assign n4321 = n4319 | n4320 ;
  assign n4322 = n66973 & n4321 ;
  assign n4323 = n66974 & n4322 ;
  assign n4324 = n4318 | n4323 ;
  assign n4325 = n66043 & n4324 ;
  assign n4326 = n3990 & n4183 ;
  assign n4104 = n3999 | n4103 ;
  assign n67000 = ~n4104 ;
  assign n4327 = n4100 & n67000 ;
  assign n67001 = ~n4105 ;
  assign n4328 = n4103 & n67001 ;
  assign n4329 = n4327 | n4328 ;
  assign n4330 = n66973 & n4329 ;
  assign n4331 = n66974 & n4330 ;
  assign n4332 = n4326 | n4331 ;
  assign n4333 = n65960 & n4332 ;
  assign n4334 = n3998 & n4183 ;
  assign n4099 = n4007 | n4098 ;
  assign n67002 = ~n4099 ;
  assign n4335 = n67002 & n4203 ;
  assign n67003 = ~n4204 ;
  assign n4336 = n4098 & n67003 ;
  assign n4337 = n4335 | n4336 ;
  assign n4338 = n66973 & n4337 ;
  assign n4339 = n66974 & n4338 ;
  assign n4340 = n4334 | n4339 ;
  assign n4341 = n65909 & n4340 ;
  assign n4342 = n4006 & n4183 ;
  assign n4092 = n4015 | n4091 ;
  assign n67004 = ~n4092 ;
  assign n4343 = n4088 & n67004 ;
  assign n67005 = ~n4093 ;
  assign n4344 = n4091 & n67005 ;
  assign n4345 = n4343 | n4344 ;
  assign n4346 = n66973 & n4345 ;
  assign n4347 = n66974 & n4346 ;
  assign n4348 = n4342 | n4347 ;
  assign n4349 = n65877 & n4348 ;
  assign n4350 = n4014 & n4183 ;
  assign n4087 = n4024 | n4086 ;
  assign n67006 = ~n4087 ;
  assign n4351 = n67006 & n4199 ;
  assign n67007 = ~n4200 ;
  assign n4352 = n4086 & n67007 ;
  assign n4353 = n4351 | n4352 ;
  assign n4354 = n66973 & n4353 ;
  assign n4355 = n66974 & n4354 ;
  assign n4356 = n4350 | n4355 ;
  assign n4357 = n65820 & n4356 ;
  assign n4358 = n4023 & n4183 ;
  assign n4186 = n4032 | n4080 ;
  assign n67008 = ~n4186 ;
  assign n4359 = n4077 & n67008 ;
  assign n67009 = ~n4081 ;
  assign n4360 = n4080 & n67009 ;
  assign n4361 = n4359 | n4360 ;
  assign n4362 = n66973 & n4361 ;
  assign n4363 = n66974 & n4362 ;
  assign n4364 = n4358 | n4363 ;
  assign n4365 = n65791 & n4364 ;
  assign n4366 = n4031 & n4183 ;
  assign n4367 = n4040 | n4076 ;
  assign n67010 = ~n4367 ;
  assign n4368 = n4195 & n67010 ;
  assign n67011 = ~n4196 ;
  assign n4369 = n4076 & n67011 ;
  assign n4370 = n4368 | n4369 ;
  assign n4371 = n66973 & n4370 ;
  assign n4372 = n66974 & n4371 ;
  assign n4373 = n4366 | n4372 ;
  assign n4374 = n65772 & n4373 ;
  assign n4375 = n4039 & n4183 ;
  assign n4376 = n4048 | n4070 ;
  assign n67012 = ~n4376 ;
  assign n4377 = n4193 & n67012 ;
  assign n67013 = ~n4071 ;
  assign n4378 = n4070 & n67013 ;
  assign n4379 = n4377 | n4378 ;
  assign n4380 = n66973 & n4379 ;
  assign n4381 = n66974 & n4380 ;
  assign n4382 = n4375 | n4381 ;
  assign n4383 = n65746 & n4382 ;
  assign n4384 = n4047 & n4183 ;
  assign n4191 = n4062 | n4066 ;
  assign n67014 = ~n4191 ;
  assign n4385 = n4060 & n67014 ;
  assign n67015 = ~n4192 ;
  assign n4386 = n4066 & n67015 ;
  assign n4387 = n4385 | n4386 ;
  assign n4388 = n66973 & n4387 ;
  assign n4389 = n66974 & n4388 ;
  assign n4390 = n4384 | n4389 ;
  assign n4391 = n65721 & n4390 ;
  assign n4185 = n4061 & n4183 ;
  assign n4189 = n4057 & n4058 ;
  assign n4392 = n66928 & n4189 ;
  assign n4393 = n4182 | n4392 ;
  assign n67016 = ~n4393 ;
  assign n4394 = n4060 & n67016 ;
  assign n4395 = n66974 & n4394 ;
  assign n4396 = n4185 | n4395 ;
  assign n4397 = n65686 & n4396 ;
  assign n67017 = ~n65579 ;
  assign n4406 = n67017 & n4058 ;
  assign n67018 = ~n65564 ;
  assign n4407 = n67018 & n4406 ;
  assign n67019 = ~n65647 ;
  assign n4408 = n67019 & n4407 ;
  assign n67020 = ~n65542 ;
  assign n4409 = n67020 & n4408 ;
  assign n67021 = ~n65429 ;
  assign n4410 = n67021 & n4409 ;
  assign n4411 = n66974 & n4410 ;
  assign n4398 = x64 & n66979 ;
  assign n67022 = ~n71642 ;
  assign n4399 = n67022 & n4398 ;
  assign n67023 = ~n74615 ;
  assign n4400 = n67023 & n4399 ;
  assign n67024 = ~n458 ;
  assign n4401 = n67024 & n4400 ;
  assign n67025 = ~n468 ;
  assign n4402 = n67025 & n4401 ;
  assign n67026 = ~n465 ;
  assign n4403 = n67026 & n4402 ;
  assign n4230 = n66968 & n4229 ;
  assign n4419 = n4175 | n4230 ;
  assign n4420 = n66969 & n4419 ;
  assign n67027 = ~n4420 ;
  assign n4421 = n4403 & n67027 ;
  assign n67028 = ~n4421 ;
  assign n4422 = x42 & n67028 ;
  assign n4423 = n4411 | n4422 ;
  assign n4424 = n65670 & n4423 ;
  assign n4404 = n66974 & n4403 ;
  assign n67029 = ~n4404 ;
  assign n4405 = x42 & n67029 ;
  assign n4412 = n4405 | n4411 ;
  assign n4413 = x65 & n4412 ;
  assign n4415 = x65 | n4411 ;
  assign n4416 = n4405 | n4415 ;
  assign n67030 = ~n4413 ;
  assign n4417 = n67030 & n4416 ;
  assign n67031 = ~x41 ;
  assign n4418 = n67031 & x64 ;
  assign n4425 = n4417 | n4418 ;
  assign n67032 = ~n4424 ;
  assign n4426 = n67032 & n4425 ;
  assign n67033 = ~n4395 ;
  assign n4427 = x66 & n67033 ;
  assign n67034 = ~n4185 ;
  assign n4428 = n67034 & n4427 ;
  assign n4429 = n4397 | n4428 ;
  assign n4430 = n4426 | n4429 ;
  assign n67035 = ~n4397 ;
  assign n4431 = n67035 & n4430 ;
  assign n67036 = ~n4389 ;
  assign n4432 = x67 & n67036 ;
  assign n67037 = ~n4384 ;
  assign n4433 = n67037 & n4432 ;
  assign n4434 = n4391 | n4433 ;
  assign n4435 = n4431 | n4434 ;
  assign n67038 = ~n4391 ;
  assign n4436 = n67038 & n4435 ;
  assign n67039 = ~n4381 ;
  assign n4437 = x68 & n67039 ;
  assign n67040 = ~n4375 ;
  assign n4438 = n67040 & n4437 ;
  assign n4439 = n4383 | n4438 ;
  assign n4440 = n4436 | n4439 ;
  assign n67041 = ~n4383 ;
  assign n4441 = n67041 & n4440 ;
  assign n67042 = ~n4372 ;
  assign n4442 = x69 & n67042 ;
  assign n67043 = ~n4366 ;
  assign n4443 = n67043 & n4442 ;
  assign n4444 = n4374 | n4443 ;
  assign n4445 = n4441 | n4444 ;
  assign n67044 = ~n4374 ;
  assign n4446 = n67044 & n4445 ;
  assign n67045 = ~n4363 ;
  assign n4447 = x70 & n67045 ;
  assign n67046 = ~n4358 ;
  assign n4448 = n67046 & n4447 ;
  assign n4449 = n4365 | n4448 ;
  assign n4451 = n4446 | n4449 ;
  assign n67047 = ~n4365 ;
  assign n4452 = n67047 & n4451 ;
  assign n67048 = ~n4355 ;
  assign n4453 = x71 & n67048 ;
  assign n67049 = ~n4350 ;
  assign n4454 = n67049 & n4453 ;
  assign n4455 = n4357 | n4454 ;
  assign n4456 = n4452 | n4455 ;
  assign n67050 = ~n4357 ;
  assign n4457 = n67050 & n4456 ;
  assign n67051 = ~n4347 ;
  assign n4458 = x72 & n67051 ;
  assign n67052 = ~n4342 ;
  assign n4459 = n67052 & n4458 ;
  assign n4460 = n4349 | n4459 ;
  assign n4462 = n4457 | n4460 ;
  assign n67053 = ~n4349 ;
  assign n4463 = n67053 & n4462 ;
  assign n67054 = ~n4339 ;
  assign n4464 = x73 & n67054 ;
  assign n67055 = ~n4334 ;
  assign n4465 = n67055 & n4464 ;
  assign n4466 = n4341 | n4465 ;
  assign n4467 = n4463 | n4466 ;
  assign n67056 = ~n4341 ;
  assign n4468 = n67056 & n4467 ;
  assign n67057 = ~n4331 ;
  assign n4469 = x74 & n67057 ;
  assign n67058 = ~n4326 ;
  assign n4470 = n67058 & n4469 ;
  assign n4471 = n4333 | n4470 ;
  assign n4473 = n4468 | n4471 ;
  assign n67059 = ~n4333 ;
  assign n4474 = n67059 & n4473 ;
  assign n67060 = ~n4323 ;
  assign n4475 = x75 & n67060 ;
  assign n67061 = ~n4318 ;
  assign n4476 = n67061 & n4475 ;
  assign n4477 = n4325 | n4476 ;
  assign n4478 = n4474 | n4477 ;
  assign n67062 = ~n4325 ;
  assign n4479 = n67062 & n4478 ;
  assign n67063 = ~n4315 ;
  assign n4480 = x76 & n67063 ;
  assign n67064 = ~n4310 ;
  assign n4481 = n67064 & n4480 ;
  assign n4482 = n4317 | n4481 ;
  assign n4484 = n4479 | n4482 ;
  assign n67065 = ~n4317 ;
  assign n4485 = n67065 & n4484 ;
  assign n67066 = ~n4307 ;
  assign n4486 = x77 & n67066 ;
  assign n67067 = ~n4302 ;
  assign n4487 = n67067 & n4486 ;
  assign n4488 = n4309 | n4487 ;
  assign n4489 = n4485 | n4488 ;
  assign n67068 = ~n4309 ;
  assign n4490 = n67068 & n4489 ;
  assign n67069 = ~n4299 ;
  assign n4491 = x78 & n67069 ;
  assign n67070 = ~n4294 ;
  assign n4492 = n67070 & n4491 ;
  assign n4493 = n4301 | n4492 ;
  assign n4495 = n4490 | n4493 ;
  assign n67071 = ~n4301 ;
  assign n4496 = n67071 & n4495 ;
  assign n67072 = ~n4291 ;
  assign n4497 = x79 & n67072 ;
  assign n67073 = ~n4286 ;
  assign n4498 = n67073 & n4497 ;
  assign n4499 = n4293 | n4498 ;
  assign n4500 = n4496 | n4499 ;
  assign n67074 = ~n4293 ;
  assign n4501 = n67074 & n4500 ;
  assign n67075 = ~n4283 ;
  assign n4502 = x80 & n67075 ;
  assign n67076 = ~n4278 ;
  assign n4503 = n67076 & n4502 ;
  assign n4504 = n4285 | n4503 ;
  assign n4506 = n4501 | n4504 ;
  assign n67077 = ~n4285 ;
  assign n4507 = n67077 & n4506 ;
  assign n67078 = ~n4275 ;
  assign n4508 = x81 & n67078 ;
  assign n67079 = ~n4270 ;
  assign n4509 = n67079 & n4508 ;
  assign n4510 = n4277 | n4509 ;
  assign n4511 = n4507 | n4510 ;
  assign n67080 = ~n4277 ;
  assign n4512 = n67080 & n4511 ;
  assign n67081 = ~n4267 ;
  assign n4513 = x82 & n67081 ;
  assign n67082 = ~n4262 ;
  assign n4514 = n67082 & n4513 ;
  assign n4515 = n4269 | n4514 ;
  assign n4517 = n4512 | n4515 ;
  assign n67083 = ~n4269 ;
  assign n4518 = n67083 & n4517 ;
  assign n67084 = ~n4259 ;
  assign n4519 = x83 & n67084 ;
  assign n67085 = ~n4254 ;
  assign n4520 = n67085 & n4519 ;
  assign n4521 = n4261 | n4520 ;
  assign n4522 = n4518 | n4521 ;
  assign n67086 = ~n4261 ;
  assign n4523 = n67086 & n4522 ;
  assign n67087 = ~n4251 ;
  assign n4524 = x84 & n67087 ;
  assign n67088 = ~n4246 ;
  assign n4525 = n67088 & n4524 ;
  assign n4526 = n4253 | n4525 ;
  assign n4528 = n4523 | n4526 ;
  assign n67089 = ~n4253 ;
  assign n4529 = n67089 & n4528 ;
  assign n67090 = ~n4243 ;
  assign n4530 = x85 & n67090 ;
  assign n67091 = ~n4238 ;
  assign n4531 = n67091 & n4530 ;
  assign n4532 = n4245 | n4531 ;
  assign n4533 = n4529 | n4532 ;
  assign n67092 = ~n4245 ;
  assign n4534 = n67092 & n4533 ;
  assign n171 = ~n4183 ;
  assign n4535 = n171 & n4234 ;
  assign n4536 = n3894 & n4183 ;
  assign n67094 = ~n4536 ;
  assign n4537 = x86 & n67094 ;
  assign n67095 = ~n4535 ;
  assign n4538 = n67095 & n4537 ;
  assign n4539 = n4237 | n4538 ;
  assign n4541 = n4534 | n4539 ;
  assign n67096 = ~n4237 ;
  assign n4542 = n67096 & n4541 ;
  assign n4543 = n71642 | n74615 ;
  assign n4544 = n458 | n4543 ;
  assign n4545 = n468 | n4544 ;
  assign n4546 = n465 | n4545 ;
  assign n4547 = n4542 | n4546 ;
  assign n4548 = n4244 & n4547 ;
  assign n4414 = n65670 & n4412 ;
  assign n4549 = x65 & n4423 ;
  assign n67097 = ~n4549 ;
  assign n4550 = n4416 & n67097 ;
  assign n4551 = n4418 | n4550 ;
  assign n67098 = ~n4414 ;
  assign n4552 = n67098 & n4551 ;
  assign n4553 = n4429 | n4552 ;
  assign n4554 = n67035 & n4553 ;
  assign n4555 = n4433 | n4554 ;
  assign n4557 = n67038 & n4555 ;
  assign n4559 = n4439 | n4557 ;
  assign n4560 = n67041 & n4559 ;
  assign n4562 = n4444 | n4560 ;
  assign n4563 = n67044 & n4562 ;
  assign n4564 = n4449 | n4563 ;
  assign n4565 = n67047 & n4564 ;
  assign n4566 = n4455 | n4565 ;
  assign n4568 = n67050 & n4566 ;
  assign n4569 = n4460 | n4568 ;
  assign n4570 = n67053 & n4569 ;
  assign n4571 = n4466 | n4570 ;
  assign n4573 = n67056 & n4571 ;
  assign n4574 = n4471 | n4573 ;
  assign n4575 = n67059 & n4574 ;
  assign n4576 = n4477 | n4575 ;
  assign n4578 = n67062 & n4576 ;
  assign n4579 = n4482 | n4578 ;
  assign n4580 = n67065 & n4579 ;
  assign n4581 = n4488 | n4580 ;
  assign n4583 = n67068 & n4581 ;
  assign n4584 = n4493 | n4583 ;
  assign n4585 = n67071 & n4584 ;
  assign n4586 = n4499 | n4585 ;
  assign n4588 = n67074 & n4586 ;
  assign n4589 = n4504 | n4588 ;
  assign n4590 = n67077 & n4589 ;
  assign n4591 = n4510 | n4590 ;
  assign n4593 = n67080 & n4591 ;
  assign n4594 = n4515 | n4593 ;
  assign n4595 = n67083 & n4594 ;
  assign n4596 = n4521 | n4595 ;
  assign n4598 = n67086 & n4596 ;
  assign n4599 = n4526 | n4598 ;
  assign n4600 = n67089 & n4599 ;
  assign n67099 = ~n4600 ;
  assign n4601 = n4532 & n67099 ;
  assign n4603 = n4253 | n4532 ;
  assign n67100 = ~n4603 ;
  assign n4604 = n4528 & n67100 ;
  assign n4605 = n4601 | n4604 ;
  assign n67101 = ~n4546 ;
  assign n4606 = n67101 & n4605 ;
  assign n67102 = ~n4542 ;
  assign n4607 = n67102 & n4606 ;
  assign n4608 = n4548 | n4607 ;
  assign n4609 = n66979 & n4608 ;
  assign n67103 = ~n4607 ;
  assign n4897 = x86 & n67103 ;
  assign n67104 = ~n4548 ;
  assign n4898 = n67104 & n4897 ;
  assign n4899 = n4609 | n4898 ;
  assign n4610 = n4252 & n4547 ;
  assign n67105 = ~n4523 ;
  assign n4527 = n67105 & n4526 ;
  assign n4611 = n4261 | n4526 ;
  assign n67106 = ~n4611 ;
  assign n4612 = n4596 & n67106 ;
  assign n4613 = n4527 | n4612 ;
  assign n4614 = n67101 & n4613 ;
  assign n4615 = n67102 & n4614 ;
  assign n4616 = n4610 | n4615 ;
  assign n4617 = n66868 & n4616 ;
  assign n4618 = n4260 & n4547 ;
  assign n67107 = ~n4595 ;
  assign n4597 = n4521 & n67107 ;
  assign n4619 = n4269 | n4521 ;
  assign n67108 = ~n4619 ;
  assign n4620 = n4517 & n67108 ;
  assign n4621 = n4597 | n4620 ;
  assign n4622 = n67101 & n4621 ;
  assign n4623 = n67102 & n4622 ;
  assign n4624 = n4618 | n4623 ;
  assign n4625 = n66797 & n4624 ;
  assign n67109 = ~n4623 ;
  assign n4886 = x84 & n67109 ;
  assign n67110 = ~n4618 ;
  assign n4887 = n67110 & n4886 ;
  assign n4888 = n4625 | n4887 ;
  assign n4626 = n4268 & n4547 ;
  assign n67111 = ~n4512 ;
  assign n4516 = n67111 & n4515 ;
  assign n4627 = n4277 | n4515 ;
  assign n67112 = ~n4627 ;
  assign n4628 = n4591 & n67112 ;
  assign n4629 = n4516 | n4628 ;
  assign n4630 = n67101 & n4629 ;
  assign n4631 = n67102 & n4630 ;
  assign n4632 = n4626 | n4631 ;
  assign n4633 = n66654 & n4632 ;
  assign n4634 = n4276 & n4547 ;
  assign n67113 = ~n4590 ;
  assign n4592 = n4510 & n67113 ;
  assign n4635 = n4285 | n4510 ;
  assign n67114 = ~n4635 ;
  assign n4636 = n4506 & n67114 ;
  assign n4637 = n4592 | n4636 ;
  assign n4638 = n67101 & n4637 ;
  assign n4639 = n67102 & n4638 ;
  assign n4640 = n4634 | n4639 ;
  assign n4641 = n66560 & n4640 ;
  assign n67115 = ~n4639 ;
  assign n4876 = x82 & n67115 ;
  assign n67116 = ~n4634 ;
  assign n4877 = n67116 & n4876 ;
  assign n4878 = n4641 | n4877 ;
  assign n4642 = n4284 & n4547 ;
  assign n67117 = ~n4501 ;
  assign n4505 = n67117 & n4504 ;
  assign n4643 = n4293 | n4504 ;
  assign n67118 = ~n4643 ;
  assign n4644 = n4586 & n67118 ;
  assign n4645 = n4505 | n4644 ;
  assign n4646 = n67101 & n4645 ;
  assign n4647 = n67102 & n4646 ;
  assign n4648 = n4642 | n4647 ;
  assign n4649 = n66505 & n4648 ;
  assign n4650 = n4292 & n4547 ;
  assign n67119 = ~n4585 ;
  assign n4587 = n4499 & n67119 ;
  assign n4651 = n4301 | n4499 ;
  assign n67120 = ~n4651 ;
  assign n4652 = n4495 & n67120 ;
  assign n4653 = n4587 | n4652 ;
  assign n4654 = n67101 & n4653 ;
  assign n4655 = n67102 & n4654 ;
  assign n4656 = n4650 | n4655 ;
  assign n4657 = n66379 & n4656 ;
  assign n67121 = ~n4655 ;
  assign n4866 = x80 & n67121 ;
  assign n67122 = ~n4650 ;
  assign n4867 = n67122 & n4866 ;
  assign n4868 = n4657 | n4867 ;
  assign n4658 = n4300 & n4547 ;
  assign n67123 = ~n4490 ;
  assign n4494 = n67123 & n4493 ;
  assign n4659 = n4309 | n4493 ;
  assign n67124 = ~n4659 ;
  assign n4660 = n4581 & n67124 ;
  assign n4661 = n4494 | n4660 ;
  assign n4662 = n67101 & n4661 ;
  assign n4663 = n67102 & n4662 ;
  assign n4664 = n4658 | n4663 ;
  assign n4665 = n66299 & n4664 ;
  assign n4666 = n4308 & n4547 ;
  assign n67125 = ~n4580 ;
  assign n4582 = n4488 & n67125 ;
  assign n4667 = n4317 | n4488 ;
  assign n67126 = ~n4667 ;
  assign n4668 = n4484 & n67126 ;
  assign n4669 = n4582 | n4668 ;
  assign n4670 = n67101 & n4669 ;
  assign n4671 = n67102 & n4670 ;
  assign n4672 = n4666 | n4671 ;
  assign n4673 = n66244 & n4672 ;
  assign n67127 = ~n4671 ;
  assign n4856 = x78 & n67127 ;
  assign n67128 = ~n4666 ;
  assign n4857 = n67128 & n4856 ;
  assign n4858 = n4673 | n4857 ;
  assign n4674 = n4316 & n4547 ;
  assign n67129 = ~n4479 ;
  assign n4483 = n67129 & n4482 ;
  assign n4675 = n4325 | n4482 ;
  assign n67130 = ~n4675 ;
  assign n4676 = n4576 & n67130 ;
  assign n4677 = n4483 | n4676 ;
  assign n4678 = n67101 & n4677 ;
  assign n4679 = n67102 & n4678 ;
  assign n4680 = n4674 | n4679 ;
  assign n4681 = n66145 & n4680 ;
  assign n4682 = n4324 & n4547 ;
  assign n67131 = ~n4575 ;
  assign n4577 = n4477 & n67131 ;
  assign n4683 = n4333 | n4477 ;
  assign n67132 = ~n4683 ;
  assign n4684 = n4473 & n67132 ;
  assign n4685 = n4577 | n4684 ;
  assign n4686 = n67101 & n4685 ;
  assign n4687 = n67102 & n4686 ;
  assign n4688 = n4682 | n4687 ;
  assign n4689 = n66081 & n4688 ;
  assign n67133 = ~n4687 ;
  assign n4846 = x76 & n67133 ;
  assign n67134 = ~n4682 ;
  assign n4847 = n67134 & n4846 ;
  assign n4848 = n4689 | n4847 ;
  assign n4690 = n4332 & n4547 ;
  assign n67135 = ~n4468 ;
  assign n4472 = n67135 & n4471 ;
  assign n4691 = n4341 | n4471 ;
  assign n67136 = ~n4691 ;
  assign n4692 = n4571 & n67136 ;
  assign n4693 = n4472 | n4692 ;
  assign n4694 = n67101 & n4693 ;
  assign n4695 = n67102 & n4694 ;
  assign n4696 = n4690 | n4695 ;
  assign n4697 = n66043 & n4696 ;
  assign n4698 = n4340 & n4547 ;
  assign n67137 = ~n4570 ;
  assign n4572 = n4466 & n67137 ;
  assign n4699 = n4349 | n4466 ;
  assign n67138 = ~n4699 ;
  assign n4700 = n4462 & n67138 ;
  assign n4701 = n4572 | n4700 ;
  assign n4702 = n67101 & n4701 ;
  assign n4703 = n67102 & n4702 ;
  assign n4704 = n4698 | n4703 ;
  assign n4705 = n65960 & n4704 ;
  assign n67139 = ~n4703 ;
  assign n4836 = x74 & n67139 ;
  assign n67140 = ~n4698 ;
  assign n4837 = n67140 & n4836 ;
  assign n4838 = n4705 | n4837 ;
  assign n4706 = n4348 & n4547 ;
  assign n67141 = ~n4457 ;
  assign n4461 = n67141 & n4460 ;
  assign n4707 = n4357 | n4460 ;
  assign n67142 = ~n4707 ;
  assign n4708 = n4566 & n67142 ;
  assign n4709 = n4461 | n4708 ;
  assign n4710 = n67101 & n4709 ;
  assign n4711 = n67102 & n4710 ;
  assign n4712 = n4706 | n4711 ;
  assign n4713 = n65909 & n4712 ;
  assign n4714 = n4356 & n4547 ;
  assign n67143 = ~n4565 ;
  assign n4567 = n4455 & n67143 ;
  assign n4715 = n4365 | n4455 ;
  assign n67144 = ~n4715 ;
  assign n4716 = n4451 & n67144 ;
  assign n4717 = n4567 | n4716 ;
  assign n4718 = n67101 & n4717 ;
  assign n4719 = n67102 & n4718 ;
  assign n4720 = n4714 | n4719 ;
  assign n4721 = n65877 & n4720 ;
  assign n67145 = ~n4719 ;
  assign n4826 = x72 & n67145 ;
  assign n67146 = ~n4714 ;
  assign n4827 = n67146 & n4826 ;
  assign n4828 = n4721 | n4827 ;
  assign n4722 = n4364 & n4547 ;
  assign n67147 = ~n4446 ;
  assign n4450 = n67147 & n4449 ;
  assign n4723 = n4374 | n4449 ;
  assign n67148 = ~n4723 ;
  assign n4724 = n4562 & n67148 ;
  assign n4725 = n4450 | n4724 ;
  assign n4726 = n67101 & n4725 ;
  assign n4727 = n67102 & n4726 ;
  assign n4728 = n4722 | n4727 ;
  assign n4729 = n65820 & n4728 ;
  assign n4730 = n4373 & n4547 ;
  assign n67149 = ~n4560 ;
  assign n4561 = n4444 & n67149 ;
  assign n4731 = n4383 | n4444 ;
  assign n67150 = ~n4731 ;
  assign n4732 = n4559 & n67150 ;
  assign n4733 = n4561 | n4732 ;
  assign n4734 = n67101 & n4733 ;
  assign n4735 = n67102 & n4734 ;
  assign n4736 = n4730 | n4735 ;
  assign n4737 = n65791 & n4736 ;
  assign n67151 = ~n4735 ;
  assign n4816 = x70 & n67151 ;
  assign n67152 = ~n4730 ;
  assign n4817 = n67152 & n4816 ;
  assign n4818 = n4737 | n4817 ;
  assign n4738 = n4382 & n4547 ;
  assign n67153 = ~n4436 ;
  assign n4558 = n67153 & n4439 ;
  assign n4739 = n4434 | n4554 ;
  assign n4740 = n4391 | n4439 ;
  assign n67154 = ~n4740 ;
  assign n4741 = n4739 & n67154 ;
  assign n4742 = n4558 | n4741 ;
  assign n4743 = n67101 & n4742 ;
  assign n4744 = n67102 & n4743 ;
  assign n4745 = n4738 | n4744 ;
  assign n4746 = n65772 & n4745 ;
  assign n4747 = n4390 & n4547 ;
  assign n67155 = ~n4554 ;
  assign n4556 = n4434 & n67155 ;
  assign n4748 = n4397 | n4434 ;
  assign n67156 = ~n4748 ;
  assign n4749 = n4553 & n67156 ;
  assign n4750 = n4556 | n4749 ;
  assign n4751 = n67101 & n4750 ;
  assign n4752 = n67102 & n4751 ;
  assign n4753 = n4747 | n4752 ;
  assign n4754 = n65746 & n4753 ;
  assign n67157 = ~n4752 ;
  assign n4806 = x68 & n67157 ;
  assign n67158 = ~n4747 ;
  assign n4807 = n67158 & n4806 ;
  assign n4808 = n4754 | n4807 ;
  assign n4755 = n4396 & n4547 ;
  assign n4756 = n4424 | n4429 ;
  assign n67159 = ~n4756 ;
  assign n4757 = n4551 & n67159 ;
  assign n67160 = ~n4426 ;
  assign n4758 = n67160 & n4429 ;
  assign n4759 = n4757 | n4758 ;
  assign n4760 = n67101 & n4759 ;
  assign n4761 = n67102 & n4760 ;
  assign n4762 = n4755 | n4761 ;
  assign n4764 = n65721 & n4762 ;
  assign n4765 = n4412 & n4547 ;
  assign n4766 = n4416 & n4418 ;
  assign n4767 = n67097 & n4766 ;
  assign n4768 = n4546 | n4767 ;
  assign n67161 = ~n4768 ;
  assign n4769 = n4551 & n67161 ;
  assign n4770 = n67102 & n4769 ;
  assign n4771 = n4765 | n4770 ;
  assign n4772 = n65686 & n4771 ;
  assign n67162 = ~n4770 ;
  assign n4797 = x66 & n67162 ;
  assign n67163 = ~n4765 ;
  assign n4798 = n67163 & n4797 ;
  assign n4799 = n4772 | n4798 ;
  assign n4602 = n4532 | n4600 ;
  assign n4773 = n67092 & n4602 ;
  assign n4774 = n4539 | n4773 ;
  assign n4775 = n67096 & n4774 ;
  assign n67164 = ~x87 ;
  assign n4776 = x64 & n67164 ;
  assign n4777 = n67018 & n4776 ;
  assign n4778 = n67019 & n4777 ;
  assign n4779 = n67020 & n4778 ;
  assign n4780 = n67021 & n4779 ;
  assign n67165 = ~n4775 ;
  assign n4781 = n67165 & n4780 ;
  assign n67166 = ~n4781 ;
  assign n4782 = x41 & n67166 ;
  assign n4783 = n67022 & n4418 ;
  assign n4784 = n67023 & n4783 ;
  assign n4785 = n67024 & n4784 ;
  assign n4786 = n67025 & n4785 ;
  assign n4787 = n67026 & n4786 ;
  assign n4788 = n67102 & n4787 ;
  assign n4789 = n4782 | n4788 ;
  assign n4790 = x65 & n4789 ;
  assign n4791 = x65 | n4788 ;
  assign n4792 = n4782 | n4791 ;
  assign n67167 = ~n4790 ;
  assign n4793 = n67167 & n4792 ;
  assign n67168 = ~x40 ;
  assign n4794 = n67168 & x64 ;
  assign n4795 = n4793 | n4794 ;
  assign n4796 = n65670 & n4789 ;
  assign n67169 = ~n4796 ;
  assign n4800 = n4795 & n67169 ;
  assign n4801 = n4799 | n4800 ;
  assign n67170 = ~n4772 ;
  assign n4802 = n67170 & n4801 ;
  assign n67171 = ~n4761 ;
  assign n4763 = x67 & n67171 ;
  assign n67172 = ~n4755 ;
  assign n4803 = n67172 & n4763 ;
  assign n4804 = n4764 | n4803 ;
  assign n4805 = n4802 | n4804 ;
  assign n67173 = ~n4764 ;
  assign n4809 = n67173 & n4805 ;
  assign n4810 = n4808 | n4809 ;
  assign n67174 = ~n4754 ;
  assign n4811 = n67174 & n4810 ;
  assign n67175 = ~n4744 ;
  assign n4812 = x69 & n67175 ;
  assign n67176 = ~n4738 ;
  assign n4813 = n67176 & n4812 ;
  assign n4814 = n4746 | n4813 ;
  assign n4815 = n4811 | n4814 ;
  assign n67177 = ~n4746 ;
  assign n4819 = n67177 & n4815 ;
  assign n4820 = n4818 | n4819 ;
  assign n67178 = ~n4737 ;
  assign n4821 = n67178 & n4820 ;
  assign n67179 = ~n4727 ;
  assign n4822 = x71 & n67179 ;
  assign n67180 = ~n4722 ;
  assign n4823 = n67180 & n4822 ;
  assign n4824 = n4729 | n4823 ;
  assign n4825 = n4821 | n4824 ;
  assign n67181 = ~n4729 ;
  assign n4829 = n67181 & n4825 ;
  assign n4830 = n4828 | n4829 ;
  assign n67182 = ~n4721 ;
  assign n4831 = n67182 & n4830 ;
  assign n67183 = ~n4711 ;
  assign n4832 = x73 & n67183 ;
  assign n67184 = ~n4706 ;
  assign n4833 = n67184 & n4832 ;
  assign n4834 = n4713 | n4833 ;
  assign n4835 = n4831 | n4834 ;
  assign n67185 = ~n4713 ;
  assign n4839 = n67185 & n4835 ;
  assign n4840 = n4838 | n4839 ;
  assign n67186 = ~n4705 ;
  assign n4841 = n67186 & n4840 ;
  assign n67187 = ~n4695 ;
  assign n4842 = x75 & n67187 ;
  assign n67188 = ~n4690 ;
  assign n4843 = n67188 & n4842 ;
  assign n4844 = n4697 | n4843 ;
  assign n4845 = n4841 | n4844 ;
  assign n67189 = ~n4697 ;
  assign n4849 = n67189 & n4845 ;
  assign n4850 = n4848 | n4849 ;
  assign n67190 = ~n4689 ;
  assign n4851 = n67190 & n4850 ;
  assign n67191 = ~n4679 ;
  assign n4852 = x77 & n67191 ;
  assign n67192 = ~n4674 ;
  assign n4853 = n67192 & n4852 ;
  assign n4854 = n4681 | n4853 ;
  assign n4855 = n4851 | n4854 ;
  assign n67193 = ~n4681 ;
  assign n4859 = n67193 & n4855 ;
  assign n4860 = n4858 | n4859 ;
  assign n67194 = ~n4673 ;
  assign n4861 = n67194 & n4860 ;
  assign n67195 = ~n4663 ;
  assign n4862 = x79 & n67195 ;
  assign n67196 = ~n4658 ;
  assign n4863 = n67196 & n4862 ;
  assign n4864 = n4665 | n4863 ;
  assign n4865 = n4861 | n4864 ;
  assign n67197 = ~n4665 ;
  assign n4869 = n67197 & n4865 ;
  assign n4870 = n4868 | n4869 ;
  assign n67198 = ~n4657 ;
  assign n4871 = n67198 & n4870 ;
  assign n67199 = ~n4647 ;
  assign n4872 = x81 & n67199 ;
  assign n67200 = ~n4642 ;
  assign n4873 = n67200 & n4872 ;
  assign n4874 = n4649 | n4873 ;
  assign n4875 = n4871 | n4874 ;
  assign n67201 = ~n4649 ;
  assign n4879 = n67201 & n4875 ;
  assign n4880 = n4878 | n4879 ;
  assign n67202 = ~n4641 ;
  assign n4881 = n67202 & n4880 ;
  assign n67203 = ~n4631 ;
  assign n4882 = x83 & n67203 ;
  assign n67204 = ~n4626 ;
  assign n4883 = n67204 & n4882 ;
  assign n4884 = n4633 | n4883 ;
  assign n4885 = n4881 | n4884 ;
  assign n67205 = ~n4633 ;
  assign n4889 = n67205 & n4885 ;
  assign n4890 = n4888 | n4889 ;
  assign n67206 = ~n4625 ;
  assign n4891 = n67206 & n4890 ;
  assign n67207 = ~n4615 ;
  assign n4892 = x85 & n67207 ;
  assign n67208 = ~n4610 ;
  assign n4893 = n67208 & n4892 ;
  assign n4894 = n4617 | n4893 ;
  assign n4896 = n4891 | n4894 ;
  assign n67209 = ~n4617 ;
  assign n4900 = n67209 & n4896 ;
  assign n4901 = n4899 | n4900 ;
  assign n67210 = ~n4609 ;
  assign n4902 = n67210 & n4901 ;
  assign n67211 = ~n4534 ;
  assign n4540 = n67211 & n4539 ;
  assign n4903 = n4245 | n4539 ;
  assign n67212 = ~n4903 ;
  assign n4904 = n4602 & n67212 ;
  assign n4905 = n4540 | n4904 ;
  assign n4906 = n4547 | n4905 ;
  assign n67213 = ~n4236 ;
  assign n4907 = n67213 & n4547 ;
  assign n67214 = ~n4907 ;
  assign n4908 = n4906 & n67214 ;
  assign n4909 = n67164 & n4908 ;
  assign n170 = ~n4547 ;
  assign n4910 = n170 & n4905 ;
  assign n4911 = n4236 & n4547 ;
  assign n67216 = ~n4911 ;
  assign n4912 = x87 & n67216 ;
  assign n67217 = ~n4910 ;
  assign n4913 = n67217 & n4912 ;
  assign n4914 = n67215 | n67349 ;
  assign n4915 = n66858 | n4914 ;
  assign n4916 = n4913 | n4915 ;
  assign n4917 = n4909 | n4916 ;
  assign n4918 = n4902 | n4917 ;
  assign n4919 = n67101 & n4908 ;
  assign n67218 = ~n4919 ;
  assign n4920 = n4918 & n67218 ;
  assign n4922 = n4609 | n4913 ;
  assign n4923 = n4909 | n4922 ;
  assign n67219 = ~n4923 ;
  assign n4924 = n4901 & n67219 ;
  assign n4925 = n4909 | n4913 ;
  assign n67220 = ~n4902 ;
  assign n4926 = n67220 & n4925 ;
  assign n4927 = n4924 | n4926 ;
  assign n169 = ~n4920 ;
  assign n4928 = n169 & n4927 ;
  assign n4929 = n4546 & n4908 ;
  assign n4930 = n4918 & n4929 ;
  assign n4931 = n4928 | n4930 ;
  assign n67222 = ~x88 ;
  assign n4932 = n67222 & n4931 ;
  assign n67223 = ~n4900 ;
  assign n4981 = n4899 & n67223 ;
  assign n4933 = n67102 & n4780 ;
  assign n67224 = ~n4933 ;
  assign n4934 = x41 & n67224 ;
  assign n4935 = n4788 | n4934 ;
  assign n4936 = x65 & n4935 ;
  assign n67225 = ~n4936 ;
  assign n4937 = n4792 & n67225 ;
  assign n4938 = n4794 | n4937 ;
  assign n4939 = n67169 & n4938 ;
  assign n4941 = n4799 | n4939 ;
  assign n4942 = n67170 & n4941 ;
  assign n4943 = n4804 | n4942 ;
  assign n4944 = n67173 & n4943 ;
  assign n4945 = n4808 | n4944 ;
  assign n4946 = n67174 & n4945 ;
  assign n4947 = n4814 | n4946 ;
  assign n4948 = n67177 & n4947 ;
  assign n4949 = n4818 | n4948 ;
  assign n4950 = n67178 & n4949 ;
  assign n4951 = n4824 | n4950 ;
  assign n4952 = n67181 & n4951 ;
  assign n4953 = n4828 | n4952 ;
  assign n4954 = n67182 & n4953 ;
  assign n4955 = n4834 | n4954 ;
  assign n4956 = n67185 & n4955 ;
  assign n4957 = n4838 | n4956 ;
  assign n4958 = n67186 & n4957 ;
  assign n4959 = n4844 | n4958 ;
  assign n4960 = n67189 & n4959 ;
  assign n4961 = n4848 | n4960 ;
  assign n4962 = n67190 & n4961 ;
  assign n4963 = n4854 | n4962 ;
  assign n4964 = n67193 & n4963 ;
  assign n4965 = n4858 | n4964 ;
  assign n4966 = n67194 & n4965 ;
  assign n4967 = n4864 | n4966 ;
  assign n4968 = n67197 & n4967 ;
  assign n4969 = n4868 | n4968 ;
  assign n4970 = n67198 & n4969 ;
  assign n4971 = n4874 | n4970 ;
  assign n4972 = n67201 & n4971 ;
  assign n4973 = n4878 | n4972 ;
  assign n4974 = n67202 & n4973 ;
  assign n4975 = n4884 | n4974 ;
  assign n4976 = n67205 & n4975 ;
  assign n4977 = n4888 | n4976 ;
  assign n4978 = n67206 & n4977 ;
  assign n4979 = n4894 | n4978 ;
  assign n4982 = n4617 | n4899 ;
  assign n67226 = ~n4982 ;
  assign n4983 = n4979 & n67226 ;
  assign n4984 = n4981 | n4983 ;
  assign n4985 = n169 & n4984 ;
  assign n4986 = n4608 & n67218 ;
  assign n4987 = n4918 & n4986 ;
  assign n4988 = n4985 | n4987 ;
  assign n4989 = n67164 & n4988 ;
  assign n67227 = ~n4978 ;
  assign n4990 = n4894 & n67227 ;
  assign n4895 = n4625 | n4894 ;
  assign n67228 = ~n4895 ;
  assign n4991 = n67228 & n4977 ;
  assign n4992 = n4990 | n4991 ;
  assign n4993 = n169 & n4992 ;
  assign n4994 = n4616 & n67218 ;
  assign n4995 = n4918 & n4994 ;
  assign n4996 = n4993 | n4995 ;
  assign n4997 = n66979 & n4996 ;
  assign n67229 = ~n4889 ;
  assign n4998 = n4888 & n67229 ;
  assign n4999 = n4633 | n4888 ;
  assign n67230 = ~n4999 ;
  assign n5000 = n4975 & n67230 ;
  assign n5001 = n4998 | n5000 ;
  assign n5002 = n169 & n5001 ;
  assign n5003 = n4624 & n67218 ;
  assign n5004 = n4918 & n5003 ;
  assign n5005 = n5002 | n5004 ;
  assign n5006 = n66868 & n5005 ;
  assign n67231 = ~n4974 ;
  assign n5007 = n4884 & n67231 ;
  assign n5008 = n4641 | n4884 ;
  assign n67232 = ~n5008 ;
  assign n5009 = n4880 & n67232 ;
  assign n5010 = n5007 | n5009 ;
  assign n5011 = n169 & n5010 ;
  assign n5012 = n4632 & n67218 ;
  assign n5013 = n4918 & n5012 ;
  assign n5014 = n5011 | n5013 ;
  assign n5015 = n66797 & n5014 ;
  assign n67233 = ~n4879 ;
  assign n5016 = n4878 & n67233 ;
  assign n5017 = n4649 | n4878 ;
  assign n67234 = ~n5017 ;
  assign n5018 = n4971 & n67234 ;
  assign n5019 = n5016 | n5018 ;
  assign n5020 = n169 & n5019 ;
  assign n5021 = n4640 & n67218 ;
  assign n5022 = n4918 & n5021 ;
  assign n5023 = n5020 | n5022 ;
  assign n5024 = n66654 & n5023 ;
  assign n67235 = ~n4970 ;
  assign n5025 = n4874 & n67235 ;
  assign n5026 = n4657 | n4874 ;
  assign n67236 = ~n5026 ;
  assign n5027 = n4870 & n67236 ;
  assign n5028 = n5025 | n5027 ;
  assign n5029 = n169 & n5028 ;
  assign n5030 = n4648 & n67218 ;
  assign n5031 = n4918 & n5030 ;
  assign n5032 = n5029 | n5031 ;
  assign n5033 = n66560 & n5032 ;
  assign n67237 = ~n4869 ;
  assign n5034 = n4868 & n67237 ;
  assign n5035 = n4665 | n4868 ;
  assign n67238 = ~n5035 ;
  assign n5036 = n4967 & n67238 ;
  assign n5037 = n5034 | n5036 ;
  assign n5038 = n169 & n5037 ;
  assign n5039 = n4656 & n67218 ;
  assign n5040 = n4918 & n5039 ;
  assign n5041 = n5038 | n5040 ;
  assign n5042 = n66505 & n5041 ;
  assign n67239 = ~n4966 ;
  assign n5043 = n4864 & n67239 ;
  assign n5044 = n4673 | n4864 ;
  assign n67240 = ~n5044 ;
  assign n5045 = n4860 & n67240 ;
  assign n5046 = n5043 | n5045 ;
  assign n5047 = n169 & n5046 ;
  assign n5048 = n4664 & n67218 ;
  assign n5049 = n4918 & n5048 ;
  assign n5050 = n5047 | n5049 ;
  assign n5051 = n66379 & n5050 ;
  assign n67241 = ~n4859 ;
  assign n5052 = n4858 & n67241 ;
  assign n5053 = n4681 | n4858 ;
  assign n67242 = ~n5053 ;
  assign n5054 = n4963 & n67242 ;
  assign n5055 = n5052 | n5054 ;
  assign n5056 = n169 & n5055 ;
  assign n5057 = n4672 & n67218 ;
  assign n5058 = n4918 & n5057 ;
  assign n5059 = n5056 | n5058 ;
  assign n5060 = n66299 & n5059 ;
  assign n67243 = ~n4962 ;
  assign n5061 = n4854 & n67243 ;
  assign n5062 = n4689 | n4854 ;
  assign n67244 = ~n5062 ;
  assign n5063 = n4850 & n67244 ;
  assign n5064 = n5061 | n5063 ;
  assign n5065 = n169 & n5064 ;
  assign n5066 = n4680 & n67218 ;
  assign n5067 = n4918 & n5066 ;
  assign n5068 = n5065 | n5067 ;
  assign n5069 = n66244 & n5068 ;
  assign n67245 = ~n4849 ;
  assign n5070 = n4848 & n67245 ;
  assign n5071 = n4697 | n4848 ;
  assign n67246 = ~n5071 ;
  assign n5072 = n4959 & n67246 ;
  assign n5073 = n5070 | n5072 ;
  assign n5074 = n169 & n5073 ;
  assign n5075 = n4688 & n67218 ;
  assign n5076 = n4918 & n5075 ;
  assign n5077 = n5074 | n5076 ;
  assign n5078 = n66145 & n5077 ;
  assign n67247 = ~n4958 ;
  assign n5079 = n4844 & n67247 ;
  assign n5080 = n4705 | n4844 ;
  assign n67248 = ~n5080 ;
  assign n5081 = n4840 & n67248 ;
  assign n5082 = n5079 | n5081 ;
  assign n5083 = n169 & n5082 ;
  assign n5084 = n4696 & n67218 ;
  assign n5085 = n4918 & n5084 ;
  assign n5086 = n5083 | n5085 ;
  assign n5087 = n66081 & n5086 ;
  assign n67249 = ~n4839 ;
  assign n5088 = n4838 & n67249 ;
  assign n5089 = n4713 | n4838 ;
  assign n67250 = ~n5089 ;
  assign n5090 = n4955 & n67250 ;
  assign n5091 = n5088 | n5090 ;
  assign n5092 = n169 & n5091 ;
  assign n5093 = n4704 & n67218 ;
  assign n5094 = n4918 & n5093 ;
  assign n5095 = n5092 | n5094 ;
  assign n5096 = n66043 & n5095 ;
  assign n67251 = ~n4954 ;
  assign n5097 = n4834 & n67251 ;
  assign n5098 = n4721 | n4834 ;
  assign n67252 = ~n5098 ;
  assign n5099 = n4830 & n67252 ;
  assign n5100 = n5097 | n5099 ;
  assign n5101 = n169 & n5100 ;
  assign n5102 = n4712 & n67218 ;
  assign n5103 = n4918 & n5102 ;
  assign n5104 = n5101 | n5103 ;
  assign n5105 = n65960 & n5104 ;
  assign n67253 = ~n4829 ;
  assign n5106 = n4828 & n67253 ;
  assign n5107 = n4729 | n4828 ;
  assign n67254 = ~n5107 ;
  assign n5108 = n4951 & n67254 ;
  assign n5109 = n5106 | n5108 ;
  assign n5110 = n169 & n5109 ;
  assign n5111 = n4720 & n67218 ;
  assign n5112 = n4918 & n5111 ;
  assign n5113 = n5110 | n5112 ;
  assign n5114 = n65909 & n5113 ;
  assign n67255 = ~n4950 ;
  assign n5115 = n4824 & n67255 ;
  assign n5116 = n4737 | n4824 ;
  assign n67256 = ~n5116 ;
  assign n5117 = n4820 & n67256 ;
  assign n5118 = n5115 | n5117 ;
  assign n5119 = n169 & n5118 ;
  assign n5120 = n4728 & n67218 ;
  assign n5121 = n4918 & n5120 ;
  assign n5122 = n5119 | n5121 ;
  assign n5123 = n65877 & n5122 ;
  assign n67257 = ~n4819 ;
  assign n5124 = n4818 & n67257 ;
  assign n5125 = n4746 | n4818 ;
  assign n67258 = ~n5125 ;
  assign n5126 = n4947 & n67258 ;
  assign n5127 = n5124 | n5126 ;
  assign n5128 = n169 & n5127 ;
  assign n5129 = n4736 & n67218 ;
  assign n5130 = n4918 & n5129 ;
  assign n5131 = n5128 | n5130 ;
  assign n5132 = n65820 & n5131 ;
  assign n67259 = ~n4946 ;
  assign n5133 = n4814 & n67259 ;
  assign n5134 = n4754 | n4814 ;
  assign n67260 = ~n5134 ;
  assign n5135 = n4810 & n67260 ;
  assign n5136 = n5133 | n5135 ;
  assign n5137 = n169 & n5136 ;
  assign n5138 = n4745 & n67218 ;
  assign n5139 = n4918 & n5138 ;
  assign n5140 = n5137 | n5139 ;
  assign n5141 = n65791 & n5140 ;
  assign n67261 = ~n4809 ;
  assign n5142 = n4808 & n67261 ;
  assign n5143 = n4764 | n4808 ;
  assign n67262 = ~n5143 ;
  assign n5144 = n4943 & n67262 ;
  assign n5145 = n5142 | n5144 ;
  assign n5146 = n169 & n5145 ;
  assign n5147 = n4753 & n67218 ;
  assign n5148 = n4918 & n5147 ;
  assign n5149 = n5146 | n5148 ;
  assign n5150 = n65772 & n5149 ;
  assign n67263 = ~n4942 ;
  assign n5152 = n4804 & n67263 ;
  assign n5151 = n4772 | n4804 ;
  assign n67264 = ~n5151 ;
  assign n5153 = n4941 & n67264 ;
  assign n5154 = n5152 | n5153 ;
  assign n5155 = n169 & n5154 ;
  assign n5156 = n4762 & n67218 ;
  assign n5157 = n4918 & n5156 ;
  assign n5158 = n5155 | n5157 ;
  assign n5159 = n65746 & n5158 ;
  assign n67265 = ~n4800 ;
  assign n5160 = n4799 & n67265 ;
  assign n4940 = n4796 | n4799 ;
  assign n67266 = ~n4940 ;
  assign n5161 = n4795 & n67266 ;
  assign n5162 = n5160 | n5161 ;
  assign n5163 = n169 & n5162 ;
  assign n5164 = n4771 & n67218 ;
  assign n5165 = n4918 & n5164 ;
  assign n5166 = n5163 | n5165 ;
  assign n5167 = n65721 & n5166 ;
  assign n5168 = n4792 & n4794 ;
  assign n5169 = n67167 & n5168 ;
  assign n67267 = ~n5169 ;
  assign n5170 = n4795 & n67267 ;
  assign n5171 = n169 & n5170 ;
  assign n5172 = n4789 & n67218 ;
  assign n5173 = n4918 & n5172 ;
  assign n5174 = n5171 | n5173 ;
  assign n5175 = n65686 & n5174 ;
  assign n4921 = n4794 & n169 ;
  assign n5176 = x64 & n169 ;
  assign n67268 = ~n5176 ;
  assign n5177 = x40 & n67268 ;
  assign n5178 = n4921 | n5177 ;
  assign n5191 = n65670 & n5178 ;
  assign n4980 = n67209 & n4979 ;
  assign n5179 = n4899 | n4980 ;
  assign n5180 = n67210 & n5179 ;
  assign n5181 = n4917 | n5180 ;
  assign n5182 = n67218 & n5181 ;
  assign n67269 = ~n5182 ;
  assign n5183 = x64 & n67269 ;
  assign n67270 = ~n5183 ;
  assign n5184 = x40 & n67270 ;
  assign n5185 = n4921 | n5184 ;
  assign n5186 = x65 & n5185 ;
  assign n5187 = x65 | n4921 ;
  assign n5188 = n5184 | n5187 ;
  assign n67271 = ~n5186 ;
  assign n5189 = n67271 & n5188 ;
  assign n67272 = ~x39 ;
  assign n5190 = n67272 & x64 ;
  assign n5192 = n5189 | n5190 ;
  assign n67273 = ~n5191 ;
  assign n5193 = n67273 & n5192 ;
  assign n67274 = ~n5173 ;
  assign n5194 = x66 & n67274 ;
  assign n67275 = ~n5171 ;
  assign n5195 = n67275 & n5194 ;
  assign n5196 = n5175 | n5195 ;
  assign n5197 = n5193 | n5196 ;
  assign n67276 = ~n5175 ;
  assign n5198 = n67276 & n5197 ;
  assign n67277 = ~n5165 ;
  assign n5199 = x67 & n67277 ;
  assign n67278 = ~n5163 ;
  assign n5200 = n67278 & n5199 ;
  assign n5201 = n5167 | n5200 ;
  assign n5202 = n5198 | n5201 ;
  assign n67279 = ~n5167 ;
  assign n5203 = n67279 & n5202 ;
  assign n67280 = ~n5157 ;
  assign n5204 = x68 & n67280 ;
  assign n67281 = ~n5155 ;
  assign n5205 = n67281 & n5204 ;
  assign n5206 = n5159 | n5205 ;
  assign n5207 = n5203 | n5206 ;
  assign n67282 = ~n5159 ;
  assign n5208 = n67282 & n5207 ;
  assign n67283 = ~n5148 ;
  assign n5209 = x69 & n67283 ;
  assign n67284 = ~n5146 ;
  assign n5210 = n67284 & n5209 ;
  assign n5211 = n5150 | n5210 ;
  assign n5212 = n5208 | n5211 ;
  assign n67285 = ~n5150 ;
  assign n5213 = n67285 & n5212 ;
  assign n67286 = ~n5139 ;
  assign n5214 = x70 & n67286 ;
  assign n67287 = ~n5137 ;
  assign n5215 = n67287 & n5214 ;
  assign n5216 = n5141 | n5215 ;
  assign n5218 = n5213 | n5216 ;
  assign n67288 = ~n5141 ;
  assign n5219 = n67288 & n5218 ;
  assign n67289 = ~n5130 ;
  assign n5220 = x71 & n67289 ;
  assign n67290 = ~n5128 ;
  assign n5221 = n67290 & n5220 ;
  assign n5222 = n5132 | n5221 ;
  assign n5223 = n5219 | n5222 ;
  assign n67291 = ~n5132 ;
  assign n5224 = n67291 & n5223 ;
  assign n67292 = ~n5121 ;
  assign n5225 = x72 & n67292 ;
  assign n67293 = ~n5119 ;
  assign n5226 = n67293 & n5225 ;
  assign n5227 = n5123 | n5226 ;
  assign n5229 = n5224 | n5227 ;
  assign n67294 = ~n5123 ;
  assign n5230 = n67294 & n5229 ;
  assign n67295 = ~n5112 ;
  assign n5231 = x73 & n67295 ;
  assign n67296 = ~n5110 ;
  assign n5232 = n67296 & n5231 ;
  assign n5233 = n5114 | n5232 ;
  assign n5234 = n5230 | n5233 ;
  assign n67297 = ~n5114 ;
  assign n5235 = n67297 & n5234 ;
  assign n67298 = ~n5103 ;
  assign n5236 = x74 & n67298 ;
  assign n67299 = ~n5101 ;
  assign n5237 = n67299 & n5236 ;
  assign n5238 = n5105 | n5237 ;
  assign n5240 = n5235 | n5238 ;
  assign n67300 = ~n5105 ;
  assign n5241 = n67300 & n5240 ;
  assign n67301 = ~n5094 ;
  assign n5242 = x75 & n67301 ;
  assign n67302 = ~n5092 ;
  assign n5243 = n67302 & n5242 ;
  assign n5244 = n5096 | n5243 ;
  assign n5245 = n5241 | n5244 ;
  assign n67303 = ~n5096 ;
  assign n5246 = n67303 & n5245 ;
  assign n67304 = ~n5085 ;
  assign n5247 = x76 & n67304 ;
  assign n67305 = ~n5083 ;
  assign n5248 = n67305 & n5247 ;
  assign n5249 = n5087 | n5248 ;
  assign n5251 = n5246 | n5249 ;
  assign n67306 = ~n5087 ;
  assign n5252 = n67306 & n5251 ;
  assign n67307 = ~n5076 ;
  assign n5253 = x77 & n67307 ;
  assign n67308 = ~n5074 ;
  assign n5254 = n67308 & n5253 ;
  assign n5255 = n5078 | n5254 ;
  assign n5256 = n5252 | n5255 ;
  assign n67309 = ~n5078 ;
  assign n5257 = n67309 & n5256 ;
  assign n67310 = ~n5067 ;
  assign n5258 = x78 & n67310 ;
  assign n67311 = ~n5065 ;
  assign n5259 = n67311 & n5258 ;
  assign n5260 = n5069 | n5259 ;
  assign n5262 = n5257 | n5260 ;
  assign n67312 = ~n5069 ;
  assign n5263 = n67312 & n5262 ;
  assign n67313 = ~n5058 ;
  assign n5264 = x79 & n67313 ;
  assign n67314 = ~n5056 ;
  assign n5265 = n67314 & n5264 ;
  assign n5266 = n5060 | n5265 ;
  assign n5267 = n5263 | n5266 ;
  assign n67315 = ~n5060 ;
  assign n5268 = n67315 & n5267 ;
  assign n67316 = ~n5049 ;
  assign n5269 = x80 & n67316 ;
  assign n67317 = ~n5047 ;
  assign n5270 = n67317 & n5269 ;
  assign n5271 = n5051 | n5270 ;
  assign n5273 = n5268 | n5271 ;
  assign n67318 = ~n5051 ;
  assign n5274 = n67318 & n5273 ;
  assign n67319 = ~n5040 ;
  assign n5275 = x81 & n67319 ;
  assign n67320 = ~n5038 ;
  assign n5276 = n67320 & n5275 ;
  assign n5277 = n5042 | n5276 ;
  assign n5278 = n5274 | n5277 ;
  assign n67321 = ~n5042 ;
  assign n5279 = n67321 & n5278 ;
  assign n67322 = ~n5031 ;
  assign n5280 = x82 & n67322 ;
  assign n67323 = ~n5029 ;
  assign n5281 = n67323 & n5280 ;
  assign n5282 = n5033 | n5281 ;
  assign n5284 = n5279 | n5282 ;
  assign n67324 = ~n5033 ;
  assign n5285 = n67324 & n5284 ;
  assign n67325 = ~n5022 ;
  assign n5286 = x83 & n67325 ;
  assign n67326 = ~n5020 ;
  assign n5287 = n67326 & n5286 ;
  assign n5288 = n5024 | n5287 ;
  assign n5289 = n5285 | n5288 ;
  assign n67327 = ~n5024 ;
  assign n5290 = n67327 & n5289 ;
  assign n67328 = ~n5013 ;
  assign n5291 = x84 & n67328 ;
  assign n67329 = ~n5011 ;
  assign n5292 = n67329 & n5291 ;
  assign n5293 = n5015 | n5292 ;
  assign n5295 = n5290 | n5293 ;
  assign n67330 = ~n5015 ;
  assign n5296 = n67330 & n5295 ;
  assign n67331 = ~n5004 ;
  assign n5297 = x85 & n67331 ;
  assign n67332 = ~n5002 ;
  assign n5298 = n67332 & n5297 ;
  assign n5299 = n5006 | n5298 ;
  assign n5300 = n5296 | n5299 ;
  assign n67333 = ~n5006 ;
  assign n5301 = n67333 & n5300 ;
  assign n67334 = ~n4995 ;
  assign n5302 = x86 & n67334 ;
  assign n67335 = ~n4993 ;
  assign n5303 = n67335 & n5302 ;
  assign n5304 = n4997 | n5303 ;
  assign n5306 = n5301 | n5304 ;
  assign n67336 = ~n4997 ;
  assign n5307 = n67336 & n5306 ;
  assign n67337 = ~n4987 ;
  assign n5308 = x87 & n67337 ;
  assign n67338 = ~n4985 ;
  assign n5309 = n67338 & n5308 ;
  assign n5310 = n4989 | n5309 ;
  assign n5311 = n5307 | n5310 ;
  assign n67339 = ~n4989 ;
  assign n5312 = n67339 & n5311 ;
  assign n67340 = ~n4930 ;
  assign n5313 = x88 & n67340 ;
  assign n67341 = ~n4928 ;
  assign n5314 = n67341 & n5313 ;
  assign n5315 = n4932 | n5314 ;
  assign n5317 = n5312 | n5315 ;
  assign n67342 = ~n4932 ;
  assign n5318 = n67342 & n5317 ;
  assign n5319 = n74914 | n294 ;
  assign n5320 = n279 | n5319 ;
  assign n5321 = n5318 | n5320 ;
  assign n67343 = ~n5312 ;
  assign n5316 = n67343 & n5315 ;
  assign n5322 = x65 & n5178 ;
  assign n67344 = ~n5322 ;
  assign n5323 = n5188 & n67344 ;
  assign n5324 = n5190 | n5323 ;
  assign n5325 = n67273 & n5324 ;
  assign n5326 = n5196 | n5325 ;
  assign n5327 = n67276 & n5326 ;
  assign n5329 = n5201 | n5327 ;
  assign n5330 = n67279 & n5329 ;
  assign n5332 = n5206 | n5330 ;
  assign n5333 = n67282 & n5332 ;
  assign n5334 = n5211 | n5333 ;
  assign n5336 = n67285 & n5334 ;
  assign n5337 = n5216 | n5336 ;
  assign n5338 = n67288 & n5337 ;
  assign n5339 = n5222 | n5338 ;
  assign n5341 = n67291 & n5339 ;
  assign n5342 = n5227 | n5341 ;
  assign n5343 = n67294 & n5342 ;
  assign n5344 = n5233 | n5343 ;
  assign n5346 = n67297 & n5344 ;
  assign n5347 = n5238 | n5346 ;
  assign n5348 = n67300 & n5347 ;
  assign n5349 = n5244 | n5348 ;
  assign n5351 = n67303 & n5349 ;
  assign n5352 = n5249 | n5351 ;
  assign n5353 = n67306 & n5352 ;
  assign n5354 = n5255 | n5353 ;
  assign n5356 = n67309 & n5354 ;
  assign n5357 = n5260 | n5356 ;
  assign n5358 = n67312 & n5357 ;
  assign n5359 = n5266 | n5358 ;
  assign n5361 = n67315 & n5359 ;
  assign n5362 = n5271 | n5361 ;
  assign n5363 = n67318 & n5362 ;
  assign n5364 = n5277 | n5363 ;
  assign n5366 = n67321 & n5364 ;
  assign n5367 = n5282 | n5366 ;
  assign n5368 = n67324 & n5367 ;
  assign n5369 = n5288 | n5368 ;
  assign n5371 = n67327 & n5369 ;
  assign n5372 = n5293 | n5371 ;
  assign n5373 = n67330 & n5372 ;
  assign n5374 = n5299 | n5373 ;
  assign n5376 = n67333 & n5374 ;
  assign n5377 = n5304 | n5376 ;
  assign n5378 = n67336 & n5377 ;
  assign n5380 = n5310 | n5378 ;
  assign n5381 = n4989 | n5315 ;
  assign n67345 = ~n5381 ;
  assign n5382 = n5380 & n67345 ;
  assign n5383 = n5316 | n5382 ;
  assign n5384 = n5321 | n5383 ;
  assign n67346 = ~n4931 ;
  assign n5385 = n67346 & n5321 ;
  assign n67347 = ~n5385 ;
  assign n5386 = n5384 & n67347 ;
  assign n67348 = ~x89 ;
  assign n5387 = n67348 & n5386 ;
  assign n168 = ~n5321 ;
  assign n5733 = n168 & n5383 ;
  assign n5734 = n4931 & n5321 ;
  assign n67350 = ~n5734 ;
  assign n5735 = x89 & n67350 ;
  assign n67351 = ~n5733 ;
  assign n5736 = n67351 & n5735 ;
  assign n5737 = n5387 | n5736 ;
  assign n5388 = n4988 & n5321 ;
  assign n67352 = ~n5378 ;
  assign n5379 = n5310 & n67352 ;
  assign n5389 = n4997 | n5310 ;
  assign n67353 = ~n5389 ;
  assign n5390 = n5306 & n67353 ;
  assign n5391 = n5379 | n5390 ;
  assign n67354 = ~n5320 ;
  assign n5392 = n67354 & n5391 ;
  assign n67355 = ~n5318 ;
  assign n5393 = n67355 & n5392 ;
  assign n5394 = n5388 | n5393 ;
  assign n5395 = n67222 & n5394 ;
  assign n5396 = n4996 & n5321 ;
  assign n67356 = ~n5301 ;
  assign n5305 = n67356 & n5304 ;
  assign n5397 = n5006 | n5304 ;
  assign n67357 = ~n5397 ;
  assign n5398 = n5374 & n67357 ;
  assign n5399 = n5305 | n5398 ;
  assign n5400 = n67354 & n5399 ;
  assign n5401 = n67355 & n5400 ;
  assign n5402 = n5396 | n5401 ;
  assign n5403 = n67164 & n5402 ;
  assign n67358 = ~n5401 ;
  assign n5721 = x87 & n67358 ;
  assign n67359 = ~n5396 ;
  assign n5722 = n67359 & n5721 ;
  assign n5723 = n5403 | n5722 ;
  assign n5404 = n5005 & n5321 ;
  assign n67360 = ~n5373 ;
  assign n5375 = n5299 & n67360 ;
  assign n5405 = n5015 | n5299 ;
  assign n67361 = ~n5405 ;
  assign n5406 = n5295 & n67361 ;
  assign n5407 = n5375 | n5406 ;
  assign n5408 = n67354 & n5407 ;
  assign n5409 = n67355 & n5408 ;
  assign n5410 = n5404 | n5409 ;
  assign n5411 = n66979 & n5410 ;
  assign n5412 = n5014 & n5321 ;
  assign n67362 = ~n5290 ;
  assign n5294 = n67362 & n5293 ;
  assign n5413 = n5024 | n5293 ;
  assign n67363 = ~n5413 ;
  assign n5414 = n5369 & n67363 ;
  assign n5415 = n5294 | n5414 ;
  assign n5416 = n67354 & n5415 ;
  assign n5417 = n67355 & n5416 ;
  assign n5418 = n5412 | n5417 ;
  assign n5419 = n66868 & n5418 ;
  assign n67364 = ~n5417 ;
  assign n5709 = x85 & n67364 ;
  assign n67365 = ~n5412 ;
  assign n5710 = n67365 & n5709 ;
  assign n5711 = n5419 | n5710 ;
  assign n5420 = n5023 & n5321 ;
  assign n67366 = ~n5368 ;
  assign n5370 = n5288 & n67366 ;
  assign n5421 = n5033 | n5288 ;
  assign n67367 = ~n5421 ;
  assign n5422 = n5284 & n67367 ;
  assign n5423 = n5370 | n5422 ;
  assign n5424 = n67354 & n5423 ;
  assign n5425 = n67355 & n5424 ;
  assign n5426 = n5420 | n5425 ;
  assign n5427 = n66797 & n5426 ;
  assign n5428 = n5032 & n5321 ;
  assign n67368 = ~n5279 ;
  assign n5283 = n67368 & n5282 ;
  assign n5429 = n5042 | n5282 ;
  assign n67369 = ~n5429 ;
  assign n5430 = n5364 & n67369 ;
  assign n5431 = n5283 | n5430 ;
  assign n5432 = n67354 & n5431 ;
  assign n5433 = n67355 & n5432 ;
  assign n5434 = n5428 | n5433 ;
  assign n5435 = n66654 & n5434 ;
  assign n67370 = ~n5433 ;
  assign n5697 = x83 & n67370 ;
  assign n67371 = ~n5428 ;
  assign n5698 = n67371 & n5697 ;
  assign n5699 = n5435 | n5698 ;
  assign n5436 = n5041 & n5321 ;
  assign n67372 = ~n5363 ;
  assign n5365 = n5277 & n67372 ;
  assign n5437 = n5051 | n5277 ;
  assign n67373 = ~n5437 ;
  assign n5438 = n5273 & n67373 ;
  assign n5439 = n5365 | n5438 ;
  assign n5440 = n67354 & n5439 ;
  assign n5441 = n67355 & n5440 ;
  assign n5442 = n5436 | n5441 ;
  assign n5443 = n66560 & n5442 ;
  assign n5444 = n5050 & n5321 ;
  assign n67374 = ~n5268 ;
  assign n5272 = n67374 & n5271 ;
  assign n5445 = n5060 | n5271 ;
  assign n67375 = ~n5445 ;
  assign n5446 = n5359 & n67375 ;
  assign n5447 = n5272 | n5446 ;
  assign n5448 = n67354 & n5447 ;
  assign n5449 = n67355 & n5448 ;
  assign n5450 = n5444 | n5449 ;
  assign n5451 = n66505 & n5450 ;
  assign n67376 = ~n5449 ;
  assign n5685 = x81 & n67376 ;
  assign n67377 = ~n5444 ;
  assign n5686 = n67377 & n5685 ;
  assign n5687 = n5451 | n5686 ;
  assign n5452 = n5059 & n5321 ;
  assign n67378 = ~n5358 ;
  assign n5360 = n5266 & n67378 ;
  assign n5453 = n5069 | n5266 ;
  assign n67379 = ~n5453 ;
  assign n5454 = n5262 & n67379 ;
  assign n5455 = n5360 | n5454 ;
  assign n5456 = n67354 & n5455 ;
  assign n5457 = n67355 & n5456 ;
  assign n5458 = n5452 | n5457 ;
  assign n5459 = n66379 & n5458 ;
  assign n5460 = n5068 & n5321 ;
  assign n67380 = ~n5257 ;
  assign n5261 = n67380 & n5260 ;
  assign n5461 = n5078 | n5260 ;
  assign n67381 = ~n5461 ;
  assign n5462 = n5354 & n67381 ;
  assign n5463 = n5261 | n5462 ;
  assign n5464 = n67354 & n5463 ;
  assign n5465 = n67355 & n5464 ;
  assign n5466 = n5460 | n5465 ;
  assign n5467 = n66299 & n5466 ;
  assign n67382 = ~n5465 ;
  assign n5673 = x79 & n67382 ;
  assign n67383 = ~n5460 ;
  assign n5674 = n67383 & n5673 ;
  assign n5675 = n5467 | n5674 ;
  assign n5468 = n5077 & n5321 ;
  assign n67384 = ~n5353 ;
  assign n5355 = n5255 & n67384 ;
  assign n5469 = n5087 | n5255 ;
  assign n67385 = ~n5469 ;
  assign n5470 = n5251 & n67385 ;
  assign n5471 = n5355 | n5470 ;
  assign n5472 = n67354 & n5471 ;
  assign n5473 = n67355 & n5472 ;
  assign n5474 = n5468 | n5473 ;
  assign n5475 = n66244 & n5474 ;
  assign n5476 = n5086 & n5321 ;
  assign n67386 = ~n5246 ;
  assign n5250 = n67386 & n5249 ;
  assign n5477 = n5096 | n5249 ;
  assign n67387 = ~n5477 ;
  assign n5478 = n5349 & n67387 ;
  assign n5479 = n5250 | n5478 ;
  assign n5480 = n67354 & n5479 ;
  assign n5481 = n67355 & n5480 ;
  assign n5482 = n5476 | n5481 ;
  assign n5483 = n66145 & n5482 ;
  assign n67388 = ~n5481 ;
  assign n5661 = x77 & n67388 ;
  assign n67389 = ~n5476 ;
  assign n5662 = n67389 & n5661 ;
  assign n5663 = n5483 | n5662 ;
  assign n5484 = n5095 & n5321 ;
  assign n67390 = ~n5348 ;
  assign n5350 = n5244 & n67390 ;
  assign n5485 = n5105 | n5244 ;
  assign n67391 = ~n5485 ;
  assign n5486 = n5240 & n67391 ;
  assign n5487 = n5350 | n5486 ;
  assign n5488 = n67354 & n5487 ;
  assign n5489 = n67355 & n5488 ;
  assign n5490 = n5484 | n5489 ;
  assign n5491 = n66081 & n5490 ;
  assign n5492 = n5104 & n5321 ;
  assign n67392 = ~n5235 ;
  assign n5239 = n67392 & n5238 ;
  assign n5493 = n5114 | n5238 ;
  assign n67393 = ~n5493 ;
  assign n5494 = n5344 & n67393 ;
  assign n5495 = n5239 | n5494 ;
  assign n5496 = n67354 & n5495 ;
  assign n5497 = n67355 & n5496 ;
  assign n5498 = n5492 | n5497 ;
  assign n5499 = n66043 & n5498 ;
  assign n67394 = ~n5497 ;
  assign n5649 = x75 & n67394 ;
  assign n67395 = ~n5492 ;
  assign n5650 = n67395 & n5649 ;
  assign n5651 = n5499 | n5650 ;
  assign n5500 = n5113 & n5321 ;
  assign n67396 = ~n5343 ;
  assign n5345 = n5233 & n67396 ;
  assign n5501 = n5123 | n5233 ;
  assign n67397 = ~n5501 ;
  assign n5502 = n5229 & n67397 ;
  assign n5503 = n5345 | n5502 ;
  assign n5504 = n67354 & n5503 ;
  assign n5505 = n67355 & n5504 ;
  assign n5506 = n5500 | n5505 ;
  assign n5507 = n65960 & n5506 ;
  assign n5508 = n5122 & n5321 ;
  assign n67398 = ~n5224 ;
  assign n5228 = n67398 & n5227 ;
  assign n5509 = n5132 | n5227 ;
  assign n67399 = ~n5509 ;
  assign n5510 = n5339 & n67399 ;
  assign n5511 = n5228 | n5510 ;
  assign n5512 = n67354 & n5511 ;
  assign n5513 = n67355 & n5512 ;
  assign n5514 = n5508 | n5513 ;
  assign n5515 = n65909 & n5514 ;
  assign n67400 = ~n5513 ;
  assign n5637 = x73 & n67400 ;
  assign n67401 = ~n5508 ;
  assign n5638 = n67401 & n5637 ;
  assign n5639 = n5515 | n5638 ;
  assign n5516 = n5131 & n5321 ;
  assign n67402 = ~n5338 ;
  assign n5340 = n5222 & n67402 ;
  assign n5517 = n5141 | n5222 ;
  assign n67403 = ~n5517 ;
  assign n5518 = n5218 & n67403 ;
  assign n5519 = n5340 | n5518 ;
  assign n5520 = n67354 & n5519 ;
  assign n5521 = n67355 & n5520 ;
  assign n5522 = n5516 | n5521 ;
  assign n5523 = n65877 & n5522 ;
  assign n5524 = n5140 & n5321 ;
  assign n67404 = ~n5213 ;
  assign n5217 = n67404 & n5216 ;
  assign n5525 = n5150 | n5216 ;
  assign n67405 = ~n5525 ;
  assign n5526 = n5334 & n67405 ;
  assign n5527 = n5217 | n5526 ;
  assign n5528 = n67354 & n5527 ;
  assign n5529 = n67355 & n5528 ;
  assign n5530 = n5524 | n5529 ;
  assign n5531 = n65820 & n5530 ;
  assign n67406 = ~n5529 ;
  assign n5625 = x71 & n67406 ;
  assign n67407 = ~n5524 ;
  assign n5626 = n67407 & n5625 ;
  assign n5627 = n5531 | n5626 ;
  assign n5532 = n5149 & n5321 ;
  assign n67408 = ~n5333 ;
  assign n5335 = n5211 & n67408 ;
  assign n5533 = n5159 | n5211 ;
  assign n67409 = ~n5533 ;
  assign n5534 = n5207 & n67409 ;
  assign n5535 = n5335 | n5534 ;
  assign n5536 = n67354 & n5535 ;
  assign n5537 = n67355 & n5536 ;
  assign n5538 = n5532 | n5537 ;
  assign n5539 = n65791 & n5538 ;
  assign n5540 = n5158 & n5321 ;
  assign n67410 = ~n5203 ;
  assign n5331 = n67410 & n5206 ;
  assign n5541 = n5167 | n5206 ;
  assign n67411 = ~n5541 ;
  assign n5542 = n5329 & n67411 ;
  assign n5543 = n5331 | n5542 ;
  assign n5544 = n67354 & n5543 ;
  assign n5545 = n67355 & n5544 ;
  assign n5546 = n5540 | n5545 ;
  assign n5547 = n65772 & n5546 ;
  assign n67412 = ~n5545 ;
  assign n5614 = x69 & n67412 ;
  assign n67413 = ~n5540 ;
  assign n5615 = n67413 & n5614 ;
  assign n5616 = n5547 | n5615 ;
  assign n5548 = n5166 & n5321 ;
  assign n67414 = ~n5327 ;
  assign n5328 = n5201 & n67414 ;
  assign n5549 = n5175 | n5201 ;
  assign n67415 = ~n5549 ;
  assign n5550 = n5326 & n67415 ;
  assign n5551 = n5328 | n5550 ;
  assign n5552 = n67354 & n5551 ;
  assign n5553 = n67355 & n5552 ;
  assign n5554 = n5548 | n5553 ;
  assign n5555 = n65746 & n5554 ;
  assign n5556 = n5174 & n5321 ;
  assign n5557 = n5191 | n5196 ;
  assign n67416 = ~n5557 ;
  assign n5558 = n5324 & n67416 ;
  assign n67417 = ~n5193 ;
  assign n5559 = n67417 & n5196 ;
  assign n5560 = n5558 | n5559 ;
  assign n5561 = n67354 & n5560 ;
  assign n5562 = n67355 & n5561 ;
  assign n5563 = n5556 | n5562 ;
  assign n5564 = n65721 & n5563 ;
  assign n67418 = ~n5562 ;
  assign n5604 = x67 & n67418 ;
  assign n67419 = ~n5556 ;
  assign n5605 = n67419 & n5604 ;
  assign n5606 = n5564 | n5605 ;
  assign n5565 = n5185 & n5321 ;
  assign n5566 = n5188 & n5190 ;
  assign n5567 = n67344 & n5566 ;
  assign n5568 = n5320 | n5567 ;
  assign n67420 = ~n5568 ;
  assign n5569 = n5324 & n67420 ;
  assign n5570 = n67355 & n5569 ;
  assign n5571 = n5565 | n5570 ;
  assign n5572 = n65686 & n5571 ;
  assign n67421 = ~x38 ;
  assign n5594 = n67421 & x64 ;
  assign n5573 = x64 & n67348 ;
  assign n67422 = ~n65557 ;
  assign n5574 = n67422 & n5573 ;
  assign n67423 = ~n65639 ;
  assign n5575 = n67423 & n5574 ;
  assign n5576 = n66509 & n5575 ;
  assign n5577 = n66510 & n5576 ;
  assign n5578 = n67355 & n5577 ;
  assign n67424 = ~n5578 ;
  assign n5579 = x39 & n67424 ;
  assign n5580 = n67023 & n5190 ;
  assign n5581 = n67024 & n5580 ;
  assign n5582 = n67025 & n5581 ;
  assign n5583 = n67026 & n5582 ;
  assign n5584 = n67355 & n5583 ;
  assign n5585 = n5579 | n5584 ;
  assign n5586 = x65 & n5585 ;
  assign n5587 = n67339 & n5380 ;
  assign n5588 = n5315 | n5587 ;
  assign n5589 = n67342 & n5588 ;
  assign n67425 = ~n5589 ;
  assign n5590 = n5577 & n67425 ;
  assign n67426 = ~n5590 ;
  assign n5591 = x39 & n67426 ;
  assign n5592 = x65 | n5584 ;
  assign n5593 = n5591 | n5592 ;
  assign n67427 = ~n5586 ;
  assign n5595 = n67427 & n5593 ;
  assign n5596 = n5594 | n5595 ;
  assign n5597 = n5584 | n5591 ;
  assign n5598 = n65670 & n5597 ;
  assign n67428 = ~n5598 ;
  assign n5599 = n5596 & n67428 ;
  assign n67429 = ~n5570 ;
  assign n5600 = x66 & n67429 ;
  assign n67430 = ~n5565 ;
  assign n5601 = n67430 & n5600 ;
  assign n5602 = n5572 | n5601 ;
  assign n5603 = n5599 | n5602 ;
  assign n67431 = ~n5572 ;
  assign n5607 = n67431 & n5603 ;
  assign n5608 = n5606 | n5607 ;
  assign n67432 = ~n5564 ;
  assign n5609 = n67432 & n5608 ;
  assign n67433 = ~n5553 ;
  assign n5610 = x68 & n67433 ;
  assign n67434 = ~n5548 ;
  assign n5611 = n67434 & n5610 ;
  assign n5612 = n5555 | n5611 ;
  assign n5613 = n5609 | n5612 ;
  assign n67435 = ~n5555 ;
  assign n5617 = n67435 & n5613 ;
  assign n5618 = n5616 | n5617 ;
  assign n67436 = ~n5547 ;
  assign n5619 = n67436 & n5618 ;
  assign n67437 = ~n5537 ;
  assign n5620 = x70 & n67437 ;
  assign n67438 = ~n5532 ;
  assign n5621 = n67438 & n5620 ;
  assign n5622 = n5539 | n5621 ;
  assign n5624 = n5619 | n5622 ;
  assign n67439 = ~n5539 ;
  assign n5629 = n67439 & n5624 ;
  assign n5630 = n5627 | n5629 ;
  assign n67440 = ~n5531 ;
  assign n5631 = n67440 & n5630 ;
  assign n67441 = ~n5521 ;
  assign n5632 = x72 & n67441 ;
  assign n67442 = ~n5516 ;
  assign n5633 = n67442 & n5632 ;
  assign n5634 = n5523 | n5633 ;
  assign n5636 = n5631 | n5634 ;
  assign n67443 = ~n5523 ;
  assign n5641 = n67443 & n5636 ;
  assign n5642 = n5639 | n5641 ;
  assign n67444 = ~n5515 ;
  assign n5643 = n67444 & n5642 ;
  assign n67445 = ~n5505 ;
  assign n5644 = x74 & n67445 ;
  assign n67446 = ~n5500 ;
  assign n5645 = n67446 & n5644 ;
  assign n5646 = n5507 | n5645 ;
  assign n5648 = n5643 | n5646 ;
  assign n67447 = ~n5507 ;
  assign n5653 = n67447 & n5648 ;
  assign n5654 = n5651 | n5653 ;
  assign n67448 = ~n5499 ;
  assign n5655 = n67448 & n5654 ;
  assign n67449 = ~n5489 ;
  assign n5656 = x76 & n67449 ;
  assign n67450 = ~n5484 ;
  assign n5657 = n67450 & n5656 ;
  assign n5658 = n5491 | n5657 ;
  assign n5660 = n5655 | n5658 ;
  assign n67451 = ~n5491 ;
  assign n5665 = n67451 & n5660 ;
  assign n5666 = n5663 | n5665 ;
  assign n67452 = ~n5483 ;
  assign n5667 = n67452 & n5666 ;
  assign n67453 = ~n5473 ;
  assign n5668 = x78 & n67453 ;
  assign n67454 = ~n5468 ;
  assign n5669 = n67454 & n5668 ;
  assign n5670 = n5475 | n5669 ;
  assign n5672 = n5667 | n5670 ;
  assign n67455 = ~n5475 ;
  assign n5677 = n67455 & n5672 ;
  assign n5678 = n5675 | n5677 ;
  assign n67456 = ~n5467 ;
  assign n5679 = n67456 & n5678 ;
  assign n67457 = ~n5457 ;
  assign n5680 = x80 & n67457 ;
  assign n67458 = ~n5452 ;
  assign n5681 = n67458 & n5680 ;
  assign n5682 = n5459 | n5681 ;
  assign n5684 = n5679 | n5682 ;
  assign n67459 = ~n5459 ;
  assign n5689 = n67459 & n5684 ;
  assign n5690 = n5687 | n5689 ;
  assign n67460 = ~n5451 ;
  assign n5691 = n67460 & n5690 ;
  assign n67461 = ~n5441 ;
  assign n5692 = x82 & n67461 ;
  assign n67462 = ~n5436 ;
  assign n5693 = n67462 & n5692 ;
  assign n5694 = n5443 | n5693 ;
  assign n5696 = n5691 | n5694 ;
  assign n67463 = ~n5443 ;
  assign n5701 = n67463 & n5696 ;
  assign n5702 = n5699 | n5701 ;
  assign n67464 = ~n5435 ;
  assign n5703 = n67464 & n5702 ;
  assign n67465 = ~n5425 ;
  assign n5704 = x84 & n67465 ;
  assign n67466 = ~n5420 ;
  assign n5705 = n67466 & n5704 ;
  assign n5706 = n5427 | n5705 ;
  assign n5708 = n5703 | n5706 ;
  assign n67467 = ~n5427 ;
  assign n5713 = n67467 & n5708 ;
  assign n5714 = n5711 | n5713 ;
  assign n67468 = ~n5419 ;
  assign n5715 = n67468 & n5714 ;
  assign n67469 = ~n5409 ;
  assign n5716 = x86 & n67469 ;
  assign n67470 = ~n5404 ;
  assign n5717 = n67470 & n5716 ;
  assign n5718 = n5411 | n5717 ;
  assign n5720 = n5715 | n5718 ;
  assign n67471 = ~n5411 ;
  assign n5725 = n67471 & n5720 ;
  assign n5726 = n5723 | n5725 ;
  assign n67472 = ~n5403 ;
  assign n5727 = n67472 & n5726 ;
  assign n67473 = ~n5393 ;
  assign n5728 = x88 & n67473 ;
  assign n67474 = ~n5388 ;
  assign n5729 = n67474 & n5728 ;
  assign n5730 = n5395 | n5729 ;
  assign n5732 = n5727 | n5730 ;
  assign n67475 = ~n5395 ;
  assign n5738 = n67475 & n5732 ;
  assign n5739 = n5737 | n5738 ;
  assign n67476 = ~n5387 ;
  assign n5740 = n67476 & n5739 ;
  assign n5744 = n5740 | n5743 ;
  assign n67477 = ~n5386 ;
  assign n5746 = n67477 & n5744 ;
  assign n67478 = ~n5738 ;
  assign n6146 = n5737 & n67478 ;
  assign n5748 = x65 & n5597 ;
  assign n67479 = ~n5748 ;
  assign n5749 = n5593 & n67479 ;
  assign n5751 = n5594 | n5749 ;
  assign n5752 = n67428 & n5751 ;
  assign n5753 = n5602 | n5752 ;
  assign n5754 = n67431 & n5753 ;
  assign n5755 = n5606 | n5754 ;
  assign n5756 = n67432 & n5755 ;
  assign n5757 = n5612 | n5756 ;
  assign n5758 = n67435 & n5757 ;
  assign n5759 = n5616 | n5758 ;
  assign n5760 = n67436 & n5759 ;
  assign n5761 = n5622 | n5760 ;
  assign n5762 = n67439 & n5761 ;
  assign n5763 = n5627 | n5762 ;
  assign n5764 = n67440 & n5763 ;
  assign n5765 = n5634 | n5764 ;
  assign n5766 = n67443 & n5765 ;
  assign n5767 = n5639 | n5766 ;
  assign n5768 = n67444 & n5767 ;
  assign n5769 = n5646 | n5768 ;
  assign n5770 = n67447 & n5769 ;
  assign n5771 = n5651 | n5770 ;
  assign n5772 = n67448 & n5771 ;
  assign n5773 = n5658 | n5772 ;
  assign n5774 = n67451 & n5773 ;
  assign n5775 = n5663 | n5774 ;
  assign n5776 = n67452 & n5775 ;
  assign n5777 = n5670 | n5776 ;
  assign n5778 = n67455 & n5777 ;
  assign n5779 = n5675 | n5778 ;
  assign n5780 = n67456 & n5779 ;
  assign n5781 = n5682 | n5780 ;
  assign n5782 = n67459 & n5781 ;
  assign n5783 = n5687 | n5782 ;
  assign n5784 = n67460 & n5783 ;
  assign n5785 = n5694 | n5784 ;
  assign n5786 = n67463 & n5785 ;
  assign n5787 = n5699 | n5786 ;
  assign n5788 = n67464 & n5787 ;
  assign n5789 = n5706 | n5788 ;
  assign n5790 = n67467 & n5789 ;
  assign n5791 = n5711 | n5790 ;
  assign n5792 = n67468 & n5791 ;
  assign n5793 = n5718 | n5792 ;
  assign n5794 = n67471 & n5793 ;
  assign n5795 = n5723 | n5794 ;
  assign n5797 = n67472 & n5795 ;
  assign n5997 = n5730 | n5797 ;
  assign n6147 = n5395 | n5737 ;
  assign n67480 = ~n6147 ;
  assign n6148 = n5997 & n67480 ;
  assign n6149 = n6146 | n6148 ;
  assign n6150 = n5744 | n6149 ;
  assign n67481 = ~n5746 ;
  assign n6151 = n67481 & n6150 ;
  assign n67482 = ~n5743 ;
  assign n6162 = n67482 & n6151 ;
  assign n5747 = n5394 & n5744 ;
  assign n5731 = n5403 | n5730 ;
  assign n67483 = ~n5731 ;
  assign n5796 = n67483 & n5795 ;
  assign n67484 = ~n5797 ;
  assign n5798 = n5730 & n67484 ;
  assign n5799 = n5796 | n5798 ;
  assign n5800 = n67482 & n5799 ;
  assign n67485 = ~n5740 ;
  assign n5801 = n67485 & n5800 ;
  assign n5802 = n5747 | n5801 ;
  assign n5803 = n67348 & n5802 ;
  assign n5804 = n5402 & n5744 ;
  assign n5724 = n5411 | n5723 ;
  assign n67486 = ~n5724 ;
  assign n5805 = n5720 & n67486 ;
  assign n67487 = ~n5725 ;
  assign n5806 = n5723 & n67487 ;
  assign n5807 = n5805 | n5806 ;
  assign n5808 = n67482 & n5807 ;
  assign n5809 = n67485 & n5808 ;
  assign n5810 = n5804 | n5809 ;
  assign n5811 = n67222 & n5810 ;
  assign n5812 = n5410 & n5744 ;
  assign n5719 = n5419 | n5718 ;
  assign n67488 = ~n5719 ;
  assign n5813 = n67488 & n5791 ;
  assign n67489 = ~n5792 ;
  assign n5814 = n5718 & n67489 ;
  assign n5815 = n5813 | n5814 ;
  assign n5816 = n67482 & n5815 ;
  assign n5817 = n67485 & n5816 ;
  assign n5818 = n5812 | n5817 ;
  assign n5819 = n67164 & n5818 ;
  assign n5820 = n5418 & n5744 ;
  assign n5712 = n5427 | n5711 ;
  assign n67490 = ~n5712 ;
  assign n5821 = n5708 & n67490 ;
  assign n67491 = ~n5713 ;
  assign n5822 = n5711 & n67491 ;
  assign n5823 = n5821 | n5822 ;
  assign n5824 = n67482 & n5823 ;
  assign n5825 = n67485 & n5824 ;
  assign n5826 = n5820 | n5825 ;
  assign n5827 = n66979 & n5826 ;
  assign n5828 = n5426 & n5744 ;
  assign n5707 = n5435 | n5706 ;
  assign n67492 = ~n5707 ;
  assign n5829 = n67492 & n5787 ;
  assign n67493 = ~n5788 ;
  assign n5830 = n5706 & n67493 ;
  assign n5831 = n5829 | n5830 ;
  assign n5832 = n67482 & n5831 ;
  assign n5833 = n67485 & n5832 ;
  assign n5834 = n5828 | n5833 ;
  assign n5835 = n66868 & n5834 ;
  assign n5836 = n5434 & n5744 ;
  assign n5700 = n5443 | n5699 ;
  assign n67494 = ~n5700 ;
  assign n5837 = n5696 & n67494 ;
  assign n67495 = ~n5701 ;
  assign n5838 = n5699 & n67495 ;
  assign n5839 = n5837 | n5838 ;
  assign n5840 = n67482 & n5839 ;
  assign n5841 = n67485 & n5840 ;
  assign n5842 = n5836 | n5841 ;
  assign n5843 = n66797 & n5842 ;
  assign n5844 = n5442 & n5744 ;
  assign n5695 = n5451 | n5694 ;
  assign n67496 = ~n5695 ;
  assign n5845 = n67496 & n5783 ;
  assign n67497 = ~n5784 ;
  assign n5846 = n5694 & n67497 ;
  assign n5847 = n5845 | n5846 ;
  assign n5848 = n67482 & n5847 ;
  assign n5849 = n67485 & n5848 ;
  assign n5850 = n5844 | n5849 ;
  assign n5851 = n66654 & n5850 ;
  assign n5852 = n5450 & n5744 ;
  assign n5688 = n5459 | n5687 ;
  assign n67498 = ~n5688 ;
  assign n5853 = n5684 & n67498 ;
  assign n67499 = ~n5689 ;
  assign n5854 = n5687 & n67499 ;
  assign n5855 = n5853 | n5854 ;
  assign n5856 = n67482 & n5855 ;
  assign n5857 = n67485 & n5856 ;
  assign n5858 = n5852 | n5857 ;
  assign n5859 = n66560 & n5858 ;
  assign n5860 = n5458 & n5744 ;
  assign n5683 = n5467 | n5682 ;
  assign n67500 = ~n5683 ;
  assign n5861 = n67500 & n5779 ;
  assign n67501 = ~n5780 ;
  assign n5862 = n5682 & n67501 ;
  assign n5863 = n5861 | n5862 ;
  assign n5864 = n67482 & n5863 ;
  assign n5865 = n67485 & n5864 ;
  assign n5866 = n5860 | n5865 ;
  assign n5867 = n66505 & n5866 ;
  assign n5868 = n5466 & n5744 ;
  assign n5676 = n5475 | n5675 ;
  assign n67502 = ~n5676 ;
  assign n5869 = n5672 & n67502 ;
  assign n67503 = ~n5677 ;
  assign n5870 = n5675 & n67503 ;
  assign n5871 = n5869 | n5870 ;
  assign n5872 = n67482 & n5871 ;
  assign n5873 = n67485 & n5872 ;
  assign n5874 = n5868 | n5873 ;
  assign n5875 = n66379 & n5874 ;
  assign n5876 = n5474 & n5744 ;
  assign n5671 = n5483 | n5670 ;
  assign n67504 = ~n5671 ;
  assign n5877 = n67504 & n5775 ;
  assign n67505 = ~n5776 ;
  assign n5878 = n5670 & n67505 ;
  assign n5879 = n5877 | n5878 ;
  assign n5880 = n67482 & n5879 ;
  assign n5881 = n67485 & n5880 ;
  assign n5882 = n5876 | n5881 ;
  assign n5883 = n66299 & n5882 ;
  assign n5884 = n5482 & n5744 ;
  assign n5664 = n5491 | n5663 ;
  assign n67506 = ~n5664 ;
  assign n5885 = n5660 & n67506 ;
  assign n67507 = ~n5665 ;
  assign n5886 = n5663 & n67507 ;
  assign n5887 = n5885 | n5886 ;
  assign n5888 = n67482 & n5887 ;
  assign n5889 = n67485 & n5888 ;
  assign n5890 = n5884 | n5889 ;
  assign n5891 = n66244 & n5890 ;
  assign n5892 = n5490 & n5744 ;
  assign n5659 = n5499 | n5658 ;
  assign n67508 = ~n5659 ;
  assign n5893 = n67508 & n5771 ;
  assign n67509 = ~n5772 ;
  assign n5894 = n5658 & n67509 ;
  assign n5895 = n5893 | n5894 ;
  assign n5896 = n67482 & n5895 ;
  assign n5897 = n67485 & n5896 ;
  assign n5898 = n5892 | n5897 ;
  assign n5899 = n66145 & n5898 ;
  assign n5900 = n5498 & n5744 ;
  assign n5652 = n5507 | n5651 ;
  assign n67510 = ~n5652 ;
  assign n5901 = n5648 & n67510 ;
  assign n67511 = ~n5653 ;
  assign n5902 = n5651 & n67511 ;
  assign n5903 = n5901 | n5902 ;
  assign n5904 = n67482 & n5903 ;
  assign n5905 = n67485 & n5904 ;
  assign n5906 = n5900 | n5905 ;
  assign n5907 = n66081 & n5906 ;
  assign n5908 = n5506 & n5744 ;
  assign n5647 = n5515 | n5646 ;
  assign n67512 = ~n5647 ;
  assign n5909 = n67512 & n5767 ;
  assign n67513 = ~n5768 ;
  assign n5910 = n5646 & n67513 ;
  assign n5911 = n5909 | n5910 ;
  assign n5912 = n67482 & n5911 ;
  assign n5913 = n67485 & n5912 ;
  assign n5914 = n5908 | n5913 ;
  assign n5915 = n66043 & n5914 ;
  assign n5916 = n5514 & n5744 ;
  assign n5640 = n5523 | n5639 ;
  assign n67514 = ~n5640 ;
  assign n5917 = n5636 & n67514 ;
  assign n67515 = ~n5641 ;
  assign n5918 = n5639 & n67515 ;
  assign n5919 = n5917 | n5918 ;
  assign n5920 = n67482 & n5919 ;
  assign n5921 = n67485 & n5920 ;
  assign n5922 = n5916 | n5921 ;
  assign n5923 = n65960 & n5922 ;
  assign n5924 = n5522 & n5744 ;
  assign n5635 = n5531 | n5634 ;
  assign n67516 = ~n5635 ;
  assign n5925 = n67516 & n5763 ;
  assign n67517 = ~n5764 ;
  assign n5926 = n5634 & n67517 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = n67482 & n5927 ;
  assign n5929 = n67485 & n5928 ;
  assign n5930 = n5924 | n5929 ;
  assign n5931 = n65909 & n5930 ;
  assign n5932 = n5530 & n5744 ;
  assign n5628 = n5539 | n5627 ;
  assign n67518 = ~n5628 ;
  assign n5933 = n5624 & n67518 ;
  assign n67519 = ~n5629 ;
  assign n5934 = n5627 & n67519 ;
  assign n5935 = n5933 | n5934 ;
  assign n5936 = n67482 & n5935 ;
  assign n5937 = n67485 & n5936 ;
  assign n5938 = n5932 | n5937 ;
  assign n5939 = n65877 & n5938 ;
  assign n5940 = n5538 & n5744 ;
  assign n5623 = n5547 | n5622 ;
  assign n67520 = ~n5623 ;
  assign n5941 = n5618 & n67520 ;
  assign n67521 = ~n5760 ;
  assign n5942 = n5622 & n67521 ;
  assign n5943 = n5941 | n5942 ;
  assign n5944 = n67482 & n5943 ;
  assign n5945 = n67485 & n5944 ;
  assign n5946 = n5940 | n5945 ;
  assign n5947 = n65820 & n5946 ;
  assign n5948 = n5546 & n5744 ;
  assign n5949 = n5555 | n5616 ;
  assign n67522 = ~n5949 ;
  assign n5950 = n5613 & n67522 ;
  assign n67523 = ~n5617 ;
  assign n5951 = n5616 & n67523 ;
  assign n5952 = n5950 | n5951 ;
  assign n5953 = n67482 & n5952 ;
  assign n5954 = n67485 & n5953 ;
  assign n5955 = n5948 | n5954 ;
  assign n5956 = n65791 & n5955 ;
  assign n5957 = n5554 & n5744 ;
  assign n5958 = n5564 | n5612 ;
  assign n67524 = ~n5958 ;
  assign n5959 = n5608 & n67524 ;
  assign n67525 = ~n5756 ;
  assign n5960 = n5612 & n67525 ;
  assign n5961 = n5959 | n5960 ;
  assign n5962 = n67482 & n5961 ;
  assign n5963 = n67485 & n5962 ;
  assign n5964 = n5957 | n5963 ;
  assign n5965 = n65772 & n5964 ;
  assign n5966 = n5563 & n5744 ;
  assign n5967 = n5572 | n5606 ;
  assign n67526 = ~n5967 ;
  assign n5968 = n5603 & n67526 ;
  assign n67527 = ~n5607 ;
  assign n5969 = n5606 & n67527 ;
  assign n5970 = n5968 | n5969 ;
  assign n5971 = n67482 & n5970 ;
  assign n5972 = n67485 & n5971 ;
  assign n5973 = n5966 | n5972 ;
  assign n5974 = n65746 & n5973 ;
  assign n5975 = n5571 & n5744 ;
  assign n67528 = ~n5599 ;
  assign n5976 = n67528 & n5602 ;
  assign n5977 = n5598 | n5602 ;
  assign n67529 = ~n5977 ;
  assign n5978 = n5596 & n67529 ;
  assign n5979 = n5976 | n5978 ;
  assign n5980 = n67482 & n5979 ;
  assign n5981 = n67485 & n5980 ;
  assign n5982 = n5975 | n5981 ;
  assign n5983 = n65721 & n5982 ;
  assign n5745 = n5597 & n5744 ;
  assign n5750 = n5593 & n5594 ;
  assign n5984 = n67427 & n5750 ;
  assign n5985 = n5743 | n5984 ;
  assign n67530 = ~n5985 ;
  assign n5986 = n5596 & n67530 ;
  assign n5987 = n67485 & n5986 ;
  assign n5988 = n5745 | n5987 ;
  assign n5989 = n65686 & n5988 ;
  assign n67531 = ~x90 ;
  assign n5990 = x64 & n67531 ;
  assign n67532 = ~n74608 ;
  assign n5991 = n67532 & n5990 ;
  assign n67533 = ~n73745 ;
  assign n5992 = n67533 & n5991 ;
  assign n5993 = n66714 & n5992 ;
  assign n5994 = n66715 & n5993 ;
  assign n5998 = n67475 & n5997 ;
  assign n5999 = n5737 | n5998 ;
  assign n6000 = n67476 & n5999 ;
  assign n67534 = ~n6000 ;
  assign n6001 = n5994 & n67534 ;
  assign n67535 = ~n6001 ;
  assign n6002 = x38 & n67535 ;
  assign n6003 = n67422 & n5594 ;
  assign n6004 = n67423 & n6003 ;
  assign n6005 = n66509 & n6004 ;
  assign n6006 = n66510 & n6005 ;
  assign n6007 = n67485 & n6006 ;
  assign n6008 = n6002 | n6007 ;
  assign n6010 = x65 & n6008 ;
  assign n5995 = n67485 & n5994 ;
  assign n67536 = ~n5995 ;
  assign n5996 = x38 & n67536 ;
  assign n6009 = x65 | n6007 ;
  assign n6011 = n5996 | n6009 ;
  assign n67537 = ~n6010 ;
  assign n6012 = n67537 & n6011 ;
  assign n67538 = ~x37 ;
  assign n6013 = n67538 & x64 ;
  assign n6014 = n6012 | n6013 ;
  assign n6015 = n65670 & n6008 ;
  assign n67539 = ~n6015 ;
  assign n6016 = n6014 & n67539 ;
  assign n67540 = ~n5987 ;
  assign n6017 = x66 & n67540 ;
  assign n67541 = ~n5745 ;
  assign n6018 = n67541 & n6017 ;
  assign n6019 = n5989 | n6018 ;
  assign n6020 = n6016 | n6019 ;
  assign n67542 = ~n5989 ;
  assign n6021 = n67542 & n6020 ;
  assign n67543 = ~n5981 ;
  assign n6022 = x67 & n67543 ;
  assign n67544 = ~n5975 ;
  assign n6023 = n67544 & n6022 ;
  assign n6024 = n6021 | n6023 ;
  assign n67545 = ~n5983 ;
  assign n6025 = n67545 & n6024 ;
  assign n67546 = ~n5972 ;
  assign n6026 = x68 & n67546 ;
  assign n67547 = ~n5966 ;
  assign n6027 = n67547 & n6026 ;
  assign n6028 = n5974 | n6027 ;
  assign n6029 = n6025 | n6028 ;
  assign n67548 = ~n5974 ;
  assign n6030 = n67548 & n6029 ;
  assign n67549 = ~n5963 ;
  assign n6031 = x69 & n67549 ;
  assign n67550 = ~n5957 ;
  assign n6032 = n67550 & n6031 ;
  assign n6033 = n5965 | n6032 ;
  assign n6034 = n6030 | n6033 ;
  assign n67551 = ~n5965 ;
  assign n6035 = n67551 & n6034 ;
  assign n67552 = ~n5954 ;
  assign n6036 = x70 & n67552 ;
  assign n67553 = ~n5948 ;
  assign n6037 = n67553 & n6036 ;
  assign n6038 = n5956 | n6037 ;
  assign n6039 = n6035 | n6038 ;
  assign n67554 = ~n5956 ;
  assign n6040 = n67554 & n6039 ;
  assign n67555 = ~n5945 ;
  assign n6041 = x71 & n67555 ;
  assign n67556 = ~n5940 ;
  assign n6042 = n67556 & n6041 ;
  assign n6043 = n5947 | n6042 ;
  assign n6045 = n6040 | n6043 ;
  assign n67557 = ~n5947 ;
  assign n6046 = n67557 & n6045 ;
  assign n67558 = ~n5937 ;
  assign n6047 = x72 & n67558 ;
  assign n67559 = ~n5932 ;
  assign n6048 = n67559 & n6047 ;
  assign n6049 = n5939 | n6048 ;
  assign n6050 = n6046 | n6049 ;
  assign n67560 = ~n5939 ;
  assign n6051 = n67560 & n6050 ;
  assign n67561 = ~n5929 ;
  assign n6052 = x73 & n67561 ;
  assign n67562 = ~n5924 ;
  assign n6053 = n67562 & n6052 ;
  assign n6054 = n5931 | n6053 ;
  assign n6056 = n6051 | n6054 ;
  assign n67563 = ~n5931 ;
  assign n6057 = n67563 & n6056 ;
  assign n67564 = ~n5921 ;
  assign n6058 = x74 & n67564 ;
  assign n67565 = ~n5916 ;
  assign n6059 = n67565 & n6058 ;
  assign n6060 = n5923 | n6059 ;
  assign n6061 = n6057 | n6060 ;
  assign n67566 = ~n5923 ;
  assign n6062 = n67566 & n6061 ;
  assign n67567 = ~n5913 ;
  assign n6063 = x75 & n67567 ;
  assign n67568 = ~n5908 ;
  assign n6064 = n67568 & n6063 ;
  assign n6065 = n5915 | n6064 ;
  assign n6067 = n6062 | n6065 ;
  assign n67569 = ~n5915 ;
  assign n6068 = n67569 & n6067 ;
  assign n67570 = ~n5905 ;
  assign n6069 = x76 & n67570 ;
  assign n67571 = ~n5900 ;
  assign n6070 = n67571 & n6069 ;
  assign n6071 = n5907 | n6070 ;
  assign n6072 = n6068 | n6071 ;
  assign n67572 = ~n5907 ;
  assign n6073 = n67572 & n6072 ;
  assign n67573 = ~n5897 ;
  assign n6074 = x77 & n67573 ;
  assign n67574 = ~n5892 ;
  assign n6075 = n67574 & n6074 ;
  assign n6076 = n5899 | n6075 ;
  assign n6078 = n6073 | n6076 ;
  assign n67575 = ~n5899 ;
  assign n6079 = n67575 & n6078 ;
  assign n67576 = ~n5889 ;
  assign n6080 = x78 & n67576 ;
  assign n67577 = ~n5884 ;
  assign n6081 = n67577 & n6080 ;
  assign n6082 = n5891 | n6081 ;
  assign n6083 = n6079 | n6082 ;
  assign n67578 = ~n5891 ;
  assign n6084 = n67578 & n6083 ;
  assign n67579 = ~n5881 ;
  assign n6085 = x79 & n67579 ;
  assign n67580 = ~n5876 ;
  assign n6086 = n67580 & n6085 ;
  assign n6087 = n5883 | n6086 ;
  assign n6089 = n6084 | n6087 ;
  assign n67581 = ~n5883 ;
  assign n6090 = n67581 & n6089 ;
  assign n67582 = ~n5873 ;
  assign n6091 = x80 & n67582 ;
  assign n67583 = ~n5868 ;
  assign n6092 = n67583 & n6091 ;
  assign n6093 = n5875 | n6092 ;
  assign n6094 = n6090 | n6093 ;
  assign n67584 = ~n5875 ;
  assign n6095 = n67584 & n6094 ;
  assign n67585 = ~n5865 ;
  assign n6096 = x81 & n67585 ;
  assign n67586 = ~n5860 ;
  assign n6097 = n67586 & n6096 ;
  assign n6098 = n5867 | n6097 ;
  assign n6100 = n6095 | n6098 ;
  assign n67587 = ~n5867 ;
  assign n6101 = n67587 & n6100 ;
  assign n67588 = ~n5857 ;
  assign n6102 = x82 & n67588 ;
  assign n67589 = ~n5852 ;
  assign n6103 = n67589 & n6102 ;
  assign n6104 = n5859 | n6103 ;
  assign n6105 = n6101 | n6104 ;
  assign n67590 = ~n5859 ;
  assign n6106 = n67590 & n6105 ;
  assign n67591 = ~n5849 ;
  assign n6107 = x83 & n67591 ;
  assign n67592 = ~n5844 ;
  assign n6108 = n67592 & n6107 ;
  assign n6109 = n5851 | n6108 ;
  assign n6111 = n6106 | n6109 ;
  assign n67593 = ~n5851 ;
  assign n6112 = n67593 & n6111 ;
  assign n67594 = ~n5841 ;
  assign n6113 = x84 & n67594 ;
  assign n67595 = ~n5836 ;
  assign n6114 = n67595 & n6113 ;
  assign n6115 = n5843 | n6114 ;
  assign n6116 = n6112 | n6115 ;
  assign n67596 = ~n5843 ;
  assign n6117 = n67596 & n6116 ;
  assign n67597 = ~n5833 ;
  assign n6118 = x85 & n67597 ;
  assign n67598 = ~n5828 ;
  assign n6119 = n67598 & n6118 ;
  assign n6120 = n5835 | n6119 ;
  assign n6122 = n6117 | n6120 ;
  assign n67599 = ~n5835 ;
  assign n6123 = n67599 & n6122 ;
  assign n67600 = ~n5825 ;
  assign n6124 = x86 & n67600 ;
  assign n67601 = ~n5820 ;
  assign n6125 = n67601 & n6124 ;
  assign n6126 = n5827 | n6125 ;
  assign n6127 = n6123 | n6126 ;
  assign n67602 = ~n5827 ;
  assign n6128 = n67602 & n6127 ;
  assign n67603 = ~n5817 ;
  assign n6129 = x87 & n67603 ;
  assign n67604 = ~n5812 ;
  assign n6130 = n67604 & n6129 ;
  assign n6131 = n5819 | n6130 ;
  assign n6133 = n6128 | n6131 ;
  assign n67605 = ~n5819 ;
  assign n6134 = n67605 & n6133 ;
  assign n67606 = ~n5809 ;
  assign n6135 = x88 & n67606 ;
  assign n67607 = ~n5804 ;
  assign n6136 = n67607 & n6135 ;
  assign n6137 = n5811 | n6136 ;
  assign n6138 = n6134 | n6137 ;
  assign n67608 = ~n5811 ;
  assign n6139 = n67608 & n6138 ;
  assign n67609 = ~n5801 ;
  assign n6140 = x89 & n67609 ;
  assign n67610 = ~n5747 ;
  assign n6141 = n67610 & n6140 ;
  assign n6142 = n5803 | n6141 ;
  assign n6144 = n6139 | n6142 ;
  assign n67611 = ~n5803 ;
  assign n6145 = n67611 & n6144 ;
  assign n6152 = n67531 & n6151 ;
  assign n167 = ~n5744 ;
  assign n6153 = n167 & n6149 ;
  assign n6154 = n5386 & n5744 ;
  assign n67613 = ~n6154 ;
  assign n6155 = x90 & n67613 ;
  assign n67614 = ~n6153 ;
  assign n6156 = n67614 & n6155 ;
  assign n6157 = n73745 | n74608 ;
  assign n6158 = n294 | n6157 ;
  assign n6159 = n279 | n6158 ;
  assign n6160 = n6156 | n6159 ;
  assign n6161 = n6152 | n6160 ;
  assign n6163 = n6145 | n6161 ;
  assign n67615 = ~n6162 ;
  assign n6164 = n67615 & n6163 ;
  assign n67616 = ~n6139 ;
  assign n6143 = n67616 & n6142 ;
  assign n6167 = n5996 | n6007 ;
  assign n6168 = x65 & n6167 ;
  assign n67617 = ~n6168 ;
  assign n6169 = n6011 & n67617 ;
  assign n6170 = n6013 | n6169 ;
  assign n6171 = n67539 & n6170 ;
  assign n6173 = n6018 | n6171 ;
  assign n6174 = n67542 & n6173 ;
  assign n6175 = n5983 | n6023 ;
  assign n6177 = n6174 | n6175 ;
  assign n6178 = n67545 & n6177 ;
  assign n6180 = n6028 | n6178 ;
  assign n6181 = n67548 & n6180 ;
  assign n6183 = n6033 | n6181 ;
  assign n6184 = n67551 & n6183 ;
  assign n6185 = n6038 | n6184 ;
  assign n6187 = n67554 & n6185 ;
  assign n6188 = n6043 | n6187 ;
  assign n6189 = n67557 & n6188 ;
  assign n6190 = n6049 | n6189 ;
  assign n6192 = n67560 & n6190 ;
  assign n6193 = n6054 | n6192 ;
  assign n6194 = n67563 & n6193 ;
  assign n6195 = n6060 | n6194 ;
  assign n6197 = n67566 & n6195 ;
  assign n6198 = n6065 | n6197 ;
  assign n6199 = n67569 & n6198 ;
  assign n6200 = n6071 | n6199 ;
  assign n6202 = n67572 & n6200 ;
  assign n6203 = n6076 | n6202 ;
  assign n6204 = n67575 & n6203 ;
  assign n6205 = n6082 | n6204 ;
  assign n6207 = n67578 & n6205 ;
  assign n6208 = n6087 | n6207 ;
  assign n6209 = n67581 & n6208 ;
  assign n6210 = n6093 | n6209 ;
  assign n6212 = n67584 & n6210 ;
  assign n6213 = n6098 | n6212 ;
  assign n6214 = n67587 & n6213 ;
  assign n6215 = n6104 | n6214 ;
  assign n6217 = n67590 & n6215 ;
  assign n6218 = n6109 | n6217 ;
  assign n6219 = n67593 & n6218 ;
  assign n6220 = n6115 | n6219 ;
  assign n6222 = n67596 & n6220 ;
  assign n6223 = n6120 | n6222 ;
  assign n6224 = n67599 & n6223 ;
  assign n6225 = n6126 | n6224 ;
  assign n6227 = n67602 & n6225 ;
  assign n6228 = n6131 | n6227 ;
  assign n6229 = n67605 & n6228 ;
  assign n6230 = n6137 | n6229 ;
  assign n6247 = n5811 | n6142 ;
  assign n67618 = ~n6247 ;
  assign n6248 = n6230 & n67618 ;
  assign n6249 = n6143 | n6248 ;
  assign n166 = ~n6164 ;
  assign n6250 = n166 & n6249 ;
  assign n6232 = n67608 & n6230 ;
  assign n6233 = n6142 | n6232 ;
  assign n6234 = n67611 & n6233 ;
  assign n6235 = n6161 | n6234 ;
  assign n6251 = n5802 & n67615 ;
  assign n6252 = n6235 & n6251 ;
  assign n6253 = n6250 | n6252 ;
  assign n6236 = n5803 | n6156 ;
  assign n6237 = n6152 | n6236 ;
  assign n67620 = ~n6237 ;
  assign n6238 = n6144 & n67620 ;
  assign n6239 = n6152 | n6156 ;
  assign n67621 = ~n6234 ;
  assign n6240 = n67621 & n6239 ;
  assign n6241 = n6238 | n6240 ;
  assign n6242 = n166 & n6241 ;
  assign n6243 = n5743 & n6151 ;
  assign n6244 = n6235 & n6243 ;
  assign n6245 = n6242 | n6244 ;
  assign n67622 = ~x91 ;
  assign n6246 = n67622 & n6245 ;
  assign n67623 = ~n6244 ;
  assign n6608 = x91 & n67623 ;
  assign n67624 = ~n6242 ;
  assign n6609 = n67624 & n6608 ;
  assign n6610 = n6246 | n6609 ;
  assign n6254 = n67531 & n6253 ;
  assign n67625 = ~n6229 ;
  assign n6231 = n6137 & n67625 ;
  assign n6255 = n5819 | n6137 ;
  assign n67626 = ~n6255 ;
  assign n6256 = n6133 & n67626 ;
  assign n6257 = n6231 | n6256 ;
  assign n6258 = n166 & n6257 ;
  assign n6259 = n5810 & n67615 ;
  assign n6260 = n6235 & n6259 ;
  assign n6261 = n6258 | n6260 ;
  assign n6262 = n67348 & n6261 ;
  assign n67627 = ~n6260 ;
  assign n6596 = x89 & n67627 ;
  assign n67628 = ~n6258 ;
  assign n6597 = n67628 & n6596 ;
  assign n6598 = n6262 | n6597 ;
  assign n67629 = ~n6128 ;
  assign n6132 = n67629 & n6131 ;
  assign n6263 = n5827 | n6131 ;
  assign n67630 = ~n6263 ;
  assign n6264 = n6225 & n67630 ;
  assign n6265 = n6132 | n6264 ;
  assign n6266 = n166 & n6265 ;
  assign n6267 = n5818 & n67615 ;
  assign n6268 = n6235 & n6267 ;
  assign n6269 = n6266 | n6268 ;
  assign n6270 = n67222 & n6269 ;
  assign n67631 = ~n6224 ;
  assign n6226 = n6126 & n67631 ;
  assign n6271 = n5835 | n6126 ;
  assign n67632 = ~n6271 ;
  assign n6272 = n6122 & n67632 ;
  assign n6273 = n6226 | n6272 ;
  assign n6274 = n166 & n6273 ;
  assign n6275 = n5826 & n67615 ;
  assign n6276 = n6235 & n6275 ;
  assign n6277 = n6274 | n6276 ;
  assign n6278 = n67164 & n6277 ;
  assign n67633 = ~n6276 ;
  assign n6584 = x87 & n67633 ;
  assign n67634 = ~n6274 ;
  assign n6585 = n67634 & n6584 ;
  assign n6586 = n6278 | n6585 ;
  assign n67635 = ~n6117 ;
  assign n6121 = n67635 & n6120 ;
  assign n6279 = n5843 | n6120 ;
  assign n67636 = ~n6279 ;
  assign n6280 = n6220 & n67636 ;
  assign n6281 = n6121 | n6280 ;
  assign n6282 = n166 & n6281 ;
  assign n6283 = n5834 & n67615 ;
  assign n6284 = n6235 & n6283 ;
  assign n6285 = n6282 | n6284 ;
  assign n6286 = n66979 & n6285 ;
  assign n67637 = ~n6219 ;
  assign n6221 = n6115 & n67637 ;
  assign n6287 = n5851 | n6115 ;
  assign n67638 = ~n6287 ;
  assign n6288 = n6111 & n67638 ;
  assign n6289 = n6221 | n6288 ;
  assign n6290 = n166 & n6289 ;
  assign n6291 = n5842 & n67615 ;
  assign n6292 = n6235 & n6291 ;
  assign n6293 = n6290 | n6292 ;
  assign n6294 = n66868 & n6293 ;
  assign n67639 = ~n6292 ;
  assign n6572 = x85 & n67639 ;
  assign n67640 = ~n6290 ;
  assign n6573 = n67640 & n6572 ;
  assign n6574 = n6294 | n6573 ;
  assign n67641 = ~n6106 ;
  assign n6110 = n67641 & n6109 ;
  assign n6295 = n5859 | n6109 ;
  assign n67642 = ~n6295 ;
  assign n6296 = n6215 & n67642 ;
  assign n6297 = n6110 | n6296 ;
  assign n6298 = n166 & n6297 ;
  assign n6299 = n5850 & n67615 ;
  assign n6300 = n6235 & n6299 ;
  assign n6301 = n6298 | n6300 ;
  assign n6302 = n66797 & n6301 ;
  assign n67643 = ~n6214 ;
  assign n6216 = n6104 & n67643 ;
  assign n6303 = n5867 | n6104 ;
  assign n67644 = ~n6303 ;
  assign n6304 = n6100 & n67644 ;
  assign n6305 = n6216 | n6304 ;
  assign n6306 = n166 & n6305 ;
  assign n6307 = n5858 & n67615 ;
  assign n6308 = n6235 & n6307 ;
  assign n6309 = n6306 | n6308 ;
  assign n6310 = n66654 & n6309 ;
  assign n67645 = ~n6308 ;
  assign n6560 = x83 & n67645 ;
  assign n67646 = ~n6306 ;
  assign n6561 = n67646 & n6560 ;
  assign n6562 = n6310 | n6561 ;
  assign n67647 = ~n6095 ;
  assign n6099 = n67647 & n6098 ;
  assign n6311 = n5875 | n6098 ;
  assign n67648 = ~n6311 ;
  assign n6312 = n6210 & n67648 ;
  assign n6313 = n6099 | n6312 ;
  assign n6314 = n166 & n6313 ;
  assign n6315 = n5866 & n67615 ;
  assign n6316 = n6235 & n6315 ;
  assign n6317 = n6314 | n6316 ;
  assign n6318 = n66560 & n6317 ;
  assign n67649 = ~n6209 ;
  assign n6211 = n6093 & n67649 ;
  assign n6319 = n5883 | n6093 ;
  assign n67650 = ~n6319 ;
  assign n6320 = n6089 & n67650 ;
  assign n6321 = n6211 | n6320 ;
  assign n6322 = n166 & n6321 ;
  assign n6323 = n5874 & n67615 ;
  assign n6324 = n6235 & n6323 ;
  assign n6325 = n6322 | n6324 ;
  assign n6326 = n66505 & n6325 ;
  assign n67651 = ~n6324 ;
  assign n6548 = x81 & n67651 ;
  assign n67652 = ~n6322 ;
  assign n6549 = n67652 & n6548 ;
  assign n6550 = n6326 | n6549 ;
  assign n67653 = ~n6084 ;
  assign n6088 = n67653 & n6087 ;
  assign n6327 = n5891 | n6087 ;
  assign n67654 = ~n6327 ;
  assign n6328 = n6205 & n67654 ;
  assign n6329 = n6088 | n6328 ;
  assign n6330 = n166 & n6329 ;
  assign n6331 = n5882 & n67615 ;
  assign n6332 = n6235 & n6331 ;
  assign n6333 = n6330 | n6332 ;
  assign n6334 = n66379 & n6333 ;
  assign n67655 = ~n6204 ;
  assign n6206 = n6082 & n67655 ;
  assign n6335 = n5899 | n6082 ;
  assign n67656 = ~n6335 ;
  assign n6336 = n6078 & n67656 ;
  assign n6337 = n6206 | n6336 ;
  assign n6338 = n166 & n6337 ;
  assign n6339 = n5890 & n67615 ;
  assign n6340 = n6235 & n6339 ;
  assign n6341 = n6338 | n6340 ;
  assign n6342 = n66299 & n6341 ;
  assign n67657 = ~n6340 ;
  assign n6536 = x79 & n67657 ;
  assign n67658 = ~n6338 ;
  assign n6537 = n67658 & n6536 ;
  assign n6538 = n6342 | n6537 ;
  assign n67659 = ~n6073 ;
  assign n6077 = n67659 & n6076 ;
  assign n6343 = n5907 | n6076 ;
  assign n67660 = ~n6343 ;
  assign n6344 = n6200 & n67660 ;
  assign n6345 = n6077 | n6344 ;
  assign n6346 = n166 & n6345 ;
  assign n6347 = n5898 & n67615 ;
  assign n6348 = n6235 & n6347 ;
  assign n6349 = n6346 | n6348 ;
  assign n6350 = n66244 & n6349 ;
  assign n67661 = ~n6199 ;
  assign n6201 = n6071 & n67661 ;
  assign n6351 = n5915 | n6071 ;
  assign n67662 = ~n6351 ;
  assign n6352 = n6067 & n67662 ;
  assign n6353 = n6201 | n6352 ;
  assign n6354 = n166 & n6353 ;
  assign n6355 = n5906 & n67615 ;
  assign n6356 = n6235 & n6355 ;
  assign n6357 = n6354 | n6356 ;
  assign n6358 = n66145 & n6357 ;
  assign n67663 = ~n6356 ;
  assign n6524 = x77 & n67663 ;
  assign n67664 = ~n6354 ;
  assign n6525 = n67664 & n6524 ;
  assign n6526 = n6358 | n6525 ;
  assign n67665 = ~n6062 ;
  assign n6066 = n67665 & n6065 ;
  assign n6359 = n5923 | n6065 ;
  assign n67666 = ~n6359 ;
  assign n6360 = n6195 & n67666 ;
  assign n6361 = n6066 | n6360 ;
  assign n6362 = n166 & n6361 ;
  assign n6363 = n5914 & n67615 ;
  assign n6364 = n6235 & n6363 ;
  assign n6365 = n6362 | n6364 ;
  assign n6366 = n66081 & n6365 ;
  assign n67667 = ~n6194 ;
  assign n6196 = n6060 & n67667 ;
  assign n6367 = n5931 | n6060 ;
  assign n67668 = ~n6367 ;
  assign n6368 = n6056 & n67668 ;
  assign n6369 = n6196 | n6368 ;
  assign n6370 = n166 & n6369 ;
  assign n6371 = n5922 & n67615 ;
  assign n6372 = n6235 & n6371 ;
  assign n6373 = n6370 | n6372 ;
  assign n6374 = n66043 & n6373 ;
  assign n67669 = ~n6372 ;
  assign n6512 = x75 & n67669 ;
  assign n67670 = ~n6370 ;
  assign n6513 = n67670 & n6512 ;
  assign n6514 = n6374 | n6513 ;
  assign n67671 = ~n6051 ;
  assign n6055 = n67671 & n6054 ;
  assign n6375 = n5939 | n6054 ;
  assign n67672 = ~n6375 ;
  assign n6376 = n6190 & n67672 ;
  assign n6377 = n6055 | n6376 ;
  assign n6378 = n166 & n6377 ;
  assign n6379 = n5930 & n67615 ;
  assign n6380 = n6235 & n6379 ;
  assign n6381 = n6378 | n6380 ;
  assign n6382 = n65960 & n6381 ;
  assign n67673 = ~n6189 ;
  assign n6191 = n6049 & n67673 ;
  assign n6383 = n5947 | n6049 ;
  assign n67674 = ~n6383 ;
  assign n6384 = n6045 & n67674 ;
  assign n6385 = n6191 | n6384 ;
  assign n6386 = n166 & n6385 ;
  assign n6387 = n5938 & n67615 ;
  assign n6388 = n6235 & n6387 ;
  assign n6389 = n6386 | n6388 ;
  assign n6390 = n65909 & n6389 ;
  assign n67675 = ~n6388 ;
  assign n6500 = x73 & n67675 ;
  assign n67676 = ~n6386 ;
  assign n6501 = n67676 & n6500 ;
  assign n6502 = n6390 | n6501 ;
  assign n67677 = ~n6040 ;
  assign n6044 = n67677 & n6043 ;
  assign n6391 = n5956 | n6043 ;
  assign n67678 = ~n6391 ;
  assign n6392 = n6185 & n67678 ;
  assign n6393 = n6044 | n6392 ;
  assign n6394 = n166 & n6393 ;
  assign n6395 = n5946 & n67615 ;
  assign n6396 = n6235 & n6395 ;
  assign n6397 = n6394 | n6396 ;
  assign n6398 = n65877 & n6397 ;
  assign n67679 = ~n6184 ;
  assign n6186 = n6038 & n67679 ;
  assign n6399 = n5965 | n6038 ;
  assign n67680 = ~n6399 ;
  assign n6400 = n6034 & n67680 ;
  assign n6401 = n6186 | n6400 ;
  assign n6402 = n166 & n6401 ;
  assign n6403 = n5955 & n67615 ;
  assign n6404 = n6235 & n6403 ;
  assign n6405 = n6402 | n6404 ;
  assign n6406 = n65820 & n6405 ;
  assign n67681 = ~n6404 ;
  assign n6488 = x71 & n67681 ;
  assign n67682 = ~n6402 ;
  assign n6489 = n67682 & n6488 ;
  assign n6490 = n6406 | n6489 ;
  assign n67683 = ~n6030 ;
  assign n6182 = n67683 & n6033 ;
  assign n6407 = n5974 | n6033 ;
  assign n67684 = ~n6407 ;
  assign n6408 = n6180 & n67684 ;
  assign n6409 = n6182 | n6408 ;
  assign n6410 = n166 & n6409 ;
  assign n6411 = n5964 & n67615 ;
  assign n6412 = n6235 & n6411 ;
  assign n6413 = n6410 | n6412 ;
  assign n6414 = n65791 & n6413 ;
  assign n67685 = ~n6178 ;
  assign n6179 = n6028 & n67685 ;
  assign n6415 = n6021 | n6175 ;
  assign n6416 = n5983 | n6028 ;
  assign n67686 = ~n6416 ;
  assign n6417 = n6415 & n67686 ;
  assign n6418 = n6179 | n6417 ;
  assign n6419 = n166 & n6418 ;
  assign n6420 = n5973 & n67615 ;
  assign n6421 = n6235 & n6420 ;
  assign n6422 = n6419 | n6421 ;
  assign n6423 = n65772 & n6422 ;
  assign n67687 = ~n6421 ;
  assign n6477 = x69 & n67687 ;
  assign n67688 = ~n6419 ;
  assign n6478 = n67688 & n6477 ;
  assign n6479 = n6423 | n6478 ;
  assign n67689 = ~n6021 ;
  assign n6176 = n67689 & n6175 ;
  assign n6424 = n5989 | n6175 ;
  assign n67690 = ~n6424 ;
  assign n6425 = n6020 & n67690 ;
  assign n6426 = n6176 | n6425 ;
  assign n6427 = n166 & n6426 ;
  assign n6428 = n5982 & n67615 ;
  assign n6429 = n6235 & n6428 ;
  assign n6430 = n6427 | n6429 ;
  assign n6431 = n65746 & n6430 ;
  assign n67691 = ~n6171 ;
  assign n6172 = n6019 & n67691 ;
  assign n6432 = n6015 | n6019 ;
  assign n67692 = ~n6432 ;
  assign n6433 = n6014 & n67692 ;
  assign n6434 = n6172 | n6433 ;
  assign n6435 = n166 & n6434 ;
  assign n6436 = n5988 & n67615 ;
  assign n6437 = n6235 & n6436 ;
  assign n6438 = n6435 | n6437 ;
  assign n6439 = n65721 & n6438 ;
  assign n67693 = ~n6437 ;
  assign n6467 = x67 & n67693 ;
  assign n67694 = ~n6435 ;
  assign n6468 = n67694 & n6467 ;
  assign n6469 = n6439 | n6468 ;
  assign n6440 = n6011 & n6013 ;
  assign n6441 = n67537 & n6440 ;
  assign n67695 = ~n6441 ;
  assign n6442 = n6170 & n67695 ;
  assign n6443 = n166 & n6442 ;
  assign n6444 = n6008 & n67615 ;
  assign n6445 = n6235 & n6444 ;
  assign n6446 = n6443 | n6445 ;
  assign n6447 = n65686 & n6446 ;
  assign n67696 = ~x36 ;
  assign n6457 = n67696 & x64 ;
  assign n6166 = n6013 & n166 ;
  assign n6448 = n67615 & n6235 ;
  assign n67697 = ~n6448 ;
  assign n6449 = x64 & n67697 ;
  assign n67698 = ~n6449 ;
  assign n6450 = x37 & n67698 ;
  assign n6451 = n6166 | n6450 ;
  assign n6452 = x65 & n6451 ;
  assign n6165 = x64 & n166 ;
  assign n67699 = ~n6165 ;
  assign n6453 = x37 & n67699 ;
  assign n6454 = n6013 & n67697 ;
  assign n6455 = x65 | n6454 ;
  assign n6456 = n6453 | n6455 ;
  assign n67700 = ~n6452 ;
  assign n6458 = n67700 & n6456 ;
  assign n6459 = n6457 | n6458 ;
  assign n6460 = n6166 | n6453 ;
  assign n6461 = n65670 & n6460 ;
  assign n67701 = ~n6461 ;
  assign n6462 = n6459 & n67701 ;
  assign n67702 = ~n6445 ;
  assign n6463 = x66 & n67702 ;
  assign n67703 = ~n6443 ;
  assign n6464 = n67703 & n6463 ;
  assign n6465 = n6447 | n6464 ;
  assign n6466 = n6462 | n6465 ;
  assign n67704 = ~n6447 ;
  assign n6470 = n67704 & n6466 ;
  assign n6471 = n6469 | n6470 ;
  assign n67705 = ~n6439 ;
  assign n6472 = n67705 & n6471 ;
  assign n67706 = ~n6429 ;
  assign n6473 = x68 & n67706 ;
  assign n67707 = ~n6427 ;
  assign n6474 = n67707 & n6473 ;
  assign n6475 = n6431 | n6474 ;
  assign n6476 = n6472 | n6475 ;
  assign n67708 = ~n6431 ;
  assign n6480 = n67708 & n6476 ;
  assign n6481 = n6479 | n6480 ;
  assign n67709 = ~n6423 ;
  assign n6482 = n67709 & n6481 ;
  assign n67710 = ~n6412 ;
  assign n6483 = x70 & n67710 ;
  assign n67711 = ~n6410 ;
  assign n6484 = n67711 & n6483 ;
  assign n6485 = n6414 | n6484 ;
  assign n6487 = n6482 | n6485 ;
  assign n67712 = ~n6414 ;
  assign n6492 = n67712 & n6487 ;
  assign n6493 = n6490 | n6492 ;
  assign n67713 = ~n6406 ;
  assign n6494 = n67713 & n6493 ;
  assign n67714 = ~n6396 ;
  assign n6495 = x72 & n67714 ;
  assign n67715 = ~n6394 ;
  assign n6496 = n67715 & n6495 ;
  assign n6497 = n6398 | n6496 ;
  assign n6499 = n6494 | n6497 ;
  assign n67716 = ~n6398 ;
  assign n6504 = n67716 & n6499 ;
  assign n6505 = n6502 | n6504 ;
  assign n67717 = ~n6390 ;
  assign n6506 = n67717 & n6505 ;
  assign n67718 = ~n6380 ;
  assign n6507 = x74 & n67718 ;
  assign n67719 = ~n6378 ;
  assign n6508 = n67719 & n6507 ;
  assign n6509 = n6382 | n6508 ;
  assign n6511 = n6506 | n6509 ;
  assign n67720 = ~n6382 ;
  assign n6516 = n67720 & n6511 ;
  assign n6517 = n6514 | n6516 ;
  assign n67721 = ~n6374 ;
  assign n6518 = n67721 & n6517 ;
  assign n67722 = ~n6364 ;
  assign n6519 = x76 & n67722 ;
  assign n67723 = ~n6362 ;
  assign n6520 = n67723 & n6519 ;
  assign n6521 = n6366 | n6520 ;
  assign n6523 = n6518 | n6521 ;
  assign n67724 = ~n6366 ;
  assign n6528 = n67724 & n6523 ;
  assign n6529 = n6526 | n6528 ;
  assign n67725 = ~n6358 ;
  assign n6530 = n67725 & n6529 ;
  assign n67726 = ~n6348 ;
  assign n6531 = x78 & n67726 ;
  assign n67727 = ~n6346 ;
  assign n6532 = n67727 & n6531 ;
  assign n6533 = n6350 | n6532 ;
  assign n6535 = n6530 | n6533 ;
  assign n67728 = ~n6350 ;
  assign n6540 = n67728 & n6535 ;
  assign n6541 = n6538 | n6540 ;
  assign n67729 = ~n6342 ;
  assign n6542 = n67729 & n6541 ;
  assign n67730 = ~n6332 ;
  assign n6543 = x80 & n67730 ;
  assign n67731 = ~n6330 ;
  assign n6544 = n67731 & n6543 ;
  assign n6545 = n6334 | n6544 ;
  assign n6547 = n6542 | n6545 ;
  assign n67732 = ~n6334 ;
  assign n6552 = n67732 & n6547 ;
  assign n6553 = n6550 | n6552 ;
  assign n67733 = ~n6326 ;
  assign n6554 = n67733 & n6553 ;
  assign n67734 = ~n6316 ;
  assign n6555 = x82 & n67734 ;
  assign n67735 = ~n6314 ;
  assign n6556 = n67735 & n6555 ;
  assign n6557 = n6318 | n6556 ;
  assign n6559 = n6554 | n6557 ;
  assign n67736 = ~n6318 ;
  assign n6564 = n67736 & n6559 ;
  assign n6565 = n6562 | n6564 ;
  assign n67737 = ~n6310 ;
  assign n6566 = n67737 & n6565 ;
  assign n67738 = ~n6300 ;
  assign n6567 = x84 & n67738 ;
  assign n67739 = ~n6298 ;
  assign n6568 = n67739 & n6567 ;
  assign n6569 = n6302 | n6568 ;
  assign n6571 = n6566 | n6569 ;
  assign n67740 = ~n6302 ;
  assign n6576 = n67740 & n6571 ;
  assign n6577 = n6574 | n6576 ;
  assign n67741 = ~n6294 ;
  assign n6578 = n67741 & n6577 ;
  assign n67742 = ~n6284 ;
  assign n6579 = x86 & n67742 ;
  assign n67743 = ~n6282 ;
  assign n6580 = n67743 & n6579 ;
  assign n6581 = n6286 | n6580 ;
  assign n6583 = n6578 | n6581 ;
  assign n67744 = ~n6286 ;
  assign n6588 = n67744 & n6583 ;
  assign n6589 = n6586 | n6588 ;
  assign n67745 = ~n6278 ;
  assign n6590 = n67745 & n6589 ;
  assign n67746 = ~n6268 ;
  assign n6591 = x88 & n67746 ;
  assign n67747 = ~n6266 ;
  assign n6592 = n67747 & n6591 ;
  assign n6593 = n6270 | n6592 ;
  assign n6595 = n6590 | n6593 ;
  assign n67748 = ~n6270 ;
  assign n6600 = n67748 & n6595 ;
  assign n6601 = n6598 | n6600 ;
  assign n67749 = ~n6262 ;
  assign n6602 = n67749 & n6601 ;
  assign n67750 = ~n6252 ;
  assign n6603 = x90 & n67750 ;
  assign n67751 = ~n6250 ;
  assign n6604 = n67751 & n6603 ;
  assign n6605 = n6254 | n6604 ;
  assign n6607 = n6602 | n6605 ;
  assign n67752 = ~n6254 ;
  assign n6611 = n67752 & n6607 ;
  assign n6612 = n6610 | n6611 ;
  assign n67753 = ~n6246 ;
  assign n6613 = n67753 & n6612 ;
  assign n6614 = n65542 | n65647 ;
  assign n6615 = n65429 | n6614 ;
  assign n6616 = n6613 | n6615 ;
  assign n6683 = n6253 & n6616 ;
  assign n6606 = n6262 | n6605 ;
  assign n6620 = x65 & n6460 ;
  assign n67754 = ~n6620 ;
  assign n6621 = n6456 & n67754 ;
  assign n6623 = n6457 | n6621 ;
  assign n6625 = n67701 & n6623 ;
  assign n6626 = n6465 | n6625 ;
  assign n6627 = n67704 & n6626 ;
  assign n6628 = n6469 | n6627 ;
  assign n6629 = n67705 & n6628 ;
  assign n6630 = n6475 | n6629 ;
  assign n6631 = n67708 & n6630 ;
  assign n6632 = n6479 | n6631 ;
  assign n6633 = n67709 & n6632 ;
  assign n6634 = n6485 | n6633 ;
  assign n6635 = n67712 & n6634 ;
  assign n6636 = n6490 | n6635 ;
  assign n6637 = n67713 & n6636 ;
  assign n6638 = n6497 | n6637 ;
  assign n6639 = n67716 & n6638 ;
  assign n6640 = n6502 | n6639 ;
  assign n6641 = n67717 & n6640 ;
  assign n6642 = n6509 | n6641 ;
  assign n6643 = n67720 & n6642 ;
  assign n6644 = n6514 | n6643 ;
  assign n6645 = n67721 & n6644 ;
  assign n6646 = n6521 | n6645 ;
  assign n6647 = n67724 & n6646 ;
  assign n6648 = n6526 | n6647 ;
  assign n6649 = n67725 & n6648 ;
  assign n6650 = n6533 | n6649 ;
  assign n6651 = n67728 & n6650 ;
  assign n6652 = n6538 | n6651 ;
  assign n6653 = n67729 & n6652 ;
  assign n6654 = n6545 | n6653 ;
  assign n6655 = n67732 & n6654 ;
  assign n6656 = n6550 | n6655 ;
  assign n6657 = n67733 & n6656 ;
  assign n6658 = n6557 | n6657 ;
  assign n6659 = n67736 & n6658 ;
  assign n6660 = n6562 | n6659 ;
  assign n6661 = n67737 & n6660 ;
  assign n6662 = n6569 | n6661 ;
  assign n6663 = n67740 & n6662 ;
  assign n6664 = n6574 | n6663 ;
  assign n6665 = n67741 & n6664 ;
  assign n6666 = n6581 | n6665 ;
  assign n6667 = n67744 & n6666 ;
  assign n6668 = n6586 | n6667 ;
  assign n6669 = n67745 & n6668 ;
  assign n6670 = n6593 | n6669 ;
  assign n6671 = n67748 & n6670 ;
  assign n6672 = n6598 | n6671 ;
  assign n67755 = ~n6606 ;
  assign n6684 = n67755 & n6672 ;
  assign n6673 = n67749 & n6672 ;
  assign n67756 = ~n6673 ;
  assign n6685 = n6605 & n67756 ;
  assign n6686 = n6684 | n6685 ;
  assign n67757 = ~n6615 ;
  assign n6687 = n67757 & n6686 ;
  assign n67758 = ~n6613 ;
  assign n6688 = n67758 & n6687 ;
  assign n6689 = n6683 | n6688 ;
  assign n67759 = ~n6245 ;
  assign n6618 = n67759 & n6616 ;
  assign n67760 = ~n6611 ;
  assign n6676 = n6610 & n67760 ;
  assign n6674 = n6605 | n6673 ;
  assign n6677 = n6254 | n6610 ;
  assign n67761 = ~n6677 ;
  assign n6678 = n6674 & n67761 ;
  assign n6679 = n6676 | n6678 ;
  assign n6680 = n6616 | n6679 ;
  assign n67762 = ~n6618 ;
  assign n6681 = n67762 & n6680 ;
  assign n67763 = ~x92 ;
  assign n6682 = n67763 & n6681 ;
  assign n6690 = n67622 & n6689 ;
  assign n6691 = n6261 & n6616 ;
  assign n6599 = n6270 | n6598 ;
  assign n67764 = ~n6599 ;
  assign n6692 = n6595 & n67764 ;
  assign n67765 = ~n6600 ;
  assign n6693 = n6598 & n67765 ;
  assign n6694 = n6692 | n6693 ;
  assign n6695 = n67757 & n6694 ;
  assign n6696 = n67758 & n6695 ;
  assign n6697 = n6691 | n6696 ;
  assign n6698 = n67531 & n6697 ;
  assign n6699 = n6269 & n6616 ;
  assign n6594 = n6278 | n6593 ;
  assign n67766 = ~n6594 ;
  assign n6700 = n67766 & n6668 ;
  assign n67767 = ~n6669 ;
  assign n6701 = n6593 & n67767 ;
  assign n6702 = n6700 | n6701 ;
  assign n6703 = n67757 & n6702 ;
  assign n6704 = n67758 & n6703 ;
  assign n6705 = n6699 | n6704 ;
  assign n6706 = n67348 & n6705 ;
  assign n6707 = n6277 & n6616 ;
  assign n6587 = n6286 | n6586 ;
  assign n67768 = ~n6587 ;
  assign n6708 = n6583 & n67768 ;
  assign n67769 = ~n6588 ;
  assign n6709 = n6586 & n67769 ;
  assign n6710 = n6708 | n6709 ;
  assign n6711 = n67757 & n6710 ;
  assign n6712 = n67758 & n6711 ;
  assign n6713 = n6707 | n6712 ;
  assign n6714 = n67222 & n6713 ;
  assign n6715 = n6285 & n6616 ;
  assign n6582 = n6294 | n6581 ;
  assign n67770 = ~n6582 ;
  assign n6716 = n67770 & n6664 ;
  assign n67771 = ~n6665 ;
  assign n6717 = n6581 & n67771 ;
  assign n6718 = n6716 | n6717 ;
  assign n6719 = n67757 & n6718 ;
  assign n6720 = n67758 & n6719 ;
  assign n6721 = n6715 | n6720 ;
  assign n6722 = n67164 & n6721 ;
  assign n6723 = n6293 & n6616 ;
  assign n6575 = n6302 | n6574 ;
  assign n67772 = ~n6575 ;
  assign n6724 = n6571 & n67772 ;
  assign n67773 = ~n6576 ;
  assign n6725 = n6574 & n67773 ;
  assign n6726 = n6724 | n6725 ;
  assign n6727 = n67757 & n6726 ;
  assign n6728 = n67758 & n6727 ;
  assign n6729 = n6723 | n6728 ;
  assign n6730 = n66979 & n6729 ;
  assign n6731 = n6301 & n6616 ;
  assign n6570 = n6310 | n6569 ;
  assign n67774 = ~n6570 ;
  assign n6732 = n67774 & n6660 ;
  assign n67775 = ~n6661 ;
  assign n6733 = n6569 & n67775 ;
  assign n6734 = n6732 | n6733 ;
  assign n6735 = n67757 & n6734 ;
  assign n6736 = n67758 & n6735 ;
  assign n6737 = n6731 | n6736 ;
  assign n6738 = n66868 & n6737 ;
  assign n6739 = n6309 & n6616 ;
  assign n6563 = n6318 | n6562 ;
  assign n67776 = ~n6563 ;
  assign n6740 = n6559 & n67776 ;
  assign n67777 = ~n6564 ;
  assign n6741 = n6562 & n67777 ;
  assign n6742 = n6740 | n6741 ;
  assign n6743 = n67757 & n6742 ;
  assign n6744 = n67758 & n6743 ;
  assign n6745 = n6739 | n6744 ;
  assign n6746 = n66797 & n6745 ;
  assign n6747 = n6317 & n6616 ;
  assign n6558 = n6326 | n6557 ;
  assign n67778 = ~n6558 ;
  assign n6748 = n67778 & n6656 ;
  assign n67779 = ~n6657 ;
  assign n6749 = n6557 & n67779 ;
  assign n6750 = n6748 | n6749 ;
  assign n6751 = n67757 & n6750 ;
  assign n6752 = n67758 & n6751 ;
  assign n6753 = n6747 | n6752 ;
  assign n6754 = n66654 & n6753 ;
  assign n6755 = n6325 & n6616 ;
  assign n6551 = n6334 | n6550 ;
  assign n67780 = ~n6551 ;
  assign n6756 = n6547 & n67780 ;
  assign n67781 = ~n6552 ;
  assign n6757 = n6550 & n67781 ;
  assign n6758 = n6756 | n6757 ;
  assign n6759 = n67757 & n6758 ;
  assign n6760 = n67758 & n6759 ;
  assign n6761 = n6755 | n6760 ;
  assign n6762 = n66560 & n6761 ;
  assign n6763 = n6333 & n6616 ;
  assign n6546 = n6342 | n6545 ;
  assign n67782 = ~n6546 ;
  assign n6764 = n67782 & n6652 ;
  assign n67783 = ~n6653 ;
  assign n6765 = n6545 & n67783 ;
  assign n6766 = n6764 | n6765 ;
  assign n6767 = n67757 & n6766 ;
  assign n6768 = n67758 & n6767 ;
  assign n6769 = n6763 | n6768 ;
  assign n6770 = n66505 & n6769 ;
  assign n6771 = n6341 & n6616 ;
  assign n6539 = n6350 | n6538 ;
  assign n67784 = ~n6539 ;
  assign n6772 = n6535 & n67784 ;
  assign n67785 = ~n6540 ;
  assign n6773 = n6538 & n67785 ;
  assign n6774 = n6772 | n6773 ;
  assign n6775 = n67757 & n6774 ;
  assign n6776 = n67758 & n6775 ;
  assign n6777 = n6771 | n6776 ;
  assign n6778 = n66379 & n6777 ;
  assign n6779 = n6349 & n6616 ;
  assign n6534 = n6358 | n6533 ;
  assign n67786 = ~n6534 ;
  assign n6780 = n67786 & n6648 ;
  assign n67787 = ~n6649 ;
  assign n6781 = n6533 & n67787 ;
  assign n6782 = n6780 | n6781 ;
  assign n6783 = n67757 & n6782 ;
  assign n6784 = n67758 & n6783 ;
  assign n6785 = n6779 | n6784 ;
  assign n6786 = n66299 & n6785 ;
  assign n6787 = n6357 & n6616 ;
  assign n6527 = n6366 | n6526 ;
  assign n67788 = ~n6527 ;
  assign n6788 = n6523 & n67788 ;
  assign n67789 = ~n6528 ;
  assign n6789 = n6526 & n67789 ;
  assign n6790 = n6788 | n6789 ;
  assign n6791 = n67757 & n6790 ;
  assign n6792 = n67758 & n6791 ;
  assign n6793 = n6787 | n6792 ;
  assign n6794 = n66244 & n6793 ;
  assign n6795 = n6365 & n6616 ;
  assign n6522 = n6374 | n6521 ;
  assign n67790 = ~n6522 ;
  assign n6796 = n67790 & n6644 ;
  assign n67791 = ~n6645 ;
  assign n6797 = n6521 & n67791 ;
  assign n6798 = n6796 | n6797 ;
  assign n6799 = n67757 & n6798 ;
  assign n6800 = n67758 & n6799 ;
  assign n6801 = n6795 | n6800 ;
  assign n6802 = n66145 & n6801 ;
  assign n6803 = n6373 & n6616 ;
  assign n6515 = n6382 | n6514 ;
  assign n67792 = ~n6515 ;
  assign n6804 = n6511 & n67792 ;
  assign n67793 = ~n6516 ;
  assign n6805 = n6514 & n67793 ;
  assign n6806 = n6804 | n6805 ;
  assign n6807 = n67757 & n6806 ;
  assign n6808 = n67758 & n6807 ;
  assign n6809 = n6803 | n6808 ;
  assign n6810 = n66081 & n6809 ;
  assign n6811 = n6381 & n6616 ;
  assign n6510 = n6390 | n6509 ;
  assign n67794 = ~n6510 ;
  assign n6812 = n67794 & n6640 ;
  assign n67795 = ~n6641 ;
  assign n6813 = n6509 & n67795 ;
  assign n6814 = n6812 | n6813 ;
  assign n6815 = n67757 & n6814 ;
  assign n6816 = n67758 & n6815 ;
  assign n6817 = n6811 | n6816 ;
  assign n6818 = n66043 & n6817 ;
  assign n6819 = n6389 & n6616 ;
  assign n6503 = n6398 | n6502 ;
  assign n67796 = ~n6503 ;
  assign n6820 = n6499 & n67796 ;
  assign n67797 = ~n6504 ;
  assign n6821 = n6502 & n67797 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = n67757 & n6822 ;
  assign n6824 = n67758 & n6823 ;
  assign n6825 = n6819 | n6824 ;
  assign n6826 = n65960 & n6825 ;
  assign n6827 = n6397 & n6616 ;
  assign n6498 = n6406 | n6497 ;
  assign n67798 = ~n6498 ;
  assign n6828 = n67798 & n6636 ;
  assign n67799 = ~n6637 ;
  assign n6829 = n6497 & n67799 ;
  assign n6830 = n6828 | n6829 ;
  assign n6831 = n67757 & n6830 ;
  assign n6832 = n67758 & n6831 ;
  assign n6833 = n6827 | n6832 ;
  assign n6834 = n65909 & n6833 ;
  assign n6835 = n6405 & n6616 ;
  assign n6491 = n6414 | n6490 ;
  assign n67800 = ~n6491 ;
  assign n6836 = n6487 & n67800 ;
  assign n67801 = ~n6492 ;
  assign n6837 = n6490 & n67801 ;
  assign n6838 = n6836 | n6837 ;
  assign n6839 = n67757 & n6838 ;
  assign n6840 = n67758 & n6839 ;
  assign n6841 = n6835 | n6840 ;
  assign n6842 = n65877 & n6841 ;
  assign n6843 = n6413 & n6616 ;
  assign n6486 = n6423 | n6485 ;
  assign n67802 = ~n6486 ;
  assign n6844 = n67802 & n6632 ;
  assign n67803 = ~n6633 ;
  assign n6845 = n6485 & n67803 ;
  assign n6846 = n6844 | n6845 ;
  assign n6847 = n67757 & n6846 ;
  assign n6848 = n67758 & n6847 ;
  assign n6849 = n6843 | n6848 ;
  assign n6850 = n65820 & n6849 ;
  assign n6851 = n6422 & n6616 ;
  assign n6619 = n6431 | n6479 ;
  assign n67804 = ~n6619 ;
  assign n6852 = n6476 & n67804 ;
  assign n67805 = ~n6480 ;
  assign n6853 = n6479 & n67805 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = n67757 & n6854 ;
  assign n6856 = n67758 & n6855 ;
  assign n6857 = n6851 | n6856 ;
  assign n6858 = n65791 & n6857 ;
  assign n6859 = n6430 & n6616 ;
  assign n6860 = n6439 | n6475 ;
  assign n67806 = ~n6860 ;
  assign n6861 = n6628 & n67806 ;
  assign n67807 = ~n6629 ;
  assign n6862 = n6475 & n67807 ;
  assign n6863 = n6861 | n6862 ;
  assign n6864 = n67757 & n6863 ;
  assign n6865 = n67758 & n6864 ;
  assign n6866 = n6859 | n6865 ;
  assign n6867 = n65772 & n6866 ;
  assign n6868 = n6438 & n6616 ;
  assign n6869 = n6447 | n6469 ;
  assign n67808 = ~n6869 ;
  assign n6870 = n6626 & n67808 ;
  assign n67809 = ~n6470 ;
  assign n6871 = n6469 & n67809 ;
  assign n6872 = n6870 | n6871 ;
  assign n6873 = n67757 & n6872 ;
  assign n6874 = n67758 & n6873 ;
  assign n6875 = n6868 | n6874 ;
  assign n6876 = n65746 & n6875 ;
  assign n6877 = n6446 & n6616 ;
  assign n6624 = n6461 | n6465 ;
  assign n67810 = ~n6624 ;
  assign n6878 = n6459 & n67810 ;
  assign n67811 = ~n6625 ;
  assign n6879 = n6465 & n67811 ;
  assign n6880 = n6878 | n6879 ;
  assign n6881 = n67757 & n6880 ;
  assign n6882 = n67758 & n6881 ;
  assign n6883 = n6877 | n6882 ;
  assign n6884 = n65721 & n6883 ;
  assign n6617 = n6460 & n6616 ;
  assign n6622 = n6456 & n6457 ;
  assign n6885 = n67700 & n6622 ;
  assign n6886 = n6615 | n6885 ;
  assign n67812 = ~n6886 ;
  assign n6887 = n6459 & n67812 ;
  assign n6888 = n67758 & n6887 ;
  assign n6889 = n6617 | n6888 ;
  assign n6890 = n65686 & n6889 ;
  assign n6897 = n67423 & n6457 ;
  assign n6898 = n66509 & n6897 ;
  assign n6899 = n66510 & n6898 ;
  assign n6900 = n67758 & n6899 ;
  assign n6891 = x64 & n67763 ;
  assign n6892 = n67533 & n6891 ;
  assign n6893 = n66714 & n6892 ;
  assign n6894 = n66715 & n6893 ;
  assign n6675 = n67752 & n6674 ;
  assign n6908 = n6610 | n6675 ;
  assign n6909 = n67753 & n6908 ;
  assign n67813 = ~n6909 ;
  assign n6910 = n6894 & n67813 ;
  assign n67814 = ~n6910 ;
  assign n6911 = x36 & n67814 ;
  assign n6912 = n6900 | n6911 ;
  assign n6913 = n65670 & n6912 ;
  assign n6895 = n67758 & n6894 ;
  assign n67815 = ~n6895 ;
  assign n6896 = x36 & n67815 ;
  assign n6901 = n6896 | n6900 ;
  assign n6902 = x65 & n6901 ;
  assign n6904 = x65 | n6900 ;
  assign n6905 = n6896 | n6904 ;
  assign n67816 = ~n6902 ;
  assign n6906 = n67816 & n6905 ;
  assign n67817 = ~x35 ;
  assign n6907 = n67817 & x64 ;
  assign n6914 = n6906 | n6907 ;
  assign n67818 = ~n6913 ;
  assign n6915 = n67818 & n6914 ;
  assign n67819 = ~n6888 ;
  assign n6916 = x66 & n67819 ;
  assign n67820 = ~n6617 ;
  assign n6917 = n67820 & n6916 ;
  assign n6918 = n6890 | n6917 ;
  assign n6919 = n6915 | n6918 ;
  assign n67821 = ~n6890 ;
  assign n6920 = n67821 & n6919 ;
  assign n67822 = ~n6882 ;
  assign n6921 = x67 & n67822 ;
  assign n67823 = ~n6877 ;
  assign n6922 = n67823 & n6921 ;
  assign n6923 = n6884 | n6922 ;
  assign n6924 = n6920 | n6923 ;
  assign n67824 = ~n6884 ;
  assign n6925 = n67824 & n6924 ;
  assign n67825 = ~n6874 ;
  assign n6926 = x68 & n67825 ;
  assign n67826 = ~n6868 ;
  assign n6927 = n67826 & n6926 ;
  assign n6928 = n6876 | n6927 ;
  assign n6929 = n6925 | n6928 ;
  assign n67827 = ~n6876 ;
  assign n6930 = n67827 & n6929 ;
  assign n67828 = ~n6865 ;
  assign n6931 = x69 & n67828 ;
  assign n67829 = ~n6859 ;
  assign n6932 = n67829 & n6931 ;
  assign n6933 = n6867 | n6932 ;
  assign n6934 = n6930 | n6933 ;
  assign n67830 = ~n6867 ;
  assign n6935 = n67830 & n6934 ;
  assign n67831 = ~n6856 ;
  assign n6936 = x70 & n67831 ;
  assign n67832 = ~n6851 ;
  assign n6937 = n67832 & n6936 ;
  assign n6938 = n6858 | n6937 ;
  assign n6940 = n6935 | n6938 ;
  assign n67833 = ~n6858 ;
  assign n6941 = n67833 & n6940 ;
  assign n67834 = ~n6848 ;
  assign n6942 = x71 & n67834 ;
  assign n67835 = ~n6843 ;
  assign n6943 = n67835 & n6942 ;
  assign n6944 = n6850 | n6943 ;
  assign n6945 = n6941 | n6944 ;
  assign n67836 = ~n6850 ;
  assign n6946 = n67836 & n6945 ;
  assign n67837 = ~n6840 ;
  assign n6947 = x72 & n67837 ;
  assign n67838 = ~n6835 ;
  assign n6948 = n67838 & n6947 ;
  assign n6949 = n6842 | n6948 ;
  assign n6951 = n6946 | n6949 ;
  assign n67839 = ~n6842 ;
  assign n6952 = n67839 & n6951 ;
  assign n67840 = ~n6832 ;
  assign n6953 = x73 & n67840 ;
  assign n67841 = ~n6827 ;
  assign n6954 = n67841 & n6953 ;
  assign n6955 = n6834 | n6954 ;
  assign n6956 = n6952 | n6955 ;
  assign n67842 = ~n6834 ;
  assign n6957 = n67842 & n6956 ;
  assign n67843 = ~n6824 ;
  assign n6958 = x74 & n67843 ;
  assign n67844 = ~n6819 ;
  assign n6959 = n67844 & n6958 ;
  assign n6960 = n6826 | n6959 ;
  assign n6962 = n6957 | n6960 ;
  assign n67845 = ~n6826 ;
  assign n6963 = n67845 & n6962 ;
  assign n67846 = ~n6816 ;
  assign n6964 = x75 & n67846 ;
  assign n67847 = ~n6811 ;
  assign n6965 = n67847 & n6964 ;
  assign n6966 = n6818 | n6965 ;
  assign n6967 = n6963 | n6966 ;
  assign n67848 = ~n6818 ;
  assign n6968 = n67848 & n6967 ;
  assign n67849 = ~n6808 ;
  assign n6969 = x76 & n67849 ;
  assign n67850 = ~n6803 ;
  assign n6970 = n67850 & n6969 ;
  assign n6971 = n6810 | n6970 ;
  assign n6973 = n6968 | n6971 ;
  assign n67851 = ~n6810 ;
  assign n6974 = n67851 & n6973 ;
  assign n67852 = ~n6800 ;
  assign n6975 = x77 & n67852 ;
  assign n67853 = ~n6795 ;
  assign n6976 = n67853 & n6975 ;
  assign n6977 = n6802 | n6976 ;
  assign n6978 = n6974 | n6977 ;
  assign n67854 = ~n6802 ;
  assign n6979 = n67854 & n6978 ;
  assign n67855 = ~n6792 ;
  assign n6980 = x78 & n67855 ;
  assign n67856 = ~n6787 ;
  assign n6981 = n67856 & n6980 ;
  assign n6982 = n6794 | n6981 ;
  assign n6984 = n6979 | n6982 ;
  assign n67857 = ~n6794 ;
  assign n6985 = n67857 & n6984 ;
  assign n67858 = ~n6784 ;
  assign n6986 = x79 & n67858 ;
  assign n67859 = ~n6779 ;
  assign n6987 = n67859 & n6986 ;
  assign n6988 = n6786 | n6987 ;
  assign n6989 = n6985 | n6988 ;
  assign n67860 = ~n6786 ;
  assign n6990 = n67860 & n6989 ;
  assign n67861 = ~n6776 ;
  assign n6991 = x80 & n67861 ;
  assign n67862 = ~n6771 ;
  assign n6992 = n67862 & n6991 ;
  assign n6993 = n6778 | n6992 ;
  assign n6995 = n6990 | n6993 ;
  assign n67863 = ~n6778 ;
  assign n6996 = n67863 & n6995 ;
  assign n67864 = ~n6768 ;
  assign n6997 = x81 & n67864 ;
  assign n67865 = ~n6763 ;
  assign n6998 = n67865 & n6997 ;
  assign n6999 = n6770 | n6998 ;
  assign n7000 = n6996 | n6999 ;
  assign n67866 = ~n6770 ;
  assign n7001 = n67866 & n7000 ;
  assign n67867 = ~n6760 ;
  assign n7002 = x82 & n67867 ;
  assign n67868 = ~n6755 ;
  assign n7003 = n67868 & n7002 ;
  assign n7004 = n6762 | n7003 ;
  assign n7006 = n7001 | n7004 ;
  assign n67869 = ~n6762 ;
  assign n7007 = n67869 & n7006 ;
  assign n67870 = ~n6752 ;
  assign n7008 = x83 & n67870 ;
  assign n67871 = ~n6747 ;
  assign n7009 = n67871 & n7008 ;
  assign n7010 = n6754 | n7009 ;
  assign n7011 = n7007 | n7010 ;
  assign n67872 = ~n6754 ;
  assign n7012 = n67872 & n7011 ;
  assign n67873 = ~n6744 ;
  assign n7013 = x84 & n67873 ;
  assign n67874 = ~n6739 ;
  assign n7014 = n67874 & n7013 ;
  assign n7015 = n6746 | n7014 ;
  assign n7017 = n7012 | n7015 ;
  assign n67875 = ~n6746 ;
  assign n7018 = n67875 & n7017 ;
  assign n67876 = ~n6736 ;
  assign n7019 = x85 & n67876 ;
  assign n67877 = ~n6731 ;
  assign n7020 = n67877 & n7019 ;
  assign n7021 = n6738 | n7020 ;
  assign n7022 = n7018 | n7021 ;
  assign n67878 = ~n6738 ;
  assign n7023 = n67878 & n7022 ;
  assign n67879 = ~n6728 ;
  assign n7024 = x86 & n67879 ;
  assign n67880 = ~n6723 ;
  assign n7025 = n67880 & n7024 ;
  assign n7026 = n6730 | n7025 ;
  assign n7028 = n7023 | n7026 ;
  assign n67881 = ~n6730 ;
  assign n7029 = n67881 & n7028 ;
  assign n67882 = ~n6720 ;
  assign n7030 = x87 & n67882 ;
  assign n67883 = ~n6715 ;
  assign n7031 = n67883 & n7030 ;
  assign n7032 = n6722 | n7031 ;
  assign n7033 = n7029 | n7032 ;
  assign n67884 = ~n6722 ;
  assign n7034 = n67884 & n7033 ;
  assign n67885 = ~n6712 ;
  assign n7035 = x88 & n67885 ;
  assign n67886 = ~n6707 ;
  assign n7036 = n67886 & n7035 ;
  assign n7037 = n6714 | n7036 ;
  assign n7039 = n7034 | n7037 ;
  assign n67887 = ~n6714 ;
  assign n7040 = n67887 & n7039 ;
  assign n67888 = ~n6704 ;
  assign n7041 = x89 & n67888 ;
  assign n67889 = ~n6699 ;
  assign n7042 = n67889 & n7041 ;
  assign n7043 = n6706 | n7042 ;
  assign n7044 = n7040 | n7043 ;
  assign n67890 = ~n6706 ;
  assign n7045 = n67890 & n7044 ;
  assign n67891 = ~n6696 ;
  assign n7046 = x90 & n67891 ;
  assign n67892 = ~n6691 ;
  assign n7047 = n67892 & n7046 ;
  assign n7048 = n6698 | n7047 ;
  assign n7050 = n7045 | n7048 ;
  assign n67893 = ~n6698 ;
  assign n7051 = n67893 & n7050 ;
  assign n67894 = ~n6688 ;
  assign n7052 = x91 & n67894 ;
  assign n67895 = ~n6683 ;
  assign n7053 = n67895 & n7052 ;
  assign n7054 = n6690 | n7053 ;
  assign n7055 = n7051 | n7054 ;
  assign n67896 = ~n6690 ;
  assign n7056 = n67896 & n7055 ;
  assign n165 = ~n6616 ;
  assign n7057 = n165 & n6679 ;
  assign n7058 = n6245 & n6616 ;
  assign n67898 = ~n7058 ;
  assign n7059 = x92 & n67898 ;
  assign n67899 = ~n7057 ;
  assign n7060 = n67899 & n7059 ;
  assign n7061 = n6682 | n7060 ;
  assign n7063 = n7056 | n7061 ;
  assign n67900 = ~n6682 ;
  assign n7064 = n67900 & n7063 ;
  assign n7065 = n458 | n468 ;
  assign n7066 = n465 | n7065 ;
  assign n7067 = n7064 | n7066 ;
  assign n7068 = n6689 & n7067 ;
  assign n6903 = n65670 & n6901 ;
  assign n7069 = x65 & n6912 ;
  assign n67901 = ~n7069 ;
  assign n7070 = n6905 & n67901 ;
  assign n7071 = n6907 | n7070 ;
  assign n67902 = ~n6903 ;
  assign n7072 = n67902 & n7071 ;
  assign n7073 = n6918 | n7072 ;
  assign n7074 = n67821 & n7073 ;
  assign n7075 = n6922 | n7074 ;
  assign n7077 = n67824 & n7075 ;
  assign n7079 = n6928 | n7077 ;
  assign n7080 = n67827 & n7079 ;
  assign n7082 = n6933 | n7080 ;
  assign n7083 = n67830 & n7082 ;
  assign n7084 = n6938 | n7083 ;
  assign n7085 = n67833 & n7084 ;
  assign n7086 = n6944 | n7085 ;
  assign n7088 = n67836 & n7086 ;
  assign n7089 = n6949 | n7088 ;
  assign n7090 = n67839 & n7089 ;
  assign n7091 = n6955 | n7090 ;
  assign n7093 = n67842 & n7091 ;
  assign n7094 = n6960 | n7093 ;
  assign n7095 = n67845 & n7094 ;
  assign n7096 = n6966 | n7095 ;
  assign n7098 = n67848 & n7096 ;
  assign n7099 = n6971 | n7098 ;
  assign n7100 = n67851 & n7099 ;
  assign n7101 = n6977 | n7100 ;
  assign n7103 = n67854 & n7101 ;
  assign n7104 = n6982 | n7103 ;
  assign n7105 = n67857 & n7104 ;
  assign n7106 = n6988 | n7105 ;
  assign n7108 = n67860 & n7106 ;
  assign n7109 = n6993 | n7108 ;
  assign n7110 = n67863 & n7109 ;
  assign n7111 = n6999 | n7110 ;
  assign n7113 = n67866 & n7111 ;
  assign n7114 = n7004 | n7113 ;
  assign n7115 = n67869 & n7114 ;
  assign n7116 = n7010 | n7115 ;
  assign n7118 = n67872 & n7116 ;
  assign n7119 = n7015 | n7118 ;
  assign n7120 = n67875 & n7119 ;
  assign n7121 = n7021 | n7120 ;
  assign n7123 = n67878 & n7121 ;
  assign n7124 = n7026 | n7123 ;
  assign n7125 = n67881 & n7124 ;
  assign n7126 = n7032 | n7125 ;
  assign n7128 = n67884 & n7126 ;
  assign n7129 = n7037 | n7128 ;
  assign n7130 = n67887 & n7129 ;
  assign n7131 = n7043 | n7130 ;
  assign n7133 = n67890 & n7131 ;
  assign n7134 = n7048 | n7133 ;
  assign n7135 = n67893 & n7134 ;
  assign n67903 = ~n7135 ;
  assign n7136 = n7054 & n67903 ;
  assign n7138 = n6698 | n7054 ;
  assign n67904 = ~n7138 ;
  assign n7139 = n7050 & n67904 ;
  assign n7140 = n7136 | n7139 ;
  assign n67905 = ~n7066 ;
  assign n7141 = n67905 & n7140 ;
  assign n67906 = ~n7064 ;
  assign n7142 = n67906 & n7141 ;
  assign n7143 = n7068 | n7142 ;
  assign n7144 = n67763 & n7143 ;
  assign n67907 = ~n7142 ;
  assign n7508 = x92 & n67907 ;
  assign n67908 = ~n7068 ;
  assign n7509 = n67908 & n7508 ;
  assign n7510 = n7144 | n7509 ;
  assign n7145 = n6697 & n7067 ;
  assign n67909 = ~n7045 ;
  assign n7049 = n67909 & n7048 ;
  assign n7146 = n6706 | n7048 ;
  assign n67910 = ~n7146 ;
  assign n7147 = n7131 & n67910 ;
  assign n7148 = n7049 | n7147 ;
  assign n7149 = n67905 & n7148 ;
  assign n7150 = n67906 & n7149 ;
  assign n7151 = n7145 | n7150 ;
  assign n7152 = n67622 & n7151 ;
  assign n7153 = n6705 & n7067 ;
  assign n67911 = ~n7130 ;
  assign n7132 = n7043 & n67911 ;
  assign n7154 = n6714 | n7043 ;
  assign n67912 = ~n7154 ;
  assign n7155 = n7039 & n67912 ;
  assign n7156 = n7132 | n7155 ;
  assign n7157 = n67905 & n7156 ;
  assign n7158 = n67906 & n7157 ;
  assign n7159 = n7153 | n7158 ;
  assign n7160 = n67531 & n7159 ;
  assign n67913 = ~n7158 ;
  assign n7498 = x90 & n67913 ;
  assign n67914 = ~n7153 ;
  assign n7499 = n67914 & n7498 ;
  assign n7500 = n7160 | n7499 ;
  assign n7161 = n6713 & n7067 ;
  assign n67915 = ~n7034 ;
  assign n7038 = n67915 & n7037 ;
  assign n7162 = n6722 | n7037 ;
  assign n67916 = ~n7162 ;
  assign n7163 = n7126 & n67916 ;
  assign n7164 = n7038 | n7163 ;
  assign n7165 = n67905 & n7164 ;
  assign n7166 = n67906 & n7165 ;
  assign n7167 = n7161 | n7166 ;
  assign n7168 = n67348 & n7167 ;
  assign n7169 = n6721 & n7067 ;
  assign n67917 = ~n7125 ;
  assign n7127 = n7032 & n67917 ;
  assign n7170 = n6730 | n7032 ;
  assign n67918 = ~n7170 ;
  assign n7171 = n7028 & n67918 ;
  assign n7172 = n7127 | n7171 ;
  assign n7173 = n67905 & n7172 ;
  assign n7174 = n67906 & n7173 ;
  assign n7175 = n7169 | n7174 ;
  assign n7176 = n67222 & n7175 ;
  assign n67919 = ~n7174 ;
  assign n7488 = x88 & n67919 ;
  assign n67920 = ~n7169 ;
  assign n7489 = n67920 & n7488 ;
  assign n7490 = n7176 | n7489 ;
  assign n7177 = n6729 & n7067 ;
  assign n67921 = ~n7023 ;
  assign n7027 = n67921 & n7026 ;
  assign n7178 = n6738 | n7026 ;
  assign n67922 = ~n7178 ;
  assign n7179 = n7121 & n67922 ;
  assign n7180 = n7027 | n7179 ;
  assign n7181 = n67905 & n7180 ;
  assign n7182 = n67906 & n7181 ;
  assign n7183 = n7177 | n7182 ;
  assign n7184 = n67164 & n7183 ;
  assign n7185 = n6737 & n7067 ;
  assign n67923 = ~n7120 ;
  assign n7122 = n7021 & n67923 ;
  assign n7186 = n6746 | n7021 ;
  assign n67924 = ~n7186 ;
  assign n7187 = n7017 & n67924 ;
  assign n7188 = n7122 | n7187 ;
  assign n7189 = n67905 & n7188 ;
  assign n7190 = n67906 & n7189 ;
  assign n7191 = n7185 | n7190 ;
  assign n7192 = n66979 & n7191 ;
  assign n67925 = ~n7190 ;
  assign n7478 = x86 & n67925 ;
  assign n67926 = ~n7185 ;
  assign n7479 = n67926 & n7478 ;
  assign n7480 = n7192 | n7479 ;
  assign n7193 = n6745 & n7067 ;
  assign n67927 = ~n7012 ;
  assign n7016 = n67927 & n7015 ;
  assign n7194 = n6754 | n7015 ;
  assign n67928 = ~n7194 ;
  assign n7195 = n7116 & n67928 ;
  assign n7196 = n7016 | n7195 ;
  assign n7197 = n67905 & n7196 ;
  assign n7198 = n67906 & n7197 ;
  assign n7199 = n7193 | n7198 ;
  assign n7200 = n66868 & n7199 ;
  assign n7201 = n6753 & n7067 ;
  assign n67929 = ~n7115 ;
  assign n7117 = n7010 & n67929 ;
  assign n7202 = n6762 | n7010 ;
  assign n67930 = ~n7202 ;
  assign n7203 = n7006 & n67930 ;
  assign n7204 = n7117 | n7203 ;
  assign n7205 = n67905 & n7204 ;
  assign n7206 = n67906 & n7205 ;
  assign n7207 = n7201 | n7206 ;
  assign n7208 = n66797 & n7207 ;
  assign n67931 = ~n7206 ;
  assign n7468 = x84 & n67931 ;
  assign n67932 = ~n7201 ;
  assign n7469 = n67932 & n7468 ;
  assign n7470 = n7208 | n7469 ;
  assign n7209 = n6761 & n7067 ;
  assign n67933 = ~n7001 ;
  assign n7005 = n67933 & n7004 ;
  assign n7210 = n6770 | n7004 ;
  assign n67934 = ~n7210 ;
  assign n7211 = n7111 & n67934 ;
  assign n7212 = n7005 | n7211 ;
  assign n7213 = n67905 & n7212 ;
  assign n7214 = n67906 & n7213 ;
  assign n7215 = n7209 | n7214 ;
  assign n7216 = n66654 & n7215 ;
  assign n7217 = n6769 & n7067 ;
  assign n67935 = ~n7110 ;
  assign n7112 = n6999 & n67935 ;
  assign n7218 = n6778 | n6999 ;
  assign n67936 = ~n7218 ;
  assign n7219 = n6995 & n67936 ;
  assign n7220 = n7112 | n7219 ;
  assign n7221 = n67905 & n7220 ;
  assign n7222 = n67906 & n7221 ;
  assign n7223 = n7217 | n7222 ;
  assign n7224 = n66560 & n7223 ;
  assign n67937 = ~n7222 ;
  assign n7458 = x82 & n67937 ;
  assign n67938 = ~n7217 ;
  assign n7459 = n67938 & n7458 ;
  assign n7460 = n7224 | n7459 ;
  assign n7225 = n6777 & n7067 ;
  assign n67939 = ~n6990 ;
  assign n6994 = n67939 & n6993 ;
  assign n7226 = n6786 | n6993 ;
  assign n67940 = ~n7226 ;
  assign n7227 = n7106 & n67940 ;
  assign n7228 = n6994 | n7227 ;
  assign n7229 = n67905 & n7228 ;
  assign n7230 = n67906 & n7229 ;
  assign n7231 = n7225 | n7230 ;
  assign n7232 = n66505 & n7231 ;
  assign n7233 = n6785 & n7067 ;
  assign n67941 = ~n7105 ;
  assign n7107 = n6988 & n67941 ;
  assign n7234 = n6794 | n6988 ;
  assign n67942 = ~n7234 ;
  assign n7235 = n6984 & n67942 ;
  assign n7236 = n7107 | n7235 ;
  assign n7237 = n67905 & n7236 ;
  assign n7238 = n67906 & n7237 ;
  assign n7239 = n7233 | n7238 ;
  assign n7240 = n66379 & n7239 ;
  assign n67943 = ~n7238 ;
  assign n7448 = x80 & n67943 ;
  assign n67944 = ~n7233 ;
  assign n7449 = n67944 & n7448 ;
  assign n7450 = n7240 | n7449 ;
  assign n7241 = n6793 & n7067 ;
  assign n67945 = ~n6979 ;
  assign n6983 = n67945 & n6982 ;
  assign n7242 = n6802 | n6982 ;
  assign n67946 = ~n7242 ;
  assign n7243 = n7101 & n67946 ;
  assign n7244 = n6983 | n7243 ;
  assign n7245 = n67905 & n7244 ;
  assign n7246 = n67906 & n7245 ;
  assign n7247 = n7241 | n7246 ;
  assign n7248 = n66299 & n7247 ;
  assign n7249 = n6801 & n7067 ;
  assign n67947 = ~n7100 ;
  assign n7102 = n6977 & n67947 ;
  assign n7250 = n6810 | n6977 ;
  assign n67948 = ~n7250 ;
  assign n7251 = n6973 & n67948 ;
  assign n7252 = n7102 | n7251 ;
  assign n7253 = n67905 & n7252 ;
  assign n7254 = n67906 & n7253 ;
  assign n7255 = n7249 | n7254 ;
  assign n7256 = n66244 & n7255 ;
  assign n67949 = ~n7254 ;
  assign n7437 = x78 & n67949 ;
  assign n67950 = ~n7249 ;
  assign n7438 = n67950 & n7437 ;
  assign n7439 = n7256 | n7438 ;
  assign n7257 = n6809 & n7067 ;
  assign n67951 = ~n6968 ;
  assign n6972 = n67951 & n6971 ;
  assign n7258 = n6818 | n6971 ;
  assign n67952 = ~n7258 ;
  assign n7259 = n7096 & n67952 ;
  assign n7260 = n6972 | n7259 ;
  assign n7261 = n67905 & n7260 ;
  assign n7262 = n67906 & n7261 ;
  assign n7263 = n7257 | n7262 ;
  assign n7264 = n66145 & n7263 ;
  assign n7265 = n6817 & n7067 ;
  assign n67953 = ~n7095 ;
  assign n7097 = n6966 & n67953 ;
  assign n7266 = n6826 | n6966 ;
  assign n67954 = ~n7266 ;
  assign n7267 = n6962 & n67954 ;
  assign n7268 = n7097 | n7267 ;
  assign n7269 = n67905 & n7268 ;
  assign n7270 = n67906 & n7269 ;
  assign n7271 = n7265 | n7270 ;
  assign n7272 = n66081 & n7271 ;
  assign n67955 = ~n7270 ;
  assign n7427 = x76 & n67955 ;
  assign n67956 = ~n7265 ;
  assign n7428 = n67956 & n7427 ;
  assign n7429 = n7272 | n7428 ;
  assign n7273 = n6825 & n7067 ;
  assign n67957 = ~n6957 ;
  assign n6961 = n67957 & n6960 ;
  assign n7274 = n6834 | n6960 ;
  assign n67958 = ~n7274 ;
  assign n7275 = n7091 & n67958 ;
  assign n7276 = n6961 | n7275 ;
  assign n7277 = n67905 & n7276 ;
  assign n7278 = n67906 & n7277 ;
  assign n7279 = n7273 | n7278 ;
  assign n7280 = n66043 & n7279 ;
  assign n7281 = n6833 & n7067 ;
  assign n67959 = ~n7090 ;
  assign n7092 = n6955 & n67959 ;
  assign n7282 = n6842 | n6955 ;
  assign n67960 = ~n7282 ;
  assign n7283 = n6951 & n67960 ;
  assign n7284 = n7092 | n7283 ;
  assign n7285 = n67905 & n7284 ;
  assign n7286 = n67906 & n7285 ;
  assign n7287 = n7281 | n7286 ;
  assign n7288 = n65960 & n7287 ;
  assign n67961 = ~n7286 ;
  assign n7417 = x74 & n67961 ;
  assign n67962 = ~n7281 ;
  assign n7418 = n67962 & n7417 ;
  assign n7419 = n7288 | n7418 ;
  assign n7289 = n6841 & n7067 ;
  assign n67963 = ~n6946 ;
  assign n6950 = n67963 & n6949 ;
  assign n7290 = n6850 | n6949 ;
  assign n67964 = ~n7290 ;
  assign n7291 = n7086 & n67964 ;
  assign n7292 = n6950 | n7291 ;
  assign n7293 = n67905 & n7292 ;
  assign n7294 = n67906 & n7293 ;
  assign n7295 = n7289 | n7294 ;
  assign n7296 = n65909 & n7295 ;
  assign n7297 = n6849 & n7067 ;
  assign n67965 = ~n7085 ;
  assign n7087 = n6944 & n67965 ;
  assign n7298 = n6858 | n6944 ;
  assign n67966 = ~n7298 ;
  assign n7299 = n6940 & n67966 ;
  assign n7300 = n7087 | n7299 ;
  assign n7301 = n67905 & n7300 ;
  assign n7302 = n67906 & n7301 ;
  assign n7303 = n7297 | n7302 ;
  assign n7304 = n65877 & n7303 ;
  assign n67967 = ~n7302 ;
  assign n7407 = x72 & n67967 ;
  assign n67968 = ~n7297 ;
  assign n7408 = n67968 & n7407 ;
  assign n7409 = n7304 | n7408 ;
  assign n7305 = n6857 & n7067 ;
  assign n67969 = ~n6935 ;
  assign n6939 = n67969 & n6938 ;
  assign n7306 = n6867 | n6938 ;
  assign n67970 = ~n7306 ;
  assign n7307 = n7082 & n67970 ;
  assign n7308 = n6939 | n7307 ;
  assign n7309 = n67905 & n7308 ;
  assign n7310 = n67906 & n7309 ;
  assign n7311 = n7305 | n7310 ;
  assign n7312 = n65820 & n7311 ;
  assign n7313 = n6866 & n7067 ;
  assign n67971 = ~n7080 ;
  assign n7081 = n6933 & n67971 ;
  assign n7314 = n6876 | n6933 ;
  assign n67972 = ~n7314 ;
  assign n7315 = n7079 & n67972 ;
  assign n7316 = n7081 | n7315 ;
  assign n7317 = n67905 & n7316 ;
  assign n7318 = n67906 & n7317 ;
  assign n7319 = n7313 | n7318 ;
  assign n7320 = n65791 & n7319 ;
  assign n67973 = ~n7318 ;
  assign n7397 = x70 & n67973 ;
  assign n67974 = ~n7313 ;
  assign n7398 = n67974 & n7397 ;
  assign n7399 = n7320 | n7398 ;
  assign n7321 = n6875 & n7067 ;
  assign n67975 = ~n6925 ;
  assign n7078 = n67975 & n6928 ;
  assign n7322 = n6923 | n7074 ;
  assign n7323 = n6884 | n6928 ;
  assign n67976 = ~n7323 ;
  assign n7324 = n7322 & n67976 ;
  assign n7325 = n7078 | n7324 ;
  assign n7326 = n67905 & n7325 ;
  assign n7327 = n67906 & n7326 ;
  assign n7328 = n7321 | n7327 ;
  assign n7329 = n65772 & n7328 ;
  assign n7330 = n6883 & n7067 ;
  assign n67977 = ~n7074 ;
  assign n7076 = n6923 & n67977 ;
  assign n7331 = n6890 | n6923 ;
  assign n67978 = ~n7331 ;
  assign n7332 = n7073 & n67978 ;
  assign n7333 = n7076 | n7332 ;
  assign n7334 = n67905 & n7333 ;
  assign n7335 = n67906 & n7334 ;
  assign n7336 = n7330 | n7335 ;
  assign n7337 = n65746 & n7336 ;
  assign n67979 = ~n7335 ;
  assign n7387 = x68 & n67979 ;
  assign n67980 = ~n7330 ;
  assign n7388 = n67980 & n7387 ;
  assign n7389 = n7337 | n7388 ;
  assign n7338 = n6889 & n7067 ;
  assign n7339 = n6913 | n6918 ;
  assign n67981 = ~n7339 ;
  assign n7340 = n7071 & n67981 ;
  assign n67982 = ~n6915 ;
  assign n7341 = n67982 & n6918 ;
  assign n7342 = n7340 | n7341 ;
  assign n7343 = n67905 & n7342 ;
  assign n7344 = n67906 & n7343 ;
  assign n7345 = n7338 | n7344 ;
  assign n7347 = n65721 & n7345 ;
  assign n7348 = n6901 & n7067 ;
  assign n7349 = n6905 & n6907 ;
  assign n7350 = n67901 & n7349 ;
  assign n7351 = n7066 | n7350 ;
  assign n67983 = ~n7351 ;
  assign n7352 = n7071 & n67983 ;
  assign n7353 = n67906 & n7352 ;
  assign n7354 = n7348 | n7353 ;
  assign n7355 = n65686 & n7354 ;
  assign n67984 = ~n7353 ;
  assign n7378 = x66 & n67984 ;
  assign n67985 = ~n7348 ;
  assign n7379 = n67985 & n7378 ;
  assign n7380 = n7355 | n7379 ;
  assign n7137 = n7054 | n7135 ;
  assign n7356 = n67896 & n7137 ;
  assign n7357 = n7061 | n7356 ;
  assign n7358 = n67900 & n7357 ;
  assign n67986 = ~x93 ;
  assign n7359 = x64 & n67986 ;
  assign n67987 = ~n65632 ;
  assign n7360 = n67987 & n7359 ;
  assign n67988 = ~n65617 ;
  assign n7361 = n67988 & n7360 ;
  assign n7362 = n67020 & n7361 ;
  assign n7363 = n67021 & n7362 ;
  assign n67989 = ~n7358 ;
  assign n7364 = n67989 & n7363 ;
  assign n67990 = ~n7364 ;
  assign n7365 = x35 & n67990 ;
  assign n7366 = n67533 & n6907 ;
  assign n7367 = n66714 & n7366 ;
  assign n7368 = n66715 & n7367 ;
  assign n7369 = n67906 & n7368 ;
  assign n7370 = n7365 | n7369 ;
  assign n7371 = x65 & n7370 ;
  assign n7372 = x65 | n7369 ;
  assign n7373 = n7365 | n7372 ;
  assign n67991 = ~n7371 ;
  assign n7374 = n67991 & n7373 ;
  assign n67992 = ~x34 ;
  assign n7375 = n67992 & x64 ;
  assign n7376 = n7374 | n7375 ;
  assign n7377 = n65670 & n7370 ;
  assign n67993 = ~n7377 ;
  assign n7381 = n7376 & n67993 ;
  assign n7382 = n7380 | n7381 ;
  assign n67994 = ~n7355 ;
  assign n7383 = n67994 & n7382 ;
  assign n67995 = ~n7344 ;
  assign n7346 = x67 & n67995 ;
  assign n67996 = ~n7338 ;
  assign n7384 = n67996 & n7346 ;
  assign n7385 = n7347 | n7384 ;
  assign n7386 = n7383 | n7385 ;
  assign n67997 = ~n7347 ;
  assign n7390 = n67997 & n7386 ;
  assign n7391 = n7389 | n7390 ;
  assign n67998 = ~n7337 ;
  assign n7392 = n67998 & n7391 ;
  assign n67999 = ~n7327 ;
  assign n7393 = x69 & n67999 ;
  assign n68000 = ~n7321 ;
  assign n7394 = n68000 & n7393 ;
  assign n7395 = n7329 | n7394 ;
  assign n7396 = n7392 | n7395 ;
  assign n68001 = ~n7329 ;
  assign n7400 = n68001 & n7396 ;
  assign n7401 = n7399 | n7400 ;
  assign n68002 = ~n7320 ;
  assign n7402 = n68002 & n7401 ;
  assign n68003 = ~n7310 ;
  assign n7403 = x71 & n68003 ;
  assign n68004 = ~n7305 ;
  assign n7404 = n68004 & n7403 ;
  assign n7405 = n7312 | n7404 ;
  assign n7406 = n7402 | n7405 ;
  assign n68005 = ~n7312 ;
  assign n7410 = n68005 & n7406 ;
  assign n7411 = n7409 | n7410 ;
  assign n68006 = ~n7304 ;
  assign n7412 = n68006 & n7411 ;
  assign n68007 = ~n7294 ;
  assign n7413 = x73 & n68007 ;
  assign n68008 = ~n7289 ;
  assign n7414 = n68008 & n7413 ;
  assign n7415 = n7296 | n7414 ;
  assign n7416 = n7412 | n7415 ;
  assign n68009 = ~n7296 ;
  assign n7420 = n68009 & n7416 ;
  assign n7421 = n7419 | n7420 ;
  assign n68010 = ~n7288 ;
  assign n7422 = n68010 & n7421 ;
  assign n68011 = ~n7278 ;
  assign n7423 = x75 & n68011 ;
  assign n68012 = ~n7273 ;
  assign n7424 = n68012 & n7423 ;
  assign n7425 = n7280 | n7424 ;
  assign n7426 = n7422 | n7425 ;
  assign n68013 = ~n7280 ;
  assign n7430 = n68013 & n7426 ;
  assign n7431 = n7429 | n7430 ;
  assign n68014 = ~n7272 ;
  assign n7432 = n68014 & n7431 ;
  assign n68015 = ~n7262 ;
  assign n7433 = x77 & n68015 ;
  assign n68016 = ~n7257 ;
  assign n7434 = n68016 & n7433 ;
  assign n7435 = n7264 | n7434 ;
  assign n7436 = n7432 | n7435 ;
  assign n68017 = ~n7264 ;
  assign n7441 = n68017 & n7436 ;
  assign n7442 = n7439 | n7441 ;
  assign n68018 = ~n7256 ;
  assign n7443 = n68018 & n7442 ;
  assign n68019 = ~n7246 ;
  assign n7444 = x79 & n68019 ;
  assign n68020 = ~n7241 ;
  assign n7445 = n68020 & n7444 ;
  assign n7446 = n7248 | n7445 ;
  assign n7447 = n7443 | n7446 ;
  assign n68021 = ~n7248 ;
  assign n7451 = n68021 & n7447 ;
  assign n7452 = n7450 | n7451 ;
  assign n68022 = ~n7240 ;
  assign n7453 = n68022 & n7452 ;
  assign n68023 = ~n7230 ;
  assign n7454 = x81 & n68023 ;
  assign n68024 = ~n7225 ;
  assign n7455 = n68024 & n7454 ;
  assign n7456 = n7232 | n7455 ;
  assign n7457 = n7453 | n7456 ;
  assign n68025 = ~n7232 ;
  assign n7461 = n68025 & n7457 ;
  assign n7462 = n7460 | n7461 ;
  assign n68026 = ~n7224 ;
  assign n7463 = n68026 & n7462 ;
  assign n68027 = ~n7214 ;
  assign n7464 = x83 & n68027 ;
  assign n68028 = ~n7209 ;
  assign n7465 = n68028 & n7464 ;
  assign n7466 = n7216 | n7465 ;
  assign n7467 = n7463 | n7466 ;
  assign n68029 = ~n7216 ;
  assign n7471 = n68029 & n7467 ;
  assign n7472 = n7470 | n7471 ;
  assign n68030 = ~n7208 ;
  assign n7473 = n68030 & n7472 ;
  assign n68031 = ~n7198 ;
  assign n7474 = x85 & n68031 ;
  assign n68032 = ~n7193 ;
  assign n7475 = n68032 & n7474 ;
  assign n7476 = n7200 | n7475 ;
  assign n7477 = n7473 | n7476 ;
  assign n68033 = ~n7200 ;
  assign n7481 = n68033 & n7477 ;
  assign n7482 = n7480 | n7481 ;
  assign n68034 = ~n7192 ;
  assign n7483 = n68034 & n7482 ;
  assign n68035 = ~n7182 ;
  assign n7484 = x87 & n68035 ;
  assign n68036 = ~n7177 ;
  assign n7485 = n68036 & n7484 ;
  assign n7486 = n7184 | n7485 ;
  assign n7487 = n7483 | n7486 ;
  assign n68037 = ~n7184 ;
  assign n7491 = n68037 & n7487 ;
  assign n7492 = n7490 | n7491 ;
  assign n68038 = ~n7176 ;
  assign n7493 = n68038 & n7492 ;
  assign n68039 = ~n7166 ;
  assign n7494 = x89 & n68039 ;
  assign n68040 = ~n7161 ;
  assign n7495 = n68040 & n7494 ;
  assign n7496 = n7168 | n7495 ;
  assign n7497 = n7493 | n7496 ;
  assign n68041 = ~n7168 ;
  assign n7501 = n68041 & n7497 ;
  assign n7502 = n7500 | n7501 ;
  assign n68042 = ~n7160 ;
  assign n7503 = n68042 & n7502 ;
  assign n68043 = ~n7150 ;
  assign n7504 = x91 & n68043 ;
  assign n68044 = ~n7145 ;
  assign n7505 = n68044 & n7504 ;
  assign n7506 = n7152 | n7505 ;
  assign n7507 = n7503 | n7506 ;
  assign n68045 = ~n7152 ;
  assign n7511 = n68045 & n7507 ;
  assign n7512 = n7510 | n7511 ;
  assign n68046 = ~n7144 ;
  assign n7513 = n68046 & n7512 ;
  assign n68047 = ~n7056 ;
  assign n7062 = n68047 & n7061 ;
  assign n7514 = n6690 | n7061 ;
  assign n68048 = ~n7514 ;
  assign n7515 = n7137 & n68048 ;
  assign n7516 = n7062 | n7515 ;
  assign n7517 = n7067 | n7516 ;
  assign n68049 = ~n6681 ;
  assign n7518 = n68049 & n7067 ;
  assign n68050 = ~n7518 ;
  assign n7519 = n7517 & n68050 ;
  assign n7520 = n67986 & n7519 ;
  assign n164 = ~n7067 ;
  assign n7521 = n164 & n7516 ;
  assign n7522 = n6681 & n7067 ;
  assign n68052 = ~n7522 ;
  assign n7523 = x93 & n68052 ;
  assign n68053 = ~n7521 ;
  assign n7524 = n68053 & n7523 ;
  assign n7525 = n65617 | n65632 ;
  assign n7526 = n65542 | n7525 ;
  assign n7527 = n65429 | n7526 ;
  assign n7528 = n7524 | n7527 ;
  assign n7529 = n7520 | n7528 ;
  assign n7530 = n7513 | n7529 ;
  assign n7531 = n67905 & n7519 ;
  assign n68054 = ~n7531 ;
  assign n7532 = n7530 & n68054 ;
  assign n7534 = n7144 | n7524 ;
  assign n7535 = n7520 | n7534 ;
  assign n68055 = ~n7535 ;
  assign n7536 = n7512 & n68055 ;
  assign n7537 = n7520 | n7524 ;
  assign n68056 = ~n7513 ;
  assign n7538 = n68056 & n7537 ;
  assign n7539 = n7536 | n7538 ;
  assign n163 = ~n7532 ;
  assign n7540 = n163 & n7539 ;
  assign n7541 = n7066 & n7519 ;
  assign n7542 = n7530 & n7541 ;
  assign n7543 = n7540 | n7542 ;
  assign n68058 = ~x94 ;
  assign n7544 = n68058 & n7543 ;
  assign n68059 = ~n7511 ;
  assign n7604 = n7510 & n68059 ;
  assign n7545 = n67906 & n7363 ;
  assign n68060 = ~n7545 ;
  assign n7546 = x35 & n68060 ;
  assign n7547 = n7369 | n7546 ;
  assign n7548 = x65 & n7547 ;
  assign n68061 = ~n7548 ;
  assign n7549 = n7373 & n68061 ;
  assign n7550 = n7375 | n7549 ;
  assign n7551 = n67993 & n7550 ;
  assign n7552 = n7380 | n7551 ;
  assign n7553 = n67994 & n7552 ;
  assign n7554 = n7385 | n7553 ;
  assign n7555 = n67997 & n7554 ;
  assign n7556 = n7389 | n7555 ;
  assign n7557 = n67998 & n7556 ;
  assign n7558 = n7395 | n7557 ;
  assign n7559 = n68001 & n7558 ;
  assign n7560 = n7399 | n7559 ;
  assign n7561 = n68002 & n7560 ;
  assign n7562 = n7405 | n7561 ;
  assign n7563 = n68005 & n7562 ;
  assign n7564 = n7409 | n7563 ;
  assign n7565 = n68006 & n7564 ;
  assign n7566 = n7415 | n7565 ;
  assign n7567 = n68009 & n7566 ;
  assign n7568 = n7419 | n7567 ;
  assign n7569 = n68010 & n7568 ;
  assign n7570 = n7425 | n7569 ;
  assign n7571 = n68013 & n7570 ;
  assign n7572 = n7429 | n7571 ;
  assign n7573 = n68014 & n7572 ;
  assign n7574 = n7435 | n7573 ;
  assign n7575 = n68017 & n7574 ;
  assign n7576 = n7439 | n7575 ;
  assign n7577 = n68018 & n7576 ;
  assign n7578 = n7446 | n7577 ;
  assign n7579 = n68021 & n7578 ;
  assign n7580 = n7450 | n7579 ;
  assign n7581 = n68022 & n7580 ;
  assign n7582 = n7456 | n7581 ;
  assign n7583 = n68025 & n7582 ;
  assign n7584 = n7460 | n7583 ;
  assign n7585 = n68026 & n7584 ;
  assign n7586 = n7466 | n7585 ;
  assign n7587 = n68029 & n7586 ;
  assign n7588 = n7470 | n7587 ;
  assign n7589 = n68030 & n7588 ;
  assign n7590 = n7476 | n7589 ;
  assign n7591 = n68033 & n7590 ;
  assign n7592 = n7480 | n7591 ;
  assign n7593 = n68034 & n7592 ;
  assign n7594 = n7486 | n7593 ;
  assign n7595 = n68037 & n7594 ;
  assign n7596 = n7490 | n7595 ;
  assign n7597 = n68038 & n7596 ;
  assign n7598 = n7496 | n7597 ;
  assign n7599 = n68041 & n7598 ;
  assign n7600 = n7500 | n7599 ;
  assign n7601 = n68042 & n7600 ;
  assign n7602 = n7506 | n7601 ;
  assign n7605 = n7152 | n7510 ;
  assign n68062 = ~n7605 ;
  assign n7606 = n7602 & n68062 ;
  assign n7607 = n7604 | n7606 ;
  assign n7608 = n163 & n7607 ;
  assign n7609 = n7143 & n68054 ;
  assign n7610 = n7530 & n7609 ;
  assign n7611 = n7608 | n7610 ;
  assign n7612 = n67986 & n7611 ;
  assign n68063 = ~n7601 ;
  assign n7613 = n7506 & n68063 ;
  assign n7614 = n7160 | n7506 ;
  assign n68064 = ~n7614 ;
  assign n7615 = n7502 & n68064 ;
  assign n7616 = n7613 | n7615 ;
  assign n7617 = n163 & n7616 ;
  assign n7618 = n7151 & n68054 ;
  assign n7619 = n7530 & n7618 ;
  assign n7620 = n7617 | n7619 ;
  assign n7621 = n67763 & n7620 ;
  assign n68065 = ~n7501 ;
  assign n7622 = n7500 & n68065 ;
  assign n7623 = n7168 | n7500 ;
  assign n68066 = ~n7623 ;
  assign n7624 = n7598 & n68066 ;
  assign n7625 = n7622 | n7624 ;
  assign n7626 = n163 & n7625 ;
  assign n7627 = n7159 & n68054 ;
  assign n7628 = n7530 & n7627 ;
  assign n7629 = n7626 | n7628 ;
  assign n7630 = n67622 & n7629 ;
  assign n68067 = ~n7597 ;
  assign n7631 = n7496 & n68067 ;
  assign n7632 = n7176 | n7496 ;
  assign n68068 = ~n7632 ;
  assign n7633 = n7492 & n68068 ;
  assign n7634 = n7631 | n7633 ;
  assign n7635 = n163 & n7634 ;
  assign n7636 = n7167 & n68054 ;
  assign n7637 = n7530 & n7636 ;
  assign n7638 = n7635 | n7637 ;
  assign n7639 = n67531 & n7638 ;
  assign n68069 = ~n7491 ;
  assign n7640 = n7490 & n68069 ;
  assign n7641 = n7184 | n7490 ;
  assign n68070 = ~n7641 ;
  assign n7642 = n7594 & n68070 ;
  assign n7643 = n7640 | n7642 ;
  assign n7644 = n163 & n7643 ;
  assign n7645 = n7175 & n68054 ;
  assign n7646 = n7530 & n7645 ;
  assign n7647 = n7644 | n7646 ;
  assign n7648 = n67348 & n7647 ;
  assign n68071 = ~n7593 ;
  assign n7649 = n7486 & n68071 ;
  assign n7650 = n7192 | n7486 ;
  assign n68072 = ~n7650 ;
  assign n7651 = n7482 & n68072 ;
  assign n7652 = n7649 | n7651 ;
  assign n7653 = n163 & n7652 ;
  assign n7654 = n7183 & n68054 ;
  assign n7655 = n7530 & n7654 ;
  assign n7656 = n7653 | n7655 ;
  assign n7657 = n67222 & n7656 ;
  assign n68073 = ~n7481 ;
  assign n7658 = n7480 & n68073 ;
  assign n7659 = n7200 | n7480 ;
  assign n68074 = ~n7659 ;
  assign n7660 = n7590 & n68074 ;
  assign n7661 = n7658 | n7660 ;
  assign n7662 = n163 & n7661 ;
  assign n7663 = n7191 & n68054 ;
  assign n7664 = n7530 & n7663 ;
  assign n7665 = n7662 | n7664 ;
  assign n7666 = n67164 & n7665 ;
  assign n68075 = ~n7589 ;
  assign n7667 = n7476 & n68075 ;
  assign n7668 = n7208 | n7476 ;
  assign n68076 = ~n7668 ;
  assign n7669 = n7472 & n68076 ;
  assign n7670 = n7667 | n7669 ;
  assign n7671 = n163 & n7670 ;
  assign n7672 = n7199 & n68054 ;
  assign n7673 = n7530 & n7672 ;
  assign n7674 = n7671 | n7673 ;
  assign n7675 = n66979 & n7674 ;
  assign n68077 = ~n7471 ;
  assign n7676 = n7470 & n68077 ;
  assign n7677 = n7216 | n7470 ;
  assign n68078 = ~n7677 ;
  assign n7678 = n7586 & n68078 ;
  assign n7679 = n7676 | n7678 ;
  assign n7680 = n163 & n7679 ;
  assign n7681 = n7207 & n68054 ;
  assign n7682 = n7530 & n7681 ;
  assign n7683 = n7680 | n7682 ;
  assign n7684 = n66868 & n7683 ;
  assign n68079 = ~n7585 ;
  assign n7685 = n7466 & n68079 ;
  assign n7686 = n7224 | n7466 ;
  assign n68080 = ~n7686 ;
  assign n7687 = n7462 & n68080 ;
  assign n7688 = n7685 | n7687 ;
  assign n7689 = n163 & n7688 ;
  assign n7690 = n7215 & n68054 ;
  assign n7691 = n7530 & n7690 ;
  assign n7692 = n7689 | n7691 ;
  assign n7693 = n66797 & n7692 ;
  assign n68081 = ~n7461 ;
  assign n7694 = n7460 & n68081 ;
  assign n7695 = n7232 | n7460 ;
  assign n68082 = ~n7695 ;
  assign n7696 = n7582 & n68082 ;
  assign n7697 = n7694 | n7696 ;
  assign n7698 = n163 & n7697 ;
  assign n7699 = n7223 & n68054 ;
  assign n7700 = n7530 & n7699 ;
  assign n7701 = n7698 | n7700 ;
  assign n7702 = n66654 & n7701 ;
  assign n68083 = ~n7581 ;
  assign n7703 = n7456 & n68083 ;
  assign n7704 = n7240 | n7456 ;
  assign n68084 = ~n7704 ;
  assign n7705 = n7452 & n68084 ;
  assign n7706 = n7703 | n7705 ;
  assign n7707 = n163 & n7706 ;
  assign n7708 = n7231 & n68054 ;
  assign n7709 = n7530 & n7708 ;
  assign n7710 = n7707 | n7709 ;
  assign n7711 = n66560 & n7710 ;
  assign n68085 = ~n7451 ;
  assign n7712 = n7450 & n68085 ;
  assign n7713 = n7248 | n7450 ;
  assign n68086 = ~n7713 ;
  assign n7714 = n7578 & n68086 ;
  assign n7715 = n7712 | n7714 ;
  assign n7716 = n163 & n7715 ;
  assign n7717 = n7239 & n68054 ;
  assign n7718 = n7530 & n7717 ;
  assign n7719 = n7716 | n7718 ;
  assign n7720 = n66505 & n7719 ;
  assign n68087 = ~n7577 ;
  assign n7721 = n7446 & n68087 ;
  assign n7722 = n7256 | n7446 ;
  assign n68088 = ~n7722 ;
  assign n7723 = n7442 & n68088 ;
  assign n7724 = n7721 | n7723 ;
  assign n7725 = n163 & n7724 ;
  assign n7726 = n7247 & n68054 ;
  assign n7727 = n7530 & n7726 ;
  assign n7728 = n7725 | n7727 ;
  assign n7729 = n66379 & n7728 ;
  assign n68089 = ~n7441 ;
  assign n7730 = n7439 & n68089 ;
  assign n7440 = n7264 | n7439 ;
  assign n68090 = ~n7440 ;
  assign n7731 = n7436 & n68090 ;
  assign n7732 = n7730 | n7731 ;
  assign n7733 = n163 & n7732 ;
  assign n7734 = n7255 & n68054 ;
  assign n7735 = n7530 & n7734 ;
  assign n7736 = n7733 | n7735 ;
  assign n7737 = n66299 & n7736 ;
  assign n68091 = ~n7573 ;
  assign n7738 = n7435 & n68091 ;
  assign n7739 = n7272 | n7435 ;
  assign n68092 = ~n7739 ;
  assign n7740 = n7431 & n68092 ;
  assign n7741 = n7738 | n7740 ;
  assign n7742 = n163 & n7741 ;
  assign n7743 = n7263 & n68054 ;
  assign n7744 = n7530 & n7743 ;
  assign n7745 = n7742 | n7744 ;
  assign n7746 = n66244 & n7745 ;
  assign n68093 = ~n7430 ;
  assign n7747 = n7429 & n68093 ;
  assign n7748 = n7280 | n7429 ;
  assign n68094 = ~n7748 ;
  assign n7749 = n7570 & n68094 ;
  assign n7750 = n7747 | n7749 ;
  assign n7751 = n163 & n7750 ;
  assign n7752 = n7271 & n68054 ;
  assign n7753 = n7530 & n7752 ;
  assign n7754 = n7751 | n7753 ;
  assign n7755 = n66145 & n7754 ;
  assign n68095 = ~n7569 ;
  assign n7756 = n7425 & n68095 ;
  assign n7757 = n7288 | n7425 ;
  assign n68096 = ~n7757 ;
  assign n7758 = n7421 & n68096 ;
  assign n7759 = n7756 | n7758 ;
  assign n7760 = n163 & n7759 ;
  assign n7761 = n7279 & n68054 ;
  assign n7762 = n7530 & n7761 ;
  assign n7763 = n7760 | n7762 ;
  assign n7764 = n66081 & n7763 ;
  assign n68097 = ~n7420 ;
  assign n7765 = n7419 & n68097 ;
  assign n7766 = n7296 | n7419 ;
  assign n68098 = ~n7766 ;
  assign n7767 = n7566 & n68098 ;
  assign n7768 = n7765 | n7767 ;
  assign n7769 = n163 & n7768 ;
  assign n7770 = n7287 & n68054 ;
  assign n7771 = n7530 & n7770 ;
  assign n7772 = n7769 | n7771 ;
  assign n7773 = n66043 & n7772 ;
  assign n68099 = ~n7565 ;
  assign n7774 = n7415 & n68099 ;
  assign n7775 = n7304 | n7415 ;
  assign n68100 = ~n7775 ;
  assign n7776 = n7411 & n68100 ;
  assign n7777 = n7774 | n7776 ;
  assign n7778 = n163 & n7777 ;
  assign n7779 = n7295 & n68054 ;
  assign n7780 = n7530 & n7779 ;
  assign n7781 = n7778 | n7780 ;
  assign n7782 = n65960 & n7781 ;
  assign n68101 = ~n7410 ;
  assign n7783 = n7409 & n68101 ;
  assign n7784 = n7312 | n7409 ;
  assign n68102 = ~n7784 ;
  assign n7785 = n7562 & n68102 ;
  assign n7786 = n7783 | n7785 ;
  assign n7787 = n163 & n7786 ;
  assign n7788 = n7303 & n68054 ;
  assign n7789 = n7530 & n7788 ;
  assign n7790 = n7787 | n7789 ;
  assign n7791 = n65909 & n7790 ;
  assign n68103 = ~n7561 ;
  assign n7792 = n7405 & n68103 ;
  assign n7793 = n7320 | n7405 ;
  assign n68104 = ~n7793 ;
  assign n7794 = n7401 & n68104 ;
  assign n7795 = n7792 | n7794 ;
  assign n7796 = n163 & n7795 ;
  assign n7797 = n7311 & n68054 ;
  assign n7798 = n7530 & n7797 ;
  assign n7799 = n7796 | n7798 ;
  assign n7800 = n65877 & n7799 ;
  assign n68105 = ~n7400 ;
  assign n7801 = n7399 & n68105 ;
  assign n7802 = n7329 | n7399 ;
  assign n68106 = ~n7802 ;
  assign n7803 = n7558 & n68106 ;
  assign n7804 = n7801 | n7803 ;
  assign n7805 = n163 & n7804 ;
  assign n7806 = n7319 & n68054 ;
  assign n7807 = n7530 & n7806 ;
  assign n7808 = n7805 | n7807 ;
  assign n7809 = n65820 & n7808 ;
  assign n68107 = ~n7557 ;
  assign n7810 = n7395 & n68107 ;
  assign n7811 = n7337 | n7395 ;
  assign n68108 = ~n7811 ;
  assign n7812 = n7391 & n68108 ;
  assign n7813 = n7810 | n7812 ;
  assign n7814 = n163 & n7813 ;
  assign n7815 = n7328 & n68054 ;
  assign n7816 = n7530 & n7815 ;
  assign n7817 = n7814 | n7816 ;
  assign n7818 = n65791 & n7817 ;
  assign n68109 = ~n7390 ;
  assign n7820 = n7389 & n68109 ;
  assign n7819 = n7347 | n7389 ;
  assign n68110 = ~n7819 ;
  assign n7821 = n7386 & n68110 ;
  assign n7822 = n7820 | n7821 ;
  assign n7823 = n163 & n7822 ;
  assign n7824 = n7336 & n68054 ;
  assign n7825 = n7530 & n7824 ;
  assign n7826 = n7823 | n7825 ;
  assign n7827 = n65772 & n7826 ;
  assign n68111 = ~n7553 ;
  assign n7829 = n7385 & n68111 ;
  assign n7828 = n7355 | n7385 ;
  assign n68112 = ~n7828 ;
  assign n7830 = n7552 & n68112 ;
  assign n7831 = n7829 | n7830 ;
  assign n7832 = n163 & n7831 ;
  assign n7833 = n7345 & n68054 ;
  assign n7834 = n7530 & n7833 ;
  assign n7835 = n7832 | n7834 ;
  assign n7836 = n65746 & n7835 ;
  assign n68113 = ~n7381 ;
  assign n7838 = n7380 & n68113 ;
  assign n7837 = n7377 | n7380 ;
  assign n68114 = ~n7837 ;
  assign n7839 = n7376 & n68114 ;
  assign n7840 = n7838 | n7839 ;
  assign n7841 = n163 & n7840 ;
  assign n7842 = n7354 & n68054 ;
  assign n7843 = n7530 & n7842 ;
  assign n7844 = n7841 | n7843 ;
  assign n7845 = n65721 & n7844 ;
  assign n7846 = n7373 & n7375 ;
  assign n7847 = n67991 & n7846 ;
  assign n68115 = ~n7847 ;
  assign n7848 = n7376 & n68115 ;
  assign n7849 = n163 & n7848 ;
  assign n7850 = n7370 & n68054 ;
  assign n7851 = n7530 & n7850 ;
  assign n7852 = n7849 | n7851 ;
  assign n7853 = n65686 & n7852 ;
  assign n7533 = n7375 & n163 ;
  assign n7854 = x64 & n163 ;
  assign n68116 = ~n7854 ;
  assign n7855 = x34 & n68116 ;
  assign n7856 = n7533 | n7855 ;
  assign n7869 = n65670 & n7856 ;
  assign n7603 = n68045 & n7602 ;
  assign n7857 = n7510 | n7603 ;
  assign n7858 = n68046 & n7857 ;
  assign n7859 = n7529 | n7858 ;
  assign n7860 = n68054 & n7859 ;
  assign n68117 = ~n7860 ;
  assign n7861 = x64 & n68117 ;
  assign n68118 = ~n7861 ;
  assign n7862 = x34 & n68118 ;
  assign n7863 = n7533 | n7862 ;
  assign n7864 = x65 & n7863 ;
  assign n7865 = x65 | n7533 ;
  assign n7866 = n7862 | n7865 ;
  assign n68119 = ~n7864 ;
  assign n7867 = n68119 & n7866 ;
  assign n68120 = ~x33 ;
  assign n7868 = n68120 & x64 ;
  assign n7870 = n7867 | n7868 ;
  assign n68121 = ~n7869 ;
  assign n7871 = n68121 & n7870 ;
  assign n68122 = ~n7851 ;
  assign n7872 = x66 & n68122 ;
  assign n68123 = ~n7849 ;
  assign n7873 = n68123 & n7872 ;
  assign n7874 = n7853 | n7873 ;
  assign n7875 = n7871 | n7874 ;
  assign n68124 = ~n7853 ;
  assign n7876 = n68124 & n7875 ;
  assign n68125 = ~n7843 ;
  assign n7877 = x67 & n68125 ;
  assign n68126 = ~n7841 ;
  assign n7878 = n68126 & n7877 ;
  assign n7879 = n7845 | n7878 ;
  assign n7880 = n7876 | n7879 ;
  assign n68127 = ~n7845 ;
  assign n7881 = n68127 & n7880 ;
  assign n68128 = ~n7834 ;
  assign n7882 = x68 & n68128 ;
  assign n68129 = ~n7832 ;
  assign n7883 = n68129 & n7882 ;
  assign n7884 = n7836 | n7883 ;
  assign n7885 = n7881 | n7884 ;
  assign n68130 = ~n7836 ;
  assign n7886 = n68130 & n7885 ;
  assign n68131 = ~n7825 ;
  assign n7887 = x69 & n68131 ;
  assign n68132 = ~n7823 ;
  assign n7888 = n68132 & n7887 ;
  assign n7889 = n7827 | n7888 ;
  assign n7890 = n7886 | n7889 ;
  assign n68133 = ~n7827 ;
  assign n7891 = n68133 & n7890 ;
  assign n68134 = ~n7816 ;
  assign n7892 = x70 & n68134 ;
  assign n68135 = ~n7814 ;
  assign n7893 = n68135 & n7892 ;
  assign n7894 = n7818 | n7893 ;
  assign n7896 = n7891 | n7894 ;
  assign n68136 = ~n7818 ;
  assign n7897 = n68136 & n7896 ;
  assign n68137 = ~n7807 ;
  assign n7898 = x71 & n68137 ;
  assign n68138 = ~n7805 ;
  assign n7899 = n68138 & n7898 ;
  assign n7900 = n7809 | n7899 ;
  assign n7901 = n7897 | n7900 ;
  assign n68139 = ~n7809 ;
  assign n7902 = n68139 & n7901 ;
  assign n68140 = ~n7798 ;
  assign n7903 = x72 & n68140 ;
  assign n68141 = ~n7796 ;
  assign n7904 = n68141 & n7903 ;
  assign n7905 = n7800 | n7904 ;
  assign n7907 = n7902 | n7905 ;
  assign n68142 = ~n7800 ;
  assign n7908 = n68142 & n7907 ;
  assign n68143 = ~n7789 ;
  assign n7909 = x73 & n68143 ;
  assign n68144 = ~n7787 ;
  assign n7910 = n68144 & n7909 ;
  assign n7911 = n7791 | n7910 ;
  assign n7912 = n7908 | n7911 ;
  assign n68145 = ~n7791 ;
  assign n7913 = n68145 & n7912 ;
  assign n68146 = ~n7780 ;
  assign n7914 = x74 & n68146 ;
  assign n68147 = ~n7778 ;
  assign n7915 = n68147 & n7914 ;
  assign n7916 = n7782 | n7915 ;
  assign n7918 = n7913 | n7916 ;
  assign n68148 = ~n7782 ;
  assign n7919 = n68148 & n7918 ;
  assign n68149 = ~n7771 ;
  assign n7920 = x75 & n68149 ;
  assign n68150 = ~n7769 ;
  assign n7921 = n68150 & n7920 ;
  assign n7922 = n7773 | n7921 ;
  assign n7923 = n7919 | n7922 ;
  assign n68151 = ~n7773 ;
  assign n7924 = n68151 & n7923 ;
  assign n68152 = ~n7762 ;
  assign n7925 = x76 & n68152 ;
  assign n68153 = ~n7760 ;
  assign n7926 = n68153 & n7925 ;
  assign n7927 = n7764 | n7926 ;
  assign n7929 = n7924 | n7927 ;
  assign n68154 = ~n7764 ;
  assign n7930 = n68154 & n7929 ;
  assign n68155 = ~n7753 ;
  assign n7931 = x77 & n68155 ;
  assign n68156 = ~n7751 ;
  assign n7932 = n68156 & n7931 ;
  assign n7933 = n7755 | n7932 ;
  assign n7934 = n7930 | n7933 ;
  assign n68157 = ~n7755 ;
  assign n7935 = n68157 & n7934 ;
  assign n68158 = ~n7744 ;
  assign n7936 = x78 & n68158 ;
  assign n68159 = ~n7742 ;
  assign n7937 = n68159 & n7936 ;
  assign n7938 = n7746 | n7937 ;
  assign n7940 = n7935 | n7938 ;
  assign n68160 = ~n7746 ;
  assign n7941 = n68160 & n7940 ;
  assign n68161 = ~n7735 ;
  assign n7942 = x79 & n68161 ;
  assign n68162 = ~n7733 ;
  assign n7943 = n68162 & n7942 ;
  assign n7944 = n7737 | n7943 ;
  assign n7945 = n7941 | n7944 ;
  assign n68163 = ~n7737 ;
  assign n7946 = n68163 & n7945 ;
  assign n68164 = ~n7727 ;
  assign n7947 = x80 & n68164 ;
  assign n68165 = ~n7725 ;
  assign n7948 = n68165 & n7947 ;
  assign n7949 = n7729 | n7948 ;
  assign n7951 = n7946 | n7949 ;
  assign n68166 = ~n7729 ;
  assign n7952 = n68166 & n7951 ;
  assign n68167 = ~n7718 ;
  assign n7953 = x81 & n68167 ;
  assign n68168 = ~n7716 ;
  assign n7954 = n68168 & n7953 ;
  assign n7955 = n7720 | n7954 ;
  assign n7956 = n7952 | n7955 ;
  assign n68169 = ~n7720 ;
  assign n7957 = n68169 & n7956 ;
  assign n68170 = ~n7709 ;
  assign n7958 = x82 & n68170 ;
  assign n68171 = ~n7707 ;
  assign n7959 = n68171 & n7958 ;
  assign n7960 = n7711 | n7959 ;
  assign n7962 = n7957 | n7960 ;
  assign n68172 = ~n7711 ;
  assign n7963 = n68172 & n7962 ;
  assign n68173 = ~n7700 ;
  assign n7964 = x83 & n68173 ;
  assign n68174 = ~n7698 ;
  assign n7965 = n68174 & n7964 ;
  assign n7966 = n7702 | n7965 ;
  assign n7967 = n7963 | n7966 ;
  assign n68175 = ~n7702 ;
  assign n7968 = n68175 & n7967 ;
  assign n68176 = ~n7691 ;
  assign n7969 = x84 & n68176 ;
  assign n68177 = ~n7689 ;
  assign n7970 = n68177 & n7969 ;
  assign n7971 = n7693 | n7970 ;
  assign n7973 = n7968 | n7971 ;
  assign n68178 = ~n7693 ;
  assign n7974 = n68178 & n7973 ;
  assign n68179 = ~n7682 ;
  assign n7975 = x85 & n68179 ;
  assign n68180 = ~n7680 ;
  assign n7976 = n68180 & n7975 ;
  assign n7977 = n7684 | n7976 ;
  assign n7978 = n7974 | n7977 ;
  assign n68181 = ~n7684 ;
  assign n7979 = n68181 & n7978 ;
  assign n68182 = ~n7673 ;
  assign n7980 = x86 & n68182 ;
  assign n68183 = ~n7671 ;
  assign n7981 = n68183 & n7980 ;
  assign n7982 = n7675 | n7981 ;
  assign n7984 = n7979 | n7982 ;
  assign n68184 = ~n7675 ;
  assign n7985 = n68184 & n7984 ;
  assign n68185 = ~n7664 ;
  assign n7986 = x87 & n68185 ;
  assign n68186 = ~n7662 ;
  assign n7987 = n68186 & n7986 ;
  assign n7988 = n7666 | n7987 ;
  assign n7989 = n7985 | n7988 ;
  assign n68187 = ~n7666 ;
  assign n7990 = n68187 & n7989 ;
  assign n68188 = ~n7655 ;
  assign n7991 = x88 & n68188 ;
  assign n68189 = ~n7653 ;
  assign n7992 = n68189 & n7991 ;
  assign n7993 = n7657 | n7992 ;
  assign n7995 = n7990 | n7993 ;
  assign n68190 = ~n7657 ;
  assign n7996 = n68190 & n7995 ;
  assign n68191 = ~n7646 ;
  assign n7997 = x89 & n68191 ;
  assign n68192 = ~n7644 ;
  assign n7998 = n68192 & n7997 ;
  assign n7999 = n7648 | n7998 ;
  assign n8000 = n7996 | n7999 ;
  assign n68193 = ~n7648 ;
  assign n8001 = n68193 & n8000 ;
  assign n68194 = ~n7637 ;
  assign n8002 = x90 & n68194 ;
  assign n68195 = ~n7635 ;
  assign n8003 = n68195 & n8002 ;
  assign n8004 = n7639 | n8003 ;
  assign n8006 = n8001 | n8004 ;
  assign n68196 = ~n7639 ;
  assign n8007 = n68196 & n8006 ;
  assign n68197 = ~n7628 ;
  assign n8008 = x91 & n68197 ;
  assign n68198 = ~n7626 ;
  assign n8009 = n68198 & n8008 ;
  assign n8010 = n7630 | n8009 ;
  assign n8011 = n8007 | n8010 ;
  assign n68199 = ~n7630 ;
  assign n8012 = n68199 & n8011 ;
  assign n68200 = ~n7619 ;
  assign n8013 = x92 & n68200 ;
  assign n68201 = ~n7617 ;
  assign n8014 = n68201 & n8013 ;
  assign n8015 = n7621 | n8014 ;
  assign n8017 = n8012 | n8015 ;
  assign n68202 = ~n7621 ;
  assign n8018 = n68202 & n8017 ;
  assign n68203 = ~n7610 ;
  assign n8019 = x93 & n68203 ;
  assign n68204 = ~n7608 ;
  assign n8020 = n68204 & n8019 ;
  assign n8021 = n7612 | n8020 ;
  assign n8022 = n8018 | n8021 ;
  assign n68205 = ~n7612 ;
  assign n8023 = n68205 & n8022 ;
  assign n68206 = ~n7542 ;
  assign n8024 = x94 & n68206 ;
  assign n68207 = ~n7540 ;
  assign n8025 = n68207 & n8024 ;
  assign n8026 = n7544 | n8025 ;
  assign n8028 = n8023 | n8026 ;
  assign n68208 = ~n7544 ;
  assign n8029 = n68208 & n8028 ;
  assign n8030 = n73737 | n285 ;
  assign n8031 = n468 | n8030 ;
  assign n8032 = n465 | n8031 ;
  assign n8033 = n8029 | n8032 ;
  assign n68209 = ~n8023 ;
  assign n8027 = n68209 & n8026 ;
  assign n8034 = x65 & n7856 ;
  assign n68210 = ~n8034 ;
  assign n8035 = n7866 & n68210 ;
  assign n8036 = n7868 | n8035 ;
  assign n8037 = n68121 & n8036 ;
  assign n8038 = n7874 | n8037 ;
  assign n8039 = n68124 & n8038 ;
  assign n8041 = n7879 | n8039 ;
  assign n8042 = n68127 & n8041 ;
  assign n8044 = n7884 | n8042 ;
  assign n8045 = n68130 & n8044 ;
  assign n8046 = n7889 | n8045 ;
  assign n8048 = n68133 & n8046 ;
  assign n8049 = n7894 | n8048 ;
  assign n8050 = n68136 & n8049 ;
  assign n8051 = n7900 | n8050 ;
  assign n8053 = n68139 & n8051 ;
  assign n8054 = n7905 | n8053 ;
  assign n8055 = n68142 & n8054 ;
  assign n8056 = n7911 | n8055 ;
  assign n8058 = n68145 & n8056 ;
  assign n8059 = n7916 | n8058 ;
  assign n8060 = n68148 & n8059 ;
  assign n8061 = n7922 | n8060 ;
  assign n8063 = n68151 & n8061 ;
  assign n8064 = n7927 | n8063 ;
  assign n8065 = n68154 & n8064 ;
  assign n8066 = n7933 | n8065 ;
  assign n8068 = n68157 & n8066 ;
  assign n8069 = n7938 | n8068 ;
  assign n8070 = n68160 & n8069 ;
  assign n8071 = n7944 | n8070 ;
  assign n8073 = n68163 & n8071 ;
  assign n8074 = n7949 | n8073 ;
  assign n8075 = n68166 & n8074 ;
  assign n8076 = n7955 | n8075 ;
  assign n8078 = n68169 & n8076 ;
  assign n8079 = n7960 | n8078 ;
  assign n8080 = n68172 & n8079 ;
  assign n8081 = n7966 | n8080 ;
  assign n8083 = n68175 & n8081 ;
  assign n8084 = n7971 | n8083 ;
  assign n8085 = n68178 & n8084 ;
  assign n8086 = n7977 | n8085 ;
  assign n8088 = n68181 & n8086 ;
  assign n8089 = n7982 | n8088 ;
  assign n8090 = n68184 & n8089 ;
  assign n8091 = n7988 | n8090 ;
  assign n8093 = n68187 & n8091 ;
  assign n8094 = n7993 | n8093 ;
  assign n8095 = n68190 & n8094 ;
  assign n8096 = n7999 | n8095 ;
  assign n8098 = n68193 & n8096 ;
  assign n8099 = n8004 | n8098 ;
  assign n8100 = n68196 & n8099 ;
  assign n8101 = n8010 | n8100 ;
  assign n8103 = n68199 & n8101 ;
  assign n8104 = n8015 | n8103 ;
  assign n8105 = n68202 & n8104 ;
  assign n8107 = n8021 | n8105 ;
  assign n8108 = n7612 | n8026 ;
  assign n68211 = ~n8108 ;
  assign n8109 = n8107 & n68211 ;
  assign n8110 = n8027 | n8109 ;
  assign n8111 = n8033 | n8110 ;
  assign n68212 = ~n7543 ;
  assign n8112 = n68212 & n8033 ;
  assign n68213 = ~n8112 ;
  assign n8113 = n8111 & n68213 ;
  assign n68214 = ~x95 ;
  assign n8114 = n68214 & n8113 ;
  assign n162 = ~n8033 ;
  assign n8543 = n162 & n8110 ;
  assign n8544 = n7543 & n8033 ;
  assign n68216 = ~n8544 ;
  assign n8545 = x95 & n68216 ;
  assign n68217 = ~n8543 ;
  assign n8546 = n68217 & n8545 ;
  assign n8547 = n8114 | n8546 ;
  assign n8115 = n7611 & n8033 ;
  assign n68218 = ~n8105 ;
  assign n8106 = n8021 & n68218 ;
  assign n8116 = n7621 | n8021 ;
  assign n68219 = ~n8116 ;
  assign n8117 = n8017 & n68219 ;
  assign n8118 = n8106 | n8117 ;
  assign n68220 = ~n8032 ;
  assign n8119 = n68220 & n8118 ;
  assign n68221 = ~n8029 ;
  assign n8120 = n68221 & n8119 ;
  assign n8121 = n8115 | n8120 ;
  assign n8122 = n68058 & n8121 ;
  assign n8123 = n7620 & n8033 ;
  assign n68222 = ~n8012 ;
  assign n8016 = n68222 & n8015 ;
  assign n8124 = n7630 | n8015 ;
  assign n68223 = ~n8124 ;
  assign n8125 = n8101 & n68223 ;
  assign n8126 = n8016 | n8125 ;
  assign n8127 = n68220 & n8126 ;
  assign n8128 = n68221 & n8127 ;
  assign n8129 = n8123 | n8128 ;
  assign n8130 = n67986 & n8129 ;
  assign n68224 = ~n8128 ;
  assign n8531 = x93 & n68224 ;
  assign n68225 = ~n8123 ;
  assign n8532 = n68225 & n8531 ;
  assign n8533 = n8130 | n8532 ;
  assign n8131 = n7629 & n8033 ;
  assign n68226 = ~n8100 ;
  assign n8102 = n8010 & n68226 ;
  assign n8132 = n7639 | n8010 ;
  assign n68227 = ~n8132 ;
  assign n8133 = n8006 & n68227 ;
  assign n8134 = n8102 | n8133 ;
  assign n8135 = n68220 & n8134 ;
  assign n8136 = n68221 & n8135 ;
  assign n8137 = n8131 | n8136 ;
  assign n8138 = n67763 & n8137 ;
  assign n8139 = n7638 & n8033 ;
  assign n68228 = ~n8001 ;
  assign n8005 = n68228 & n8004 ;
  assign n8140 = n7648 | n8004 ;
  assign n68229 = ~n8140 ;
  assign n8141 = n8096 & n68229 ;
  assign n8142 = n8005 | n8141 ;
  assign n8143 = n68220 & n8142 ;
  assign n8144 = n68221 & n8143 ;
  assign n8145 = n8139 | n8144 ;
  assign n8146 = n67622 & n8145 ;
  assign n68230 = ~n8144 ;
  assign n8519 = x91 & n68230 ;
  assign n68231 = ~n8139 ;
  assign n8520 = n68231 & n8519 ;
  assign n8521 = n8146 | n8520 ;
  assign n8147 = n7647 & n8033 ;
  assign n68232 = ~n8095 ;
  assign n8097 = n7999 & n68232 ;
  assign n8148 = n7657 | n7999 ;
  assign n68233 = ~n8148 ;
  assign n8149 = n7995 & n68233 ;
  assign n8150 = n8097 | n8149 ;
  assign n8151 = n68220 & n8150 ;
  assign n8152 = n68221 & n8151 ;
  assign n8153 = n8147 | n8152 ;
  assign n8154 = n67531 & n8153 ;
  assign n8155 = n7656 & n8033 ;
  assign n68234 = ~n7990 ;
  assign n7994 = n68234 & n7993 ;
  assign n8156 = n7666 | n7993 ;
  assign n68235 = ~n8156 ;
  assign n8157 = n8091 & n68235 ;
  assign n8158 = n7994 | n8157 ;
  assign n8159 = n68220 & n8158 ;
  assign n8160 = n68221 & n8159 ;
  assign n8161 = n8155 | n8160 ;
  assign n8162 = n67348 & n8161 ;
  assign n68236 = ~n8160 ;
  assign n8507 = x89 & n68236 ;
  assign n68237 = ~n8155 ;
  assign n8508 = n68237 & n8507 ;
  assign n8509 = n8162 | n8508 ;
  assign n8163 = n7665 & n8033 ;
  assign n68238 = ~n8090 ;
  assign n8092 = n7988 & n68238 ;
  assign n8164 = n7675 | n7988 ;
  assign n68239 = ~n8164 ;
  assign n8165 = n7984 & n68239 ;
  assign n8166 = n8092 | n8165 ;
  assign n8167 = n68220 & n8166 ;
  assign n8168 = n68221 & n8167 ;
  assign n8169 = n8163 | n8168 ;
  assign n8170 = n67222 & n8169 ;
  assign n8171 = n7674 & n8033 ;
  assign n68240 = ~n7979 ;
  assign n7983 = n68240 & n7982 ;
  assign n8172 = n7684 | n7982 ;
  assign n68241 = ~n8172 ;
  assign n8173 = n8086 & n68241 ;
  assign n8174 = n7983 | n8173 ;
  assign n8175 = n68220 & n8174 ;
  assign n8176 = n68221 & n8175 ;
  assign n8177 = n8171 | n8176 ;
  assign n8178 = n67164 & n8177 ;
  assign n68242 = ~n8176 ;
  assign n8495 = x87 & n68242 ;
  assign n68243 = ~n8171 ;
  assign n8496 = n68243 & n8495 ;
  assign n8497 = n8178 | n8496 ;
  assign n8179 = n7683 & n8033 ;
  assign n68244 = ~n8085 ;
  assign n8087 = n7977 & n68244 ;
  assign n8180 = n7693 | n7977 ;
  assign n68245 = ~n8180 ;
  assign n8181 = n7973 & n68245 ;
  assign n8182 = n8087 | n8181 ;
  assign n8183 = n68220 & n8182 ;
  assign n8184 = n68221 & n8183 ;
  assign n8185 = n8179 | n8184 ;
  assign n8186 = n66979 & n8185 ;
  assign n8187 = n7692 & n8033 ;
  assign n68246 = ~n7968 ;
  assign n7972 = n68246 & n7971 ;
  assign n8188 = n7702 | n7971 ;
  assign n68247 = ~n8188 ;
  assign n8189 = n8081 & n68247 ;
  assign n8190 = n7972 | n8189 ;
  assign n8191 = n68220 & n8190 ;
  assign n8192 = n68221 & n8191 ;
  assign n8193 = n8187 | n8192 ;
  assign n8194 = n66868 & n8193 ;
  assign n68248 = ~n8192 ;
  assign n8483 = x85 & n68248 ;
  assign n68249 = ~n8187 ;
  assign n8484 = n68249 & n8483 ;
  assign n8485 = n8194 | n8484 ;
  assign n8195 = n7701 & n8033 ;
  assign n68250 = ~n8080 ;
  assign n8082 = n7966 & n68250 ;
  assign n8196 = n7711 | n7966 ;
  assign n68251 = ~n8196 ;
  assign n8197 = n7962 & n68251 ;
  assign n8198 = n8082 | n8197 ;
  assign n8199 = n68220 & n8198 ;
  assign n8200 = n68221 & n8199 ;
  assign n8201 = n8195 | n8200 ;
  assign n8202 = n66797 & n8201 ;
  assign n8203 = n7710 & n8033 ;
  assign n68252 = ~n7957 ;
  assign n7961 = n68252 & n7960 ;
  assign n8204 = n7720 | n7960 ;
  assign n68253 = ~n8204 ;
  assign n8205 = n8076 & n68253 ;
  assign n8206 = n7961 | n8205 ;
  assign n8207 = n68220 & n8206 ;
  assign n8208 = n68221 & n8207 ;
  assign n8209 = n8203 | n8208 ;
  assign n8210 = n66654 & n8209 ;
  assign n68254 = ~n8208 ;
  assign n8471 = x83 & n68254 ;
  assign n68255 = ~n8203 ;
  assign n8472 = n68255 & n8471 ;
  assign n8473 = n8210 | n8472 ;
  assign n8211 = n7719 & n8033 ;
  assign n68256 = ~n8075 ;
  assign n8077 = n7955 & n68256 ;
  assign n8212 = n7729 | n7955 ;
  assign n68257 = ~n8212 ;
  assign n8213 = n7951 & n68257 ;
  assign n8214 = n8077 | n8213 ;
  assign n8215 = n68220 & n8214 ;
  assign n8216 = n68221 & n8215 ;
  assign n8217 = n8211 | n8216 ;
  assign n8218 = n66560 & n8217 ;
  assign n8219 = n7728 & n8033 ;
  assign n68258 = ~n7946 ;
  assign n7950 = n68258 & n7949 ;
  assign n8220 = n7737 | n7949 ;
  assign n68259 = ~n8220 ;
  assign n8221 = n8071 & n68259 ;
  assign n8222 = n7950 | n8221 ;
  assign n8223 = n68220 & n8222 ;
  assign n8224 = n68221 & n8223 ;
  assign n8225 = n8219 | n8224 ;
  assign n8226 = n66505 & n8225 ;
  assign n68260 = ~n8224 ;
  assign n8459 = x81 & n68260 ;
  assign n68261 = ~n8219 ;
  assign n8460 = n68261 & n8459 ;
  assign n8461 = n8226 | n8460 ;
  assign n8227 = n7736 & n8033 ;
  assign n68262 = ~n8070 ;
  assign n8072 = n7944 & n68262 ;
  assign n8228 = n7746 | n7944 ;
  assign n68263 = ~n8228 ;
  assign n8229 = n7940 & n68263 ;
  assign n8230 = n8072 | n8229 ;
  assign n8231 = n68220 & n8230 ;
  assign n8232 = n68221 & n8231 ;
  assign n8233 = n8227 | n8232 ;
  assign n8234 = n66379 & n8233 ;
  assign n8235 = n7745 & n8033 ;
  assign n68264 = ~n7935 ;
  assign n7939 = n68264 & n7938 ;
  assign n8236 = n7755 | n7938 ;
  assign n68265 = ~n8236 ;
  assign n8237 = n8066 & n68265 ;
  assign n8238 = n7939 | n8237 ;
  assign n8239 = n68220 & n8238 ;
  assign n8240 = n68221 & n8239 ;
  assign n8241 = n8235 | n8240 ;
  assign n8242 = n66299 & n8241 ;
  assign n68266 = ~n8240 ;
  assign n8447 = x79 & n68266 ;
  assign n68267 = ~n8235 ;
  assign n8448 = n68267 & n8447 ;
  assign n8449 = n8242 | n8448 ;
  assign n8243 = n7754 & n8033 ;
  assign n68268 = ~n8065 ;
  assign n8067 = n7933 & n68268 ;
  assign n8244 = n7764 | n7933 ;
  assign n68269 = ~n8244 ;
  assign n8245 = n7929 & n68269 ;
  assign n8246 = n8067 | n8245 ;
  assign n8247 = n68220 & n8246 ;
  assign n8248 = n68221 & n8247 ;
  assign n8249 = n8243 | n8248 ;
  assign n8250 = n66244 & n8249 ;
  assign n8251 = n7763 & n8033 ;
  assign n68270 = ~n7924 ;
  assign n7928 = n68270 & n7927 ;
  assign n8252 = n7773 | n7927 ;
  assign n68271 = ~n8252 ;
  assign n8253 = n8061 & n68271 ;
  assign n8254 = n7928 | n8253 ;
  assign n8255 = n68220 & n8254 ;
  assign n8256 = n68221 & n8255 ;
  assign n8257 = n8251 | n8256 ;
  assign n8258 = n66145 & n8257 ;
  assign n68272 = ~n8256 ;
  assign n8435 = x77 & n68272 ;
  assign n68273 = ~n8251 ;
  assign n8436 = n68273 & n8435 ;
  assign n8437 = n8258 | n8436 ;
  assign n8259 = n7772 & n8033 ;
  assign n68274 = ~n8060 ;
  assign n8062 = n7922 & n68274 ;
  assign n8260 = n7782 | n7922 ;
  assign n68275 = ~n8260 ;
  assign n8261 = n7918 & n68275 ;
  assign n8262 = n8062 | n8261 ;
  assign n8263 = n68220 & n8262 ;
  assign n8264 = n68221 & n8263 ;
  assign n8265 = n8259 | n8264 ;
  assign n8266 = n66081 & n8265 ;
  assign n8267 = n7781 & n8033 ;
  assign n68276 = ~n7913 ;
  assign n7917 = n68276 & n7916 ;
  assign n8268 = n7791 | n7916 ;
  assign n68277 = ~n8268 ;
  assign n8269 = n8056 & n68277 ;
  assign n8270 = n7917 | n8269 ;
  assign n8271 = n68220 & n8270 ;
  assign n8272 = n68221 & n8271 ;
  assign n8273 = n8267 | n8272 ;
  assign n8274 = n66043 & n8273 ;
  assign n68278 = ~n8272 ;
  assign n8423 = x75 & n68278 ;
  assign n68279 = ~n8267 ;
  assign n8424 = n68279 & n8423 ;
  assign n8425 = n8274 | n8424 ;
  assign n8275 = n7790 & n8033 ;
  assign n68280 = ~n8055 ;
  assign n8057 = n7911 & n68280 ;
  assign n8276 = n7800 | n7911 ;
  assign n68281 = ~n8276 ;
  assign n8277 = n7907 & n68281 ;
  assign n8278 = n8057 | n8277 ;
  assign n8279 = n68220 & n8278 ;
  assign n8280 = n68221 & n8279 ;
  assign n8281 = n8275 | n8280 ;
  assign n8282 = n65960 & n8281 ;
  assign n8283 = n7799 & n8033 ;
  assign n68282 = ~n7902 ;
  assign n7906 = n68282 & n7905 ;
  assign n8284 = n7809 | n7905 ;
  assign n68283 = ~n8284 ;
  assign n8285 = n8051 & n68283 ;
  assign n8286 = n7906 | n8285 ;
  assign n8287 = n68220 & n8286 ;
  assign n8288 = n68221 & n8287 ;
  assign n8289 = n8283 | n8288 ;
  assign n8290 = n65909 & n8289 ;
  assign n68284 = ~n8288 ;
  assign n8411 = x73 & n68284 ;
  assign n68285 = ~n8283 ;
  assign n8412 = n68285 & n8411 ;
  assign n8413 = n8290 | n8412 ;
  assign n8291 = n7808 & n8033 ;
  assign n68286 = ~n8050 ;
  assign n8052 = n7900 & n68286 ;
  assign n8292 = n7818 | n7900 ;
  assign n68287 = ~n8292 ;
  assign n8293 = n7896 & n68287 ;
  assign n8294 = n8052 | n8293 ;
  assign n8295 = n68220 & n8294 ;
  assign n8296 = n68221 & n8295 ;
  assign n8297 = n8291 | n8296 ;
  assign n8298 = n65877 & n8297 ;
  assign n8299 = n7817 & n8033 ;
  assign n68288 = ~n7891 ;
  assign n7895 = n68288 & n7894 ;
  assign n8300 = n7827 | n7894 ;
  assign n68289 = ~n8300 ;
  assign n8301 = n8046 & n68289 ;
  assign n8302 = n7895 | n8301 ;
  assign n8303 = n68220 & n8302 ;
  assign n8304 = n68221 & n8303 ;
  assign n8305 = n8299 | n8304 ;
  assign n8306 = n65820 & n8305 ;
  assign n68290 = ~n8304 ;
  assign n8399 = x71 & n68290 ;
  assign n68291 = ~n8299 ;
  assign n8400 = n68291 & n8399 ;
  assign n8401 = n8306 | n8400 ;
  assign n8307 = n7826 & n8033 ;
  assign n68292 = ~n8045 ;
  assign n8047 = n7889 & n68292 ;
  assign n8308 = n7836 | n7889 ;
  assign n68293 = ~n8308 ;
  assign n8309 = n7885 & n68293 ;
  assign n8310 = n8047 | n8309 ;
  assign n8311 = n68220 & n8310 ;
  assign n8312 = n68221 & n8311 ;
  assign n8313 = n8307 | n8312 ;
  assign n8314 = n65791 & n8313 ;
  assign n8315 = n7835 & n8033 ;
  assign n68294 = ~n7881 ;
  assign n8043 = n68294 & n7884 ;
  assign n8316 = n7845 | n7884 ;
  assign n68295 = ~n8316 ;
  assign n8317 = n8041 & n68295 ;
  assign n8318 = n8043 | n8317 ;
  assign n8319 = n68220 & n8318 ;
  assign n8320 = n68221 & n8319 ;
  assign n8321 = n8315 | n8320 ;
  assign n8322 = n65772 & n8321 ;
  assign n68296 = ~n8320 ;
  assign n8388 = x69 & n68296 ;
  assign n68297 = ~n8315 ;
  assign n8389 = n68297 & n8388 ;
  assign n8390 = n8322 | n8389 ;
  assign n8323 = n7844 & n8033 ;
  assign n68298 = ~n8039 ;
  assign n8040 = n7879 & n68298 ;
  assign n8324 = n7853 | n7879 ;
  assign n68299 = ~n8324 ;
  assign n8325 = n8038 & n68299 ;
  assign n8326 = n8040 | n8325 ;
  assign n8327 = n68220 & n8326 ;
  assign n8328 = n68221 & n8327 ;
  assign n8329 = n8323 | n8328 ;
  assign n8330 = n65746 & n8329 ;
  assign n8331 = n7852 & n8033 ;
  assign n8332 = n7869 | n7874 ;
  assign n68300 = ~n8332 ;
  assign n8333 = n8036 & n68300 ;
  assign n68301 = ~n7871 ;
  assign n8334 = n68301 & n7874 ;
  assign n8335 = n8333 | n8334 ;
  assign n8336 = n68220 & n8335 ;
  assign n8337 = n68221 & n8336 ;
  assign n8338 = n8331 | n8337 ;
  assign n8339 = n65721 & n8338 ;
  assign n68302 = ~n8337 ;
  assign n8378 = x67 & n68302 ;
  assign n68303 = ~n8331 ;
  assign n8379 = n68303 & n8378 ;
  assign n8380 = n8339 | n8379 ;
  assign n8340 = n7863 & n8033 ;
  assign n8341 = n7866 & n7868 ;
  assign n8342 = n68210 & n8341 ;
  assign n8343 = n8032 | n8342 ;
  assign n68304 = ~n8343 ;
  assign n8344 = n8036 & n68304 ;
  assign n8345 = n68221 & n8344 ;
  assign n8346 = n8340 | n8345 ;
  assign n8347 = n65686 & n8346 ;
  assign n68305 = ~x32 ;
  assign n8368 = n68305 & x64 ;
  assign n8348 = x64 & n68214 ;
  assign n8349 = n67988 & n8348 ;
  assign n8350 = n67020 & n8349 ;
  assign n8351 = n67021 & n8350 ;
  assign n8352 = n68221 & n8351 ;
  assign n68306 = ~n8352 ;
  assign n8353 = x33 & n68306 ;
  assign n68307 = ~n73737 ;
  assign n8354 = n68307 & n7868 ;
  assign n68308 = ~n285 ;
  assign n8355 = n68308 & n8354 ;
  assign n8356 = n67025 & n8355 ;
  assign n8357 = n67026 & n8356 ;
  assign n8358 = n68221 & n8357 ;
  assign n8359 = n8353 | n8358 ;
  assign n8360 = x65 & n8359 ;
  assign n8361 = n68205 & n8107 ;
  assign n8362 = n8026 | n8361 ;
  assign n8363 = n68208 & n8362 ;
  assign n68309 = ~n8363 ;
  assign n8364 = n8351 & n68309 ;
  assign n68310 = ~n8364 ;
  assign n8365 = x33 & n68310 ;
  assign n8366 = x65 | n8358 ;
  assign n8367 = n8365 | n8366 ;
  assign n68311 = ~n8360 ;
  assign n8369 = n68311 & n8367 ;
  assign n8370 = n8368 | n8369 ;
  assign n8371 = n8358 | n8365 ;
  assign n8372 = n65670 & n8371 ;
  assign n68312 = ~n8372 ;
  assign n8373 = n8370 & n68312 ;
  assign n68313 = ~n8345 ;
  assign n8374 = x66 & n68313 ;
  assign n68314 = ~n8340 ;
  assign n8375 = n68314 & n8374 ;
  assign n8376 = n8347 | n8375 ;
  assign n8377 = n8373 | n8376 ;
  assign n68315 = ~n8347 ;
  assign n8381 = n68315 & n8377 ;
  assign n8382 = n8380 | n8381 ;
  assign n68316 = ~n8339 ;
  assign n8383 = n68316 & n8382 ;
  assign n68317 = ~n8328 ;
  assign n8384 = x68 & n68317 ;
  assign n68318 = ~n8323 ;
  assign n8385 = n68318 & n8384 ;
  assign n8386 = n8330 | n8385 ;
  assign n8387 = n8383 | n8386 ;
  assign n68319 = ~n8330 ;
  assign n8391 = n68319 & n8387 ;
  assign n8392 = n8390 | n8391 ;
  assign n68320 = ~n8322 ;
  assign n8393 = n68320 & n8392 ;
  assign n68321 = ~n8312 ;
  assign n8394 = x70 & n68321 ;
  assign n68322 = ~n8307 ;
  assign n8395 = n68322 & n8394 ;
  assign n8396 = n8314 | n8395 ;
  assign n8398 = n8393 | n8396 ;
  assign n68323 = ~n8314 ;
  assign n8403 = n68323 & n8398 ;
  assign n8404 = n8401 | n8403 ;
  assign n68324 = ~n8306 ;
  assign n8405 = n68324 & n8404 ;
  assign n68325 = ~n8296 ;
  assign n8406 = x72 & n68325 ;
  assign n68326 = ~n8291 ;
  assign n8407 = n68326 & n8406 ;
  assign n8408 = n8298 | n8407 ;
  assign n8410 = n8405 | n8408 ;
  assign n68327 = ~n8298 ;
  assign n8415 = n68327 & n8410 ;
  assign n8416 = n8413 | n8415 ;
  assign n68328 = ~n8290 ;
  assign n8417 = n68328 & n8416 ;
  assign n68329 = ~n8280 ;
  assign n8418 = x74 & n68329 ;
  assign n68330 = ~n8275 ;
  assign n8419 = n68330 & n8418 ;
  assign n8420 = n8282 | n8419 ;
  assign n8422 = n8417 | n8420 ;
  assign n68331 = ~n8282 ;
  assign n8427 = n68331 & n8422 ;
  assign n8428 = n8425 | n8427 ;
  assign n68332 = ~n8274 ;
  assign n8429 = n68332 & n8428 ;
  assign n68333 = ~n8264 ;
  assign n8430 = x76 & n68333 ;
  assign n68334 = ~n8259 ;
  assign n8431 = n68334 & n8430 ;
  assign n8432 = n8266 | n8431 ;
  assign n8434 = n8429 | n8432 ;
  assign n68335 = ~n8266 ;
  assign n8439 = n68335 & n8434 ;
  assign n8440 = n8437 | n8439 ;
  assign n68336 = ~n8258 ;
  assign n8441 = n68336 & n8440 ;
  assign n68337 = ~n8248 ;
  assign n8442 = x78 & n68337 ;
  assign n68338 = ~n8243 ;
  assign n8443 = n68338 & n8442 ;
  assign n8444 = n8250 | n8443 ;
  assign n8446 = n8441 | n8444 ;
  assign n68339 = ~n8250 ;
  assign n8451 = n68339 & n8446 ;
  assign n8452 = n8449 | n8451 ;
  assign n68340 = ~n8242 ;
  assign n8453 = n68340 & n8452 ;
  assign n68341 = ~n8232 ;
  assign n8454 = x80 & n68341 ;
  assign n68342 = ~n8227 ;
  assign n8455 = n68342 & n8454 ;
  assign n8456 = n8234 | n8455 ;
  assign n8458 = n8453 | n8456 ;
  assign n68343 = ~n8234 ;
  assign n8463 = n68343 & n8458 ;
  assign n8464 = n8461 | n8463 ;
  assign n68344 = ~n8226 ;
  assign n8465 = n68344 & n8464 ;
  assign n68345 = ~n8216 ;
  assign n8466 = x82 & n68345 ;
  assign n68346 = ~n8211 ;
  assign n8467 = n68346 & n8466 ;
  assign n8468 = n8218 | n8467 ;
  assign n8470 = n8465 | n8468 ;
  assign n68347 = ~n8218 ;
  assign n8475 = n68347 & n8470 ;
  assign n8476 = n8473 | n8475 ;
  assign n68348 = ~n8210 ;
  assign n8477 = n68348 & n8476 ;
  assign n68349 = ~n8200 ;
  assign n8478 = x84 & n68349 ;
  assign n68350 = ~n8195 ;
  assign n8479 = n68350 & n8478 ;
  assign n8480 = n8202 | n8479 ;
  assign n8482 = n8477 | n8480 ;
  assign n68351 = ~n8202 ;
  assign n8487 = n68351 & n8482 ;
  assign n8488 = n8485 | n8487 ;
  assign n68352 = ~n8194 ;
  assign n8489 = n68352 & n8488 ;
  assign n68353 = ~n8184 ;
  assign n8490 = x86 & n68353 ;
  assign n68354 = ~n8179 ;
  assign n8491 = n68354 & n8490 ;
  assign n8492 = n8186 | n8491 ;
  assign n8494 = n8489 | n8492 ;
  assign n68355 = ~n8186 ;
  assign n8499 = n68355 & n8494 ;
  assign n8500 = n8497 | n8499 ;
  assign n68356 = ~n8178 ;
  assign n8501 = n68356 & n8500 ;
  assign n68357 = ~n8168 ;
  assign n8502 = x88 & n68357 ;
  assign n68358 = ~n8163 ;
  assign n8503 = n68358 & n8502 ;
  assign n8504 = n8170 | n8503 ;
  assign n8506 = n8501 | n8504 ;
  assign n68359 = ~n8170 ;
  assign n8511 = n68359 & n8506 ;
  assign n8512 = n8509 | n8511 ;
  assign n68360 = ~n8162 ;
  assign n8513 = n68360 & n8512 ;
  assign n68361 = ~n8152 ;
  assign n8514 = x90 & n68361 ;
  assign n68362 = ~n8147 ;
  assign n8515 = n68362 & n8514 ;
  assign n8516 = n8154 | n8515 ;
  assign n8518 = n8513 | n8516 ;
  assign n68363 = ~n8154 ;
  assign n8523 = n68363 & n8518 ;
  assign n8524 = n8521 | n8523 ;
  assign n68364 = ~n8146 ;
  assign n8525 = n68364 & n8524 ;
  assign n68365 = ~n8136 ;
  assign n8526 = x92 & n68365 ;
  assign n68366 = ~n8131 ;
  assign n8527 = n68366 & n8526 ;
  assign n8528 = n8138 | n8527 ;
  assign n8530 = n8525 | n8528 ;
  assign n68367 = ~n8138 ;
  assign n8535 = n68367 & n8530 ;
  assign n8536 = n8533 | n8535 ;
  assign n68368 = ~n8130 ;
  assign n8537 = n68368 & n8536 ;
  assign n68369 = ~n8120 ;
  assign n8538 = x94 & n68369 ;
  assign n68370 = ~n8115 ;
  assign n8539 = n68370 & n8538 ;
  assign n8540 = n8122 | n8539 ;
  assign n8542 = n8537 | n8540 ;
  assign n68371 = ~n8122 ;
  assign n8548 = n68371 & n8542 ;
  assign n8549 = n8547 | n8548 ;
  assign n68372 = ~n8114 ;
  assign n8550 = n68372 & n8549 ;
  assign n8551 = n303 | n8550 ;
  assign n68373 = ~n8113 ;
  assign n8553 = n68373 & n8551 ;
  assign n68374 = ~n8548 ;
  assign n9044 = n8547 & n68374 ;
  assign n8555 = x65 & n8371 ;
  assign n68375 = ~n8555 ;
  assign n8556 = n8367 & n68375 ;
  assign n8558 = n8368 | n8556 ;
  assign n8559 = n68312 & n8558 ;
  assign n8560 = n8376 | n8559 ;
  assign n8561 = n68315 & n8560 ;
  assign n8562 = n8380 | n8561 ;
  assign n8563 = n68316 & n8562 ;
  assign n8564 = n8386 | n8563 ;
  assign n8565 = n68319 & n8564 ;
  assign n8566 = n8390 | n8565 ;
  assign n8567 = n68320 & n8566 ;
  assign n8568 = n8396 | n8567 ;
  assign n8569 = n68323 & n8568 ;
  assign n8570 = n8401 | n8569 ;
  assign n8571 = n68324 & n8570 ;
  assign n8572 = n8408 | n8571 ;
  assign n8573 = n68327 & n8572 ;
  assign n8574 = n8413 | n8573 ;
  assign n8575 = n68328 & n8574 ;
  assign n8576 = n8420 | n8575 ;
  assign n8577 = n68331 & n8576 ;
  assign n8578 = n8425 | n8577 ;
  assign n8579 = n68332 & n8578 ;
  assign n8580 = n8432 | n8579 ;
  assign n8581 = n68335 & n8580 ;
  assign n8582 = n8437 | n8581 ;
  assign n8583 = n68336 & n8582 ;
  assign n8584 = n8444 | n8583 ;
  assign n8585 = n68339 & n8584 ;
  assign n8586 = n8449 | n8585 ;
  assign n8587 = n68340 & n8586 ;
  assign n8588 = n8456 | n8587 ;
  assign n8589 = n68343 & n8588 ;
  assign n8590 = n8461 | n8589 ;
  assign n8591 = n68344 & n8590 ;
  assign n8592 = n8468 | n8591 ;
  assign n8593 = n68347 & n8592 ;
  assign n8594 = n8473 | n8593 ;
  assign n8595 = n68348 & n8594 ;
  assign n8596 = n8480 | n8595 ;
  assign n8597 = n68351 & n8596 ;
  assign n8598 = n8485 | n8597 ;
  assign n8599 = n68352 & n8598 ;
  assign n8600 = n8492 | n8599 ;
  assign n8601 = n68355 & n8600 ;
  assign n8602 = n8497 | n8601 ;
  assign n8603 = n68356 & n8602 ;
  assign n8604 = n8504 | n8603 ;
  assign n8605 = n68359 & n8604 ;
  assign n8606 = n8509 | n8605 ;
  assign n8607 = n68360 & n8606 ;
  assign n8608 = n8516 | n8607 ;
  assign n8609 = n68363 & n8608 ;
  assign n8610 = n8521 | n8609 ;
  assign n8611 = n68364 & n8610 ;
  assign n8612 = n8528 | n8611 ;
  assign n8613 = n68367 & n8612 ;
  assign n8614 = n8533 | n8613 ;
  assign n8616 = n68368 & n8614 ;
  assign n8863 = n8540 | n8616 ;
  assign n9045 = n8122 | n8547 ;
  assign n68376 = ~n9045 ;
  assign n9046 = n8863 & n68376 ;
  assign n9047 = n9044 | n9046 ;
  assign n9048 = n8551 | n9047 ;
  assign n68377 = ~n8553 ;
  assign n9049 = n68377 & n9048 ;
  assign n9057 = n65696 & n9049 ;
  assign n8554 = n8121 & n8551 ;
  assign n8541 = n8130 | n8540 ;
  assign n68378 = ~n8541 ;
  assign n8615 = n68378 & n8614 ;
  assign n68379 = ~n8616 ;
  assign n8617 = n8540 & n68379 ;
  assign n8618 = n8615 | n8617 ;
  assign n8619 = n65696 & n8618 ;
  assign n68380 = ~n8550 ;
  assign n8620 = n68380 & n8619 ;
  assign n8621 = n8554 | n8620 ;
  assign n8622 = n68214 & n8621 ;
  assign n8623 = n8129 & n8551 ;
  assign n8534 = n8138 | n8533 ;
  assign n68381 = ~n8534 ;
  assign n8624 = n8530 & n68381 ;
  assign n68382 = ~n8535 ;
  assign n8625 = n8533 & n68382 ;
  assign n8626 = n8624 | n8625 ;
  assign n8627 = n65696 & n8626 ;
  assign n8628 = n68380 & n8627 ;
  assign n8629 = n8623 | n8628 ;
  assign n8630 = n68058 & n8629 ;
  assign n8631 = n8137 & n8551 ;
  assign n8529 = n8146 | n8528 ;
  assign n68383 = ~n8529 ;
  assign n8632 = n68383 & n8610 ;
  assign n68384 = ~n8611 ;
  assign n8633 = n8528 & n68384 ;
  assign n8634 = n8632 | n8633 ;
  assign n8635 = n65696 & n8634 ;
  assign n8636 = n68380 & n8635 ;
  assign n8637 = n8631 | n8636 ;
  assign n8638 = n67986 & n8637 ;
  assign n8639 = n8145 & n8551 ;
  assign n8522 = n8154 | n8521 ;
  assign n68385 = ~n8522 ;
  assign n8640 = n8518 & n68385 ;
  assign n68386 = ~n8523 ;
  assign n8641 = n8521 & n68386 ;
  assign n8642 = n8640 | n8641 ;
  assign n8643 = n65696 & n8642 ;
  assign n8644 = n68380 & n8643 ;
  assign n8645 = n8639 | n8644 ;
  assign n8646 = n67763 & n8645 ;
  assign n8647 = n8153 & n8551 ;
  assign n8517 = n8162 | n8516 ;
  assign n68387 = ~n8517 ;
  assign n8648 = n68387 & n8606 ;
  assign n68388 = ~n8607 ;
  assign n8649 = n8516 & n68388 ;
  assign n8650 = n8648 | n8649 ;
  assign n8651 = n65696 & n8650 ;
  assign n8652 = n68380 & n8651 ;
  assign n8653 = n8647 | n8652 ;
  assign n8654 = n67622 & n8653 ;
  assign n8655 = n8161 & n8551 ;
  assign n8510 = n8170 | n8509 ;
  assign n68389 = ~n8510 ;
  assign n8656 = n8506 & n68389 ;
  assign n68390 = ~n8511 ;
  assign n8657 = n8509 & n68390 ;
  assign n8658 = n8656 | n8657 ;
  assign n8659 = n65696 & n8658 ;
  assign n8660 = n68380 & n8659 ;
  assign n8661 = n8655 | n8660 ;
  assign n8662 = n67531 & n8661 ;
  assign n8663 = n8169 & n8551 ;
  assign n8505 = n8178 | n8504 ;
  assign n68391 = ~n8505 ;
  assign n8664 = n68391 & n8602 ;
  assign n68392 = ~n8603 ;
  assign n8665 = n8504 & n68392 ;
  assign n8666 = n8664 | n8665 ;
  assign n8667 = n65696 & n8666 ;
  assign n8668 = n68380 & n8667 ;
  assign n8669 = n8663 | n8668 ;
  assign n8670 = n67348 & n8669 ;
  assign n8671 = n8177 & n8551 ;
  assign n8498 = n8186 | n8497 ;
  assign n68393 = ~n8498 ;
  assign n8672 = n8494 & n68393 ;
  assign n68394 = ~n8499 ;
  assign n8673 = n8497 & n68394 ;
  assign n8674 = n8672 | n8673 ;
  assign n8675 = n65696 & n8674 ;
  assign n8676 = n68380 & n8675 ;
  assign n8677 = n8671 | n8676 ;
  assign n8678 = n67222 & n8677 ;
  assign n8679 = n8185 & n8551 ;
  assign n8493 = n8194 | n8492 ;
  assign n68395 = ~n8493 ;
  assign n8680 = n68395 & n8598 ;
  assign n68396 = ~n8599 ;
  assign n8681 = n8492 & n68396 ;
  assign n8682 = n8680 | n8681 ;
  assign n8683 = n65696 & n8682 ;
  assign n8684 = n68380 & n8683 ;
  assign n8685 = n8679 | n8684 ;
  assign n8686 = n67164 & n8685 ;
  assign n8687 = n8193 & n8551 ;
  assign n8486 = n8202 | n8485 ;
  assign n68397 = ~n8486 ;
  assign n8688 = n8482 & n68397 ;
  assign n68398 = ~n8487 ;
  assign n8689 = n8485 & n68398 ;
  assign n8690 = n8688 | n8689 ;
  assign n8691 = n65696 & n8690 ;
  assign n8692 = n68380 & n8691 ;
  assign n8693 = n8687 | n8692 ;
  assign n8694 = n66979 & n8693 ;
  assign n8695 = n8201 & n8551 ;
  assign n8481 = n8210 | n8480 ;
  assign n68399 = ~n8481 ;
  assign n8696 = n68399 & n8594 ;
  assign n68400 = ~n8595 ;
  assign n8697 = n8480 & n68400 ;
  assign n8698 = n8696 | n8697 ;
  assign n8699 = n65696 & n8698 ;
  assign n8700 = n68380 & n8699 ;
  assign n8701 = n8695 | n8700 ;
  assign n8702 = n66868 & n8701 ;
  assign n8703 = n8209 & n8551 ;
  assign n8474 = n8218 | n8473 ;
  assign n68401 = ~n8474 ;
  assign n8704 = n8470 & n68401 ;
  assign n68402 = ~n8475 ;
  assign n8705 = n8473 & n68402 ;
  assign n8706 = n8704 | n8705 ;
  assign n8707 = n65696 & n8706 ;
  assign n8708 = n68380 & n8707 ;
  assign n8709 = n8703 | n8708 ;
  assign n8710 = n66797 & n8709 ;
  assign n8711 = n8217 & n8551 ;
  assign n8469 = n8226 | n8468 ;
  assign n68403 = ~n8469 ;
  assign n8712 = n68403 & n8590 ;
  assign n68404 = ~n8591 ;
  assign n8713 = n8468 & n68404 ;
  assign n8714 = n8712 | n8713 ;
  assign n8715 = n65696 & n8714 ;
  assign n8716 = n68380 & n8715 ;
  assign n8717 = n8711 | n8716 ;
  assign n8718 = n66654 & n8717 ;
  assign n8719 = n8225 & n8551 ;
  assign n8462 = n8234 | n8461 ;
  assign n68405 = ~n8462 ;
  assign n8720 = n8458 & n68405 ;
  assign n68406 = ~n8463 ;
  assign n8721 = n8461 & n68406 ;
  assign n8722 = n8720 | n8721 ;
  assign n8723 = n65696 & n8722 ;
  assign n8724 = n68380 & n8723 ;
  assign n8725 = n8719 | n8724 ;
  assign n8726 = n66560 & n8725 ;
  assign n8727 = n8233 & n8551 ;
  assign n8457 = n8242 | n8456 ;
  assign n68407 = ~n8457 ;
  assign n8728 = n68407 & n8586 ;
  assign n68408 = ~n8587 ;
  assign n8729 = n8456 & n68408 ;
  assign n8730 = n8728 | n8729 ;
  assign n8731 = n65696 & n8730 ;
  assign n8732 = n68380 & n8731 ;
  assign n8733 = n8727 | n8732 ;
  assign n8734 = n66505 & n8733 ;
  assign n8735 = n8241 & n8551 ;
  assign n8450 = n8250 | n8449 ;
  assign n68409 = ~n8450 ;
  assign n8736 = n8446 & n68409 ;
  assign n68410 = ~n8451 ;
  assign n8737 = n8449 & n68410 ;
  assign n8738 = n8736 | n8737 ;
  assign n8739 = n65696 & n8738 ;
  assign n8740 = n68380 & n8739 ;
  assign n8741 = n8735 | n8740 ;
  assign n8742 = n66379 & n8741 ;
  assign n8743 = n8249 & n8551 ;
  assign n8445 = n8258 | n8444 ;
  assign n68411 = ~n8445 ;
  assign n8744 = n68411 & n8582 ;
  assign n68412 = ~n8583 ;
  assign n8745 = n8444 & n68412 ;
  assign n8746 = n8744 | n8745 ;
  assign n8747 = n65696 & n8746 ;
  assign n8748 = n68380 & n8747 ;
  assign n8749 = n8743 | n8748 ;
  assign n8750 = n66299 & n8749 ;
  assign n8751 = n8257 & n8551 ;
  assign n8438 = n8266 | n8437 ;
  assign n68413 = ~n8438 ;
  assign n8752 = n8434 & n68413 ;
  assign n68414 = ~n8439 ;
  assign n8753 = n8437 & n68414 ;
  assign n8754 = n8752 | n8753 ;
  assign n8755 = n65696 & n8754 ;
  assign n8756 = n68380 & n8755 ;
  assign n8757 = n8751 | n8756 ;
  assign n8758 = n66244 & n8757 ;
  assign n8759 = n8265 & n8551 ;
  assign n8433 = n8274 | n8432 ;
  assign n68415 = ~n8433 ;
  assign n8760 = n68415 & n8578 ;
  assign n68416 = ~n8579 ;
  assign n8761 = n8432 & n68416 ;
  assign n8762 = n8760 | n8761 ;
  assign n8763 = n65696 & n8762 ;
  assign n8764 = n68380 & n8763 ;
  assign n8765 = n8759 | n8764 ;
  assign n8766 = n66145 & n8765 ;
  assign n8767 = n8273 & n8551 ;
  assign n8426 = n8282 | n8425 ;
  assign n68417 = ~n8426 ;
  assign n8768 = n8422 & n68417 ;
  assign n68418 = ~n8427 ;
  assign n8769 = n8425 & n68418 ;
  assign n8770 = n8768 | n8769 ;
  assign n8771 = n65696 & n8770 ;
  assign n8772 = n68380 & n8771 ;
  assign n8773 = n8767 | n8772 ;
  assign n8774 = n66081 & n8773 ;
  assign n8775 = n8281 & n8551 ;
  assign n8421 = n8290 | n8420 ;
  assign n68419 = ~n8421 ;
  assign n8776 = n68419 & n8574 ;
  assign n68420 = ~n8575 ;
  assign n8777 = n8420 & n68420 ;
  assign n8778 = n8776 | n8777 ;
  assign n8779 = n65696 & n8778 ;
  assign n8780 = n68380 & n8779 ;
  assign n8781 = n8775 | n8780 ;
  assign n8782 = n66043 & n8781 ;
  assign n8783 = n8289 & n8551 ;
  assign n8414 = n8298 | n8413 ;
  assign n68421 = ~n8414 ;
  assign n8784 = n8410 & n68421 ;
  assign n68422 = ~n8415 ;
  assign n8785 = n8413 & n68422 ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = n65696 & n8786 ;
  assign n8788 = n68380 & n8787 ;
  assign n8789 = n8783 | n8788 ;
  assign n8790 = n65960 & n8789 ;
  assign n8791 = n8297 & n8551 ;
  assign n8409 = n8306 | n8408 ;
  assign n68423 = ~n8409 ;
  assign n8792 = n68423 & n8570 ;
  assign n68424 = ~n8571 ;
  assign n8793 = n8408 & n68424 ;
  assign n8794 = n8792 | n8793 ;
  assign n8795 = n65696 & n8794 ;
  assign n8796 = n68380 & n8795 ;
  assign n8797 = n8791 | n8796 ;
  assign n8798 = n65909 & n8797 ;
  assign n8799 = n8305 & n8551 ;
  assign n8402 = n8314 | n8401 ;
  assign n68425 = ~n8402 ;
  assign n8800 = n8398 & n68425 ;
  assign n68426 = ~n8403 ;
  assign n8801 = n8401 & n68426 ;
  assign n8802 = n8800 | n8801 ;
  assign n8803 = n65696 & n8802 ;
  assign n8804 = n68380 & n8803 ;
  assign n8805 = n8799 | n8804 ;
  assign n8806 = n65877 & n8805 ;
  assign n8807 = n8313 & n8551 ;
  assign n8397 = n8322 | n8396 ;
  assign n68427 = ~n8397 ;
  assign n8808 = n8392 & n68427 ;
  assign n68428 = ~n8567 ;
  assign n8809 = n8396 & n68428 ;
  assign n8810 = n8808 | n8809 ;
  assign n8811 = n65696 & n8810 ;
  assign n8812 = n68380 & n8811 ;
  assign n8813 = n8807 | n8812 ;
  assign n8814 = n65820 & n8813 ;
  assign n8815 = n8321 & n8551 ;
  assign n8816 = n8330 | n8390 ;
  assign n68429 = ~n8816 ;
  assign n8817 = n8387 & n68429 ;
  assign n68430 = ~n8391 ;
  assign n8818 = n8390 & n68430 ;
  assign n8819 = n8817 | n8818 ;
  assign n8820 = n65696 & n8819 ;
  assign n8821 = n68380 & n8820 ;
  assign n8822 = n8815 | n8821 ;
  assign n8823 = n65791 & n8822 ;
  assign n8824 = n8329 & n8551 ;
  assign n8825 = n8339 | n8386 ;
  assign n68431 = ~n8825 ;
  assign n8826 = n8382 & n68431 ;
  assign n68432 = ~n8563 ;
  assign n8827 = n8386 & n68432 ;
  assign n8828 = n8826 | n8827 ;
  assign n8829 = n65696 & n8828 ;
  assign n8830 = n68380 & n8829 ;
  assign n8831 = n8824 | n8830 ;
  assign n8832 = n65772 & n8831 ;
  assign n8833 = n8338 & n8551 ;
  assign n8834 = n8347 | n8380 ;
  assign n68433 = ~n8834 ;
  assign n8835 = n8377 & n68433 ;
  assign n68434 = ~n8381 ;
  assign n8836 = n8380 & n68434 ;
  assign n8837 = n8835 | n8836 ;
  assign n8838 = n65696 & n8837 ;
  assign n8839 = n68380 & n8838 ;
  assign n8840 = n8833 | n8839 ;
  assign n8841 = n65746 & n8840 ;
  assign n8842 = n8346 & n8551 ;
  assign n68435 = ~n8373 ;
  assign n8843 = n68435 & n8376 ;
  assign n8844 = n8372 | n8376 ;
  assign n68436 = ~n8844 ;
  assign n8845 = n8370 & n68436 ;
  assign n8846 = n8843 | n8845 ;
  assign n8847 = n65696 & n8846 ;
  assign n8848 = n68380 & n8847 ;
  assign n8849 = n8842 | n8848 ;
  assign n8850 = n65721 & n8849 ;
  assign n8552 = n8371 & n8551 ;
  assign n8557 = n8367 & n8368 ;
  assign n8851 = n68311 & n8557 ;
  assign n8852 = n303 | n8851 ;
  assign n68437 = ~n8852 ;
  assign n8853 = n8370 & n68437 ;
  assign n8854 = n68380 & n8853 ;
  assign n8855 = n8552 | n8854 ;
  assign n8856 = n65686 & n8855 ;
  assign n68438 = ~x96 ;
  assign n8857 = x64 & n68438 ;
  assign n8858 = n68308 & n8857 ;
  assign n8859 = n67025 & n8858 ;
  assign n8860 = n67026 & n8859 ;
  assign n8864 = n68371 & n8863 ;
  assign n8865 = n8547 | n8864 ;
  assign n8866 = n68372 & n8865 ;
  assign n68439 = ~n8866 ;
  assign n8867 = n8860 & n68439 ;
  assign n68440 = ~n8867 ;
  assign n8868 = x32 & n68440 ;
  assign n8869 = n67988 & n8368 ;
  assign n8870 = n67020 & n8869 ;
  assign n8871 = n67021 & n8870 ;
  assign n8872 = n68380 & n8871 ;
  assign n8873 = n8868 | n8872 ;
  assign n8875 = x65 & n8873 ;
  assign n8861 = n68380 & n8860 ;
  assign n68441 = ~n8861 ;
  assign n8862 = x32 & n68441 ;
  assign n8874 = x65 | n8872 ;
  assign n8876 = n8862 | n8874 ;
  assign n68442 = ~n8875 ;
  assign n8877 = n68442 & n8876 ;
  assign n68443 = ~x31 ;
  assign n8878 = n68443 & x64 ;
  assign n8879 = n8877 | n8878 ;
  assign n8880 = n65670 & n8873 ;
  assign n68444 = ~n8880 ;
  assign n8881 = n8879 & n68444 ;
  assign n68445 = ~n8854 ;
  assign n8882 = x66 & n68445 ;
  assign n68446 = ~n8552 ;
  assign n8883 = n68446 & n8882 ;
  assign n8884 = n8856 | n8883 ;
  assign n8885 = n8881 | n8884 ;
  assign n68447 = ~n8856 ;
  assign n8886 = n68447 & n8885 ;
  assign n68448 = ~n8848 ;
  assign n8887 = x67 & n68448 ;
  assign n68449 = ~n8842 ;
  assign n8888 = n68449 & n8887 ;
  assign n8889 = n8886 | n8888 ;
  assign n68450 = ~n8850 ;
  assign n8890 = n68450 & n8889 ;
  assign n68451 = ~n8839 ;
  assign n8891 = x68 & n68451 ;
  assign n68452 = ~n8833 ;
  assign n8892 = n68452 & n8891 ;
  assign n8893 = n8841 | n8892 ;
  assign n8894 = n8890 | n8893 ;
  assign n68453 = ~n8841 ;
  assign n8895 = n68453 & n8894 ;
  assign n68454 = ~n8830 ;
  assign n8896 = x69 & n68454 ;
  assign n68455 = ~n8824 ;
  assign n8897 = n68455 & n8896 ;
  assign n8898 = n8832 | n8897 ;
  assign n8899 = n8895 | n8898 ;
  assign n68456 = ~n8832 ;
  assign n8900 = n68456 & n8899 ;
  assign n68457 = ~n8821 ;
  assign n8901 = x70 & n68457 ;
  assign n68458 = ~n8815 ;
  assign n8902 = n68458 & n8901 ;
  assign n8903 = n8823 | n8902 ;
  assign n8904 = n8900 | n8903 ;
  assign n68459 = ~n8823 ;
  assign n8905 = n68459 & n8904 ;
  assign n68460 = ~n8812 ;
  assign n8906 = x71 & n68460 ;
  assign n68461 = ~n8807 ;
  assign n8907 = n68461 & n8906 ;
  assign n8908 = n8814 | n8907 ;
  assign n8910 = n8905 | n8908 ;
  assign n68462 = ~n8814 ;
  assign n8911 = n68462 & n8910 ;
  assign n68463 = ~n8804 ;
  assign n8912 = x72 & n68463 ;
  assign n68464 = ~n8799 ;
  assign n8913 = n68464 & n8912 ;
  assign n8914 = n8806 | n8913 ;
  assign n8915 = n8911 | n8914 ;
  assign n68465 = ~n8806 ;
  assign n8916 = n68465 & n8915 ;
  assign n68466 = ~n8796 ;
  assign n8917 = x73 & n68466 ;
  assign n68467 = ~n8791 ;
  assign n8918 = n68467 & n8917 ;
  assign n8919 = n8798 | n8918 ;
  assign n8921 = n8916 | n8919 ;
  assign n68468 = ~n8798 ;
  assign n8922 = n68468 & n8921 ;
  assign n68469 = ~n8788 ;
  assign n8923 = x74 & n68469 ;
  assign n68470 = ~n8783 ;
  assign n8924 = n68470 & n8923 ;
  assign n8925 = n8790 | n8924 ;
  assign n8926 = n8922 | n8925 ;
  assign n68471 = ~n8790 ;
  assign n8927 = n68471 & n8926 ;
  assign n68472 = ~n8780 ;
  assign n8928 = x75 & n68472 ;
  assign n68473 = ~n8775 ;
  assign n8929 = n68473 & n8928 ;
  assign n8930 = n8782 | n8929 ;
  assign n8932 = n8927 | n8930 ;
  assign n68474 = ~n8782 ;
  assign n8933 = n68474 & n8932 ;
  assign n68475 = ~n8772 ;
  assign n8934 = x76 & n68475 ;
  assign n68476 = ~n8767 ;
  assign n8935 = n68476 & n8934 ;
  assign n8936 = n8774 | n8935 ;
  assign n8937 = n8933 | n8936 ;
  assign n68477 = ~n8774 ;
  assign n8938 = n68477 & n8937 ;
  assign n68478 = ~n8764 ;
  assign n8939 = x77 & n68478 ;
  assign n68479 = ~n8759 ;
  assign n8940 = n68479 & n8939 ;
  assign n8941 = n8766 | n8940 ;
  assign n8943 = n8938 | n8941 ;
  assign n68480 = ~n8766 ;
  assign n8944 = n68480 & n8943 ;
  assign n68481 = ~n8756 ;
  assign n8945 = x78 & n68481 ;
  assign n68482 = ~n8751 ;
  assign n8946 = n68482 & n8945 ;
  assign n8947 = n8758 | n8946 ;
  assign n8948 = n8944 | n8947 ;
  assign n68483 = ~n8758 ;
  assign n8949 = n68483 & n8948 ;
  assign n68484 = ~n8748 ;
  assign n8950 = x79 & n68484 ;
  assign n68485 = ~n8743 ;
  assign n8951 = n68485 & n8950 ;
  assign n8952 = n8750 | n8951 ;
  assign n8954 = n8949 | n8952 ;
  assign n68486 = ~n8750 ;
  assign n8955 = n68486 & n8954 ;
  assign n68487 = ~n8740 ;
  assign n8956 = x80 & n68487 ;
  assign n68488 = ~n8735 ;
  assign n8957 = n68488 & n8956 ;
  assign n8958 = n8742 | n8957 ;
  assign n8959 = n8955 | n8958 ;
  assign n68489 = ~n8742 ;
  assign n8960 = n68489 & n8959 ;
  assign n68490 = ~n8732 ;
  assign n8961 = x81 & n68490 ;
  assign n68491 = ~n8727 ;
  assign n8962 = n68491 & n8961 ;
  assign n8963 = n8734 | n8962 ;
  assign n8965 = n8960 | n8963 ;
  assign n68492 = ~n8734 ;
  assign n8966 = n68492 & n8965 ;
  assign n68493 = ~n8724 ;
  assign n8967 = x82 & n68493 ;
  assign n68494 = ~n8719 ;
  assign n8968 = n68494 & n8967 ;
  assign n8969 = n8726 | n8968 ;
  assign n8970 = n8966 | n8969 ;
  assign n68495 = ~n8726 ;
  assign n8971 = n68495 & n8970 ;
  assign n68496 = ~n8716 ;
  assign n8972 = x83 & n68496 ;
  assign n68497 = ~n8711 ;
  assign n8973 = n68497 & n8972 ;
  assign n8974 = n8718 | n8973 ;
  assign n8976 = n8971 | n8974 ;
  assign n68498 = ~n8718 ;
  assign n8977 = n68498 & n8976 ;
  assign n68499 = ~n8708 ;
  assign n8978 = x84 & n68499 ;
  assign n68500 = ~n8703 ;
  assign n8979 = n68500 & n8978 ;
  assign n8980 = n8710 | n8979 ;
  assign n8981 = n8977 | n8980 ;
  assign n68501 = ~n8710 ;
  assign n8982 = n68501 & n8981 ;
  assign n68502 = ~n8700 ;
  assign n8983 = x85 & n68502 ;
  assign n68503 = ~n8695 ;
  assign n8984 = n68503 & n8983 ;
  assign n8985 = n8702 | n8984 ;
  assign n8987 = n8982 | n8985 ;
  assign n68504 = ~n8702 ;
  assign n8988 = n68504 & n8987 ;
  assign n68505 = ~n8692 ;
  assign n8989 = x86 & n68505 ;
  assign n68506 = ~n8687 ;
  assign n8990 = n68506 & n8989 ;
  assign n8991 = n8694 | n8990 ;
  assign n8992 = n8988 | n8991 ;
  assign n68507 = ~n8694 ;
  assign n8993 = n68507 & n8992 ;
  assign n68508 = ~n8684 ;
  assign n8994 = x87 & n68508 ;
  assign n68509 = ~n8679 ;
  assign n8995 = n68509 & n8994 ;
  assign n8996 = n8686 | n8995 ;
  assign n8998 = n8993 | n8996 ;
  assign n68510 = ~n8686 ;
  assign n8999 = n68510 & n8998 ;
  assign n68511 = ~n8676 ;
  assign n9000 = x88 & n68511 ;
  assign n68512 = ~n8671 ;
  assign n9001 = n68512 & n9000 ;
  assign n9002 = n8678 | n9001 ;
  assign n9003 = n8999 | n9002 ;
  assign n68513 = ~n8678 ;
  assign n9004 = n68513 & n9003 ;
  assign n68514 = ~n8668 ;
  assign n9005 = x89 & n68514 ;
  assign n68515 = ~n8663 ;
  assign n9006 = n68515 & n9005 ;
  assign n9007 = n8670 | n9006 ;
  assign n9009 = n9004 | n9007 ;
  assign n68516 = ~n8670 ;
  assign n9010 = n68516 & n9009 ;
  assign n68517 = ~n8660 ;
  assign n9011 = x90 & n68517 ;
  assign n68518 = ~n8655 ;
  assign n9012 = n68518 & n9011 ;
  assign n9013 = n8662 | n9012 ;
  assign n9014 = n9010 | n9013 ;
  assign n68519 = ~n8662 ;
  assign n9015 = n68519 & n9014 ;
  assign n68520 = ~n8652 ;
  assign n9016 = x91 & n68520 ;
  assign n68521 = ~n8647 ;
  assign n9017 = n68521 & n9016 ;
  assign n9018 = n8654 | n9017 ;
  assign n9020 = n9015 | n9018 ;
  assign n68522 = ~n8654 ;
  assign n9021 = n68522 & n9020 ;
  assign n68523 = ~n8644 ;
  assign n9022 = x92 & n68523 ;
  assign n68524 = ~n8639 ;
  assign n9023 = n68524 & n9022 ;
  assign n9024 = n8646 | n9023 ;
  assign n9025 = n9021 | n9024 ;
  assign n68525 = ~n8646 ;
  assign n9026 = n68525 & n9025 ;
  assign n68526 = ~n8636 ;
  assign n9027 = x93 & n68526 ;
  assign n68527 = ~n8631 ;
  assign n9028 = n68527 & n9027 ;
  assign n9029 = n8638 | n9028 ;
  assign n9031 = n9026 | n9029 ;
  assign n68528 = ~n8638 ;
  assign n9032 = n68528 & n9031 ;
  assign n68529 = ~n8628 ;
  assign n9033 = x94 & n68529 ;
  assign n68530 = ~n8623 ;
  assign n9034 = n68530 & n9033 ;
  assign n9035 = n8630 | n9034 ;
  assign n9036 = n9032 | n9035 ;
  assign n68531 = ~n8630 ;
  assign n9037 = n68531 & n9036 ;
  assign n68532 = ~n8620 ;
  assign n9038 = x95 & n68532 ;
  assign n68533 = ~n8554 ;
  assign n9039 = n68533 & n9038 ;
  assign n9040 = n8622 | n9039 ;
  assign n9042 = n9037 | n9040 ;
  assign n68534 = ~n8622 ;
  assign n9043 = n68534 & n9042 ;
  assign n9050 = n68438 & n9049 ;
  assign n161 = ~n8551 ;
  assign n9051 = n161 & n9047 ;
  assign n9052 = n8113 & n8551 ;
  assign n68536 = ~n9052 ;
  assign n9053 = x96 & n68536 ;
  assign n68537 = ~n9051 ;
  assign n9054 = n68537 & n9053 ;
  assign n9055 = n295 | n9054 ;
  assign n9056 = n9050 | n9055 ;
  assign n9058 = n9043 | n9056 ;
  assign n68538 = ~n9057 ;
  assign n9059 = n68538 & n9058 ;
  assign n68539 = ~n9037 ;
  assign n9041 = n68539 & n9040 ;
  assign n9062 = n8862 | n8872 ;
  assign n9063 = x65 & n9062 ;
  assign n68540 = ~n9063 ;
  assign n9064 = n8876 & n68540 ;
  assign n9065 = n8878 | n9064 ;
  assign n9066 = n68444 & n9065 ;
  assign n9068 = n8883 | n9066 ;
  assign n9069 = n68447 & n9068 ;
  assign n9070 = n8850 | n8888 ;
  assign n9072 = n9069 | n9070 ;
  assign n9073 = n68450 & n9072 ;
  assign n9075 = n8893 | n9073 ;
  assign n9076 = n68453 & n9075 ;
  assign n9078 = n8898 | n9076 ;
  assign n9079 = n68456 & n9078 ;
  assign n9080 = n8903 | n9079 ;
  assign n9082 = n68459 & n9080 ;
  assign n9083 = n8908 | n9082 ;
  assign n9084 = n68462 & n9083 ;
  assign n9085 = n8914 | n9084 ;
  assign n9087 = n68465 & n9085 ;
  assign n9088 = n8919 | n9087 ;
  assign n9089 = n68468 & n9088 ;
  assign n9090 = n8925 | n9089 ;
  assign n9092 = n68471 & n9090 ;
  assign n9093 = n8930 | n9092 ;
  assign n9094 = n68474 & n9093 ;
  assign n9095 = n8936 | n9094 ;
  assign n9097 = n68477 & n9095 ;
  assign n9098 = n8941 | n9097 ;
  assign n9099 = n68480 & n9098 ;
  assign n9100 = n8947 | n9099 ;
  assign n9102 = n68483 & n9100 ;
  assign n9103 = n8952 | n9102 ;
  assign n9104 = n68486 & n9103 ;
  assign n9105 = n8958 | n9104 ;
  assign n9107 = n68489 & n9105 ;
  assign n9108 = n8963 | n9107 ;
  assign n9109 = n68492 & n9108 ;
  assign n9110 = n8969 | n9109 ;
  assign n9112 = n68495 & n9110 ;
  assign n9113 = n8974 | n9112 ;
  assign n9114 = n68498 & n9113 ;
  assign n9115 = n8980 | n9114 ;
  assign n9117 = n68501 & n9115 ;
  assign n9118 = n8985 | n9117 ;
  assign n9119 = n68504 & n9118 ;
  assign n9120 = n8991 | n9119 ;
  assign n9122 = n68507 & n9120 ;
  assign n9123 = n8996 | n9122 ;
  assign n9124 = n68510 & n9123 ;
  assign n9125 = n9002 | n9124 ;
  assign n9127 = n68513 & n9125 ;
  assign n9128 = n9007 | n9127 ;
  assign n9129 = n68516 & n9128 ;
  assign n9130 = n9013 | n9129 ;
  assign n9132 = n68519 & n9130 ;
  assign n9133 = n9018 | n9132 ;
  assign n9134 = n68522 & n9133 ;
  assign n9135 = n9024 | n9134 ;
  assign n9137 = n68525 & n9135 ;
  assign n9138 = n9029 | n9137 ;
  assign n9139 = n68528 & n9138 ;
  assign n9140 = n9035 | n9139 ;
  assign n9157 = n8630 | n9040 ;
  assign n68541 = ~n9157 ;
  assign n9158 = n9140 & n68541 ;
  assign n9159 = n9041 | n9158 ;
  assign n160 = ~n9059 ;
  assign n9160 = n160 & n9159 ;
  assign n9142 = n68531 & n9140 ;
  assign n9143 = n9040 | n9142 ;
  assign n9144 = n68534 & n9143 ;
  assign n9145 = n9056 | n9144 ;
  assign n9161 = n8621 & n68538 ;
  assign n9162 = n9145 & n9161 ;
  assign n9163 = n9160 | n9162 ;
  assign n9146 = n8622 | n9054 ;
  assign n9147 = n9050 | n9146 ;
  assign n68543 = ~n9147 ;
  assign n9148 = n9042 & n68543 ;
  assign n9149 = n9050 | n9054 ;
  assign n68544 = ~n9144 ;
  assign n9150 = n68544 & n9149 ;
  assign n9151 = n9148 | n9150 ;
  assign n9152 = n160 & n9151 ;
  assign n9153 = n303 & n8113 ;
  assign n9154 = n9145 & n9153 ;
  assign n9155 = n9152 | n9154 ;
  assign n68545 = ~x97 ;
  assign n9156 = n68545 & n9155 ;
  assign n68546 = ~n9154 ;
  assign n9602 = x97 & n68546 ;
  assign n68547 = ~n9152 ;
  assign n9603 = n68547 & n9602 ;
  assign n9604 = n9156 | n9603 ;
  assign n9164 = n68438 & n9163 ;
  assign n68548 = ~n9139 ;
  assign n9141 = n9035 & n68548 ;
  assign n9165 = n8638 | n9035 ;
  assign n68549 = ~n9165 ;
  assign n9166 = n9031 & n68549 ;
  assign n9167 = n9141 | n9166 ;
  assign n9168 = n160 & n9167 ;
  assign n9169 = n8629 & n68538 ;
  assign n9170 = n9145 & n9169 ;
  assign n9171 = n9168 | n9170 ;
  assign n9172 = n68214 & n9171 ;
  assign n68550 = ~n9170 ;
  assign n9590 = x95 & n68550 ;
  assign n68551 = ~n9168 ;
  assign n9591 = n68551 & n9590 ;
  assign n9592 = n9172 | n9591 ;
  assign n68552 = ~n9026 ;
  assign n9030 = n68552 & n9029 ;
  assign n9173 = n8646 | n9029 ;
  assign n68553 = ~n9173 ;
  assign n9174 = n9135 & n68553 ;
  assign n9175 = n9030 | n9174 ;
  assign n9176 = n160 & n9175 ;
  assign n9177 = n8637 & n68538 ;
  assign n9178 = n9145 & n9177 ;
  assign n9179 = n9176 | n9178 ;
  assign n9180 = n68058 & n9179 ;
  assign n68554 = ~n9134 ;
  assign n9136 = n9024 & n68554 ;
  assign n9181 = n8654 | n9024 ;
  assign n68555 = ~n9181 ;
  assign n9182 = n9020 & n68555 ;
  assign n9183 = n9136 | n9182 ;
  assign n9184 = n160 & n9183 ;
  assign n9185 = n8645 & n68538 ;
  assign n9186 = n9145 & n9185 ;
  assign n9187 = n9184 | n9186 ;
  assign n9188 = n67986 & n9187 ;
  assign n68556 = ~n9186 ;
  assign n9578 = x93 & n68556 ;
  assign n68557 = ~n9184 ;
  assign n9579 = n68557 & n9578 ;
  assign n9580 = n9188 | n9579 ;
  assign n68558 = ~n9015 ;
  assign n9019 = n68558 & n9018 ;
  assign n9189 = n8662 | n9018 ;
  assign n68559 = ~n9189 ;
  assign n9190 = n9130 & n68559 ;
  assign n9191 = n9019 | n9190 ;
  assign n9192 = n160 & n9191 ;
  assign n9193 = n8653 & n68538 ;
  assign n9194 = n9145 & n9193 ;
  assign n9195 = n9192 | n9194 ;
  assign n9196 = n67763 & n9195 ;
  assign n68560 = ~n9129 ;
  assign n9131 = n9013 & n68560 ;
  assign n9197 = n8670 | n9013 ;
  assign n68561 = ~n9197 ;
  assign n9198 = n9009 & n68561 ;
  assign n9199 = n9131 | n9198 ;
  assign n9200 = n160 & n9199 ;
  assign n9201 = n8661 & n68538 ;
  assign n9202 = n9145 & n9201 ;
  assign n9203 = n9200 | n9202 ;
  assign n9204 = n67622 & n9203 ;
  assign n68562 = ~n9202 ;
  assign n9566 = x91 & n68562 ;
  assign n68563 = ~n9200 ;
  assign n9567 = n68563 & n9566 ;
  assign n9568 = n9204 | n9567 ;
  assign n68564 = ~n9004 ;
  assign n9008 = n68564 & n9007 ;
  assign n9205 = n8678 | n9007 ;
  assign n68565 = ~n9205 ;
  assign n9206 = n9125 & n68565 ;
  assign n9207 = n9008 | n9206 ;
  assign n9208 = n160 & n9207 ;
  assign n9209 = n8669 & n68538 ;
  assign n9210 = n9145 & n9209 ;
  assign n9211 = n9208 | n9210 ;
  assign n9212 = n67531 & n9211 ;
  assign n68566 = ~n9124 ;
  assign n9126 = n9002 & n68566 ;
  assign n9213 = n8686 | n9002 ;
  assign n68567 = ~n9213 ;
  assign n9214 = n8998 & n68567 ;
  assign n9215 = n9126 | n9214 ;
  assign n9216 = n160 & n9215 ;
  assign n9217 = n8677 & n68538 ;
  assign n9218 = n9145 & n9217 ;
  assign n9219 = n9216 | n9218 ;
  assign n9220 = n67348 & n9219 ;
  assign n68568 = ~n9218 ;
  assign n9554 = x89 & n68568 ;
  assign n68569 = ~n9216 ;
  assign n9555 = n68569 & n9554 ;
  assign n9556 = n9220 | n9555 ;
  assign n68570 = ~n8993 ;
  assign n8997 = n68570 & n8996 ;
  assign n9221 = n8694 | n8996 ;
  assign n68571 = ~n9221 ;
  assign n9222 = n9120 & n68571 ;
  assign n9223 = n8997 | n9222 ;
  assign n9224 = n160 & n9223 ;
  assign n9225 = n8685 & n68538 ;
  assign n9226 = n9145 & n9225 ;
  assign n9227 = n9224 | n9226 ;
  assign n9228 = n67222 & n9227 ;
  assign n68572 = ~n9119 ;
  assign n9121 = n8991 & n68572 ;
  assign n9229 = n8702 | n8991 ;
  assign n68573 = ~n9229 ;
  assign n9230 = n8987 & n68573 ;
  assign n9231 = n9121 | n9230 ;
  assign n9232 = n160 & n9231 ;
  assign n9233 = n8693 & n68538 ;
  assign n9234 = n9145 & n9233 ;
  assign n9235 = n9232 | n9234 ;
  assign n9236 = n67164 & n9235 ;
  assign n68574 = ~n9234 ;
  assign n9542 = x87 & n68574 ;
  assign n68575 = ~n9232 ;
  assign n9543 = n68575 & n9542 ;
  assign n9544 = n9236 | n9543 ;
  assign n68576 = ~n8982 ;
  assign n8986 = n68576 & n8985 ;
  assign n9237 = n8710 | n8985 ;
  assign n68577 = ~n9237 ;
  assign n9238 = n9115 & n68577 ;
  assign n9239 = n8986 | n9238 ;
  assign n9240 = n160 & n9239 ;
  assign n9241 = n8701 & n68538 ;
  assign n9242 = n9145 & n9241 ;
  assign n9243 = n9240 | n9242 ;
  assign n9244 = n66979 & n9243 ;
  assign n68578 = ~n9114 ;
  assign n9116 = n8980 & n68578 ;
  assign n9245 = n8718 | n8980 ;
  assign n68579 = ~n9245 ;
  assign n9246 = n8976 & n68579 ;
  assign n9247 = n9116 | n9246 ;
  assign n9248 = n160 & n9247 ;
  assign n9249 = n8709 & n68538 ;
  assign n9250 = n9145 & n9249 ;
  assign n9251 = n9248 | n9250 ;
  assign n9252 = n66868 & n9251 ;
  assign n68580 = ~n9250 ;
  assign n9530 = x85 & n68580 ;
  assign n68581 = ~n9248 ;
  assign n9531 = n68581 & n9530 ;
  assign n9532 = n9252 | n9531 ;
  assign n68582 = ~n8971 ;
  assign n8975 = n68582 & n8974 ;
  assign n9253 = n8726 | n8974 ;
  assign n68583 = ~n9253 ;
  assign n9254 = n9110 & n68583 ;
  assign n9255 = n8975 | n9254 ;
  assign n9256 = n160 & n9255 ;
  assign n9257 = n8717 & n68538 ;
  assign n9258 = n9145 & n9257 ;
  assign n9259 = n9256 | n9258 ;
  assign n9260 = n66797 & n9259 ;
  assign n68584 = ~n9109 ;
  assign n9111 = n8969 & n68584 ;
  assign n9261 = n8734 | n8969 ;
  assign n68585 = ~n9261 ;
  assign n9262 = n8965 & n68585 ;
  assign n9263 = n9111 | n9262 ;
  assign n9264 = n160 & n9263 ;
  assign n9265 = n8725 & n68538 ;
  assign n9266 = n9145 & n9265 ;
  assign n9267 = n9264 | n9266 ;
  assign n9268 = n66654 & n9267 ;
  assign n68586 = ~n9266 ;
  assign n9518 = x83 & n68586 ;
  assign n68587 = ~n9264 ;
  assign n9519 = n68587 & n9518 ;
  assign n9520 = n9268 | n9519 ;
  assign n68588 = ~n8960 ;
  assign n8964 = n68588 & n8963 ;
  assign n9269 = n8742 | n8963 ;
  assign n68589 = ~n9269 ;
  assign n9270 = n9105 & n68589 ;
  assign n9271 = n8964 | n9270 ;
  assign n9272 = n160 & n9271 ;
  assign n9273 = n8733 & n68538 ;
  assign n9274 = n9145 & n9273 ;
  assign n9275 = n9272 | n9274 ;
  assign n9276 = n66560 & n9275 ;
  assign n68590 = ~n9104 ;
  assign n9106 = n8958 & n68590 ;
  assign n9277 = n8750 | n8958 ;
  assign n68591 = ~n9277 ;
  assign n9278 = n8954 & n68591 ;
  assign n9279 = n9106 | n9278 ;
  assign n9280 = n160 & n9279 ;
  assign n9281 = n8741 & n68538 ;
  assign n9282 = n9145 & n9281 ;
  assign n9283 = n9280 | n9282 ;
  assign n9284 = n66505 & n9283 ;
  assign n68592 = ~n9282 ;
  assign n9506 = x81 & n68592 ;
  assign n68593 = ~n9280 ;
  assign n9507 = n68593 & n9506 ;
  assign n9508 = n9284 | n9507 ;
  assign n68594 = ~n8949 ;
  assign n8953 = n68594 & n8952 ;
  assign n9285 = n8758 | n8952 ;
  assign n68595 = ~n9285 ;
  assign n9286 = n9100 & n68595 ;
  assign n9287 = n8953 | n9286 ;
  assign n9288 = n160 & n9287 ;
  assign n9289 = n8749 & n68538 ;
  assign n9290 = n9145 & n9289 ;
  assign n9291 = n9288 | n9290 ;
  assign n9292 = n66379 & n9291 ;
  assign n68596 = ~n9099 ;
  assign n9101 = n8947 & n68596 ;
  assign n9293 = n8766 | n8947 ;
  assign n68597 = ~n9293 ;
  assign n9294 = n8943 & n68597 ;
  assign n9295 = n9101 | n9294 ;
  assign n9296 = n160 & n9295 ;
  assign n9297 = n8757 & n68538 ;
  assign n9298 = n9145 & n9297 ;
  assign n9299 = n9296 | n9298 ;
  assign n9300 = n66299 & n9299 ;
  assign n68598 = ~n9298 ;
  assign n9494 = x79 & n68598 ;
  assign n68599 = ~n9296 ;
  assign n9495 = n68599 & n9494 ;
  assign n9496 = n9300 | n9495 ;
  assign n68600 = ~n8938 ;
  assign n8942 = n68600 & n8941 ;
  assign n9301 = n8774 | n8941 ;
  assign n68601 = ~n9301 ;
  assign n9302 = n9095 & n68601 ;
  assign n9303 = n8942 | n9302 ;
  assign n9304 = n160 & n9303 ;
  assign n9305 = n8765 & n68538 ;
  assign n9306 = n9145 & n9305 ;
  assign n9307 = n9304 | n9306 ;
  assign n9308 = n66244 & n9307 ;
  assign n68602 = ~n9094 ;
  assign n9096 = n8936 & n68602 ;
  assign n9309 = n8782 | n8936 ;
  assign n68603 = ~n9309 ;
  assign n9310 = n8932 & n68603 ;
  assign n9311 = n9096 | n9310 ;
  assign n9312 = n160 & n9311 ;
  assign n9313 = n8773 & n68538 ;
  assign n9314 = n9145 & n9313 ;
  assign n9315 = n9312 | n9314 ;
  assign n9316 = n66145 & n9315 ;
  assign n68604 = ~n9314 ;
  assign n9482 = x77 & n68604 ;
  assign n68605 = ~n9312 ;
  assign n9483 = n68605 & n9482 ;
  assign n9484 = n9316 | n9483 ;
  assign n68606 = ~n8927 ;
  assign n8931 = n68606 & n8930 ;
  assign n9317 = n8790 | n8930 ;
  assign n68607 = ~n9317 ;
  assign n9318 = n9090 & n68607 ;
  assign n9319 = n8931 | n9318 ;
  assign n9320 = n160 & n9319 ;
  assign n9321 = n8781 & n68538 ;
  assign n9322 = n9145 & n9321 ;
  assign n9323 = n9320 | n9322 ;
  assign n9324 = n66081 & n9323 ;
  assign n68608 = ~n9089 ;
  assign n9091 = n8925 & n68608 ;
  assign n9325 = n8798 | n8925 ;
  assign n68609 = ~n9325 ;
  assign n9326 = n8921 & n68609 ;
  assign n9327 = n9091 | n9326 ;
  assign n9328 = n160 & n9327 ;
  assign n9329 = n8789 & n68538 ;
  assign n9330 = n9145 & n9329 ;
  assign n9331 = n9328 | n9330 ;
  assign n9332 = n66043 & n9331 ;
  assign n68610 = ~n9330 ;
  assign n9470 = x75 & n68610 ;
  assign n68611 = ~n9328 ;
  assign n9471 = n68611 & n9470 ;
  assign n9472 = n9332 | n9471 ;
  assign n68612 = ~n8916 ;
  assign n8920 = n68612 & n8919 ;
  assign n9333 = n8806 | n8919 ;
  assign n68613 = ~n9333 ;
  assign n9334 = n9085 & n68613 ;
  assign n9335 = n8920 | n9334 ;
  assign n9336 = n160 & n9335 ;
  assign n9337 = n8797 & n68538 ;
  assign n9338 = n9145 & n9337 ;
  assign n9339 = n9336 | n9338 ;
  assign n9340 = n65960 & n9339 ;
  assign n68614 = ~n9084 ;
  assign n9086 = n8914 & n68614 ;
  assign n9341 = n8814 | n8914 ;
  assign n68615 = ~n9341 ;
  assign n9342 = n8910 & n68615 ;
  assign n9343 = n9086 | n9342 ;
  assign n9344 = n160 & n9343 ;
  assign n9345 = n8805 & n68538 ;
  assign n9346 = n9145 & n9345 ;
  assign n9347 = n9344 | n9346 ;
  assign n9348 = n65909 & n9347 ;
  assign n68616 = ~n9346 ;
  assign n9458 = x73 & n68616 ;
  assign n68617 = ~n9344 ;
  assign n9459 = n68617 & n9458 ;
  assign n9460 = n9348 | n9459 ;
  assign n68618 = ~n8905 ;
  assign n8909 = n68618 & n8908 ;
  assign n9349 = n8823 | n8908 ;
  assign n68619 = ~n9349 ;
  assign n9350 = n9080 & n68619 ;
  assign n9351 = n8909 | n9350 ;
  assign n9352 = n160 & n9351 ;
  assign n9353 = n8813 & n68538 ;
  assign n9354 = n9145 & n9353 ;
  assign n9355 = n9352 | n9354 ;
  assign n9356 = n65877 & n9355 ;
  assign n68620 = ~n9079 ;
  assign n9081 = n8903 & n68620 ;
  assign n9357 = n8832 | n8903 ;
  assign n68621 = ~n9357 ;
  assign n9358 = n8899 & n68621 ;
  assign n9359 = n9081 | n9358 ;
  assign n9360 = n160 & n9359 ;
  assign n9361 = n8822 & n68538 ;
  assign n9362 = n9145 & n9361 ;
  assign n9363 = n9360 | n9362 ;
  assign n9364 = n65820 & n9363 ;
  assign n68622 = ~n9362 ;
  assign n9446 = x71 & n68622 ;
  assign n68623 = ~n9360 ;
  assign n9447 = n68623 & n9446 ;
  assign n9448 = n9364 | n9447 ;
  assign n68624 = ~n8895 ;
  assign n9077 = n68624 & n8898 ;
  assign n9365 = n8841 | n8898 ;
  assign n68625 = ~n9365 ;
  assign n9366 = n9075 & n68625 ;
  assign n9367 = n9077 | n9366 ;
  assign n9368 = n160 & n9367 ;
  assign n9369 = n8831 & n68538 ;
  assign n9370 = n9145 & n9369 ;
  assign n9371 = n9368 | n9370 ;
  assign n9372 = n65791 & n9371 ;
  assign n68626 = ~n9073 ;
  assign n9074 = n8893 & n68626 ;
  assign n9373 = n8886 | n9070 ;
  assign n9374 = n8850 | n8893 ;
  assign n68627 = ~n9374 ;
  assign n9375 = n9373 & n68627 ;
  assign n9376 = n9074 | n9375 ;
  assign n9377 = n160 & n9376 ;
  assign n9378 = n8840 & n68538 ;
  assign n9379 = n9145 & n9378 ;
  assign n9380 = n9377 | n9379 ;
  assign n9381 = n65772 & n9380 ;
  assign n68628 = ~n9379 ;
  assign n9435 = x69 & n68628 ;
  assign n68629 = ~n9377 ;
  assign n9436 = n68629 & n9435 ;
  assign n9437 = n9381 | n9436 ;
  assign n68630 = ~n8886 ;
  assign n9071 = n68630 & n9070 ;
  assign n9382 = n8856 | n9070 ;
  assign n68631 = ~n9382 ;
  assign n9383 = n8885 & n68631 ;
  assign n9384 = n9071 | n9383 ;
  assign n9385 = n160 & n9384 ;
  assign n9386 = n8849 & n68538 ;
  assign n9387 = n9145 & n9386 ;
  assign n9388 = n9385 | n9387 ;
  assign n9389 = n65746 & n9388 ;
  assign n68632 = ~n9066 ;
  assign n9067 = n8884 & n68632 ;
  assign n9390 = n8880 | n8884 ;
  assign n68633 = ~n9390 ;
  assign n9391 = n8879 & n68633 ;
  assign n9392 = n9067 | n9391 ;
  assign n9393 = n160 & n9392 ;
  assign n9394 = n8855 & n68538 ;
  assign n9395 = n9145 & n9394 ;
  assign n9396 = n9393 | n9395 ;
  assign n9397 = n65721 & n9396 ;
  assign n68634 = ~n9395 ;
  assign n9425 = x67 & n68634 ;
  assign n68635 = ~n9393 ;
  assign n9426 = n68635 & n9425 ;
  assign n9427 = n9397 | n9426 ;
  assign n9398 = n8876 & n8878 ;
  assign n9399 = n68442 & n9398 ;
  assign n68636 = ~n9399 ;
  assign n9400 = n9065 & n68636 ;
  assign n9401 = n160 & n9400 ;
  assign n9402 = n8873 & n68538 ;
  assign n9403 = n9145 & n9402 ;
  assign n9404 = n9401 | n9403 ;
  assign n9405 = n65686 & n9404 ;
  assign n68637 = ~x30 ;
  assign n9415 = n68637 & x64 ;
  assign n9061 = n8878 & n160 ;
  assign n9406 = n68538 & n9145 ;
  assign n68638 = ~n9406 ;
  assign n9407 = x64 & n68638 ;
  assign n68639 = ~n9407 ;
  assign n9408 = x31 & n68639 ;
  assign n9409 = n9061 | n9408 ;
  assign n9410 = x65 & n9409 ;
  assign n9060 = x64 & n160 ;
  assign n68640 = ~n9060 ;
  assign n9411 = x31 & n68640 ;
  assign n9412 = n8878 & n68638 ;
  assign n9413 = x65 | n9412 ;
  assign n9414 = n9411 | n9413 ;
  assign n68641 = ~n9410 ;
  assign n9416 = n68641 & n9414 ;
  assign n9417 = n9415 | n9416 ;
  assign n9418 = n9061 | n9411 ;
  assign n9419 = n65670 & n9418 ;
  assign n68642 = ~n9419 ;
  assign n9420 = n9417 & n68642 ;
  assign n68643 = ~n9403 ;
  assign n9421 = x66 & n68643 ;
  assign n68644 = ~n9401 ;
  assign n9422 = n68644 & n9421 ;
  assign n9423 = n9405 | n9422 ;
  assign n9424 = n9420 | n9423 ;
  assign n68645 = ~n9405 ;
  assign n9428 = n68645 & n9424 ;
  assign n9429 = n9427 | n9428 ;
  assign n68646 = ~n9397 ;
  assign n9430 = n68646 & n9429 ;
  assign n68647 = ~n9387 ;
  assign n9431 = x68 & n68647 ;
  assign n68648 = ~n9385 ;
  assign n9432 = n68648 & n9431 ;
  assign n9433 = n9389 | n9432 ;
  assign n9434 = n9430 | n9433 ;
  assign n68649 = ~n9389 ;
  assign n9438 = n68649 & n9434 ;
  assign n9439 = n9437 | n9438 ;
  assign n68650 = ~n9381 ;
  assign n9440 = n68650 & n9439 ;
  assign n68651 = ~n9370 ;
  assign n9441 = x70 & n68651 ;
  assign n68652 = ~n9368 ;
  assign n9442 = n68652 & n9441 ;
  assign n9443 = n9372 | n9442 ;
  assign n9445 = n9440 | n9443 ;
  assign n68653 = ~n9372 ;
  assign n9450 = n68653 & n9445 ;
  assign n9451 = n9448 | n9450 ;
  assign n68654 = ~n9364 ;
  assign n9452 = n68654 & n9451 ;
  assign n68655 = ~n9354 ;
  assign n9453 = x72 & n68655 ;
  assign n68656 = ~n9352 ;
  assign n9454 = n68656 & n9453 ;
  assign n9455 = n9356 | n9454 ;
  assign n9457 = n9452 | n9455 ;
  assign n68657 = ~n9356 ;
  assign n9462 = n68657 & n9457 ;
  assign n9463 = n9460 | n9462 ;
  assign n68658 = ~n9348 ;
  assign n9464 = n68658 & n9463 ;
  assign n68659 = ~n9338 ;
  assign n9465 = x74 & n68659 ;
  assign n68660 = ~n9336 ;
  assign n9466 = n68660 & n9465 ;
  assign n9467 = n9340 | n9466 ;
  assign n9469 = n9464 | n9467 ;
  assign n68661 = ~n9340 ;
  assign n9474 = n68661 & n9469 ;
  assign n9475 = n9472 | n9474 ;
  assign n68662 = ~n9332 ;
  assign n9476 = n68662 & n9475 ;
  assign n68663 = ~n9322 ;
  assign n9477 = x76 & n68663 ;
  assign n68664 = ~n9320 ;
  assign n9478 = n68664 & n9477 ;
  assign n9479 = n9324 | n9478 ;
  assign n9481 = n9476 | n9479 ;
  assign n68665 = ~n9324 ;
  assign n9486 = n68665 & n9481 ;
  assign n9487 = n9484 | n9486 ;
  assign n68666 = ~n9316 ;
  assign n9488 = n68666 & n9487 ;
  assign n68667 = ~n9306 ;
  assign n9489 = x78 & n68667 ;
  assign n68668 = ~n9304 ;
  assign n9490 = n68668 & n9489 ;
  assign n9491 = n9308 | n9490 ;
  assign n9493 = n9488 | n9491 ;
  assign n68669 = ~n9308 ;
  assign n9498 = n68669 & n9493 ;
  assign n9499 = n9496 | n9498 ;
  assign n68670 = ~n9300 ;
  assign n9500 = n68670 & n9499 ;
  assign n68671 = ~n9290 ;
  assign n9501 = x80 & n68671 ;
  assign n68672 = ~n9288 ;
  assign n9502 = n68672 & n9501 ;
  assign n9503 = n9292 | n9502 ;
  assign n9505 = n9500 | n9503 ;
  assign n68673 = ~n9292 ;
  assign n9510 = n68673 & n9505 ;
  assign n9511 = n9508 | n9510 ;
  assign n68674 = ~n9284 ;
  assign n9512 = n68674 & n9511 ;
  assign n68675 = ~n9274 ;
  assign n9513 = x82 & n68675 ;
  assign n68676 = ~n9272 ;
  assign n9514 = n68676 & n9513 ;
  assign n9515 = n9276 | n9514 ;
  assign n9517 = n9512 | n9515 ;
  assign n68677 = ~n9276 ;
  assign n9522 = n68677 & n9517 ;
  assign n9523 = n9520 | n9522 ;
  assign n68678 = ~n9268 ;
  assign n9524 = n68678 & n9523 ;
  assign n68679 = ~n9258 ;
  assign n9525 = x84 & n68679 ;
  assign n68680 = ~n9256 ;
  assign n9526 = n68680 & n9525 ;
  assign n9527 = n9260 | n9526 ;
  assign n9529 = n9524 | n9527 ;
  assign n68681 = ~n9260 ;
  assign n9534 = n68681 & n9529 ;
  assign n9535 = n9532 | n9534 ;
  assign n68682 = ~n9252 ;
  assign n9536 = n68682 & n9535 ;
  assign n68683 = ~n9242 ;
  assign n9537 = x86 & n68683 ;
  assign n68684 = ~n9240 ;
  assign n9538 = n68684 & n9537 ;
  assign n9539 = n9244 | n9538 ;
  assign n9541 = n9536 | n9539 ;
  assign n68685 = ~n9244 ;
  assign n9546 = n68685 & n9541 ;
  assign n9547 = n9544 | n9546 ;
  assign n68686 = ~n9236 ;
  assign n9548 = n68686 & n9547 ;
  assign n68687 = ~n9226 ;
  assign n9549 = x88 & n68687 ;
  assign n68688 = ~n9224 ;
  assign n9550 = n68688 & n9549 ;
  assign n9551 = n9228 | n9550 ;
  assign n9553 = n9548 | n9551 ;
  assign n68689 = ~n9228 ;
  assign n9558 = n68689 & n9553 ;
  assign n9559 = n9556 | n9558 ;
  assign n68690 = ~n9220 ;
  assign n9560 = n68690 & n9559 ;
  assign n68691 = ~n9210 ;
  assign n9561 = x90 & n68691 ;
  assign n68692 = ~n9208 ;
  assign n9562 = n68692 & n9561 ;
  assign n9563 = n9212 | n9562 ;
  assign n9565 = n9560 | n9563 ;
  assign n68693 = ~n9212 ;
  assign n9570 = n68693 & n9565 ;
  assign n9571 = n9568 | n9570 ;
  assign n68694 = ~n9204 ;
  assign n9572 = n68694 & n9571 ;
  assign n68695 = ~n9194 ;
  assign n9573 = x92 & n68695 ;
  assign n68696 = ~n9192 ;
  assign n9574 = n68696 & n9573 ;
  assign n9575 = n9196 | n9574 ;
  assign n9577 = n9572 | n9575 ;
  assign n68697 = ~n9196 ;
  assign n9582 = n68697 & n9577 ;
  assign n9583 = n9580 | n9582 ;
  assign n68698 = ~n9188 ;
  assign n9584 = n68698 & n9583 ;
  assign n68699 = ~n9178 ;
  assign n9585 = x94 & n68699 ;
  assign n68700 = ~n9176 ;
  assign n9586 = n68700 & n9585 ;
  assign n9587 = n9180 | n9586 ;
  assign n9589 = n9584 | n9587 ;
  assign n68701 = ~n9180 ;
  assign n9594 = n68701 & n9589 ;
  assign n9595 = n9592 | n9594 ;
  assign n68702 = ~n9172 ;
  assign n9596 = n68702 & n9595 ;
  assign n68703 = ~n9162 ;
  assign n9597 = x96 & n68703 ;
  assign n68704 = ~n9160 ;
  assign n9598 = n68704 & n9597 ;
  assign n9599 = n9164 | n9598 ;
  assign n9601 = n9596 | n9599 ;
  assign n68705 = ~n9164 ;
  assign n9605 = n68705 & n9601 ;
  assign n9606 = n9604 | n9605 ;
  assign n68706 = ~n9156 ;
  assign n9607 = n68706 & n9606 ;
  assign n9608 = n65474 | n65609 ;
  assign n9609 = n67093 | n9608 ;
  assign n9610 = n66858 | n9609 ;
  assign n9611 = n9607 | n9610 ;
  assign n9690 = n9163 & n9611 ;
  assign n9600 = n9172 | n9599 ;
  assign n9615 = x65 & n9418 ;
  assign n68707 = ~n9615 ;
  assign n9616 = n9414 & n68707 ;
  assign n9618 = n9415 | n9616 ;
  assign n9620 = n68642 & n9618 ;
  assign n9621 = n9423 | n9620 ;
  assign n9622 = n68645 & n9621 ;
  assign n9623 = n9427 | n9622 ;
  assign n9624 = n68646 & n9623 ;
  assign n9625 = n9433 | n9624 ;
  assign n9626 = n68649 & n9625 ;
  assign n9627 = n9437 | n9626 ;
  assign n9628 = n68650 & n9627 ;
  assign n9629 = n9443 | n9628 ;
  assign n9630 = n68653 & n9629 ;
  assign n9631 = n9448 | n9630 ;
  assign n9632 = n68654 & n9631 ;
  assign n9633 = n9455 | n9632 ;
  assign n9634 = n68657 & n9633 ;
  assign n9635 = n9460 | n9634 ;
  assign n9636 = n68658 & n9635 ;
  assign n9637 = n9467 | n9636 ;
  assign n9638 = n68661 & n9637 ;
  assign n9639 = n9472 | n9638 ;
  assign n9640 = n68662 & n9639 ;
  assign n9641 = n9479 | n9640 ;
  assign n9642 = n68665 & n9641 ;
  assign n9643 = n9484 | n9642 ;
  assign n9644 = n68666 & n9643 ;
  assign n9645 = n9491 | n9644 ;
  assign n9646 = n68669 & n9645 ;
  assign n9647 = n9496 | n9646 ;
  assign n9648 = n68670 & n9647 ;
  assign n9649 = n9503 | n9648 ;
  assign n9650 = n68673 & n9649 ;
  assign n9651 = n9508 | n9650 ;
  assign n9652 = n68674 & n9651 ;
  assign n9653 = n9515 | n9652 ;
  assign n9654 = n68677 & n9653 ;
  assign n9655 = n9520 | n9654 ;
  assign n9656 = n68678 & n9655 ;
  assign n9657 = n9527 | n9656 ;
  assign n9658 = n68681 & n9657 ;
  assign n9659 = n9532 | n9658 ;
  assign n9660 = n68682 & n9659 ;
  assign n9661 = n9539 | n9660 ;
  assign n9662 = n68685 & n9661 ;
  assign n9663 = n9544 | n9662 ;
  assign n9664 = n68686 & n9663 ;
  assign n9665 = n9551 | n9664 ;
  assign n9666 = n68689 & n9665 ;
  assign n9667 = n9556 | n9666 ;
  assign n9668 = n68690 & n9667 ;
  assign n9669 = n9563 | n9668 ;
  assign n9670 = n68693 & n9669 ;
  assign n9671 = n9568 | n9670 ;
  assign n9672 = n68694 & n9671 ;
  assign n9673 = n9575 | n9672 ;
  assign n9674 = n68697 & n9673 ;
  assign n9675 = n9580 | n9674 ;
  assign n9676 = n68698 & n9675 ;
  assign n9677 = n9587 | n9676 ;
  assign n9678 = n68701 & n9677 ;
  assign n9679 = n9592 | n9678 ;
  assign n68708 = ~n9600 ;
  assign n9691 = n68708 & n9679 ;
  assign n9680 = n68702 & n9679 ;
  assign n68709 = ~n9680 ;
  assign n9692 = n9599 & n68709 ;
  assign n9693 = n9691 | n9692 ;
  assign n68710 = ~n9610 ;
  assign n9694 = n68710 & n9693 ;
  assign n68711 = ~n9607 ;
  assign n9695 = n68711 & n9694 ;
  assign n9696 = n9690 | n9695 ;
  assign n68712 = ~n9155 ;
  assign n9613 = n68712 & n9611 ;
  assign n68713 = ~n9605 ;
  assign n9683 = n9604 & n68713 ;
  assign n9681 = n9599 | n9680 ;
  assign n9684 = n9164 | n9604 ;
  assign n68714 = ~n9684 ;
  assign n9685 = n9681 & n68714 ;
  assign n9686 = n9683 | n9685 ;
  assign n9687 = n9611 | n9686 ;
  assign n68715 = ~n9613 ;
  assign n9688 = n68715 & n9687 ;
  assign n68716 = ~x98 ;
  assign n9689 = n68716 & n9688 ;
  assign n9697 = n68545 & n9696 ;
  assign n9698 = n9171 & n9611 ;
  assign n9593 = n9180 | n9592 ;
  assign n68717 = ~n9593 ;
  assign n9699 = n9589 & n68717 ;
  assign n68718 = ~n9594 ;
  assign n9700 = n9592 & n68718 ;
  assign n9701 = n9699 | n9700 ;
  assign n9702 = n68710 & n9701 ;
  assign n9703 = n68711 & n9702 ;
  assign n9704 = n9698 | n9703 ;
  assign n9705 = n68438 & n9704 ;
  assign n9706 = n9179 & n9611 ;
  assign n9588 = n9188 | n9587 ;
  assign n68719 = ~n9588 ;
  assign n9707 = n68719 & n9675 ;
  assign n68720 = ~n9676 ;
  assign n9708 = n9587 & n68720 ;
  assign n9709 = n9707 | n9708 ;
  assign n9710 = n68710 & n9709 ;
  assign n9711 = n68711 & n9710 ;
  assign n9712 = n9706 | n9711 ;
  assign n9713 = n68214 & n9712 ;
  assign n9714 = n9187 & n9611 ;
  assign n9581 = n9196 | n9580 ;
  assign n68721 = ~n9581 ;
  assign n9715 = n9577 & n68721 ;
  assign n68722 = ~n9582 ;
  assign n9716 = n9580 & n68722 ;
  assign n9717 = n9715 | n9716 ;
  assign n9718 = n68710 & n9717 ;
  assign n9719 = n68711 & n9718 ;
  assign n9720 = n9714 | n9719 ;
  assign n9721 = n68058 & n9720 ;
  assign n9722 = n9195 & n9611 ;
  assign n9576 = n9204 | n9575 ;
  assign n68723 = ~n9576 ;
  assign n9723 = n68723 & n9671 ;
  assign n68724 = ~n9672 ;
  assign n9724 = n9575 & n68724 ;
  assign n9725 = n9723 | n9724 ;
  assign n9726 = n68710 & n9725 ;
  assign n9727 = n68711 & n9726 ;
  assign n9728 = n9722 | n9727 ;
  assign n9729 = n67986 & n9728 ;
  assign n9730 = n9203 & n9611 ;
  assign n9569 = n9212 | n9568 ;
  assign n68725 = ~n9569 ;
  assign n9731 = n9565 & n68725 ;
  assign n68726 = ~n9570 ;
  assign n9732 = n9568 & n68726 ;
  assign n9733 = n9731 | n9732 ;
  assign n9734 = n68710 & n9733 ;
  assign n9735 = n68711 & n9734 ;
  assign n9736 = n9730 | n9735 ;
  assign n9737 = n67763 & n9736 ;
  assign n9738 = n9211 & n9611 ;
  assign n9564 = n9220 | n9563 ;
  assign n68727 = ~n9564 ;
  assign n9739 = n68727 & n9667 ;
  assign n68728 = ~n9668 ;
  assign n9740 = n9563 & n68728 ;
  assign n9741 = n9739 | n9740 ;
  assign n9742 = n68710 & n9741 ;
  assign n9743 = n68711 & n9742 ;
  assign n9744 = n9738 | n9743 ;
  assign n9745 = n67622 & n9744 ;
  assign n9746 = n9219 & n9611 ;
  assign n9557 = n9228 | n9556 ;
  assign n68729 = ~n9557 ;
  assign n9747 = n9553 & n68729 ;
  assign n68730 = ~n9558 ;
  assign n9748 = n9556 & n68730 ;
  assign n9749 = n9747 | n9748 ;
  assign n9750 = n68710 & n9749 ;
  assign n9751 = n68711 & n9750 ;
  assign n9752 = n9746 | n9751 ;
  assign n9753 = n67531 & n9752 ;
  assign n9754 = n9227 & n9611 ;
  assign n9552 = n9236 | n9551 ;
  assign n68731 = ~n9552 ;
  assign n9755 = n68731 & n9663 ;
  assign n68732 = ~n9664 ;
  assign n9756 = n9551 & n68732 ;
  assign n9757 = n9755 | n9756 ;
  assign n9758 = n68710 & n9757 ;
  assign n9759 = n68711 & n9758 ;
  assign n9760 = n9754 | n9759 ;
  assign n9761 = n67348 & n9760 ;
  assign n9762 = n9235 & n9611 ;
  assign n9545 = n9244 | n9544 ;
  assign n68733 = ~n9545 ;
  assign n9763 = n9541 & n68733 ;
  assign n68734 = ~n9546 ;
  assign n9764 = n9544 & n68734 ;
  assign n9765 = n9763 | n9764 ;
  assign n9766 = n68710 & n9765 ;
  assign n9767 = n68711 & n9766 ;
  assign n9768 = n9762 | n9767 ;
  assign n9769 = n67222 & n9768 ;
  assign n9770 = n9243 & n9611 ;
  assign n9540 = n9252 | n9539 ;
  assign n68735 = ~n9540 ;
  assign n9771 = n68735 & n9659 ;
  assign n68736 = ~n9660 ;
  assign n9772 = n9539 & n68736 ;
  assign n9773 = n9771 | n9772 ;
  assign n9774 = n68710 & n9773 ;
  assign n9775 = n68711 & n9774 ;
  assign n9776 = n9770 | n9775 ;
  assign n9777 = n67164 & n9776 ;
  assign n9778 = n9251 & n9611 ;
  assign n9533 = n9260 | n9532 ;
  assign n68737 = ~n9533 ;
  assign n9779 = n9529 & n68737 ;
  assign n68738 = ~n9534 ;
  assign n9780 = n9532 & n68738 ;
  assign n9781 = n9779 | n9780 ;
  assign n9782 = n68710 & n9781 ;
  assign n9783 = n68711 & n9782 ;
  assign n9784 = n9778 | n9783 ;
  assign n9785 = n66979 & n9784 ;
  assign n9786 = n9259 & n9611 ;
  assign n9528 = n9268 | n9527 ;
  assign n68739 = ~n9528 ;
  assign n9787 = n68739 & n9655 ;
  assign n68740 = ~n9656 ;
  assign n9788 = n9527 & n68740 ;
  assign n9789 = n9787 | n9788 ;
  assign n9790 = n68710 & n9789 ;
  assign n9791 = n68711 & n9790 ;
  assign n9792 = n9786 | n9791 ;
  assign n9793 = n66868 & n9792 ;
  assign n9794 = n9267 & n9611 ;
  assign n9521 = n9276 | n9520 ;
  assign n68741 = ~n9521 ;
  assign n9795 = n9517 & n68741 ;
  assign n68742 = ~n9522 ;
  assign n9796 = n9520 & n68742 ;
  assign n9797 = n9795 | n9796 ;
  assign n9798 = n68710 & n9797 ;
  assign n9799 = n68711 & n9798 ;
  assign n9800 = n9794 | n9799 ;
  assign n9801 = n66797 & n9800 ;
  assign n9802 = n9275 & n9611 ;
  assign n9516 = n9284 | n9515 ;
  assign n68743 = ~n9516 ;
  assign n9803 = n68743 & n9651 ;
  assign n68744 = ~n9652 ;
  assign n9804 = n9515 & n68744 ;
  assign n9805 = n9803 | n9804 ;
  assign n9806 = n68710 & n9805 ;
  assign n9807 = n68711 & n9806 ;
  assign n9808 = n9802 | n9807 ;
  assign n9809 = n66654 & n9808 ;
  assign n9810 = n9283 & n9611 ;
  assign n9509 = n9292 | n9508 ;
  assign n68745 = ~n9509 ;
  assign n9811 = n9505 & n68745 ;
  assign n68746 = ~n9510 ;
  assign n9812 = n9508 & n68746 ;
  assign n9813 = n9811 | n9812 ;
  assign n9814 = n68710 & n9813 ;
  assign n9815 = n68711 & n9814 ;
  assign n9816 = n9810 | n9815 ;
  assign n9817 = n66560 & n9816 ;
  assign n9818 = n9291 & n9611 ;
  assign n9504 = n9300 | n9503 ;
  assign n68747 = ~n9504 ;
  assign n9819 = n68747 & n9647 ;
  assign n68748 = ~n9648 ;
  assign n9820 = n9503 & n68748 ;
  assign n9821 = n9819 | n9820 ;
  assign n9822 = n68710 & n9821 ;
  assign n9823 = n68711 & n9822 ;
  assign n9824 = n9818 | n9823 ;
  assign n9825 = n66505 & n9824 ;
  assign n9826 = n9299 & n9611 ;
  assign n9497 = n9308 | n9496 ;
  assign n68749 = ~n9497 ;
  assign n9827 = n9493 & n68749 ;
  assign n68750 = ~n9498 ;
  assign n9828 = n9496 & n68750 ;
  assign n9829 = n9827 | n9828 ;
  assign n9830 = n68710 & n9829 ;
  assign n9831 = n68711 & n9830 ;
  assign n9832 = n9826 | n9831 ;
  assign n9833 = n66379 & n9832 ;
  assign n9834 = n9307 & n9611 ;
  assign n9492 = n9316 | n9491 ;
  assign n68751 = ~n9492 ;
  assign n9835 = n68751 & n9643 ;
  assign n68752 = ~n9644 ;
  assign n9836 = n9491 & n68752 ;
  assign n9837 = n9835 | n9836 ;
  assign n9838 = n68710 & n9837 ;
  assign n9839 = n68711 & n9838 ;
  assign n9840 = n9834 | n9839 ;
  assign n9841 = n66299 & n9840 ;
  assign n9842 = n9315 & n9611 ;
  assign n9485 = n9324 | n9484 ;
  assign n68753 = ~n9485 ;
  assign n9843 = n9481 & n68753 ;
  assign n68754 = ~n9486 ;
  assign n9844 = n9484 & n68754 ;
  assign n9845 = n9843 | n9844 ;
  assign n9846 = n68710 & n9845 ;
  assign n9847 = n68711 & n9846 ;
  assign n9848 = n9842 | n9847 ;
  assign n9849 = n66244 & n9848 ;
  assign n9850 = n9323 & n9611 ;
  assign n9480 = n9332 | n9479 ;
  assign n68755 = ~n9480 ;
  assign n9851 = n68755 & n9639 ;
  assign n68756 = ~n9640 ;
  assign n9852 = n9479 & n68756 ;
  assign n9853 = n9851 | n9852 ;
  assign n9854 = n68710 & n9853 ;
  assign n9855 = n68711 & n9854 ;
  assign n9856 = n9850 | n9855 ;
  assign n9857 = n66145 & n9856 ;
  assign n9858 = n9331 & n9611 ;
  assign n9473 = n9340 | n9472 ;
  assign n68757 = ~n9473 ;
  assign n9859 = n9469 & n68757 ;
  assign n68758 = ~n9474 ;
  assign n9860 = n9472 & n68758 ;
  assign n9861 = n9859 | n9860 ;
  assign n9862 = n68710 & n9861 ;
  assign n9863 = n68711 & n9862 ;
  assign n9864 = n9858 | n9863 ;
  assign n9865 = n66081 & n9864 ;
  assign n9866 = n9339 & n9611 ;
  assign n9468 = n9348 | n9467 ;
  assign n68759 = ~n9468 ;
  assign n9867 = n68759 & n9635 ;
  assign n68760 = ~n9636 ;
  assign n9868 = n9467 & n68760 ;
  assign n9869 = n9867 | n9868 ;
  assign n9870 = n68710 & n9869 ;
  assign n9871 = n68711 & n9870 ;
  assign n9872 = n9866 | n9871 ;
  assign n9873 = n66043 & n9872 ;
  assign n9874 = n9347 & n9611 ;
  assign n9461 = n9356 | n9460 ;
  assign n68761 = ~n9461 ;
  assign n9875 = n9457 & n68761 ;
  assign n68762 = ~n9462 ;
  assign n9876 = n9460 & n68762 ;
  assign n9877 = n9875 | n9876 ;
  assign n9878 = n68710 & n9877 ;
  assign n9879 = n68711 & n9878 ;
  assign n9880 = n9874 | n9879 ;
  assign n9881 = n65960 & n9880 ;
  assign n9882 = n9355 & n9611 ;
  assign n9456 = n9364 | n9455 ;
  assign n68763 = ~n9456 ;
  assign n9883 = n68763 & n9631 ;
  assign n68764 = ~n9632 ;
  assign n9884 = n9455 & n68764 ;
  assign n9885 = n9883 | n9884 ;
  assign n9886 = n68710 & n9885 ;
  assign n9887 = n68711 & n9886 ;
  assign n9888 = n9882 | n9887 ;
  assign n9889 = n65909 & n9888 ;
  assign n9890 = n9363 & n9611 ;
  assign n9449 = n9372 | n9448 ;
  assign n68765 = ~n9449 ;
  assign n9891 = n9445 & n68765 ;
  assign n68766 = ~n9450 ;
  assign n9892 = n9448 & n68766 ;
  assign n9893 = n9891 | n9892 ;
  assign n9894 = n68710 & n9893 ;
  assign n9895 = n68711 & n9894 ;
  assign n9896 = n9890 | n9895 ;
  assign n9897 = n65877 & n9896 ;
  assign n9898 = n9371 & n9611 ;
  assign n9444 = n9381 | n9443 ;
  assign n68767 = ~n9444 ;
  assign n9899 = n68767 & n9627 ;
  assign n68768 = ~n9628 ;
  assign n9900 = n9443 & n68768 ;
  assign n9901 = n9899 | n9900 ;
  assign n9902 = n68710 & n9901 ;
  assign n9903 = n68711 & n9902 ;
  assign n9904 = n9898 | n9903 ;
  assign n9905 = n65820 & n9904 ;
  assign n9906 = n9380 & n9611 ;
  assign n9614 = n9389 | n9437 ;
  assign n68769 = ~n9614 ;
  assign n9907 = n9434 & n68769 ;
  assign n68770 = ~n9438 ;
  assign n9908 = n9437 & n68770 ;
  assign n9909 = n9907 | n9908 ;
  assign n9910 = n68710 & n9909 ;
  assign n9911 = n68711 & n9910 ;
  assign n9912 = n9906 | n9911 ;
  assign n9913 = n65791 & n9912 ;
  assign n9914 = n9388 & n9611 ;
  assign n9915 = n9397 | n9433 ;
  assign n68771 = ~n9915 ;
  assign n9916 = n9623 & n68771 ;
  assign n68772 = ~n9624 ;
  assign n9917 = n9433 & n68772 ;
  assign n9918 = n9916 | n9917 ;
  assign n9919 = n68710 & n9918 ;
  assign n9920 = n68711 & n9919 ;
  assign n9921 = n9914 | n9920 ;
  assign n9922 = n65772 & n9921 ;
  assign n9923 = n9396 & n9611 ;
  assign n9924 = n9405 | n9427 ;
  assign n68773 = ~n9924 ;
  assign n9925 = n9621 & n68773 ;
  assign n68774 = ~n9428 ;
  assign n9926 = n9427 & n68774 ;
  assign n9927 = n9925 | n9926 ;
  assign n9928 = n68710 & n9927 ;
  assign n9929 = n68711 & n9928 ;
  assign n9930 = n9923 | n9929 ;
  assign n9931 = n65746 & n9930 ;
  assign n9932 = n9404 & n9611 ;
  assign n9619 = n9419 | n9423 ;
  assign n68775 = ~n9619 ;
  assign n9933 = n9417 & n68775 ;
  assign n68776 = ~n9620 ;
  assign n9934 = n9423 & n68776 ;
  assign n9935 = n9933 | n9934 ;
  assign n9936 = n68710 & n9935 ;
  assign n9937 = n68711 & n9936 ;
  assign n9938 = n9932 | n9937 ;
  assign n9939 = n65721 & n9938 ;
  assign n9612 = n9418 & n9611 ;
  assign n9617 = n9414 & n9415 ;
  assign n9940 = n68641 & n9617 ;
  assign n9941 = n9610 | n9940 ;
  assign n68777 = ~n9941 ;
  assign n9942 = n9417 & n68777 ;
  assign n9943 = n68711 & n9942 ;
  assign n9944 = n9612 | n9943 ;
  assign n9945 = n65686 & n9944 ;
  assign n68778 = ~n65609 ;
  assign n9953 = n68778 & n9415 ;
  assign n68779 = ~n65474 ;
  assign n9954 = n68779 & n9953 ;
  assign n68780 = ~n67093 ;
  assign n9955 = n68780 & n9954 ;
  assign n9956 = n66510 & n9955 ;
  assign n9957 = n68711 & n9956 ;
  assign n9946 = x64 & n68716 ;
  assign n68781 = ~n284 ;
  assign n9947 = n68781 & n9946 ;
  assign n68782 = ~n282 ;
  assign n9948 = n68782 & n9947 ;
  assign n68783 = ~n293 ;
  assign n9949 = n68783 & n9948 ;
  assign n9950 = n66715 & n9949 ;
  assign n9682 = n68705 & n9681 ;
  assign n9965 = n9604 | n9682 ;
  assign n9966 = n68706 & n9965 ;
  assign n68784 = ~n9966 ;
  assign n9967 = n9950 & n68784 ;
  assign n68785 = ~n9967 ;
  assign n9968 = x30 & n68785 ;
  assign n9969 = n9957 | n9968 ;
  assign n9970 = n65670 & n9969 ;
  assign n9951 = n68711 & n9950 ;
  assign n68786 = ~n9951 ;
  assign n9952 = x30 & n68786 ;
  assign n9958 = n9952 | n9957 ;
  assign n9959 = x65 & n9958 ;
  assign n9961 = x65 | n9957 ;
  assign n9962 = n9952 | n9961 ;
  assign n68787 = ~n9959 ;
  assign n9963 = n68787 & n9962 ;
  assign n68788 = ~x29 ;
  assign n9964 = n68788 & x64 ;
  assign n9971 = n9963 | n9964 ;
  assign n68789 = ~n9970 ;
  assign n9972 = n68789 & n9971 ;
  assign n68790 = ~n9943 ;
  assign n9973 = x66 & n68790 ;
  assign n68791 = ~n9612 ;
  assign n9974 = n68791 & n9973 ;
  assign n9975 = n9945 | n9974 ;
  assign n9976 = n9972 | n9975 ;
  assign n68792 = ~n9945 ;
  assign n9977 = n68792 & n9976 ;
  assign n68793 = ~n9937 ;
  assign n9978 = x67 & n68793 ;
  assign n68794 = ~n9932 ;
  assign n9979 = n68794 & n9978 ;
  assign n9980 = n9939 | n9979 ;
  assign n9981 = n9977 | n9980 ;
  assign n68795 = ~n9939 ;
  assign n9982 = n68795 & n9981 ;
  assign n68796 = ~n9929 ;
  assign n9983 = x68 & n68796 ;
  assign n68797 = ~n9923 ;
  assign n9984 = n68797 & n9983 ;
  assign n9985 = n9931 | n9984 ;
  assign n9986 = n9982 | n9985 ;
  assign n68798 = ~n9931 ;
  assign n9987 = n68798 & n9986 ;
  assign n68799 = ~n9920 ;
  assign n9988 = x69 & n68799 ;
  assign n68800 = ~n9914 ;
  assign n9989 = n68800 & n9988 ;
  assign n9990 = n9922 | n9989 ;
  assign n9991 = n9987 | n9990 ;
  assign n68801 = ~n9922 ;
  assign n9992 = n68801 & n9991 ;
  assign n68802 = ~n9911 ;
  assign n9993 = x70 & n68802 ;
  assign n68803 = ~n9906 ;
  assign n9994 = n68803 & n9993 ;
  assign n9995 = n9913 | n9994 ;
  assign n9997 = n9992 | n9995 ;
  assign n68804 = ~n9913 ;
  assign n9998 = n68804 & n9997 ;
  assign n68805 = ~n9903 ;
  assign n9999 = x71 & n68805 ;
  assign n68806 = ~n9898 ;
  assign n10000 = n68806 & n9999 ;
  assign n10001 = n9905 | n10000 ;
  assign n10002 = n9998 | n10001 ;
  assign n68807 = ~n9905 ;
  assign n10003 = n68807 & n10002 ;
  assign n68808 = ~n9895 ;
  assign n10004 = x72 & n68808 ;
  assign n68809 = ~n9890 ;
  assign n10005 = n68809 & n10004 ;
  assign n10006 = n9897 | n10005 ;
  assign n10008 = n10003 | n10006 ;
  assign n68810 = ~n9897 ;
  assign n10009 = n68810 & n10008 ;
  assign n68811 = ~n9887 ;
  assign n10010 = x73 & n68811 ;
  assign n68812 = ~n9882 ;
  assign n10011 = n68812 & n10010 ;
  assign n10012 = n9889 | n10011 ;
  assign n10013 = n10009 | n10012 ;
  assign n68813 = ~n9889 ;
  assign n10014 = n68813 & n10013 ;
  assign n68814 = ~n9879 ;
  assign n10015 = x74 & n68814 ;
  assign n68815 = ~n9874 ;
  assign n10016 = n68815 & n10015 ;
  assign n10017 = n9881 | n10016 ;
  assign n10019 = n10014 | n10017 ;
  assign n68816 = ~n9881 ;
  assign n10020 = n68816 & n10019 ;
  assign n68817 = ~n9871 ;
  assign n10021 = x75 & n68817 ;
  assign n68818 = ~n9866 ;
  assign n10022 = n68818 & n10021 ;
  assign n10023 = n9873 | n10022 ;
  assign n10024 = n10020 | n10023 ;
  assign n68819 = ~n9873 ;
  assign n10025 = n68819 & n10024 ;
  assign n68820 = ~n9863 ;
  assign n10026 = x76 & n68820 ;
  assign n68821 = ~n9858 ;
  assign n10027 = n68821 & n10026 ;
  assign n10028 = n9865 | n10027 ;
  assign n10030 = n10025 | n10028 ;
  assign n68822 = ~n9865 ;
  assign n10031 = n68822 & n10030 ;
  assign n68823 = ~n9855 ;
  assign n10032 = x77 & n68823 ;
  assign n68824 = ~n9850 ;
  assign n10033 = n68824 & n10032 ;
  assign n10034 = n9857 | n10033 ;
  assign n10035 = n10031 | n10034 ;
  assign n68825 = ~n9857 ;
  assign n10036 = n68825 & n10035 ;
  assign n68826 = ~n9847 ;
  assign n10037 = x78 & n68826 ;
  assign n68827 = ~n9842 ;
  assign n10038 = n68827 & n10037 ;
  assign n10039 = n9849 | n10038 ;
  assign n10041 = n10036 | n10039 ;
  assign n68828 = ~n9849 ;
  assign n10042 = n68828 & n10041 ;
  assign n68829 = ~n9839 ;
  assign n10043 = x79 & n68829 ;
  assign n68830 = ~n9834 ;
  assign n10044 = n68830 & n10043 ;
  assign n10045 = n9841 | n10044 ;
  assign n10046 = n10042 | n10045 ;
  assign n68831 = ~n9841 ;
  assign n10047 = n68831 & n10046 ;
  assign n68832 = ~n9831 ;
  assign n10048 = x80 & n68832 ;
  assign n68833 = ~n9826 ;
  assign n10049 = n68833 & n10048 ;
  assign n10050 = n9833 | n10049 ;
  assign n10052 = n10047 | n10050 ;
  assign n68834 = ~n9833 ;
  assign n10053 = n68834 & n10052 ;
  assign n68835 = ~n9823 ;
  assign n10054 = x81 & n68835 ;
  assign n68836 = ~n9818 ;
  assign n10055 = n68836 & n10054 ;
  assign n10056 = n9825 | n10055 ;
  assign n10057 = n10053 | n10056 ;
  assign n68837 = ~n9825 ;
  assign n10058 = n68837 & n10057 ;
  assign n68838 = ~n9815 ;
  assign n10059 = x82 & n68838 ;
  assign n68839 = ~n9810 ;
  assign n10060 = n68839 & n10059 ;
  assign n10061 = n9817 | n10060 ;
  assign n10063 = n10058 | n10061 ;
  assign n68840 = ~n9817 ;
  assign n10064 = n68840 & n10063 ;
  assign n68841 = ~n9807 ;
  assign n10065 = x83 & n68841 ;
  assign n68842 = ~n9802 ;
  assign n10066 = n68842 & n10065 ;
  assign n10067 = n9809 | n10066 ;
  assign n10068 = n10064 | n10067 ;
  assign n68843 = ~n9809 ;
  assign n10069 = n68843 & n10068 ;
  assign n68844 = ~n9799 ;
  assign n10070 = x84 & n68844 ;
  assign n68845 = ~n9794 ;
  assign n10071 = n68845 & n10070 ;
  assign n10072 = n9801 | n10071 ;
  assign n10074 = n10069 | n10072 ;
  assign n68846 = ~n9801 ;
  assign n10075 = n68846 & n10074 ;
  assign n68847 = ~n9791 ;
  assign n10076 = x85 & n68847 ;
  assign n68848 = ~n9786 ;
  assign n10077 = n68848 & n10076 ;
  assign n10078 = n9793 | n10077 ;
  assign n10079 = n10075 | n10078 ;
  assign n68849 = ~n9793 ;
  assign n10080 = n68849 & n10079 ;
  assign n68850 = ~n9783 ;
  assign n10081 = x86 & n68850 ;
  assign n68851 = ~n9778 ;
  assign n10082 = n68851 & n10081 ;
  assign n10083 = n9785 | n10082 ;
  assign n10085 = n10080 | n10083 ;
  assign n68852 = ~n9785 ;
  assign n10086 = n68852 & n10085 ;
  assign n68853 = ~n9775 ;
  assign n10087 = x87 & n68853 ;
  assign n68854 = ~n9770 ;
  assign n10088 = n68854 & n10087 ;
  assign n10089 = n9777 | n10088 ;
  assign n10090 = n10086 | n10089 ;
  assign n68855 = ~n9777 ;
  assign n10091 = n68855 & n10090 ;
  assign n68856 = ~n9767 ;
  assign n10092 = x88 & n68856 ;
  assign n68857 = ~n9762 ;
  assign n10093 = n68857 & n10092 ;
  assign n10094 = n9769 | n10093 ;
  assign n10096 = n10091 | n10094 ;
  assign n68858 = ~n9769 ;
  assign n10097 = n68858 & n10096 ;
  assign n68859 = ~n9759 ;
  assign n10098 = x89 & n68859 ;
  assign n68860 = ~n9754 ;
  assign n10099 = n68860 & n10098 ;
  assign n10100 = n9761 | n10099 ;
  assign n10101 = n10097 | n10100 ;
  assign n68861 = ~n9761 ;
  assign n10102 = n68861 & n10101 ;
  assign n68862 = ~n9751 ;
  assign n10103 = x90 & n68862 ;
  assign n68863 = ~n9746 ;
  assign n10104 = n68863 & n10103 ;
  assign n10105 = n9753 | n10104 ;
  assign n10107 = n10102 | n10105 ;
  assign n68864 = ~n9753 ;
  assign n10108 = n68864 & n10107 ;
  assign n68865 = ~n9743 ;
  assign n10109 = x91 & n68865 ;
  assign n68866 = ~n9738 ;
  assign n10110 = n68866 & n10109 ;
  assign n10111 = n9745 | n10110 ;
  assign n10112 = n10108 | n10111 ;
  assign n68867 = ~n9745 ;
  assign n10113 = n68867 & n10112 ;
  assign n68868 = ~n9735 ;
  assign n10114 = x92 & n68868 ;
  assign n68869 = ~n9730 ;
  assign n10115 = n68869 & n10114 ;
  assign n10116 = n9737 | n10115 ;
  assign n10118 = n10113 | n10116 ;
  assign n68870 = ~n9737 ;
  assign n10119 = n68870 & n10118 ;
  assign n68871 = ~n9727 ;
  assign n10120 = x93 & n68871 ;
  assign n68872 = ~n9722 ;
  assign n10121 = n68872 & n10120 ;
  assign n10122 = n9729 | n10121 ;
  assign n10123 = n10119 | n10122 ;
  assign n68873 = ~n9729 ;
  assign n10124 = n68873 & n10123 ;
  assign n68874 = ~n9719 ;
  assign n10125 = x94 & n68874 ;
  assign n68875 = ~n9714 ;
  assign n10126 = n68875 & n10125 ;
  assign n10127 = n9721 | n10126 ;
  assign n10129 = n10124 | n10127 ;
  assign n68876 = ~n9721 ;
  assign n10130 = n68876 & n10129 ;
  assign n68877 = ~n9711 ;
  assign n10131 = x95 & n68877 ;
  assign n68878 = ~n9706 ;
  assign n10132 = n68878 & n10131 ;
  assign n10133 = n9713 | n10132 ;
  assign n10134 = n10130 | n10133 ;
  assign n68879 = ~n9713 ;
  assign n10135 = n68879 & n10134 ;
  assign n68880 = ~n9703 ;
  assign n10136 = x96 & n68880 ;
  assign n68881 = ~n9698 ;
  assign n10137 = n68881 & n10136 ;
  assign n10138 = n9705 | n10137 ;
  assign n10140 = n10135 | n10138 ;
  assign n68882 = ~n9705 ;
  assign n10141 = n68882 & n10140 ;
  assign n68883 = ~n9695 ;
  assign n10142 = x97 & n68883 ;
  assign n68884 = ~n9690 ;
  assign n10143 = n68884 & n10142 ;
  assign n10144 = n9697 | n10143 ;
  assign n10145 = n10141 | n10144 ;
  assign n68885 = ~n9697 ;
  assign n10146 = n68885 & n10145 ;
  assign n159 = ~n9611 ;
  assign n10147 = n159 & n9686 ;
  assign n10148 = n9155 & n9611 ;
  assign n68887 = ~n10148 ;
  assign n10149 = x98 & n68887 ;
  assign n68888 = ~n10147 ;
  assign n10150 = n68888 & n10149 ;
  assign n10151 = n9689 | n10150 ;
  assign n10153 = n10146 | n10151 ;
  assign n68889 = ~n9689 ;
  assign n10154 = n68889 & n10153 ;
  assign n10155 = n282 | n284 ;
  assign n10156 = n293 | n10155 ;
  assign n10157 = n279 | n10156 ;
  assign n10158 = n10154 | n10157 ;
  assign n10159 = n9696 & n10158 ;
  assign n9960 = n65670 & n9958 ;
  assign n10160 = x65 & n9969 ;
  assign n68890 = ~n10160 ;
  assign n10161 = n9962 & n68890 ;
  assign n10162 = n9964 | n10161 ;
  assign n68891 = ~n9960 ;
  assign n10163 = n68891 & n10162 ;
  assign n10164 = n9975 | n10163 ;
  assign n10165 = n68792 & n10164 ;
  assign n10166 = n9979 | n10165 ;
  assign n10168 = n68795 & n10166 ;
  assign n10170 = n9985 | n10168 ;
  assign n10171 = n68798 & n10170 ;
  assign n10173 = n9990 | n10171 ;
  assign n10174 = n68801 & n10173 ;
  assign n10175 = n9995 | n10174 ;
  assign n10176 = n68804 & n10175 ;
  assign n10177 = n10001 | n10176 ;
  assign n10179 = n68807 & n10177 ;
  assign n10180 = n10006 | n10179 ;
  assign n10181 = n68810 & n10180 ;
  assign n10182 = n10012 | n10181 ;
  assign n10184 = n68813 & n10182 ;
  assign n10185 = n10017 | n10184 ;
  assign n10186 = n68816 & n10185 ;
  assign n10187 = n10023 | n10186 ;
  assign n10189 = n68819 & n10187 ;
  assign n10190 = n10028 | n10189 ;
  assign n10191 = n68822 & n10190 ;
  assign n10192 = n10034 | n10191 ;
  assign n10194 = n68825 & n10192 ;
  assign n10195 = n10039 | n10194 ;
  assign n10196 = n68828 & n10195 ;
  assign n10197 = n10045 | n10196 ;
  assign n10199 = n68831 & n10197 ;
  assign n10200 = n10050 | n10199 ;
  assign n10201 = n68834 & n10200 ;
  assign n10202 = n10056 | n10201 ;
  assign n10204 = n68837 & n10202 ;
  assign n10205 = n10061 | n10204 ;
  assign n10206 = n68840 & n10205 ;
  assign n10207 = n10067 | n10206 ;
  assign n10209 = n68843 & n10207 ;
  assign n10210 = n10072 | n10209 ;
  assign n10211 = n68846 & n10210 ;
  assign n10212 = n10078 | n10211 ;
  assign n10214 = n68849 & n10212 ;
  assign n10215 = n10083 | n10214 ;
  assign n10216 = n68852 & n10215 ;
  assign n10217 = n10089 | n10216 ;
  assign n10219 = n68855 & n10217 ;
  assign n10220 = n10094 | n10219 ;
  assign n10221 = n68858 & n10220 ;
  assign n10222 = n10100 | n10221 ;
  assign n10224 = n68861 & n10222 ;
  assign n10225 = n10105 | n10224 ;
  assign n10226 = n68864 & n10225 ;
  assign n10227 = n10111 | n10226 ;
  assign n10229 = n68867 & n10227 ;
  assign n10230 = n10116 | n10229 ;
  assign n10231 = n68870 & n10230 ;
  assign n10232 = n10122 | n10231 ;
  assign n10234 = n68873 & n10232 ;
  assign n10235 = n10127 | n10234 ;
  assign n10236 = n68876 & n10235 ;
  assign n10237 = n10133 | n10236 ;
  assign n10239 = n68879 & n10237 ;
  assign n10240 = n10138 | n10239 ;
  assign n10241 = n68882 & n10240 ;
  assign n68892 = ~n10241 ;
  assign n10242 = n10144 & n68892 ;
  assign n10244 = n9705 | n10144 ;
  assign n68893 = ~n10244 ;
  assign n10245 = n10140 & n68893 ;
  assign n10246 = n10242 | n10245 ;
  assign n68894 = ~n10157 ;
  assign n10247 = n68894 & n10246 ;
  assign n68895 = ~n10154 ;
  assign n10248 = n68895 & n10247 ;
  assign n10249 = n10159 | n10248 ;
  assign n10250 = n68716 & n10249 ;
  assign n68896 = ~n10248 ;
  assign n10691 = x98 & n68896 ;
  assign n68897 = ~n10159 ;
  assign n10692 = n68897 & n10691 ;
  assign n10693 = n10250 | n10692 ;
  assign n10251 = n9704 & n10158 ;
  assign n68898 = ~n10135 ;
  assign n10139 = n68898 & n10138 ;
  assign n10252 = n9713 | n10138 ;
  assign n68899 = ~n10252 ;
  assign n10253 = n10237 & n68899 ;
  assign n10254 = n10139 | n10253 ;
  assign n10255 = n68894 & n10254 ;
  assign n10256 = n68895 & n10255 ;
  assign n10257 = n10251 | n10256 ;
  assign n10258 = n68545 & n10257 ;
  assign n10259 = n9712 & n10158 ;
  assign n68900 = ~n10236 ;
  assign n10238 = n10133 & n68900 ;
  assign n10260 = n9721 | n10133 ;
  assign n68901 = ~n10260 ;
  assign n10261 = n10129 & n68901 ;
  assign n10262 = n10238 | n10261 ;
  assign n10263 = n68894 & n10262 ;
  assign n10264 = n68895 & n10263 ;
  assign n10265 = n10259 | n10264 ;
  assign n10266 = n68438 & n10265 ;
  assign n68902 = ~n10264 ;
  assign n10681 = x96 & n68902 ;
  assign n68903 = ~n10259 ;
  assign n10682 = n68903 & n10681 ;
  assign n10683 = n10266 | n10682 ;
  assign n10267 = n9720 & n10158 ;
  assign n68904 = ~n10124 ;
  assign n10128 = n68904 & n10127 ;
  assign n10268 = n9729 | n10127 ;
  assign n68905 = ~n10268 ;
  assign n10269 = n10232 & n68905 ;
  assign n10270 = n10128 | n10269 ;
  assign n10271 = n68894 & n10270 ;
  assign n10272 = n68895 & n10271 ;
  assign n10273 = n10267 | n10272 ;
  assign n10274 = n68214 & n10273 ;
  assign n10275 = n9728 & n10158 ;
  assign n68906 = ~n10231 ;
  assign n10233 = n10122 & n68906 ;
  assign n10276 = n9737 | n10122 ;
  assign n68907 = ~n10276 ;
  assign n10277 = n10118 & n68907 ;
  assign n10278 = n10233 | n10277 ;
  assign n10279 = n68894 & n10278 ;
  assign n10280 = n68895 & n10279 ;
  assign n10281 = n10275 | n10280 ;
  assign n10282 = n68058 & n10281 ;
  assign n68908 = ~n10280 ;
  assign n10671 = x94 & n68908 ;
  assign n68909 = ~n10275 ;
  assign n10672 = n68909 & n10671 ;
  assign n10673 = n10282 | n10672 ;
  assign n10283 = n9736 & n10158 ;
  assign n68910 = ~n10113 ;
  assign n10117 = n68910 & n10116 ;
  assign n10284 = n9745 | n10116 ;
  assign n68911 = ~n10284 ;
  assign n10285 = n10227 & n68911 ;
  assign n10286 = n10117 | n10285 ;
  assign n10287 = n68894 & n10286 ;
  assign n10288 = n68895 & n10287 ;
  assign n10289 = n10283 | n10288 ;
  assign n10290 = n67986 & n10289 ;
  assign n10291 = n9744 & n10158 ;
  assign n68912 = ~n10226 ;
  assign n10228 = n10111 & n68912 ;
  assign n10292 = n9753 | n10111 ;
  assign n68913 = ~n10292 ;
  assign n10293 = n10107 & n68913 ;
  assign n10294 = n10228 | n10293 ;
  assign n10295 = n68894 & n10294 ;
  assign n10296 = n68895 & n10295 ;
  assign n10297 = n10291 | n10296 ;
  assign n10298 = n67763 & n10297 ;
  assign n68914 = ~n10296 ;
  assign n10661 = x92 & n68914 ;
  assign n68915 = ~n10291 ;
  assign n10662 = n68915 & n10661 ;
  assign n10663 = n10298 | n10662 ;
  assign n10299 = n9752 & n10158 ;
  assign n68916 = ~n10102 ;
  assign n10106 = n68916 & n10105 ;
  assign n10300 = n9761 | n10105 ;
  assign n68917 = ~n10300 ;
  assign n10301 = n10222 & n68917 ;
  assign n10302 = n10106 | n10301 ;
  assign n10303 = n68894 & n10302 ;
  assign n10304 = n68895 & n10303 ;
  assign n10305 = n10299 | n10304 ;
  assign n10306 = n67622 & n10305 ;
  assign n10307 = n9760 & n10158 ;
  assign n68918 = ~n10221 ;
  assign n10223 = n10100 & n68918 ;
  assign n10308 = n9769 | n10100 ;
  assign n68919 = ~n10308 ;
  assign n10309 = n10096 & n68919 ;
  assign n10310 = n10223 | n10309 ;
  assign n10311 = n68894 & n10310 ;
  assign n10312 = n68895 & n10311 ;
  assign n10313 = n10307 | n10312 ;
  assign n10314 = n67531 & n10313 ;
  assign n68920 = ~n10312 ;
  assign n10651 = x90 & n68920 ;
  assign n68921 = ~n10307 ;
  assign n10652 = n68921 & n10651 ;
  assign n10653 = n10314 | n10652 ;
  assign n10315 = n9768 & n10158 ;
  assign n68922 = ~n10091 ;
  assign n10095 = n68922 & n10094 ;
  assign n10316 = n9777 | n10094 ;
  assign n68923 = ~n10316 ;
  assign n10317 = n10217 & n68923 ;
  assign n10318 = n10095 | n10317 ;
  assign n10319 = n68894 & n10318 ;
  assign n10320 = n68895 & n10319 ;
  assign n10321 = n10315 | n10320 ;
  assign n10322 = n67348 & n10321 ;
  assign n10323 = n9776 & n10158 ;
  assign n68924 = ~n10216 ;
  assign n10218 = n10089 & n68924 ;
  assign n10324 = n9785 | n10089 ;
  assign n68925 = ~n10324 ;
  assign n10325 = n10085 & n68925 ;
  assign n10326 = n10218 | n10325 ;
  assign n10327 = n68894 & n10326 ;
  assign n10328 = n68895 & n10327 ;
  assign n10329 = n10323 | n10328 ;
  assign n10330 = n67222 & n10329 ;
  assign n68926 = ~n10328 ;
  assign n10641 = x88 & n68926 ;
  assign n68927 = ~n10323 ;
  assign n10642 = n68927 & n10641 ;
  assign n10643 = n10330 | n10642 ;
  assign n10331 = n9784 & n10158 ;
  assign n68928 = ~n10080 ;
  assign n10084 = n68928 & n10083 ;
  assign n10332 = n9793 | n10083 ;
  assign n68929 = ~n10332 ;
  assign n10333 = n10212 & n68929 ;
  assign n10334 = n10084 | n10333 ;
  assign n10335 = n68894 & n10334 ;
  assign n10336 = n68895 & n10335 ;
  assign n10337 = n10331 | n10336 ;
  assign n10338 = n67164 & n10337 ;
  assign n10339 = n9792 & n10158 ;
  assign n68930 = ~n10211 ;
  assign n10213 = n10078 & n68930 ;
  assign n10340 = n9801 | n10078 ;
  assign n68931 = ~n10340 ;
  assign n10341 = n10074 & n68931 ;
  assign n10342 = n10213 | n10341 ;
  assign n10343 = n68894 & n10342 ;
  assign n10344 = n68895 & n10343 ;
  assign n10345 = n10339 | n10344 ;
  assign n10346 = n66979 & n10345 ;
  assign n68932 = ~n10344 ;
  assign n10631 = x86 & n68932 ;
  assign n68933 = ~n10339 ;
  assign n10632 = n68933 & n10631 ;
  assign n10633 = n10346 | n10632 ;
  assign n10347 = n9800 & n10158 ;
  assign n68934 = ~n10069 ;
  assign n10073 = n68934 & n10072 ;
  assign n10348 = n9809 | n10072 ;
  assign n68935 = ~n10348 ;
  assign n10349 = n10207 & n68935 ;
  assign n10350 = n10073 | n10349 ;
  assign n10351 = n68894 & n10350 ;
  assign n10352 = n68895 & n10351 ;
  assign n10353 = n10347 | n10352 ;
  assign n10354 = n66868 & n10353 ;
  assign n10355 = n9808 & n10158 ;
  assign n68936 = ~n10206 ;
  assign n10208 = n10067 & n68936 ;
  assign n10356 = n9817 | n10067 ;
  assign n68937 = ~n10356 ;
  assign n10357 = n10063 & n68937 ;
  assign n10358 = n10208 | n10357 ;
  assign n10359 = n68894 & n10358 ;
  assign n10360 = n68895 & n10359 ;
  assign n10361 = n10355 | n10360 ;
  assign n10362 = n66797 & n10361 ;
  assign n68938 = ~n10360 ;
  assign n10621 = x84 & n68938 ;
  assign n68939 = ~n10355 ;
  assign n10622 = n68939 & n10621 ;
  assign n10623 = n10362 | n10622 ;
  assign n10363 = n9816 & n10158 ;
  assign n68940 = ~n10058 ;
  assign n10062 = n68940 & n10061 ;
  assign n10364 = n9825 | n10061 ;
  assign n68941 = ~n10364 ;
  assign n10365 = n10202 & n68941 ;
  assign n10366 = n10062 | n10365 ;
  assign n10367 = n68894 & n10366 ;
  assign n10368 = n68895 & n10367 ;
  assign n10369 = n10363 | n10368 ;
  assign n10370 = n66654 & n10369 ;
  assign n10371 = n9824 & n10158 ;
  assign n68942 = ~n10201 ;
  assign n10203 = n10056 & n68942 ;
  assign n10372 = n9833 | n10056 ;
  assign n68943 = ~n10372 ;
  assign n10373 = n10052 & n68943 ;
  assign n10374 = n10203 | n10373 ;
  assign n10375 = n68894 & n10374 ;
  assign n10376 = n68895 & n10375 ;
  assign n10377 = n10371 | n10376 ;
  assign n10378 = n66560 & n10377 ;
  assign n68944 = ~n10376 ;
  assign n10611 = x82 & n68944 ;
  assign n68945 = ~n10371 ;
  assign n10612 = n68945 & n10611 ;
  assign n10613 = n10378 | n10612 ;
  assign n10379 = n9832 & n10158 ;
  assign n68946 = ~n10047 ;
  assign n10051 = n68946 & n10050 ;
  assign n10380 = n9841 | n10050 ;
  assign n68947 = ~n10380 ;
  assign n10381 = n10197 & n68947 ;
  assign n10382 = n10051 | n10381 ;
  assign n10383 = n68894 & n10382 ;
  assign n10384 = n68895 & n10383 ;
  assign n10385 = n10379 | n10384 ;
  assign n10386 = n66505 & n10385 ;
  assign n10387 = n9840 & n10158 ;
  assign n68948 = ~n10196 ;
  assign n10198 = n10045 & n68948 ;
  assign n10388 = n9849 | n10045 ;
  assign n68949 = ~n10388 ;
  assign n10389 = n10041 & n68949 ;
  assign n10390 = n10198 | n10389 ;
  assign n10391 = n68894 & n10390 ;
  assign n10392 = n68895 & n10391 ;
  assign n10393 = n10387 | n10392 ;
  assign n10394 = n66379 & n10393 ;
  assign n68950 = ~n10392 ;
  assign n10601 = x80 & n68950 ;
  assign n68951 = ~n10387 ;
  assign n10602 = n68951 & n10601 ;
  assign n10603 = n10394 | n10602 ;
  assign n10395 = n9848 & n10158 ;
  assign n68952 = ~n10036 ;
  assign n10040 = n68952 & n10039 ;
  assign n10396 = n9857 | n10039 ;
  assign n68953 = ~n10396 ;
  assign n10397 = n10192 & n68953 ;
  assign n10398 = n10040 | n10397 ;
  assign n10399 = n68894 & n10398 ;
  assign n10400 = n68895 & n10399 ;
  assign n10401 = n10395 | n10400 ;
  assign n10402 = n66299 & n10401 ;
  assign n10403 = n9856 & n10158 ;
  assign n68954 = ~n10191 ;
  assign n10193 = n10034 & n68954 ;
  assign n10404 = n9865 | n10034 ;
  assign n68955 = ~n10404 ;
  assign n10405 = n10030 & n68955 ;
  assign n10406 = n10193 | n10405 ;
  assign n10407 = n68894 & n10406 ;
  assign n10408 = n68895 & n10407 ;
  assign n10409 = n10403 | n10408 ;
  assign n10410 = n66244 & n10409 ;
  assign n68956 = ~n10408 ;
  assign n10591 = x78 & n68956 ;
  assign n68957 = ~n10403 ;
  assign n10592 = n68957 & n10591 ;
  assign n10593 = n10410 | n10592 ;
  assign n10411 = n9864 & n10158 ;
  assign n68958 = ~n10025 ;
  assign n10029 = n68958 & n10028 ;
  assign n10412 = n9873 | n10028 ;
  assign n68959 = ~n10412 ;
  assign n10413 = n10187 & n68959 ;
  assign n10414 = n10029 | n10413 ;
  assign n10415 = n68894 & n10414 ;
  assign n10416 = n68895 & n10415 ;
  assign n10417 = n10411 | n10416 ;
  assign n10418 = n66145 & n10417 ;
  assign n10419 = n9872 & n10158 ;
  assign n68960 = ~n10186 ;
  assign n10188 = n10023 & n68960 ;
  assign n10420 = n9881 | n10023 ;
  assign n68961 = ~n10420 ;
  assign n10421 = n10019 & n68961 ;
  assign n10422 = n10188 | n10421 ;
  assign n10423 = n68894 & n10422 ;
  assign n10424 = n68895 & n10423 ;
  assign n10425 = n10419 | n10424 ;
  assign n10426 = n66081 & n10425 ;
  assign n68962 = ~n10424 ;
  assign n10581 = x76 & n68962 ;
  assign n68963 = ~n10419 ;
  assign n10582 = n68963 & n10581 ;
  assign n10583 = n10426 | n10582 ;
  assign n10427 = n9880 & n10158 ;
  assign n68964 = ~n10014 ;
  assign n10018 = n68964 & n10017 ;
  assign n10428 = n9889 | n10017 ;
  assign n68965 = ~n10428 ;
  assign n10429 = n10182 & n68965 ;
  assign n10430 = n10018 | n10429 ;
  assign n10431 = n68894 & n10430 ;
  assign n10432 = n68895 & n10431 ;
  assign n10433 = n10427 | n10432 ;
  assign n10434 = n66043 & n10433 ;
  assign n10435 = n9888 & n10158 ;
  assign n68966 = ~n10181 ;
  assign n10183 = n10012 & n68966 ;
  assign n10436 = n9897 | n10012 ;
  assign n68967 = ~n10436 ;
  assign n10437 = n10008 & n68967 ;
  assign n10438 = n10183 | n10437 ;
  assign n10439 = n68894 & n10438 ;
  assign n10440 = n68895 & n10439 ;
  assign n10441 = n10435 | n10440 ;
  assign n10442 = n65960 & n10441 ;
  assign n68968 = ~n10440 ;
  assign n10571 = x74 & n68968 ;
  assign n68969 = ~n10435 ;
  assign n10572 = n68969 & n10571 ;
  assign n10573 = n10442 | n10572 ;
  assign n10443 = n9896 & n10158 ;
  assign n68970 = ~n10003 ;
  assign n10007 = n68970 & n10006 ;
  assign n10444 = n9905 | n10006 ;
  assign n68971 = ~n10444 ;
  assign n10445 = n10177 & n68971 ;
  assign n10446 = n10007 | n10445 ;
  assign n10447 = n68894 & n10446 ;
  assign n10448 = n68895 & n10447 ;
  assign n10449 = n10443 | n10448 ;
  assign n10450 = n65909 & n10449 ;
  assign n10451 = n9904 & n10158 ;
  assign n68972 = ~n10176 ;
  assign n10178 = n10001 & n68972 ;
  assign n10452 = n9913 | n10001 ;
  assign n68973 = ~n10452 ;
  assign n10453 = n9997 & n68973 ;
  assign n10454 = n10178 | n10453 ;
  assign n10455 = n68894 & n10454 ;
  assign n10456 = n68895 & n10455 ;
  assign n10457 = n10451 | n10456 ;
  assign n10458 = n65877 & n10457 ;
  assign n68974 = ~n10456 ;
  assign n10561 = x72 & n68974 ;
  assign n68975 = ~n10451 ;
  assign n10562 = n68975 & n10561 ;
  assign n10563 = n10458 | n10562 ;
  assign n10459 = n9912 & n10158 ;
  assign n68976 = ~n9992 ;
  assign n9996 = n68976 & n9995 ;
  assign n10460 = n9922 | n9995 ;
  assign n68977 = ~n10460 ;
  assign n10461 = n10173 & n68977 ;
  assign n10462 = n9996 | n10461 ;
  assign n10463 = n68894 & n10462 ;
  assign n10464 = n68895 & n10463 ;
  assign n10465 = n10459 | n10464 ;
  assign n10466 = n65820 & n10465 ;
  assign n10467 = n9921 & n10158 ;
  assign n68978 = ~n10171 ;
  assign n10172 = n9990 & n68978 ;
  assign n10468 = n9931 | n9990 ;
  assign n68979 = ~n10468 ;
  assign n10469 = n10170 & n68979 ;
  assign n10470 = n10172 | n10469 ;
  assign n10471 = n68894 & n10470 ;
  assign n10472 = n68895 & n10471 ;
  assign n10473 = n10467 | n10472 ;
  assign n10474 = n65791 & n10473 ;
  assign n68980 = ~n10472 ;
  assign n10551 = x70 & n68980 ;
  assign n68981 = ~n10467 ;
  assign n10552 = n68981 & n10551 ;
  assign n10553 = n10474 | n10552 ;
  assign n10475 = n9930 & n10158 ;
  assign n68982 = ~n9982 ;
  assign n10169 = n68982 & n9985 ;
  assign n10476 = n9980 | n10165 ;
  assign n10477 = n9939 | n9985 ;
  assign n68983 = ~n10477 ;
  assign n10478 = n10476 & n68983 ;
  assign n10479 = n10169 | n10478 ;
  assign n10480 = n68894 & n10479 ;
  assign n10481 = n68895 & n10480 ;
  assign n10482 = n10475 | n10481 ;
  assign n10483 = n65772 & n10482 ;
  assign n10484 = n9938 & n10158 ;
  assign n68984 = ~n10165 ;
  assign n10167 = n9980 & n68984 ;
  assign n10485 = n9945 | n9980 ;
  assign n68985 = ~n10485 ;
  assign n10486 = n10164 & n68985 ;
  assign n10487 = n10167 | n10486 ;
  assign n10488 = n68894 & n10487 ;
  assign n10489 = n68895 & n10488 ;
  assign n10490 = n10484 | n10489 ;
  assign n10491 = n65746 & n10490 ;
  assign n68986 = ~n10489 ;
  assign n10541 = x68 & n68986 ;
  assign n68987 = ~n10484 ;
  assign n10542 = n68987 & n10541 ;
  assign n10543 = n10491 | n10542 ;
  assign n10492 = n9944 & n10158 ;
  assign n10493 = n9970 | n9975 ;
  assign n68988 = ~n10493 ;
  assign n10494 = n10162 & n68988 ;
  assign n68989 = ~n9972 ;
  assign n10495 = n68989 & n9975 ;
  assign n10496 = n10494 | n10495 ;
  assign n10497 = n68894 & n10496 ;
  assign n10498 = n68895 & n10497 ;
  assign n10499 = n10492 | n10498 ;
  assign n10501 = n65721 & n10499 ;
  assign n10502 = n9958 & n10158 ;
  assign n10503 = n9962 & n9964 ;
  assign n10504 = n68890 & n10503 ;
  assign n10505 = n10157 | n10504 ;
  assign n68990 = ~n10505 ;
  assign n10506 = n10162 & n68990 ;
  assign n10507 = n68895 & n10506 ;
  assign n10508 = n10502 | n10507 ;
  assign n10509 = n65686 & n10508 ;
  assign n68991 = ~n10507 ;
  assign n10532 = x66 & n68991 ;
  assign n68992 = ~n10502 ;
  assign n10533 = n68992 & n10532 ;
  assign n10534 = n10509 | n10533 ;
  assign n10243 = n10144 | n10241 ;
  assign n10510 = n68885 & n10243 ;
  assign n10511 = n10151 | n10510 ;
  assign n10512 = n68889 & n10511 ;
  assign n68993 = ~x99 ;
  assign n10513 = x64 & n68993 ;
  assign n10514 = n68779 & n10513 ;
  assign n10515 = n68780 & n10514 ;
  assign n10516 = n66510 & n10515 ;
  assign n68994 = ~n10512 ;
  assign n10517 = n68994 & n10516 ;
  assign n68995 = ~n10517 ;
  assign n10518 = x29 & n68995 ;
  assign n10519 = n68781 & n9964 ;
  assign n10520 = n68782 & n10519 ;
  assign n10521 = n68783 & n10520 ;
  assign n10522 = n66715 & n10521 ;
  assign n10523 = n68895 & n10522 ;
  assign n10524 = n10518 | n10523 ;
  assign n10525 = x65 & n10524 ;
  assign n10526 = x65 | n10523 ;
  assign n10527 = n10518 | n10526 ;
  assign n68996 = ~n10525 ;
  assign n10528 = n68996 & n10527 ;
  assign n68997 = ~x28 ;
  assign n10529 = n68997 & x64 ;
  assign n10530 = n10528 | n10529 ;
  assign n10531 = n65670 & n10524 ;
  assign n68998 = ~n10531 ;
  assign n10535 = n10530 & n68998 ;
  assign n10536 = n10534 | n10535 ;
  assign n68999 = ~n10509 ;
  assign n10537 = n68999 & n10536 ;
  assign n69000 = ~n10498 ;
  assign n10500 = x67 & n69000 ;
  assign n69001 = ~n10492 ;
  assign n10538 = n69001 & n10500 ;
  assign n10539 = n10501 | n10538 ;
  assign n10540 = n10537 | n10539 ;
  assign n69002 = ~n10501 ;
  assign n10544 = n69002 & n10540 ;
  assign n10545 = n10543 | n10544 ;
  assign n69003 = ~n10491 ;
  assign n10546 = n69003 & n10545 ;
  assign n69004 = ~n10481 ;
  assign n10547 = x69 & n69004 ;
  assign n69005 = ~n10475 ;
  assign n10548 = n69005 & n10547 ;
  assign n10549 = n10483 | n10548 ;
  assign n10550 = n10546 | n10549 ;
  assign n69006 = ~n10483 ;
  assign n10554 = n69006 & n10550 ;
  assign n10555 = n10553 | n10554 ;
  assign n69007 = ~n10474 ;
  assign n10556 = n69007 & n10555 ;
  assign n69008 = ~n10464 ;
  assign n10557 = x71 & n69008 ;
  assign n69009 = ~n10459 ;
  assign n10558 = n69009 & n10557 ;
  assign n10559 = n10466 | n10558 ;
  assign n10560 = n10556 | n10559 ;
  assign n69010 = ~n10466 ;
  assign n10564 = n69010 & n10560 ;
  assign n10565 = n10563 | n10564 ;
  assign n69011 = ~n10458 ;
  assign n10566 = n69011 & n10565 ;
  assign n69012 = ~n10448 ;
  assign n10567 = x73 & n69012 ;
  assign n69013 = ~n10443 ;
  assign n10568 = n69013 & n10567 ;
  assign n10569 = n10450 | n10568 ;
  assign n10570 = n10566 | n10569 ;
  assign n69014 = ~n10450 ;
  assign n10574 = n69014 & n10570 ;
  assign n10575 = n10573 | n10574 ;
  assign n69015 = ~n10442 ;
  assign n10576 = n69015 & n10575 ;
  assign n69016 = ~n10432 ;
  assign n10577 = x75 & n69016 ;
  assign n69017 = ~n10427 ;
  assign n10578 = n69017 & n10577 ;
  assign n10579 = n10434 | n10578 ;
  assign n10580 = n10576 | n10579 ;
  assign n69018 = ~n10434 ;
  assign n10584 = n69018 & n10580 ;
  assign n10585 = n10583 | n10584 ;
  assign n69019 = ~n10426 ;
  assign n10586 = n69019 & n10585 ;
  assign n69020 = ~n10416 ;
  assign n10587 = x77 & n69020 ;
  assign n69021 = ~n10411 ;
  assign n10588 = n69021 & n10587 ;
  assign n10589 = n10418 | n10588 ;
  assign n10590 = n10586 | n10589 ;
  assign n69022 = ~n10418 ;
  assign n10594 = n69022 & n10590 ;
  assign n10595 = n10593 | n10594 ;
  assign n69023 = ~n10410 ;
  assign n10596 = n69023 & n10595 ;
  assign n69024 = ~n10400 ;
  assign n10597 = x79 & n69024 ;
  assign n69025 = ~n10395 ;
  assign n10598 = n69025 & n10597 ;
  assign n10599 = n10402 | n10598 ;
  assign n10600 = n10596 | n10599 ;
  assign n69026 = ~n10402 ;
  assign n10604 = n69026 & n10600 ;
  assign n10605 = n10603 | n10604 ;
  assign n69027 = ~n10394 ;
  assign n10606 = n69027 & n10605 ;
  assign n69028 = ~n10384 ;
  assign n10607 = x81 & n69028 ;
  assign n69029 = ~n10379 ;
  assign n10608 = n69029 & n10607 ;
  assign n10609 = n10386 | n10608 ;
  assign n10610 = n10606 | n10609 ;
  assign n69030 = ~n10386 ;
  assign n10614 = n69030 & n10610 ;
  assign n10615 = n10613 | n10614 ;
  assign n69031 = ~n10378 ;
  assign n10616 = n69031 & n10615 ;
  assign n69032 = ~n10368 ;
  assign n10617 = x83 & n69032 ;
  assign n69033 = ~n10363 ;
  assign n10618 = n69033 & n10617 ;
  assign n10619 = n10370 | n10618 ;
  assign n10620 = n10616 | n10619 ;
  assign n69034 = ~n10370 ;
  assign n10624 = n69034 & n10620 ;
  assign n10625 = n10623 | n10624 ;
  assign n69035 = ~n10362 ;
  assign n10626 = n69035 & n10625 ;
  assign n69036 = ~n10352 ;
  assign n10627 = x85 & n69036 ;
  assign n69037 = ~n10347 ;
  assign n10628 = n69037 & n10627 ;
  assign n10629 = n10354 | n10628 ;
  assign n10630 = n10626 | n10629 ;
  assign n69038 = ~n10354 ;
  assign n10634 = n69038 & n10630 ;
  assign n10635 = n10633 | n10634 ;
  assign n69039 = ~n10346 ;
  assign n10636 = n69039 & n10635 ;
  assign n69040 = ~n10336 ;
  assign n10637 = x87 & n69040 ;
  assign n69041 = ~n10331 ;
  assign n10638 = n69041 & n10637 ;
  assign n10639 = n10338 | n10638 ;
  assign n10640 = n10636 | n10639 ;
  assign n69042 = ~n10338 ;
  assign n10644 = n69042 & n10640 ;
  assign n10645 = n10643 | n10644 ;
  assign n69043 = ~n10330 ;
  assign n10646 = n69043 & n10645 ;
  assign n69044 = ~n10320 ;
  assign n10647 = x89 & n69044 ;
  assign n69045 = ~n10315 ;
  assign n10648 = n69045 & n10647 ;
  assign n10649 = n10322 | n10648 ;
  assign n10650 = n10646 | n10649 ;
  assign n69046 = ~n10322 ;
  assign n10654 = n69046 & n10650 ;
  assign n10655 = n10653 | n10654 ;
  assign n69047 = ~n10314 ;
  assign n10656 = n69047 & n10655 ;
  assign n69048 = ~n10304 ;
  assign n10657 = x91 & n69048 ;
  assign n69049 = ~n10299 ;
  assign n10658 = n69049 & n10657 ;
  assign n10659 = n10306 | n10658 ;
  assign n10660 = n10656 | n10659 ;
  assign n69050 = ~n10306 ;
  assign n10664 = n69050 & n10660 ;
  assign n10665 = n10663 | n10664 ;
  assign n69051 = ~n10298 ;
  assign n10666 = n69051 & n10665 ;
  assign n69052 = ~n10288 ;
  assign n10667 = x93 & n69052 ;
  assign n69053 = ~n10283 ;
  assign n10668 = n69053 & n10667 ;
  assign n10669 = n10290 | n10668 ;
  assign n10670 = n10666 | n10669 ;
  assign n69054 = ~n10290 ;
  assign n10674 = n69054 & n10670 ;
  assign n10675 = n10673 | n10674 ;
  assign n69055 = ~n10282 ;
  assign n10676 = n69055 & n10675 ;
  assign n69056 = ~n10272 ;
  assign n10677 = x95 & n69056 ;
  assign n69057 = ~n10267 ;
  assign n10678 = n69057 & n10677 ;
  assign n10679 = n10274 | n10678 ;
  assign n10680 = n10676 | n10679 ;
  assign n69058 = ~n10274 ;
  assign n10684 = n69058 & n10680 ;
  assign n10685 = n10683 | n10684 ;
  assign n69059 = ~n10266 ;
  assign n10686 = n69059 & n10685 ;
  assign n69060 = ~n10256 ;
  assign n10687 = x97 & n69060 ;
  assign n69061 = ~n10251 ;
  assign n10688 = n69061 & n10687 ;
  assign n10689 = n10258 | n10688 ;
  assign n10690 = n10686 | n10689 ;
  assign n69062 = ~n10258 ;
  assign n10694 = n69062 & n10690 ;
  assign n10695 = n10693 | n10694 ;
  assign n69063 = ~n10250 ;
  assign n10696 = n69063 & n10695 ;
  assign n69064 = ~n10146 ;
  assign n10152 = n69064 & n10151 ;
  assign n10697 = n9697 | n10151 ;
  assign n69065 = ~n10697 ;
  assign n10698 = n10243 & n69065 ;
  assign n10699 = n10152 | n10698 ;
  assign n10700 = n10158 | n10699 ;
  assign n69066 = ~n9688 ;
  assign n10701 = n69066 & n10158 ;
  assign n69067 = ~n10701 ;
  assign n10702 = n10700 & n69067 ;
  assign n10703 = n68993 & n10702 ;
  assign n158 = ~n10158 ;
  assign n10704 = n158 & n10699 ;
  assign n10705 = n9688 & n10158 ;
  assign n69069 = ~n10705 ;
  assign n10706 = x99 & n69069 ;
  assign n69070 = ~n10704 ;
  assign n10707 = n69070 & n10706 ;
  assign n10708 = n380 | n10707 ;
  assign n10709 = n10703 | n10708 ;
  assign n10710 = n10696 | n10709 ;
  assign n10711 = n68894 & n10702 ;
  assign n69071 = ~n10711 ;
  assign n10712 = n10710 & n69071 ;
  assign n10714 = n10250 | n10707 ;
  assign n10715 = n10703 | n10714 ;
  assign n69072 = ~n10715 ;
  assign n10716 = n10695 & n69072 ;
  assign n10717 = n10703 | n10707 ;
  assign n69073 = ~n10696 ;
  assign n10718 = n69073 & n10717 ;
  assign n10719 = n10716 | n10718 ;
  assign n157 = ~n10712 ;
  assign n10720 = n157 & n10719 ;
  assign n10721 = n10157 & n10702 ;
  assign n10722 = n10710 & n10721 ;
  assign n10723 = n10720 | n10722 ;
  assign n69075 = ~x100 ;
  assign n10724 = n69075 & n10723 ;
  assign n69076 = ~n10694 ;
  assign n10796 = n10693 & n69076 ;
  assign n10725 = n68895 & n10516 ;
  assign n69077 = ~n10725 ;
  assign n10726 = x29 & n69077 ;
  assign n10727 = n10523 | n10726 ;
  assign n10728 = x65 & n10727 ;
  assign n69078 = ~n10728 ;
  assign n10729 = n10527 & n69078 ;
  assign n10730 = n10529 | n10729 ;
  assign n10731 = n68998 & n10730 ;
  assign n10732 = n10534 | n10731 ;
  assign n10733 = n68999 & n10732 ;
  assign n10734 = n10539 | n10733 ;
  assign n10735 = n69002 & n10734 ;
  assign n10736 = n10543 | n10735 ;
  assign n10737 = n69003 & n10736 ;
  assign n10738 = n10549 | n10737 ;
  assign n10739 = n69006 & n10738 ;
  assign n10740 = n10553 | n10739 ;
  assign n10741 = n69007 & n10740 ;
  assign n10742 = n10559 | n10741 ;
  assign n10743 = n69010 & n10742 ;
  assign n10744 = n10563 | n10743 ;
  assign n10745 = n69011 & n10744 ;
  assign n10746 = n10569 | n10745 ;
  assign n10747 = n69014 & n10746 ;
  assign n10748 = n10573 | n10747 ;
  assign n10749 = n69015 & n10748 ;
  assign n10750 = n10579 | n10749 ;
  assign n10751 = n69018 & n10750 ;
  assign n10752 = n10583 | n10751 ;
  assign n10753 = n69019 & n10752 ;
  assign n10754 = n10589 | n10753 ;
  assign n10755 = n69022 & n10754 ;
  assign n10756 = n10593 | n10755 ;
  assign n10757 = n69023 & n10756 ;
  assign n10758 = n10599 | n10757 ;
  assign n10759 = n69026 & n10758 ;
  assign n10760 = n10603 | n10759 ;
  assign n10761 = n69027 & n10760 ;
  assign n10762 = n10609 | n10761 ;
  assign n10763 = n69030 & n10762 ;
  assign n10764 = n10613 | n10763 ;
  assign n10765 = n69031 & n10764 ;
  assign n10766 = n10619 | n10765 ;
  assign n10767 = n69034 & n10766 ;
  assign n10768 = n10623 | n10767 ;
  assign n10769 = n69035 & n10768 ;
  assign n10770 = n10629 | n10769 ;
  assign n10771 = n69038 & n10770 ;
  assign n10772 = n10633 | n10771 ;
  assign n10773 = n69039 & n10772 ;
  assign n10774 = n10639 | n10773 ;
  assign n10775 = n69042 & n10774 ;
  assign n10776 = n10643 | n10775 ;
  assign n10777 = n69043 & n10776 ;
  assign n10778 = n10649 | n10777 ;
  assign n10779 = n69046 & n10778 ;
  assign n10780 = n10653 | n10779 ;
  assign n10781 = n69047 & n10780 ;
  assign n10782 = n10659 | n10781 ;
  assign n10783 = n69050 & n10782 ;
  assign n10784 = n10663 | n10783 ;
  assign n10785 = n69051 & n10784 ;
  assign n10786 = n10669 | n10785 ;
  assign n10787 = n69054 & n10786 ;
  assign n10788 = n10673 | n10787 ;
  assign n10789 = n69055 & n10788 ;
  assign n10790 = n10679 | n10789 ;
  assign n10791 = n69058 & n10790 ;
  assign n10792 = n10683 | n10791 ;
  assign n10793 = n69059 & n10792 ;
  assign n10794 = n10689 | n10793 ;
  assign n10797 = n10258 | n10693 ;
  assign n69079 = ~n10797 ;
  assign n10798 = n10794 & n69079 ;
  assign n10799 = n10796 | n10798 ;
  assign n10800 = n157 & n10799 ;
  assign n10801 = n10249 & n69071 ;
  assign n10802 = n10710 & n10801 ;
  assign n10803 = n10800 | n10802 ;
  assign n10804 = n68993 & n10803 ;
  assign n69080 = ~n10793 ;
  assign n10805 = n10689 & n69080 ;
  assign n10806 = n10266 | n10689 ;
  assign n69081 = ~n10806 ;
  assign n10807 = n10685 & n69081 ;
  assign n10808 = n10805 | n10807 ;
  assign n10809 = n157 & n10808 ;
  assign n10810 = n10257 & n69071 ;
  assign n10811 = n10710 & n10810 ;
  assign n10812 = n10809 | n10811 ;
  assign n10813 = n68716 & n10812 ;
  assign n69082 = ~n10684 ;
  assign n10814 = n10683 & n69082 ;
  assign n10815 = n10274 | n10683 ;
  assign n69083 = ~n10815 ;
  assign n10816 = n10790 & n69083 ;
  assign n10817 = n10814 | n10816 ;
  assign n10818 = n157 & n10817 ;
  assign n10819 = n10265 & n69071 ;
  assign n10820 = n10710 & n10819 ;
  assign n10821 = n10818 | n10820 ;
  assign n10822 = n68545 & n10821 ;
  assign n69084 = ~n10789 ;
  assign n10823 = n10679 & n69084 ;
  assign n10824 = n10282 | n10679 ;
  assign n69085 = ~n10824 ;
  assign n10825 = n10675 & n69085 ;
  assign n10826 = n10823 | n10825 ;
  assign n10827 = n157 & n10826 ;
  assign n10828 = n10273 & n69071 ;
  assign n10829 = n10710 & n10828 ;
  assign n10830 = n10827 | n10829 ;
  assign n10831 = n68438 & n10830 ;
  assign n69086 = ~n10674 ;
  assign n10832 = n10673 & n69086 ;
  assign n10833 = n10290 | n10673 ;
  assign n69087 = ~n10833 ;
  assign n10834 = n10786 & n69087 ;
  assign n10835 = n10832 | n10834 ;
  assign n10836 = n157 & n10835 ;
  assign n10837 = n10281 & n69071 ;
  assign n10838 = n10710 & n10837 ;
  assign n10839 = n10836 | n10838 ;
  assign n10840 = n68214 & n10839 ;
  assign n69088 = ~n10785 ;
  assign n10841 = n10669 & n69088 ;
  assign n10842 = n10298 | n10669 ;
  assign n69089 = ~n10842 ;
  assign n10843 = n10665 & n69089 ;
  assign n10844 = n10841 | n10843 ;
  assign n10845 = n157 & n10844 ;
  assign n10846 = n10289 & n69071 ;
  assign n10847 = n10710 & n10846 ;
  assign n10848 = n10845 | n10847 ;
  assign n10849 = n68058 & n10848 ;
  assign n69090 = ~n10664 ;
  assign n10850 = n10663 & n69090 ;
  assign n10851 = n10306 | n10663 ;
  assign n69091 = ~n10851 ;
  assign n10852 = n10782 & n69091 ;
  assign n10853 = n10850 | n10852 ;
  assign n10854 = n157 & n10853 ;
  assign n10855 = n10297 & n69071 ;
  assign n10856 = n10710 & n10855 ;
  assign n10857 = n10854 | n10856 ;
  assign n10858 = n67986 & n10857 ;
  assign n69092 = ~n10781 ;
  assign n10859 = n10659 & n69092 ;
  assign n10860 = n10314 | n10659 ;
  assign n69093 = ~n10860 ;
  assign n10861 = n10655 & n69093 ;
  assign n10862 = n10859 | n10861 ;
  assign n10863 = n157 & n10862 ;
  assign n10864 = n10305 & n69071 ;
  assign n10865 = n10710 & n10864 ;
  assign n10866 = n10863 | n10865 ;
  assign n10867 = n67763 & n10866 ;
  assign n69094 = ~n10654 ;
  assign n10868 = n10653 & n69094 ;
  assign n10869 = n10322 | n10653 ;
  assign n69095 = ~n10869 ;
  assign n10870 = n10778 & n69095 ;
  assign n10871 = n10868 | n10870 ;
  assign n10872 = n157 & n10871 ;
  assign n10873 = n10313 & n69071 ;
  assign n10874 = n10710 & n10873 ;
  assign n10875 = n10872 | n10874 ;
  assign n10876 = n67622 & n10875 ;
  assign n69096 = ~n10777 ;
  assign n10877 = n10649 & n69096 ;
  assign n10878 = n10330 | n10649 ;
  assign n69097 = ~n10878 ;
  assign n10879 = n10645 & n69097 ;
  assign n10880 = n10877 | n10879 ;
  assign n10881 = n157 & n10880 ;
  assign n10882 = n10321 & n69071 ;
  assign n10883 = n10710 & n10882 ;
  assign n10884 = n10881 | n10883 ;
  assign n10885 = n67531 & n10884 ;
  assign n69098 = ~n10644 ;
  assign n10886 = n10643 & n69098 ;
  assign n10887 = n10338 | n10643 ;
  assign n69099 = ~n10887 ;
  assign n10888 = n10774 & n69099 ;
  assign n10889 = n10886 | n10888 ;
  assign n10890 = n157 & n10889 ;
  assign n10891 = n10329 & n69071 ;
  assign n10892 = n10710 & n10891 ;
  assign n10893 = n10890 | n10892 ;
  assign n10894 = n67348 & n10893 ;
  assign n69100 = ~n10773 ;
  assign n10895 = n10639 & n69100 ;
  assign n10896 = n10346 | n10639 ;
  assign n69101 = ~n10896 ;
  assign n10897 = n10635 & n69101 ;
  assign n10898 = n10895 | n10897 ;
  assign n10899 = n157 & n10898 ;
  assign n10900 = n10337 & n69071 ;
  assign n10901 = n10710 & n10900 ;
  assign n10902 = n10899 | n10901 ;
  assign n10903 = n67222 & n10902 ;
  assign n69102 = ~n10634 ;
  assign n10904 = n10633 & n69102 ;
  assign n10905 = n10354 | n10633 ;
  assign n69103 = ~n10905 ;
  assign n10906 = n10770 & n69103 ;
  assign n10907 = n10904 | n10906 ;
  assign n10908 = n157 & n10907 ;
  assign n10909 = n10345 & n69071 ;
  assign n10910 = n10710 & n10909 ;
  assign n10911 = n10908 | n10910 ;
  assign n10912 = n67164 & n10911 ;
  assign n69104 = ~n10769 ;
  assign n10913 = n10629 & n69104 ;
  assign n10914 = n10362 | n10629 ;
  assign n69105 = ~n10914 ;
  assign n10915 = n10625 & n69105 ;
  assign n10916 = n10913 | n10915 ;
  assign n10917 = n157 & n10916 ;
  assign n10918 = n10353 & n69071 ;
  assign n10919 = n10710 & n10918 ;
  assign n10920 = n10917 | n10919 ;
  assign n10921 = n66979 & n10920 ;
  assign n69106 = ~n10624 ;
  assign n10922 = n10623 & n69106 ;
  assign n10923 = n10370 | n10623 ;
  assign n69107 = ~n10923 ;
  assign n10924 = n10766 & n69107 ;
  assign n10925 = n10922 | n10924 ;
  assign n10926 = n157 & n10925 ;
  assign n10927 = n10361 & n69071 ;
  assign n10928 = n10710 & n10927 ;
  assign n10929 = n10926 | n10928 ;
  assign n10930 = n66868 & n10929 ;
  assign n69108 = ~n10765 ;
  assign n10931 = n10619 & n69108 ;
  assign n10932 = n10378 | n10619 ;
  assign n69109 = ~n10932 ;
  assign n10933 = n10615 & n69109 ;
  assign n10934 = n10931 | n10933 ;
  assign n10935 = n157 & n10934 ;
  assign n10936 = n10369 & n69071 ;
  assign n10937 = n10710 & n10936 ;
  assign n10938 = n10935 | n10937 ;
  assign n10939 = n66797 & n10938 ;
  assign n69110 = ~n10614 ;
  assign n10940 = n10613 & n69110 ;
  assign n10941 = n10386 | n10613 ;
  assign n69111 = ~n10941 ;
  assign n10942 = n10762 & n69111 ;
  assign n10943 = n10940 | n10942 ;
  assign n10944 = n157 & n10943 ;
  assign n10945 = n10377 & n69071 ;
  assign n10946 = n10710 & n10945 ;
  assign n10947 = n10944 | n10946 ;
  assign n10948 = n66654 & n10947 ;
  assign n69112 = ~n10761 ;
  assign n10949 = n10609 & n69112 ;
  assign n10950 = n10394 | n10609 ;
  assign n69113 = ~n10950 ;
  assign n10951 = n10605 & n69113 ;
  assign n10952 = n10949 | n10951 ;
  assign n10953 = n157 & n10952 ;
  assign n10954 = n10385 & n69071 ;
  assign n10955 = n10710 & n10954 ;
  assign n10956 = n10953 | n10955 ;
  assign n10957 = n66560 & n10956 ;
  assign n69114 = ~n10604 ;
  assign n10958 = n10603 & n69114 ;
  assign n10959 = n10402 | n10603 ;
  assign n69115 = ~n10959 ;
  assign n10960 = n10758 & n69115 ;
  assign n10961 = n10958 | n10960 ;
  assign n10962 = n157 & n10961 ;
  assign n10963 = n10393 & n69071 ;
  assign n10964 = n10710 & n10963 ;
  assign n10965 = n10962 | n10964 ;
  assign n10966 = n66505 & n10965 ;
  assign n69116 = ~n10757 ;
  assign n10967 = n10599 & n69116 ;
  assign n10968 = n10410 | n10599 ;
  assign n69117 = ~n10968 ;
  assign n10969 = n10595 & n69117 ;
  assign n10970 = n10967 | n10969 ;
  assign n10971 = n157 & n10970 ;
  assign n10972 = n10401 & n69071 ;
  assign n10973 = n10710 & n10972 ;
  assign n10974 = n10971 | n10973 ;
  assign n10975 = n66379 & n10974 ;
  assign n69118 = ~n10594 ;
  assign n10976 = n10593 & n69118 ;
  assign n10977 = n10418 | n10593 ;
  assign n69119 = ~n10977 ;
  assign n10978 = n10754 & n69119 ;
  assign n10979 = n10976 | n10978 ;
  assign n10980 = n157 & n10979 ;
  assign n10981 = n10409 & n69071 ;
  assign n10982 = n10710 & n10981 ;
  assign n10983 = n10980 | n10982 ;
  assign n10984 = n66299 & n10983 ;
  assign n69120 = ~n10753 ;
  assign n10985 = n10589 & n69120 ;
  assign n10986 = n10426 | n10589 ;
  assign n69121 = ~n10986 ;
  assign n10987 = n10585 & n69121 ;
  assign n10988 = n10985 | n10987 ;
  assign n10989 = n157 & n10988 ;
  assign n10990 = n10417 & n69071 ;
  assign n10991 = n10710 & n10990 ;
  assign n10992 = n10989 | n10991 ;
  assign n10993 = n66244 & n10992 ;
  assign n69122 = ~n10584 ;
  assign n10994 = n10583 & n69122 ;
  assign n10995 = n10434 | n10583 ;
  assign n69123 = ~n10995 ;
  assign n10996 = n10750 & n69123 ;
  assign n10997 = n10994 | n10996 ;
  assign n10998 = n157 & n10997 ;
  assign n10999 = n10425 & n69071 ;
  assign n11000 = n10710 & n10999 ;
  assign n11001 = n10998 | n11000 ;
  assign n11002 = n66145 & n11001 ;
  assign n69124 = ~n10749 ;
  assign n11003 = n10579 & n69124 ;
  assign n11004 = n10442 | n10579 ;
  assign n69125 = ~n11004 ;
  assign n11005 = n10575 & n69125 ;
  assign n11006 = n11003 | n11005 ;
  assign n11007 = n157 & n11006 ;
  assign n11008 = n10433 & n69071 ;
  assign n11009 = n10710 & n11008 ;
  assign n11010 = n11007 | n11009 ;
  assign n11011 = n66081 & n11010 ;
  assign n69126 = ~n10574 ;
  assign n11012 = n10573 & n69126 ;
  assign n11013 = n10450 | n10573 ;
  assign n69127 = ~n11013 ;
  assign n11014 = n10746 & n69127 ;
  assign n11015 = n11012 | n11014 ;
  assign n11016 = n157 & n11015 ;
  assign n11017 = n10441 & n69071 ;
  assign n11018 = n10710 & n11017 ;
  assign n11019 = n11016 | n11018 ;
  assign n11020 = n66043 & n11019 ;
  assign n69128 = ~n10745 ;
  assign n11021 = n10569 & n69128 ;
  assign n11022 = n10458 | n10569 ;
  assign n69129 = ~n11022 ;
  assign n11023 = n10565 & n69129 ;
  assign n11024 = n11021 | n11023 ;
  assign n11025 = n157 & n11024 ;
  assign n11026 = n10449 & n69071 ;
  assign n11027 = n10710 & n11026 ;
  assign n11028 = n11025 | n11027 ;
  assign n11029 = n65960 & n11028 ;
  assign n69130 = ~n10564 ;
  assign n11030 = n10563 & n69130 ;
  assign n11031 = n10466 | n10563 ;
  assign n69131 = ~n11031 ;
  assign n11032 = n10742 & n69131 ;
  assign n11033 = n11030 | n11032 ;
  assign n11034 = n157 & n11033 ;
  assign n11035 = n10457 & n69071 ;
  assign n11036 = n10710 & n11035 ;
  assign n11037 = n11034 | n11036 ;
  assign n11038 = n65909 & n11037 ;
  assign n69132 = ~n10741 ;
  assign n11039 = n10559 & n69132 ;
  assign n11040 = n10474 | n10559 ;
  assign n69133 = ~n11040 ;
  assign n11041 = n10555 & n69133 ;
  assign n11042 = n11039 | n11041 ;
  assign n11043 = n157 & n11042 ;
  assign n11044 = n10465 & n69071 ;
  assign n11045 = n10710 & n11044 ;
  assign n11046 = n11043 | n11045 ;
  assign n11047 = n65877 & n11046 ;
  assign n69134 = ~n10554 ;
  assign n11048 = n10553 & n69134 ;
  assign n11049 = n10483 | n10553 ;
  assign n69135 = ~n11049 ;
  assign n11050 = n10738 & n69135 ;
  assign n11051 = n11048 | n11050 ;
  assign n11052 = n157 & n11051 ;
  assign n11053 = n10473 & n69071 ;
  assign n11054 = n10710 & n11053 ;
  assign n11055 = n11052 | n11054 ;
  assign n11056 = n65820 & n11055 ;
  assign n69136 = ~n10737 ;
  assign n11057 = n10549 & n69136 ;
  assign n11058 = n10491 | n10549 ;
  assign n69137 = ~n11058 ;
  assign n11059 = n10545 & n69137 ;
  assign n11060 = n11057 | n11059 ;
  assign n11061 = n157 & n11060 ;
  assign n11062 = n10482 & n69071 ;
  assign n11063 = n10710 & n11062 ;
  assign n11064 = n11061 | n11063 ;
  assign n11065 = n65791 & n11064 ;
  assign n69138 = ~n10544 ;
  assign n11066 = n10543 & n69138 ;
  assign n11067 = n10501 | n10543 ;
  assign n69139 = ~n11067 ;
  assign n11068 = n10734 & n69139 ;
  assign n11069 = n11066 | n11068 ;
  assign n11070 = n157 & n11069 ;
  assign n11071 = n10490 & n69071 ;
  assign n11072 = n10710 & n11071 ;
  assign n11073 = n11070 | n11072 ;
  assign n11074 = n65772 & n11073 ;
  assign n69140 = ~n10733 ;
  assign n11076 = n10539 & n69140 ;
  assign n11075 = n10509 | n10539 ;
  assign n69141 = ~n11075 ;
  assign n11077 = n10732 & n69141 ;
  assign n11078 = n11076 | n11077 ;
  assign n11079 = n157 & n11078 ;
  assign n11080 = n10499 & n69071 ;
  assign n11081 = n10710 & n11080 ;
  assign n11082 = n11079 | n11081 ;
  assign n11083 = n65746 & n11082 ;
  assign n69142 = ~n10535 ;
  assign n11085 = n10534 & n69142 ;
  assign n11084 = n10531 | n10534 ;
  assign n69143 = ~n11084 ;
  assign n11086 = n10530 & n69143 ;
  assign n11087 = n11085 | n11086 ;
  assign n11088 = n157 & n11087 ;
  assign n11089 = n10508 & n69071 ;
  assign n11090 = n10710 & n11089 ;
  assign n11091 = n11088 | n11090 ;
  assign n11092 = n65721 & n11091 ;
  assign n11093 = n10527 & n10529 ;
  assign n11094 = n68996 & n11093 ;
  assign n69144 = ~n11094 ;
  assign n11095 = n10530 & n69144 ;
  assign n11096 = n157 & n11095 ;
  assign n11097 = n10524 & n69071 ;
  assign n11098 = n10710 & n11097 ;
  assign n11099 = n11096 | n11098 ;
  assign n11100 = n65686 & n11099 ;
  assign n10713 = n10529 & n157 ;
  assign n11101 = x64 & n157 ;
  assign n69145 = ~n11101 ;
  assign n11102 = x28 & n69145 ;
  assign n11103 = n10713 | n11102 ;
  assign n11116 = n65670 & n11103 ;
  assign n10795 = n69062 & n10794 ;
  assign n11104 = n10693 | n10795 ;
  assign n11105 = n69063 & n11104 ;
  assign n11106 = n10709 | n11105 ;
  assign n11107 = n69071 & n11106 ;
  assign n69146 = ~n11107 ;
  assign n11108 = x64 & n69146 ;
  assign n69147 = ~n11108 ;
  assign n11109 = x28 & n69147 ;
  assign n11110 = n10713 | n11109 ;
  assign n11111 = x65 & n11110 ;
  assign n11112 = x65 | n10713 ;
  assign n11113 = n11109 | n11112 ;
  assign n69148 = ~n11111 ;
  assign n11114 = n69148 & n11113 ;
  assign n69149 = ~x27 ;
  assign n11115 = n69149 & x64 ;
  assign n11117 = n11114 | n11115 ;
  assign n69150 = ~n11116 ;
  assign n11118 = n69150 & n11117 ;
  assign n69151 = ~n11098 ;
  assign n11119 = x66 & n69151 ;
  assign n69152 = ~n11096 ;
  assign n11120 = n69152 & n11119 ;
  assign n11121 = n11100 | n11120 ;
  assign n11122 = n11118 | n11121 ;
  assign n69153 = ~n11100 ;
  assign n11123 = n69153 & n11122 ;
  assign n69154 = ~n11090 ;
  assign n11124 = x67 & n69154 ;
  assign n69155 = ~n11088 ;
  assign n11125 = n69155 & n11124 ;
  assign n11126 = n11092 | n11125 ;
  assign n11127 = n11123 | n11126 ;
  assign n69156 = ~n11092 ;
  assign n11128 = n69156 & n11127 ;
  assign n69157 = ~n11081 ;
  assign n11129 = x68 & n69157 ;
  assign n69158 = ~n11079 ;
  assign n11130 = n69158 & n11129 ;
  assign n11131 = n11083 | n11130 ;
  assign n11132 = n11128 | n11131 ;
  assign n69159 = ~n11083 ;
  assign n11133 = n69159 & n11132 ;
  assign n69160 = ~n11072 ;
  assign n11134 = x69 & n69160 ;
  assign n69161 = ~n11070 ;
  assign n11135 = n69161 & n11134 ;
  assign n11136 = n11074 | n11135 ;
  assign n11137 = n11133 | n11136 ;
  assign n69162 = ~n11074 ;
  assign n11138 = n69162 & n11137 ;
  assign n69163 = ~n11063 ;
  assign n11139 = x70 & n69163 ;
  assign n69164 = ~n11061 ;
  assign n11140 = n69164 & n11139 ;
  assign n11141 = n11065 | n11140 ;
  assign n11143 = n11138 | n11141 ;
  assign n69165 = ~n11065 ;
  assign n11144 = n69165 & n11143 ;
  assign n69166 = ~n11054 ;
  assign n11145 = x71 & n69166 ;
  assign n69167 = ~n11052 ;
  assign n11146 = n69167 & n11145 ;
  assign n11147 = n11056 | n11146 ;
  assign n11148 = n11144 | n11147 ;
  assign n69168 = ~n11056 ;
  assign n11149 = n69168 & n11148 ;
  assign n69169 = ~n11045 ;
  assign n11150 = x72 & n69169 ;
  assign n69170 = ~n11043 ;
  assign n11151 = n69170 & n11150 ;
  assign n11152 = n11047 | n11151 ;
  assign n11154 = n11149 | n11152 ;
  assign n69171 = ~n11047 ;
  assign n11155 = n69171 & n11154 ;
  assign n69172 = ~n11036 ;
  assign n11156 = x73 & n69172 ;
  assign n69173 = ~n11034 ;
  assign n11157 = n69173 & n11156 ;
  assign n11158 = n11038 | n11157 ;
  assign n11159 = n11155 | n11158 ;
  assign n69174 = ~n11038 ;
  assign n11160 = n69174 & n11159 ;
  assign n69175 = ~n11027 ;
  assign n11161 = x74 & n69175 ;
  assign n69176 = ~n11025 ;
  assign n11162 = n69176 & n11161 ;
  assign n11163 = n11029 | n11162 ;
  assign n11165 = n11160 | n11163 ;
  assign n69177 = ~n11029 ;
  assign n11166 = n69177 & n11165 ;
  assign n69178 = ~n11018 ;
  assign n11167 = x75 & n69178 ;
  assign n69179 = ~n11016 ;
  assign n11168 = n69179 & n11167 ;
  assign n11169 = n11020 | n11168 ;
  assign n11170 = n11166 | n11169 ;
  assign n69180 = ~n11020 ;
  assign n11171 = n69180 & n11170 ;
  assign n69181 = ~n11009 ;
  assign n11172 = x76 & n69181 ;
  assign n69182 = ~n11007 ;
  assign n11173 = n69182 & n11172 ;
  assign n11174 = n11011 | n11173 ;
  assign n11176 = n11171 | n11174 ;
  assign n69183 = ~n11011 ;
  assign n11177 = n69183 & n11176 ;
  assign n69184 = ~n11000 ;
  assign n11178 = x77 & n69184 ;
  assign n69185 = ~n10998 ;
  assign n11179 = n69185 & n11178 ;
  assign n11180 = n11002 | n11179 ;
  assign n11181 = n11177 | n11180 ;
  assign n69186 = ~n11002 ;
  assign n11182 = n69186 & n11181 ;
  assign n69187 = ~n10991 ;
  assign n11183 = x78 & n69187 ;
  assign n69188 = ~n10989 ;
  assign n11184 = n69188 & n11183 ;
  assign n11185 = n10993 | n11184 ;
  assign n11187 = n11182 | n11185 ;
  assign n69189 = ~n10993 ;
  assign n11188 = n69189 & n11187 ;
  assign n69190 = ~n10982 ;
  assign n11189 = x79 & n69190 ;
  assign n69191 = ~n10980 ;
  assign n11190 = n69191 & n11189 ;
  assign n11191 = n10984 | n11190 ;
  assign n11192 = n11188 | n11191 ;
  assign n69192 = ~n10984 ;
  assign n11193 = n69192 & n11192 ;
  assign n69193 = ~n10973 ;
  assign n11194 = x80 & n69193 ;
  assign n69194 = ~n10971 ;
  assign n11195 = n69194 & n11194 ;
  assign n11196 = n10975 | n11195 ;
  assign n11198 = n11193 | n11196 ;
  assign n69195 = ~n10975 ;
  assign n11199 = n69195 & n11198 ;
  assign n69196 = ~n10964 ;
  assign n11200 = x81 & n69196 ;
  assign n69197 = ~n10962 ;
  assign n11201 = n69197 & n11200 ;
  assign n11202 = n10966 | n11201 ;
  assign n11203 = n11199 | n11202 ;
  assign n69198 = ~n10966 ;
  assign n11204 = n69198 & n11203 ;
  assign n69199 = ~n10955 ;
  assign n11205 = x82 & n69199 ;
  assign n69200 = ~n10953 ;
  assign n11206 = n69200 & n11205 ;
  assign n11207 = n10957 | n11206 ;
  assign n11209 = n11204 | n11207 ;
  assign n69201 = ~n10957 ;
  assign n11210 = n69201 & n11209 ;
  assign n69202 = ~n10946 ;
  assign n11211 = x83 & n69202 ;
  assign n69203 = ~n10944 ;
  assign n11212 = n69203 & n11211 ;
  assign n11213 = n10948 | n11212 ;
  assign n11214 = n11210 | n11213 ;
  assign n69204 = ~n10948 ;
  assign n11215 = n69204 & n11214 ;
  assign n69205 = ~n10937 ;
  assign n11216 = x84 & n69205 ;
  assign n69206 = ~n10935 ;
  assign n11217 = n69206 & n11216 ;
  assign n11218 = n10939 | n11217 ;
  assign n11220 = n11215 | n11218 ;
  assign n69207 = ~n10939 ;
  assign n11221 = n69207 & n11220 ;
  assign n69208 = ~n10928 ;
  assign n11222 = x85 & n69208 ;
  assign n69209 = ~n10926 ;
  assign n11223 = n69209 & n11222 ;
  assign n11224 = n10930 | n11223 ;
  assign n11225 = n11221 | n11224 ;
  assign n69210 = ~n10930 ;
  assign n11226 = n69210 & n11225 ;
  assign n69211 = ~n10919 ;
  assign n11227 = x86 & n69211 ;
  assign n69212 = ~n10917 ;
  assign n11228 = n69212 & n11227 ;
  assign n11229 = n10921 | n11228 ;
  assign n11231 = n11226 | n11229 ;
  assign n69213 = ~n10921 ;
  assign n11232 = n69213 & n11231 ;
  assign n69214 = ~n10910 ;
  assign n11233 = x87 & n69214 ;
  assign n69215 = ~n10908 ;
  assign n11234 = n69215 & n11233 ;
  assign n11235 = n10912 | n11234 ;
  assign n11236 = n11232 | n11235 ;
  assign n69216 = ~n10912 ;
  assign n11237 = n69216 & n11236 ;
  assign n69217 = ~n10901 ;
  assign n11238 = x88 & n69217 ;
  assign n69218 = ~n10899 ;
  assign n11239 = n69218 & n11238 ;
  assign n11240 = n10903 | n11239 ;
  assign n11242 = n11237 | n11240 ;
  assign n69219 = ~n10903 ;
  assign n11243 = n69219 & n11242 ;
  assign n69220 = ~n10892 ;
  assign n11244 = x89 & n69220 ;
  assign n69221 = ~n10890 ;
  assign n11245 = n69221 & n11244 ;
  assign n11246 = n10894 | n11245 ;
  assign n11247 = n11243 | n11246 ;
  assign n69222 = ~n10894 ;
  assign n11248 = n69222 & n11247 ;
  assign n69223 = ~n10883 ;
  assign n11249 = x90 & n69223 ;
  assign n69224 = ~n10881 ;
  assign n11250 = n69224 & n11249 ;
  assign n11251 = n10885 | n11250 ;
  assign n11253 = n11248 | n11251 ;
  assign n69225 = ~n10885 ;
  assign n11254 = n69225 & n11253 ;
  assign n69226 = ~n10874 ;
  assign n11255 = x91 & n69226 ;
  assign n69227 = ~n10872 ;
  assign n11256 = n69227 & n11255 ;
  assign n11257 = n10876 | n11256 ;
  assign n11258 = n11254 | n11257 ;
  assign n69228 = ~n10876 ;
  assign n11259 = n69228 & n11258 ;
  assign n69229 = ~n10865 ;
  assign n11260 = x92 & n69229 ;
  assign n69230 = ~n10863 ;
  assign n11261 = n69230 & n11260 ;
  assign n11262 = n10867 | n11261 ;
  assign n11264 = n11259 | n11262 ;
  assign n69231 = ~n10867 ;
  assign n11265 = n69231 & n11264 ;
  assign n69232 = ~n10856 ;
  assign n11266 = x93 & n69232 ;
  assign n69233 = ~n10854 ;
  assign n11267 = n69233 & n11266 ;
  assign n11268 = n10858 | n11267 ;
  assign n11269 = n11265 | n11268 ;
  assign n69234 = ~n10858 ;
  assign n11270 = n69234 & n11269 ;
  assign n69235 = ~n10847 ;
  assign n11271 = x94 & n69235 ;
  assign n69236 = ~n10845 ;
  assign n11272 = n69236 & n11271 ;
  assign n11273 = n10849 | n11272 ;
  assign n11275 = n11270 | n11273 ;
  assign n69237 = ~n10849 ;
  assign n11276 = n69237 & n11275 ;
  assign n69238 = ~n10838 ;
  assign n11277 = x95 & n69238 ;
  assign n69239 = ~n10836 ;
  assign n11278 = n69239 & n11277 ;
  assign n11279 = n10840 | n11278 ;
  assign n11280 = n11276 | n11279 ;
  assign n69240 = ~n10840 ;
  assign n11281 = n69240 & n11280 ;
  assign n69241 = ~n10829 ;
  assign n11282 = x96 & n69241 ;
  assign n69242 = ~n10827 ;
  assign n11283 = n69242 & n11282 ;
  assign n11284 = n10831 | n11283 ;
  assign n11286 = n11281 | n11284 ;
  assign n69243 = ~n10831 ;
  assign n11287 = n69243 & n11286 ;
  assign n69244 = ~n10820 ;
  assign n11288 = x97 & n69244 ;
  assign n69245 = ~n10818 ;
  assign n11289 = n69245 & n11288 ;
  assign n11290 = n10822 | n11289 ;
  assign n11291 = n11287 | n11290 ;
  assign n69246 = ~n10822 ;
  assign n11292 = n69246 & n11291 ;
  assign n69247 = ~n10811 ;
  assign n11293 = x98 & n69247 ;
  assign n69248 = ~n10809 ;
  assign n11294 = n69248 & n11293 ;
  assign n11295 = n10813 | n11294 ;
  assign n11297 = n11292 | n11295 ;
  assign n69249 = ~n10813 ;
  assign n11298 = n69249 & n11297 ;
  assign n69250 = ~n10802 ;
  assign n11299 = x99 & n69250 ;
  assign n69251 = ~n10800 ;
  assign n11300 = n69251 & n11299 ;
  assign n11301 = n10804 | n11300 ;
  assign n11302 = n11298 | n11301 ;
  assign n69252 = ~n10804 ;
  assign n11303 = n69252 & n11302 ;
  assign n69253 = ~n10722 ;
  assign n11304 = x100 & n69253 ;
  assign n69254 = ~n10720 ;
  assign n11305 = n69254 & n11304 ;
  assign n11306 = n10724 | n11305 ;
  assign n11308 = n11303 | n11306 ;
  assign n69255 = ~n10724 ;
  assign n11309 = n69255 & n11308 ;
  assign n11310 = n469 | n11309 ;
  assign n69256 = ~n11303 ;
  assign n11307 = n69256 & n11306 ;
  assign n11311 = x65 & n11103 ;
  assign n69257 = ~n11311 ;
  assign n11312 = n11113 & n69257 ;
  assign n11313 = n11115 | n11312 ;
  assign n11314 = n69150 & n11313 ;
  assign n11315 = n11121 | n11314 ;
  assign n11316 = n69153 & n11315 ;
  assign n11318 = n11126 | n11316 ;
  assign n11319 = n69156 & n11318 ;
  assign n11321 = n11131 | n11319 ;
  assign n11322 = n69159 & n11321 ;
  assign n11323 = n11136 | n11322 ;
  assign n11325 = n69162 & n11323 ;
  assign n11326 = n11141 | n11325 ;
  assign n11327 = n69165 & n11326 ;
  assign n11328 = n11147 | n11327 ;
  assign n11330 = n69168 & n11328 ;
  assign n11331 = n11152 | n11330 ;
  assign n11332 = n69171 & n11331 ;
  assign n11333 = n11158 | n11332 ;
  assign n11335 = n69174 & n11333 ;
  assign n11336 = n11163 | n11335 ;
  assign n11337 = n69177 & n11336 ;
  assign n11338 = n11169 | n11337 ;
  assign n11340 = n69180 & n11338 ;
  assign n11341 = n11174 | n11340 ;
  assign n11342 = n69183 & n11341 ;
  assign n11343 = n11180 | n11342 ;
  assign n11345 = n69186 & n11343 ;
  assign n11346 = n11185 | n11345 ;
  assign n11347 = n69189 & n11346 ;
  assign n11348 = n11191 | n11347 ;
  assign n11350 = n69192 & n11348 ;
  assign n11351 = n11196 | n11350 ;
  assign n11352 = n69195 & n11351 ;
  assign n11353 = n11202 | n11352 ;
  assign n11355 = n69198 & n11353 ;
  assign n11356 = n11207 | n11355 ;
  assign n11357 = n69201 & n11356 ;
  assign n11358 = n11213 | n11357 ;
  assign n11360 = n69204 & n11358 ;
  assign n11361 = n11218 | n11360 ;
  assign n11362 = n69207 & n11361 ;
  assign n11363 = n11224 | n11362 ;
  assign n11365 = n69210 & n11363 ;
  assign n11366 = n11229 | n11365 ;
  assign n11367 = n69213 & n11366 ;
  assign n11368 = n11235 | n11367 ;
  assign n11370 = n69216 & n11368 ;
  assign n11371 = n11240 | n11370 ;
  assign n11372 = n69219 & n11371 ;
  assign n11373 = n11246 | n11372 ;
  assign n11375 = n69222 & n11373 ;
  assign n11376 = n11251 | n11375 ;
  assign n11377 = n69225 & n11376 ;
  assign n11378 = n11257 | n11377 ;
  assign n11380 = n69228 & n11378 ;
  assign n11381 = n11262 | n11380 ;
  assign n11382 = n69231 & n11381 ;
  assign n11383 = n11268 | n11382 ;
  assign n11385 = n69234 & n11383 ;
  assign n11386 = n11273 | n11385 ;
  assign n11387 = n69237 & n11386 ;
  assign n11388 = n11279 | n11387 ;
  assign n11390 = n69240 & n11388 ;
  assign n11391 = n11284 | n11390 ;
  assign n11392 = n69243 & n11391 ;
  assign n11393 = n11290 | n11392 ;
  assign n11395 = n69246 & n11393 ;
  assign n11396 = n11295 | n11395 ;
  assign n11397 = n69249 & n11396 ;
  assign n11399 = n11301 | n11397 ;
  assign n11400 = n10804 | n11306 ;
  assign n69258 = ~n11400 ;
  assign n11401 = n11399 & n69258 ;
  assign n11402 = n11307 | n11401 ;
  assign n11403 = n11310 | n11402 ;
  assign n69259 = ~n10723 ;
  assign n11404 = n69259 & n11310 ;
  assign n69260 = ~n11404 ;
  assign n11405 = n11403 & n69260 ;
  assign n69261 = ~x101 ;
  assign n11406 = n69261 & n11405 ;
  assign n156 = ~n11310 ;
  assign n11919 = n156 & n11402 ;
  assign n11920 = n10723 & n11310 ;
  assign n69263 = ~n11920 ;
  assign n11921 = x101 & n69263 ;
  assign n69264 = ~n11919 ;
  assign n11922 = n69264 & n11921 ;
  assign n11923 = n11406 | n11922 ;
  assign n11407 = n10803 & n11310 ;
  assign n69265 = ~n11397 ;
  assign n11398 = n11301 & n69265 ;
  assign n11408 = n10813 | n11301 ;
  assign n69266 = ~n11408 ;
  assign n11409 = n11297 & n69266 ;
  assign n11410 = n11398 | n11409 ;
  assign n11411 = n65845 & n11410 ;
  assign n69267 = ~n11309 ;
  assign n11412 = n69267 & n11411 ;
  assign n11413 = n11407 | n11412 ;
  assign n11414 = n69075 & n11413 ;
  assign n11415 = n10812 & n11310 ;
  assign n69268 = ~n11292 ;
  assign n11296 = n69268 & n11295 ;
  assign n11416 = n10822 | n11295 ;
  assign n69269 = ~n11416 ;
  assign n11417 = n11393 & n69269 ;
  assign n11418 = n11296 | n11417 ;
  assign n11419 = n65845 & n11418 ;
  assign n11420 = n69267 & n11419 ;
  assign n11421 = n11415 | n11420 ;
  assign n11422 = n68993 & n11421 ;
  assign n69270 = ~n11420 ;
  assign n11907 = x99 & n69270 ;
  assign n69271 = ~n11415 ;
  assign n11908 = n69271 & n11907 ;
  assign n11909 = n11422 | n11908 ;
  assign n11423 = n10821 & n11310 ;
  assign n69272 = ~n11392 ;
  assign n11394 = n11290 & n69272 ;
  assign n11424 = n10831 | n11290 ;
  assign n69273 = ~n11424 ;
  assign n11425 = n11286 & n69273 ;
  assign n11426 = n11394 | n11425 ;
  assign n11427 = n65845 & n11426 ;
  assign n11428 = n69267 & n11427 ;
  assign n11429 = n11423 | n11428 ;
  assign n11430 = n68716 & n11429 ;
  assign n11431 = n10830 & n11310 ;
  assign n69274 = ~n11281 ;
  assign n11285 = n69274 & n11284 ;
  assign n11432 = n10840 | n11284 ;
  assign n69275 = ~n11432 ;
  assign n11433 = n11388 & n69275 ;
  assign n11434 = n11285 | n11433 ;
  assign n11435 = n65845 & n11434 ;
  assign n11436 = n69267 & n11435 ;
  assign n11437 = n11431 | n11436 ;
  assign n11438 = n68545 & n11437 ;
  assign n69276 = ~n11436 ;
  assign n11895 = x97 & n69276 ;
  assign n69277 = ~n11431 ;
  assign n11896 = n69277 & n11895 ;
  assign n11897 = n11438 | n11896 ;
  assign n11439 = n10839 & n11310 ;
  assign n69278 = ~n11387 ;
  assign n11389 = n11279 & n69278 ;
  assign n11440 = n10849 | n11279 ;
  assign n69279 = ~n11440 ;
  assign n11441 = n11275 & n69279 ;
  assign n11442 = n11389 | n11441 ;
  assign n11443 = n65845 & n11442 ;
  assign n11444 = n69267 & n11443 ;
  assign n11445 = n11439 | n11444 ;
  assign n11446 = n68438 & n11445 ;
  assign n11447 = n10848 & n11310 ;
  assign n69280 = ~n11270 ;
  assign n11274 = n69280 & n11273 ;
  assign n11448 = n10858 | n11273 ;
  assign n69281 = ~n11448 ;
  assign n11449 = n11383 & n69281 ;
  assign n11450 = n11274 | n11449 ;
  assign n11451 = n65845 & n11450 ;
  assign n11452 = n69267 & n11451 ;
  assign n11453 = n11447 | n11452 ;
  assign n11454 = n68214 & n11453 ;
  assign n69282 = ~n11452 ;
  assign n11883 = x95 & n69282 ;
  assign n69283 = ~n11447 ;
  assign n11884 = n69283 & n11883 ;
  assign n11885 = n11454 | n11884 ;
  assign n11455 = n10857 & n11310 ;
  assign n69284 = ~n11382 ;
  assign n11384 = n11268 & n69284 ;
  assign n11456 = n10867 | n11268 ;
  assign n69285 = ~n11456 ;
  assign n11457 = n11264 & n69285 ;
  assign n11458 = n11384 | n11457 ;
  assign n11459 = n65845 & n11458 ;
  assign n11460 = n69267 & n11459 ;
  assign n11461 = n11455 | n11460 ;
  assign n11462 = n68058 & n11461 ;
  assign n11463 = n10866 & n11310 ;
  assign n69286 = ~n11259 ;
  assign n11263 = n69286 & n11262 ;
  assign n11464 = n10876 | n11262 ;
  assign n69287 = ~n11464 ;
  assign n11465 = n11378 & n69287 ;
  assign n11466 = n11263 | n11465 ;
  assign n11467 = n65845 & n11466 ;
  assign n11468 = n69267 & n11467 ;
  assign n11469 = n11463 | n11468 ;
  assign n11470 = n67986 & n11469 ;
  assign n69288 = ~n11468 ;
  assign n11871 = x93 & n69288 ;
  assign n69289 = ~n11463 ;
  assign n11872 = n69289 & n11871 ;
  assign n11873 = n11470 | n11872 ;
  assign n11471 = n10875 & n11310 ;
  assign n69290 = ~n11377 ;
  assign n11379 = n11257 & n69290 ;
  assign n11472 = n10885 | n11257 ;
  assign n69291 = ~n11472 ;
  assign n11473 = n11253 & n69291 ;
  assign n11474 = n11379 | n11473 ;
  assign n11475 = n65845 & n11474 ;
  assign n11476 = n69267 & n11475 ;
  assign n11477 = n11471 | n11476 ;
  assign n11478 = n67763 & n11477 ;
  assign n11479 = n10884 & n11310 ;
  assign n69292 = ~n11248 ;
  assign n11252 = n69292 & n11251 ;
  assign n11480 = n10894 | n11251 ;
  assign n69293 = ~n11480 ;
  assign n11481 = n11373 & n69293 ;
  assign n11482 = n11252 | n11481 ;
  assign n11483 = n65845 & n11482 ;
  assign n11484 = n69267 & n11483 ;
  assign n11485 = n11479 | n11484 ;
  assign n11486 = n67622 & n11485 ;
  assign n69294 = ~n11484 ;
  assign n11859 = x91 & n69294 ;
  assign n69295 = ~n11479 ;
  assign n11860 = n69295 & n11859 ;
  assign n11861 = n11486 | n11860 ;
  assign n11487 = n10893 & n11310 ;
  assign n69296 = ~n11372 ;
  assign n11374 = n11246 & n69296 ;
  assign n11488 = n10903 | n11246 ;
  assign n69297 = ~n11488 ;
  assign n11489 = n11242 & n69297 ;
  assign n11490 = n11374 | n11489 ;
  assign n11491 = n65845 & n11490 ;
  assign n11492 = n69267 & n11491 ;
  assign n11493 = n11487 | n11492 ;
  assign n11494 = n67531 & n11493 ;
  assign n11495 = n10902 & n11310 ;
  assign n69298 = ~n11237 ;
  assign n11241 = n69298 & n11240 ;
  assign n11496 = n10912 | n11240 ;
  assign n69299 = ~n11496 ;
  assign n11497 = n11368 & n69299 ;
  assign n11498 = n11241 | n11497 ;
  assign n11499 = n65845 & n11498 ;
  assign n11500 = n69267 & n11499 ;
  assign n11501 = n11495 | n11500 ;
  assign n11502 = n67348 & n11501 ;
  assign n69300 = ~n11500 ;
  assign n11847 = x89 & n69300 ;
  assign n69301 = ~n11495 ;
  assign n11848 = n69301 & n11847 ;
  assign n11849 = n11502 | n11848 ;
  assign n11503 = n10911 & n11310 ;
  assign n69302 = ~n11367 ;
  assign n11369 = n11235 & n69302 ;
  assign n11504 = n10921 | n11235 ;
  assign n69303 = ~n11504 ;
  assign n11505 = n11231 & n69303 ;
  assign n11506 = n11369 | n11505 ;
  assign n11507 = n65845 & n11506 ;
  assign n11508 = n69267 & n11507 ;
  assign n11509 = n11503 | n11508 ;
  assign n11510 = n67222 & n11509 ;
  assign n11511 = n10920 & n11310 ;
  assign n69304 = ~n11226 ;
  assign n11230 = n69304 & n11229 ;
  assign n11512 = n10930 | n11229 ;
  assign n69305 = ~n11512 ;
  assign n11513 = n11363 & n69305 ;
  assign n11514 = n11230 | n11513 ;
  assign n11515 = n65845 & n11514 ;
  assign n11516 = n69267 & n11515 ;
  assign n11517 = n11511 | n11516 ;
  assign n11518 = n67164 & n11517 ;
  assign n69306 = ~n11516 ;
  assign n11835 = x87 & n69306 ;
  assign n69307 = ~n11511 ;
  assign n11836 = n69307 & n11835 ;
  assign n11837 = n11518 | n11836 ;
  assign n11519 = n10929 & n11310 ;
  assign n69308 = ~n11362 ;
  assign n11364 = n11224 & n69308 ;
  assign n11520 = n10939 | n11224 ;
  assign n69309 = ~n11520 ;
  assign n11521 = n11220 & n69309 ;
  assign n11522 = n11364 | n11521 ;
  assign n11523 = n65845 & n11522 ;
  assign n11524 = n69267 & n11523 ;
  assign n11525 = n11519 | n11524 ;
  assign n11526 = n66979 & n11525 ;
  assign n11527 = n10938 & n11310 ;
  assign n69310 = ~n11215 ;
  assign n11219 = n69310 & n11218 ;
  assign n11528 = n10948 | n11218 ;
  assign n69311 = ~n11528 ;
  assign n11529 = n11358 & n69311 ;
  assign n11530 = n11219 | n11529 ;
  assign n11531 = n65845 & n11530 ;
  assign n11532 = n69267 & n11531 ;
  assign n11533 = n11527 | n11532 ;
  assign n11534 = n66868 & n11533 ;
  assign n69312 = ~n11532 ;
  assign n11823 = x85 & n69312 ;
  assign n69313 = ~n11527 ;
  assign n11824 = n69313 & n11823 ;
  assign n11825 = n11534 | n11824 ;
  assign n11535 = n10947 & n11310 ;
  assign n69314 = ~n11357 ;
  assign n11359 = n11213 & n69314 ;
  assign n11536 = n10957 | n11213 ;
  assign n69315 = ~n11536 ;
  assign n11537 = n11209 & n69315 ;
  assign n11538 = n11359 | n11537 ;
  assign n11539 = n65845 & n11538 ;
  assign n11540 = n69267 & n11539 ;
  assign n11541 = n11535 | n11540 ;
  assign n11542 = n66797 & n11541 ;
  assign n11543 = n10956 & n11310 ;
  assign n69316 = ~n11204 ;
  assign n11208 = n69316 & n11207 ;
  assign n11544 = n10966 | n11207 ;
  assign n69317 = ~n11544 ;
  assign n11545 = n11353 & n69317 ;
  assign n11546 = n11208 | n11545 ;
  assign n11547 = n65845 & n11546 ;
  assign n11548 = n69267 & n11547 ;
  assign n11549 = n11543 | n11548 ;
  assign n11550 = n66654 & n11549 ;
  assign n69318 = ~n11548 ;
  assign n11811 = x83 & n69318 ;
  assign n69319 = ~n11543 ;
  assign n11812 = n69319 & n11811 ;
  assign n11813 = n11550 | n11812 ;
  assign n11551 = n10965 & n11310 ;
  assign n69320 = ~n11352 ;
  assign n11354 = n11202 & n69320 ;
  assign n11552 = n10975 | n11202 ;
  assign n69321 = ~n11552 ;
  assign n11553 = n11198 & n69321 ;
  assign n11554 = n11354 | n11553 ;
  assign n11555 = n65845 & n11554 ;
  assign n11556 = n69267 & n11555 ;
  assign n11557 = n11551 | n11556 ;
  assign n11558 = n66560 & n11557 ;
  assign n11559 = n10974 & n11310 ;
  assign n69322 = ~n11193 ;
  assign n11197 = n69322 & n11196 ;
  assign n11560 = n10984 | n11196 ;
  assign n69323 = ~n11560 ;
  assign n11561 = n11348 & n69323 ;
  assign n11562 = n11197 | n11561 ;
  assign n11563 = n65845 & n11562 ;
  assign n11564 = n69267 & n11563 ;
  assign n11565 = n11559 | n11564 ;
  assign n11566 = n66505 & n11565 ;
  assign n69324 = ~n11564 ;
  assign n11799 = x81 & n69324 ;
  assign n69325 = ~n11559 ;
  assign n11800 = n69325 & n11799 ;
  assign n11801 = n11566 | n11800 ;
  assign n11567 = n10983 & n11310 ;
  assign n69326 = ~n11347 ;
  assign n11349 = n11191 & n69326 ;
  assign n11568 = n10993 | n11191 ;
  assign n69327 = ~n11568 ;
  assign n11569 = n11187 & n69327 ;
  assign n11570 = n11349 | n11569 ;
  assign n11571 = n65845 & n11570 ;
  assign n11572 = n69267 & n11571 ;
  assign n11573 = n11567 | n11572 ;
  assign n11574 = n66379 & n11573 ;
  assign n11575 = n10992 & n11310 ;
  assign n69328 = ~n11182 ;
  assign n11186 = n69328 & n11185 ;
  assign n11576 = n11002 | n11185 ;
  assign n69329 = ~n11576 ;
  assign n11577 = n11343 & n69329 ;
  assign n11578 = n11186 | n11577 ;
  assign n11579 = n65845 & n11578 ;
  assign n11580 = n69267 & n11579 ;
  assign n11581 = n11575 | n11580 ;
  assign n11582 = n66299 & n11581 ;
  assign n69330 = ~n11580 ;
  assign n11787 = x79 & n69330 ;
  assign n69331 = ~n11575 ;
  assign n11788 = n69331 & n11787 ;
  assign n11789 = n11582 | n11788 ;
  assign n11583 = n11001 & n11310 ;
  assign n69332 = ~n11342 ;
  assign n11344 = n11180 & n69332 ;
  assign n11584 = n11011 | n11180 ;
  assign n69333 = ~n11584 ;
  assign n11585 = n11176 & n69333 ;
  assign n11586 = n11344 | n11585 ;
  assign n11587 = n65845 & n11586 ;
  assign n11588 = n69267 & n11587 ;
  assign n11589 = n11583 | n11588 ;
  assign n11590 = n66244 & n11589 ;
  assign n11591 = n11010 & n11310 ;
  assign n69334 = ~n11171 ;
  assign n11175 = n69334 & n11174 ;
  assign n11592 = n11020 | n11174 ;
  assign n69335 = ~n11592 ;
  assign n11593 = n11338 & n69335 ;
  assign n11594 = n11175 | n11593 ;
  assign n11595 = n65845 & n11594 ;
  assign n11596 = n69267 & n11595 ;
  assign n11597 = n11591 | n11596 ;
  assign n11598 = n66145 & n11597 ;
  assign n69336 = ~n11596 ;
  assign n11775 = x77 & n69336 ;
  assign n69337 = ~n11591 ;
  assign n11776 = n69337 & n11775 ;
  assign n11777 = n11598 | n11776 ;
  assign n11599 = n11019 & n11310 ;
  assign n69338 = ~n11337 ;
  assign n11339 = n11169 & n69338 ;
  assign n11600 = n11029 | n11169 ;
  assign n69339 = ~n11600 ;
  assign n11601 = n11165 & n69339 ;
  assign n11602 = n11339 | n11601 ;
  assign n11603 = n65845 & n11602 ;
  assign n11604 = n69267 & n11603 ;
  assign n11605 = n11599 | n11604 ;
  assign n11606 = n66081 & n11605 ;
  assign n11607 = n11028 & n11310 ;
  assign n69340 = ~n11160 ;
  assign n11164 = n69340 & n11163 ;
  assign n11608 = n11038 | n11163 ;
  assign n69341 = ~n11608 ;
  assign n11609 = n11333 & n69341 ;
  assign n11610 = n11164 | n11609 ;
  assign n11611 = n65845 & n11610 ;
  assign n11612 = n69267 & n11611 ;
  assign n11613 = n11607 | n11612 ;
  assign n11614 = n66043 & n11613 ;
  assign n69342 = ~n11612 ;
  assign n11763 = x75 & n69342 ;
  assign n69343 = ~n11607 ;
  assign n11764 = n69343 & n11763 ;
  assign n11765 = n11614 | n11764 ;
  assign n11615 = n11037 & n11310 ;
  assign n69344 = ~n11332 ;
  assign n11334 = n11158 & n69344 ;
  assign n11616 = n11047 | n11158 ;
  assign n69345 = ~n11616 ;
  assign n11617 = n11154 & n69345 ;
  assign n11618 = n11334 | n11617 ;
  assign n11619 = n65845 & n11618 ;
  assign n11620 = n69267 & n11619 ;
  assign n11621 = n11615 | n11620 ;
  assign n11622 = n65960 & n11621 ;
  assign n11623 = n11046 & n11310 ;
  assign n69346 = ~n11149 ;
  assign n11153 = n69346 & n11152 ;
  assign n11624 = n11056 | n11152 ;
  assign n69347 = ~n11624 ;
  assign n11625 = n11328 & n69347 ;
  assign n11626 = n11153 | n11625 ;
  assign n11627 = n65845 & n11626 ;
  assign n11628 = n69267 & n11627 ;
  assign n11629 = n11623 | n11628 ;
  assign n11630 = n65909 & n11629 ;
  assign n69348 = ~n11628 ;
  assign n11751 = x73 & n69348 ;
  assign n69349 = ~n11623 ;
  assign n11752 = n69349 & n11751 ;
  assign n11753 = n11630 | n11752 ;
  assign n11631 = n11055 & n11310 ;
  assign n69350 = ~n11327 ;
  assign n11329 = n11147 & n69350 ;
  assign n11632 = n11065 | n11147 ;
  assign n69351 = ~n11632 ;
  assign n11633 = n11143 & n69351 ;
  assign n11634 = n11329 | n11633 ;
  assign n11635 = n65845 & n11634 ;
  assign n11636 = n69267 & n11635 ;
  assign n11637 = n11631 | n11636 ;
  assign n11638 = n65877 & n11637 ;
  assign n11639 = n11064 & n11310 ;
  assign n69352 = ~n11138 ;
  assign n11142 = n69352 & n11141 ;
  assign n11640 = n11074 | n11141 ;
  assign n69353 = ~n11640 ;
  assign n11641 = n11323 & n69353 ;
  assign n11642 = n11142 | n11641 ;
  assign n11643 = n65845 & n11642 ;
  assign n11644 = n69267 & n11643 ;
  assign n11645 = n11639 | n11644 ;
  assign n11646 = n65820 & n11645 ;
  assign n69354 = ~n11644 ;
  assign n11739 = x71 & n69354 ;
  assign n69355 = ~n11639 ;
  assign n11740 = n69355 & n11739 ;
  assign n11741 = n11646 | n11740 ;
  assign n11647 = n11073 & n11310 ;
  assign n69356 = ~n11322 ;
  assign n11324 = n11136 & n69356 ;
  assign n11648 = n11083 | n11136 ;
  assign n69357 = ~n11648 ;
  assign n11649 = n11132 & n69357 ;
  assign n11650 = n11324 | n11649 ;
  assign n11651 = n65845 & n11650 ;
  assign n11652 = n69267 & n11651 ;
  assign n11653 = n11647 | n11652 ;
  assign n11654 = n65791 & n11653 ;
  assign n11655 = n11082 & n11310 ;
  assign n69358 = ~n11128 ;
  assign n11320 = n69358 & n11131 ;
  assign n11656 = n11092 | n11131 ;
  assign n69359 = ~n11656 ;
  assign n11657 = n11318 & n69359 ;
  assign n11658 = n11320 | n11657 ;
  assign n11659 = n65845 & n11658 ;
  assign n11660 = n69267 & n11659 ;
  assign n11661 = n11655 | n11660 ;
  assign n11662 = n65772 & n11661 ;
  assign n69360 = ~n11660 ;
  assign n11728 = x69 & n69360 ;
  assign n69361 = ~n11655 ;
  assign n11729 = n69361 & n11728 ;
  assign n11730 = n11662 | n11729 ;
  assign n11663 = n11091 & n11310 ;
  assign n69362 = ~n11316 ;
  assign n11317 = n11126 & n69362 ;
  assign n11664 = n11100 | n11126 ;
  assign n69363 = ~n11664 ;
  assign n11665 = n11315 & n69363 ;
  assign n11666 = n11317 | n11665 ;
  assign n11667 = n65845 & n11666 ;
  assign n11668 = n69267 & n11667 ;
  assign n11669 = n11663 | n11668 ;
  assign n11670 = n65746 & n11669 ;
  assign n11671 = n11099 & n11310 ;
  assign n11672 = n11116 | n11121 ;
  assign n69364 = ~n11672 ;
  assign n11673 = n11313 & n69364 ;
  assign n69365 = ~n11118 ;
  assign n11674 = n69365 & n11121 ;
  assign n11675 = n11673 | n11674 ;
  assign n11676 = n65845 & n11675 ;
  assign n11677 = n69267 & n11676 ;
  assign n11678 = n11671 | n11677 ;
  assign n11679 = n65721 & n11678 ;
  assign n69366 = ~n11677 ;
  assign n11718 = x67 & n69366 ;
  assign n69367 = ~n11671 ;
  assign n11719 = n69367 & n11718 ;
  assign n11720 = n11679 | n11719 ;
  assign n11680 = n11110 & n11310 ;
  assign n11681 = n11113 & n11115 ;
  assign n11682 = n69257 & n11681 ;
  assign n11683 = n469 | n11682 ;
  assign n69368 = ~n11683 ;
  assign n11684 = n11313 & n69368 ;
  assign n11685 = n69267 & n11684 ;
  assign n11686 = n11680 | n11685 ;
  assign n11687 = n65686 & n11686 ;
  assign n69369 = ~x26 ;
  assign n11708 = n69369 & x64 ;
  assign n11688 = x64 & n69261 ;
  assign n69370 = ~n65467 ;
  assign n11689 = n69370 & n11688 ;
  assign n69371 = ~n65452 ;
  assign n11690 = n69371 & n11689 ;
  assign n69372 = ~n65534 ;
  assign n11691 = n69372 & n11690 ;
  assign n11692 = n67021 & n11691 ;
  assign n11693 = n69267 & n11692 ;
  assign n69373 = ~n11693 ;
  assign n11694 = x27 & n69373 ;
  assign n11695 = n68782 & n11115 ;
  assign n11696 = n68783 & n11695 ;
  assign n11697 = n66715 & n11696 ;
  assign n11698 = n69267 & n11697 ;
  assign n11699 = n11694 | n11698 ;
  assign n11700 = x65 & n11699 ;
  assign n11701 = n69252 & n11399 ;
  assign n11702 = n11306 | n11701 ;
  assign n11703 = n69255 & n11702 ;
  assign n69374 = ~n11703 ;
  assign n11704 = n11692 & n69374 ;
  assign n69375 = ~n11704 ;
  assign n11705 = x27 & n69375 ;
  assign n11706 = x65 | n11698 ;
  assign n11707 = n11705 | n11706 ;
  assign n69376 = ~n11700 ;
  assign n11709 = n69376 & n11707 ;
  assign n11710 = n11708 | n11709 ;
  assign n11711 = n11698 | n11705 ;
  assign n11712 = n65670 & n11711 ;
  assign n69377 = ~n11712 ;
  assign n11713 = n11710 & n69377 ;
  assign n69378 = ~n11685 ;
  assign n11714 = x66 & n69378 ;
  assign n69379 = ~n11680 ;
  assign n11715 = n69379 & n11714 ;
  assign n11716 = n11687 | n11715 ;
  assign n11717 = n11713 | n11716 ;
  assign n69380 = ~n11687 ;
  assign n11721 = n69380 & n11717 ;
  assign n11722 = n11720 | n11721 ;
  assign n69381 = ~n11679 ;
  assign n11723 = n69381 & n11722 ;
  assign n69382 = ~n11668 ;
  assign n11724 = x68 & n69382 ;
  assign n69383 = ~n11663 ;
  assign n11725 = n69383 & n11724 ;
  assign n11726 = n11670 | n11725 ;
  assign n11727 = n11723 | n11726 ;
  assign n69384 = ~n11670 ;
  assign n11731 = n69384 & n11727 ;
  assign n11732 = n11730 | n11731 ;
  assign n69385 = ~n11662 ;
  assign n11733 = n69385 & n11732 ;
  assign n69386 = ~n11652 ;
  assign n11734 = x70 & n69386 ;
  assign n69387 = ~n11647 ;
  assign n11735 = n69387 & n11734 ;
  assign n11736 = n11654 | n11735 ;
  assign n11738 = n11733 | n11736 ;
  assign n69388 = ~n11654 ;
  assign n11743 = n69388 & n11738 ;
  assign n11744 = n11741 | n11743 ;
  assign n69389 = ~n11646 ;
  assign n11745 = n69389 & n11744 ;
  assign n69390 = ~n11636 ;
  assign n11746 = x72 & n69390 ;
  assign n69391 = ~n11631 ;
  assign n11747 = n69391 & n11746 ;
  assign n11748 = n11638 | n11747 ;
  assign n11750 = n11745 | n11748 ;
  assign n69392 = ~n11638 ;
  assign n11755 = n69392 & n11750 ;
  assign n11756 = n11753 | n11755 ;
  assign n69393 = ~n11630 ;
  assign n11757 = n69393 & n11756 ;
  assign n69394 = ~n11620 ;
  assign n11758 = x74 & n69394 ;
  assign n69395 = ~n11615 ;
  assign n11759 = n69395 & n11758 ;
  assign n11760 = n11622 | n11759 ;
  assign n11762 = n11757 | n11760 ;
  assign n69396 = ~n11622 ;
  assign n11767 = n69396 & n11762 ;
  assign n11768 = n11765 | n11767 ;
  assign n69397 = ~n11614 ;
  assign n11769 = n69397 & n11768 ;
  assign n69398 = ~n11604 ;
  assign n11770 = x76 & n69398 ;
  assign n69399 = ~n11599 ;
  assign n11771 = n69399 & n11770 ;
  assign n11772 = n11606 | n11771 ;
  assign n11774 = n11769 | n11772 ;
  assign n69400 = ~n11606 ;
  assign n11779 = n69400 & n11774 ;
  assign n11780 = n11777 | n11779 ;
  assign n69401 = ~n11598 ;
  assign n11781 = n69401 & n11780 ;
  assign n69402 = ~n11588 ;
  assign n11782 = x78 & n69402 ;
  assign n69403 = ~n11583 ;
  assign n11783 = n69403 & n11782 ;
  assign n11784 = n11590 | n11783 ;
  assign n11786 = n11781 | n11784 ;
  assign n69404 = ~n11590 ;
  assign n11791 = n69404 & n11786 ;
  assign n11792 = n11789 | n11791 ;
  assign n69405 = ~n11582 ;
  assign n11793 = n69405 & n11792 ;
  assign n69406 = ~n11572 ;
  assign n11794 = x80 & n69406 ;
  assign n69407 = ~n11567 ;
  assign n11795 = n69407 & n11794 ;
  assign n11796 = n11574 | n11795 ;
  assign n11798 = n11793 | n11796 ;
  assign n69408 = ~n11574 ;
  assign n11803 = n69408 & n11798 ;
  assign n11804 = n11801 | n11803 ;
  assign n69409 = ~n11566 ;
  assign n11805 = n69409 & n11804 ;
  assign n69410 = ~n11556 ;
  assign n11806 = x82 & n69410 ;
  assign n69411 = ~n11551 ;
  assign n11807 = n69411 & n11806 ;
  assign n11808 = n11558 | n11807 ;
  assign n11810 = n11805 | n11808 ;
  assign n69412 = ~n11558 ;
  assign n11815 = n69412 & n11810 ;
  assign n11816 = n11813 | n11815 ;
  assign n69413 = ~n11550 ;
  assign n11817 = n69413 & n11816 ;
  assign n69414 = ~n11540 ;
  assign n11818 = x84 & n69414 ;
  assign n69415 = ~n11535 ;
  assign n11819 = n69415 & n11818 ;
  assign n11820 = n11542 | n11819 ;
  assign n11822 = n11817 | n11820 ;
  assign n69416 = ~n11542 ;
  assign n11827 = n69416 & n11822 ;
  assign n11828 = n11825 | n11827 ;
  assign n69417 = ~n11534 ;
  assign n11829 = n69417 & n11828 ;
  assign n69418 = ~n11524 ;
  assign n11830 = x86 & n69418 ;
  assign n69419 = ~n11519 ;
  assign n11831 = n69419 & n11830 ;
  assign n11832 = n11526 | n11831 ;
  assign n11834 = n11829 | n11832 ;
  assign n69420 = ~n11526 ;
  assign n11839 = n69420 & n11834 ;
  assign n11840 = n11837 | n11839 ;
  assign n69421 = ~n11518 ;
  assign n11841 = n69421 & n11840 ;
  assign n69422 = ~n11508 ;
  assign n11842 = x88 & n69422 ;
  assign n69423 = ~n11503 ;
  assign n11843 = n69423 & n11842 ;
  assign n11844 = n11510 | n11843 ;
  assign n11846 = n11841 | n11844 ;
  assign n69424 = ~n11510 ;
  assign n11851 = n69424 & n11846 ;
  assign n11852 = n11849 | n11851 ;
  assign n69425 = ~n11502 ;
  assign n11853 = n69425 & n11852 ;
  assign n69426 = ~n11492 ;
  assign n11854 = x90 & n69426 ;
  assign n69427 = ~n11487 ;
  assign n11855 = n69427 & n11854 ;
  assign n11856 = n11494 | n11855 ;
  assign n11858 = n11853 | n11856 ;
  assign n69428 = ~n11494 ;
  assign n11863 = n69428 & n11858 ;
  assign n11864 = n11861 | n11863 ;
  assign n69429 = ~n11486 ;
  assign n11865 = n69429 & n11864 ;
  assign n69430 = ~n11476 ;
  assign n11866 = x92 & n69430 ;
  assign n69431 = ~n11471 ;
  assign n11867 = n69431 & n11866 ;
  assign n11868 = n11478 | n11867 ;
  assign n11870 = n11865 | n11868 ;
  assign n69432 = ~n11478 ;
  assign n11875 = n69432 & n11870 ;
  assign n11876 = n11873 | n11875 ;
  assign n69433 = ~n11470 ;
  assign n11877 = n69433 & n11876 ;
  assign n69434 = ~n11460 ;
  assign n11878 = x94 & n69434 ;
  assign n69435 = ~n11455 ;
  assign n11879 = n69435 & n11878 ;
  assign n11880 = n11462 | n11879 ;
  assign n11882 = n11877 | n11880 ;
  assign n69436 = ~n11462 ;
  assign n11887 = n69436 & n11882 ;
  assign n11888 = n11885 | n11887 ;
  assign n69437 = ~n11454 ;
  assign n11889 = n69437 & n11888 ;
  assign n69438 = ~n11444 ;
  assign n11890 = x96 & n69438 ;
  assign n69439 = ~n11439 ;
  assign n11891 = n69439 & n11890 ;
  assign n11892 = n11446 | n11891 ;
  assign n11894 = n11889 | n11892 ;
  assign n69440 = ~n11446 ;
  assign n11899 = n69440 & n11894 ;
  assign n11900 = n11897 | n11899 ;
  assign n69441 = ~n11438 ;
  assign n11901 = n69441 & n11900 ;
  assign n69442 = ~n11428 ;
  assign n11902 = x98 & n69442 ;
  assign n69443 = ~n11423 ;
  assign n11903 = n69443 & n11902 ;
  assign n11904 = n11430 | n11903 ;
  assign n11906 = n11901 | n11904 ;
  assign n69444 = ~n11430 ;
  assign n11911 = n69444 & n11906 ;
  assign n11912 = n11909 | n11911 ;
  assign n69445 = ~n11422 ;
  assign n11913 = n69445 & n11912 ;
  assign n69446 = ~n11412 ;
  assign n11914 = x100 & n69446 ;
  assign n69447 = ~n11407 ;
  assign n11915 = n69447 & n11914 ;
  assign n11916 = n11414 | n11915 ;
  assign n11918 = n11913 | n11916 ;
  assign n69448 = ~n11414 ;
  assign n11924 = n69448 & n11918 ;
  assign n11925 = n11923 | n11924 ;
  assign n69449 = ~n11406 ;
  assign n11926 = n69449 & n11925 ;
  assign n11930 = n11926 | n11929 ;
  assign n69450 = ~n11405 ;
  assign n11932 = n69450 & n11930 ;
  assign n69451 = ~n11924 ;
  assign n12518 = n11923 & n69451 ;
  assign n11934 = x65 & n11711 ;
  assign n69452 = ~n11934 ;
  assign n11935 = n11707 & n69452 ;
  assign n11937 = n11708 | n11935 ;
  assign n11938 = n69377 & n11937 ;
  assign n11939 = n11716 | n11938 ;
  assign n11940 = n69380 & n11939 ;
  assign n11941 = n11720 | n11940 ;
  assign n11942 = n69381 & n11941 ;
  assign n11943 = n11726 | n11942 ;
  assign n11944 = n69384 & n11943 ;
  assign n11945 = n11730 | n11944 ;
  assign n11946 = n69385 & n11945 ;
  assign n11947 = n11736 | n11946 ;
  assign n11948 = n69388 & n11947 ;
  assign n11949 = n11741 | n11948 ;
  assign n11950 = n69389 & n11949 ;
  assign n11951 = n11748 | n11950 ;
  assign n11952 = n69392 & n11951 ;
  assign n11953 = n11753 | n11952 ;
  assign n11954 = n69393 & n11953 ;
  assign n11955 = n11760 | n11954 ;
  assign n11956 = n69396 & n11955 ;
  assign n11957 = n11765 | n11956 ;
  assign n11958 = n69397 & n11957 ;
  assign n11959 = n11772 | n11958 ;
  assign n11960 = n69400 & n11959 ;
  assign n11961 = n11777 | n11960 ;
  assign n11962 = n69401 & n11961 ;
  assign n11963 = n11784 | n11962 ;
  assign n11964 = n69404 & n11963 ;
  assign n11965 = n11789 | n11964 ;
  assign n11966 = n69405 & n11965 ;
  assign n11967 = n11796 | n11966 ;
  assign n11968 = n69408 & n11967 ;
  assign n11969 = n11801 | n11968 ;
  assign n11970 = n69409 & n11969 ;
  assign n11971 = n11808 | n11970 ;
  assign n11972 = n69412 & n11971 ;
  assign n11973 = n11813 | n11972 ;
  assign n11974 = n69413 & n11973 ;
  assign n11975 = n11820 | n11974 ;
  assign n11976 = n69416 & n11975 ;
  assign n11977 = n11825 | n11976 ;
  assign n11978 = n69417 & n11977 ;
  assign n11979 = n11832 | n11978 ;
  assign n11980 = n69420 & n11979 ;
  assign n11981 = n11837 | n11980 ;
  assign n11982 = n69421 & n11981 ;
  assign n11983 = n11844 | n11982 ;
  assign n11984 = n69424 & n11983 ;
  assign n11985 = n11849 | n11984 ;
  assign n11986 = n69425 & n11985 ;
  assign n11987 = n11856 | n11986 ;
  assign n11988 = n69428 & n11987 ;
  assign n11989 = n11861 | n11988 ;
  assign n11990 = n69429 & n11989 ;
  assign n11991 = n11868 | n11990 ;
  assign n11992 = n69432 & n11991 ;
  assign n11993 = n11873 | n11992 ;
  assign n11994 = n69433 & n11993 ;
  assign n11995 = n11880 | n11994 ;
  assign n11996 = n69436 & n11995 ;
  assign n11997 = n11885 | n11996 ;
  assign n11998 = n69437 & n11997 ;
  assign n11999 = n11892 | n11998 ;
  assign n12000 = n69440 & n11999 ;
  assign n12001 = n11897 | n12000 ;
  assign n12002 = n69441 & n12001 ;
  assign n12003 = n11904 | n12002 ;
  assign n12004 = n69444 & n12003 ;
  assign n12005 = n11909 | n12004 ;
  assign n12007 = n69445 & n12005 ;
  assign n12303 = n11916 | n12007 ;
  assign n12519 = n11414 | n11923 ;
  assign n69453 = ~n12519 ;
  assign n12520 = n12303 & n69453 ;
  assign n12521 = n12518 | n12520 ;
  assign n12522 = n11930 | n12521 ;
  assign n69454 = ~n11932 ;
  assign n12523 = n69454 & n12522 ;
  assign n69455 = ~n11929 ;
  assign n12534 = n69455 & n12523 ;
  assign n11933 = n11413 & n11930 ;
  assign n11917 = n11422 | n11916 ;
  assign n69456 = ~n11917 ;
  assign n12006 = n69456 & n12005 ;
  assign n69457 = ~n12007 ;
  assign n12008 = n11916 & n69457 ;
  assign n12009 = n12006 | n12008 ;
  assign n12010 = n69455 & n12009 ;
  assign n69458 = ~n11926 ;
  assign n12011 = n69458 & n12010 ;
  assign n12012 = n11933 | n12011 ;
  assign n12013 = n69261 & n12012 ;
  assign n12014 = n11421 & n11930 ;
  assign n11910 = n11430 | n11909 ;
  assign n69459 = ~n11910 ;
  assign n12015 = n11906 & n69459 ;
  assign n69460 = ~n11911 ;
  assign n12016 = n11909 & n69460 ;
  assign n12017 = n12015 | n12016 ;
  assign n12018 = n69455 & n12017 ;
  assign n12019 = n69458 & n12018 ;
  assign n12020 = n12014 | n12019 ;
  assign n12021 = n69075 & n12020 ;
  assign n12022 = n11429 & n11930 ;
  assign n11905 = n11438 | n11904 ;
  assign n69461 = ~n11905 ;
  assign n12023 = n69461 & n12001 ;
  assign n69462 = ~n12002 ;
  assign n12024 = n11904 & n69462 ;
  assign n12025 = n12023 | n12024 ;
  assign n12026 = n69455 & n12025 ;
  assign n12027 = n69458 & n12026 ;
  assign n12028 = n12022 | n12027 ;
  assign n12029 = n68993 & n12028 ;
  assign n12030 = n11437 & n11930 ;
  assign n11898 = n11446 | n11897 ;
  assign n69463 = ~n11898 ;
  assign n12031 = n11894 & n69463 ;
  assign n69464 = ~n11899 ;
  assign n12032 = n11897 & n69464 ;
  assign n12033 = n12031 | n12032 ;
  assign n12034 = n69455 & n12033 ;
  assign n12035 = n69458 & n12034 ;
  assign n12036 = n12030 | n12035 ;
  assign n12037 = n68716 & n12036 ;
  assign n12038 = n11445 & n11930 ;
  assign n11893 = n11454 | n11892 ;
  assign n69465 = ~n11893 ;
  assign n12039 = n69465 & n11997 ;
  assign n69466 = ~n11998 ;
  assign n12040 = n11892 & n69466 ;
  assign n12041 = n12039 | n12040 ;
  assign n12042 = n69455 & n12041 ;
  assign n12043 = n69458 & n12042 ;
  assign n12044 = n12038 | n12043 ;
  assign n12045 = n68545 & n12044 ;
  assign n12046 = n11453 & n11930 ;
  assign n11886 = n11462 | n11885 ;
  assign n69467 = ~n11886 ;
  assign n12047 = n11882 & n69467 ;
  assign n69468 = ~n11887 ;
  assign n12048 = n11885 & n69468 ;
  assign n12049 = n12047 | n12048 ;
  assign n12050 = n69455 & n12049 ;
  assign n12051 = n69458 & n12050 ;
  assign n12052 = n12046 | n12051 ;
  assign n12053 = n68438 & n12052 ;
  assign n12054 = n11461 & n11930 ;
  assign n11881 = n11470 | n11880 ;
  assign n69469 = ~n11881 ;
  assign n12055 = n69469 & n11993 ;
  assign n69470 = ~n11994 ;
  assign n12056 = n11880 & n69470 ;
  assign n12057 = n12055 | n12056 ;
  assign n12058 = n69455 & n12057 ;
  assign n12059 = n69458 & n12058 ;
  assign n12060 = n12054 | n12059 ;
  assign n12061 = n68214 & n12060 ;
  assign n12062 = n11469 & n11930 ;
  assign n11874 = n11478 | n11873 ;
  assign n69471 = ~n11874 ;
  assign n12063 = n11870 & n69471 ;
  assign n69472 = ~n11875 ;
  assign n12064 = n11873 & n69472 ;
  assign n12065 = n12063 | n12064 ;
  assign n12066 = n69455 & n12065 ;
  assign n12067 = n69458 & n12066 ;
  assign n12068 = n12062 | n12067 ;
  assign n12069 = n68058 & n12068 ;
  assign n12070 = n11477 & n11930 ;
  assign n11869 = n11486 | n11868 ;
  assign n69473 = ~n11869 ;
  assign n12071 = n69473 & n11989 ;
  assign n69474 = ~n11990 ;
  assign n12072 = n11868 & n69474 ;
  assign n12073 = n12071 | n12072 ;
  assign n12074 = n69455 & n12073 ;
  assign n12075 = n69458 & n12074 ;
  assign n12076 = n12070 | n12075 ;
  assign n12077 = n67986 & n12076 ;
  assign n12078 = n11485 & n11930 ;
  assign n11862 = n11494 | n11861 ;
  assign n69475 = ~n11862 ;
  assign n12079 = n11858 & n69475 ;
  assign n69476 = ~n11863 ;
  assign n12080 = n11861 & n69476 ;
  assign n12081 = n12079 | n12080 ;
  assign n12082 = n69455 & n12081 ;
  assign n12083 = n69458 & n12082 ;
  assign n12084 = n12078 | n12083 ;
  assign n12085 = n67763 & n12084 ;
  assign n12086 = n11493 & n11930 ;
  assign n11857 = n11502 | n11856 ;
  assign n69477 = ~n11857 ;
  assign n12087 = n69477 & n11985 ;
  assign n69478 = ~n11986 ;
  assign n12088 = n11856 & n69478 ;
  assign n12089 = n12087 | n12088 ;
  assign n12090 = n69455 & n12089 ;
  assign n12091 = n69458 & n12090 ;
  assign n12092 = n12086 | n12091 ;
  assign n12093 = n67622 & n12092 ;
  assign n12094 = n11501 & n11930 ;
  assign n11850 = n11510 | n11849 ;
  assign n69479 = ~n11850 ;
  assign n12095 = n11846 & n69479 ;
  assign n69480 = ~n11851 ;
  assign n12096 = n11849 & n69480 ;
  assign n12097 = n12095 | n12096 ;
  assign n12098 = n69455 & n12097 ;
  assign n12099 = n69458 & n12098 ;
  assign n12100 = n12094 | n12099 ;
  assign n12101 = n67531 & n12100 ;
  assign n12102 = n11509 & n11930 ;
  assign n11845 = n11518 | n11844 ;
  assign n69481 = ~n11845 ;
  assign n12103 = n69481 & n11981 ;
  assign n69482 = ~n11982 ;
  assign n12104 = n11844 & n69482 ;
  assign n12105 = n12103 | n12104 ;
  assign n12106 = n69455 & n12105 ;
  assign n12107 = n69458 & n12106 ;
  assign n12108 = n12102 | n12107 ;
  assign n12109 = n67348 & n12108 ;
  assign n12110 = n11517 & n11930 ;
  assign n11838 = n11526 | n11837 ;
  assign n69483 = ~n11838 ;
  assign n12111 = n11834 & n69483 ;
  assign n69484 = ~n11839 ;
  assign n12112 = n11837 & n69484 ;
  assign n12113 = n12111 | n12112 ;
  assign n12114 = n69455 & n12113 ;
  assign n12115 = n69458 & n12114 ;
  assign n12116 = n12110 | n12115 ;
  assign n12117 = n67222 & n12116 ;
  assign n12118 = n11525 & n11930 ;
  assign n11833 = n11534 | n11832 ;
  assign n69485 = ~n11833 ;
  assign n12119 = n69485 & n11977 ;
  assign n69486 = ~n11978 ;
  assign n12120 = n11832 & n69486 ;
  assign n12121 = n12119 | n12120 ;
  assign n12122 = n69455 & n12121 ;
  assign n12123 = n69458 & n12122 ;
  assign n12124 = n12118 | n12123 ;
  assign n12125 = n67164 & n12124 ;
  assign n12126 = n11533 & n11930 ;
  assign n11826 = n11542 | n11825 ;
  assign n69487 = ~n11826 ;
  assign n12127 = n11822 & n69487 ;
  assign n69488 = ~n11827 ;
  assign n12128 = n11825 & n69488 ;
  assign n12129 = n12127 | n12128 ;
  assign n12130 = n69455 & n12129 ;
  assign n12131 = n69458 & n12130 ;
  assign n12132 = n12126 | n12131 ;
  assign n12133 = n66979 & n12132 ;
  assign n12134 = n11541 & n11930 ;
  assign n11821 = n11550 | n11820 ;
  assign n69489 = ~n11821 ;
  assign n12135 = n69489 & n11973 ;
  assign n69490 = ~n11974 ;
  assign n12136 = n11820 & n69490 ;
  assign n12137 = n12135 | n12136 ;
  assign n12138 = n69455 & n12137 ;
  assign n12139 = n69458 & n12138 ;
  assign n12140 = n12134 | n12139 ;
  assign n12141 = n66868 & n12140 ;
  assign n12142 = n11549 & n11930 ;
  assign n11814 = n11558 | n11813 ;
  assign n69491 = ~n11814 ;
  assign n12143 = n11810 & n69491 ;
  assign n69492 = ~n11815 ;
  assign n12144 = n11813 & n69492 ;
  assign n12145 = n12143 | n12144 ;
  assign n12146 = n69455 & n12145 ;
  assign n12147 = n69458 & n12146 ;
  assign n12148 = n12142 | n12147 ;
  assign n12149 = n66797 & n12148 ;
  assign n12150 = n11557 & n11930 ;
  assign n11809 = n11566 | n11808 ;
  assign n69493 = ~n11809 ;
  assign n12151 = n69493 & n11969 ;
  assign n69494 = ~n11970 ;
  assign n12152 = n11808 & n69494 ;
  assign n12153 = n12151 | n12152 ;
  assign n12154 = n69455 & n12153 ;
  assign n12155 = n69458 & n12154 ;
  assign n12156 = n12150 | n12155 ;
  assign n12157 = n66654 & n12156 ;
  assign n12158 = n11565 & n11930 ;
  assign n11802 = n11574 | n11801 ;
  assign n69495 = ~n11802 ;
  assign n12159 = n11798 & n69495 ;
  assign n69496 = ~n11803 ;
  assign n12160 = n11801 & n69496 ;
  assign n12161 = n12159 | n12160 ;
  assign n12162 = n69455 & n12161 ;
  assign n12163 = n69458 & n12162 ;
  assign n12164 = n12158 | n12163 ;
  assign n12165 = n66560 & n12164 ;
  assign n12166 = n11573 & n11930 ;
  assign n11797 = n11582 | n11796 ;
  assign n69497 = ~n11797 ;
  assign n12167 = n69497 & n11965 ;
  assign n69498 = ~n11966 ;
  assign n12168 = n11796 & n69498 ;
  assign n12169 = n12167 | n12168 ;
  assign n12170 = n69455 & n12169 ;
  assign n12171 = n69458 & n12170 ;
  assign n12172 = n12166 | n12171 ;
  assign n12173 = n66505 & n12172 ;
  assign n12174 = n11581 & n11930 ;
  assign n11790 = n11590 | n11789 ;
  assign n69499 = ~n11790 ;
  assign n12175 = n11786 & n69499 ;
  assign n69500 = ~n11791 ;
  assign n12176 = n11789 & n69500 ;
  assign n12177 = n12175 | n12176 ;
  assign n12178 = n69455 & n12177 ;
  assign n12179 = n69458 & n12178 ;
  assign n12180 = n12174 | n12179 ;
  assign n12181 = n66379 & n12180 ;
  assign n12182 = n11589 & n11930 ;
  assign n11785 = n11598 | n11784 ;
  assign n69501 = ~n11785 ;
  assign n12183 = n69501 & n11961 ;
  assign n69502 = ~n11962 ;
  assign n12184 = n11784 & n69502 ;
  assign n12185 = n12183 | n12184 ;
  assign n12186 = n69455 & n12185 ;
  assign n12187 = n69458 & n12186 ;
  assign n12188 = n12182 | n12187 ;
  assign n12189 = n66299 & n12188 ;
  assign n12190 = n11597 & n11930 ;
  assign n11778 = n11606 | n11777 ;
  assign n69503 = ~n11778 ;
  assign n12191 = n11774 & n69503 ;
  assign n69504 = ~n11779 ;
  assign n12192 = n11777 & n69504 ;
  assign n12193 = n12191 | n12192 ;
  assign n12194 = n69455 & n12193 ;
  assign n12195 = n69458 & n12194 ;
  assign n12196 = n12190 | n12195 ;
  assign n12197 = n66244 & n12196 ;
  assign n12198 = n11605 & n11930 ;
  assign n11773 = n11614 | n11772 ;
  assign n69505 = ~n11773 ;
  assign n12199 = n69505 & n11957 ;
  assign n69506 = ~n11958 ;
  assign n12200 = n11772 & n69506 ;
  assign n12201 = n12199 | n12200 ;
  assign n12202 = n69455 & n12201 ;
  assign n12203 = n69458 & n12202 ;
  assign n12204 = n12198 | n12203 ;
  assign n12205 = n66145 & n12204 ;
  assign n12206 = n11613 & n11930 ;
  assign n11766 = n11622 | n11765 ;
  assign n69507 = ~n11766 ;
  assign n12207 = n11762 & n69507 ;
  assign n69508 = ~n11767 ;
  assign n12208 = n11765 & n69508 ;
  assign n12209 = n12207 | n12208 ;
  assign n12210 = n69455 & n12209 ;
  assign n12211 = n69458 & n12210 ;
  assign n12212 = n12206 | n12211 ;
  assign n12213 = n66081 & n12212 ;
  assign n12214 = n11621 & n11930 ;
  assign n11761 = n11630 | n11760 ;
  assign n69509 = ~n11761 ;
  assign n12215 = n69509 & n11953 ;
  assign n69510 = ~n11954 ;
  assign n12216 = n11760 & n69510 ;
  assign n12217 = n12215 | n12216 ;
  assign n12218 = n69455 & n12217 ;
  assign n12219 = n69458 & n12218 ;
  assign n12220 = n12214 | n12219 ;
  assign n12221 = n66043 & n12220 ;
  assign n12222 = n11629 & n11930 ;
  assign n11754 = n11638 | n11753 ;
  assign n69511 = ~n11754 ;
  assign n12223 = n11750 & n69511 ;
  assign n69512 = ~n11755 ;
  assign n12224 = n11753 & n69512 ;
  assign n12225 = n12223 | n12224 ;
  assign n12226 = n69455 & n12225 ;
  assign n12227 = n69458 & n12226 ;
  assign n12228 = n12222 | n12227 ;
  assign n12229 = n65960 & n12228 ;
  assign n12230 = n11637 & n11930 ;
  assign n11749 = n11646 | n11748 ;
  assign n69513 = ~n11749 ;
  assign n12231 = n69513 & n11949 ;
  assign n69514 = ~n11950 ;
  assign n12232 = n11748 & n69514 ;
  assign n12233 = n12231 | n12232 ;
  assign n12234 = n69455 & n12233 ;
  assign n12235 = n69458 & n12234 ;
  assign n12236 = n12230 | n12235 ;
  assign n12237 = n65909 & n12236 ;
  assign n12238 = n11645 & n11930 ;
  assign n11742 = n11654 | n11741 ;
  assign n69515 = ~n11742 ;
  assign n12239 = n11738 & n69515 ;
  assign n69516 = ~n11743 ;
  assign n12240 = n11741 & n69516 ;
  assign n12241 = n12239 | n12240 ;
  assign n12242 = n69455 & n12241 ;
  assign n12243 = n69458 & n12242 ;
  assign n12244 = n12238 | n12243 ;
  assign n12245 = n65877 & n12244 ;
  assign n12246 = n11653 & n11930 ;
  assign n11737 = n11662 | n11736 ;
  assign n69517 = ~n11737 ;
  assign n12247 = n11732 & n69517 ;
  assign n69518 = ~n11946 ;
  assign n12248 = n11736 & n69518 ;
  assign n12249 = n12247 | n12248 ;
  assign n12250 = n69455 & n12249 ;
  assign n12251 = n69458 & n12250 ;
  assign n12252 = n12246 | n12251 ;
  assign n12253 = n65820 & n12252 ;
  assign n12254 = n11661 & n11930 ;
  assign n12255 = n11670 | n11730 ;
  assign n69519 = ~n12255 ;
  assign n12256 = n11727 & n69519 ;
  assign n69520 = ~n11731 ;
  assign n12257 = n11730 & n69520 ;
  assign n12258 = n12256 | n12257 ;
  assign n12259 = n69455 & n12258 ;
  assign n12260 = n69458 & n12259 ;
  assign n12261 = n12254 | n12260 ;
  assign n12262 = n65791 & n12261 ;
  assign n12263 = n11669 & n11930 ;
  assign n12264 = n11679 | n11726 ;
  assign n69521 = ~n12264 ;
  assign n12265 = n11722 & n69521 ;
  assign n69522 = ~n11942 ;
  assign n12266 = n11726 & n69522 ;
  assign n12267 = n12265 | n12266 ;
  assign n12268 = n69455 & n12267 ;
  assign n12269 = n69458 & n12268 ;
  assign n12270 = n12263 | n12269 ;
  assign n12271 = n65772 & n12270 ;
  assign n12272 = n11678 & n11930 ;
  assign n12273 = n11687 | n11720 ;
  assign n69523 = ~n12273 ;
  assign n12274 = n11717 & n69523 ;
  assign n69524 = ~n11721 ;
  assign n12275 = n11720 & n69524 ;
  assign n12276 = n12274 | n12275 ;
  assign n12277 = n69455 & n12276 ;
  assign n12278 = n69458 & n12277 ;
  assign n12279 = n12272 | n12278 ;
  assign n12280 = n65746 & n12279 ;
  assign n12281 = n11686 & n11930 ;
  assign n69525 = ~n11713 ;
  assign n12282 = n69525 & n11716 ;
  assign n12283 = n11712 | n11716 ;
  assign n69526 = ~n12283 ;
  assign n12284 = n11710 & n69526 ;
  assign n12285 = n12282 | n12284 ;
  assign n12286 = n69455 & n12285 ;
  assign n12287 = n69458 & n12286 ;
  assign n12288 = n12281 | n12287 ;
  assign n12289 = n65721 & n12288 ;
  assign n11931 = n11711 & n11930 ;
  assign n11936 = n11707 & n11708 ;
  assign n12290 = n69376 & n11936 ;
  assign n12291 = n11929 | n12290 ;
  assign n69527 = ~n12291 ;
  assign n12292 = n11710 & n69527 ;
  assign n12293 = n69458 & n12292 ;
  assign n12294 = n11931 | n12293 ;
  assign n12295 = n65686 & n12294 ;
  assign n69528 = ~x102 ;
  assign n12296 = x64 & n69528 ;
  assign n69529 = ~n281 ;
  assign n12297 = n69529 & n12296 ;
  assign n69530 = ~n292 ;
  assign n12298 = n69530 & n12297 ;
  assign n69531 = ~n467 ;
  assign n12299 = n69531 & n12298 ;
  assign n12300 = n67026 & n12299 ;
  assign n12304 = n69448 & n12303 ;
  assign n12305 = n11923 | n12304 ;
  assign n12306 = n69449 & n12305 ;
  assign n69532 = ~n12306 ;
  assign n12307 = n12300 & n69532 ;
  assign n69533 = ~n12307 ;
  assign n12308 = x26 & n69533 ;
  assign n12309 = n69370 & n11708 ;
  assign n12310 = n69371 & n12309 ;
  assign n12311 = n69372 & n12310 ;
  assign n12312 = n67021 & n12311 ;
  assign n12313 = n69458 & n12312 ;
  assign n12314 = n12308 | n12313 ;
  assign n12316 = x65 & n12314 ;
  assign n12301 = n69458 & n12300 ;
  assign n69534 = ~n12301 ;
  assign n12302 = x26 & n69534 ;
  assign n12315 = x65 | n12313 ;
  assign n12317 = n12302 | n12315 ;
  assign n69535 = ~n12316 ;
  assign n12318 = n69535 & n12317 ;
  assign n69536 = ~x25 ;
  assign n12319 = n69536 & x64 ;
  assign n12320 = n12318 | n12319 ;
  assign n12321 = n65670 & n12314 ;
  assign n69537 = ~n12321 ;
  assign n12322 = n12320 & n69537 ;
  assign n69538 = ~n12293 ;
  assign n12323 = x66 & n69538 ;
  assign n69539 = ~n11931 ;
  assign n12324 = n69539 & n12323 ;
  assign n12325 = n12295 | n12324 ;
  assign n12326 = n12322 | n12325 ;
  assign n69540 = ~n12295 ;
  assign n12327 = n69540 & n12326 ;
  assign n69541 = ~n12287 ;
  assign n12328 = x67 & n69541 ;
  assign n69542 = ~n12281 ;
  assign n12329 = n69542 & n12328 ;
  assign n12330 = n12327 | n12329 ;
  assign n69543 = ~n12289 ;
  assign n12331 = n69543 & n12330 ;
  assign n69544 = ~n12278 ;
  assign n12332 = x68 & n69544 ;
  assign n69545 = ~n12272 ;
  assign n12333 = n69545 & n12332 ;
  assign n12334 = n12280 | n12333 ;
  assign n12335 = n12331 | n12334 ;
  assign n69546 = ~n12280 ;
  assign n12336 = n69546 & n12335 ;
  assign n69547 = ~n12269 ;
  assign n12337 = x69 & n69547 ;
  assign n69548 = ~n12263 ;
  assign n12338 = n69548 & n12337 ;
  assign n12339 = n12271 | n12338 ;
  assign n12340 = n12336 | n12339 ;
  assign n69549 = ~n12271 ;
  assign n12341 = n69549 & n12340 ;
  assign n69550 = ~n12260 ;
  assign n12342 = x70 & n69550 ;
  assign n69551 = ~n12254 ;
  assign n12343 = n69551 & n12342 ;
  assign n12344 = n12262 | n12343 ;
  assign n12345 = n12341 | n12344 ;
  assign n69552 = ~n12262 ;
  assign n12346 = n69552 & n12345 ;
  assign n69553 = ~n12251 ;
  assign n12347 = x71 & n69553 ;
  assign n69554 = ~n12246 ;
  assign n12348 = n69554 & n12347 ;
  assign n12349 = n12253 | n12348 ;
  assign n12351 = n12346 | n12349 ;
  assign n69555 = ~n12253 ;
  assign n12352 = n69555 & n12351 ;
  assign n69556 = ~n12243 ;
  assign n12353 = x72 & n69556 ;
  assign n69557 = ~n12238 ;
  assign n12354 = n69557 & n12353 ;
  assign n12355 = n12245 | n12354 ;
  assign n12356 = n12352 | n12355 ;
  assign n69558 = ~n12245 ;
  assign n12357 = n69558 & n12356 ;
  assign n69559 = ~n12235 ;
  assign n12358 = x73 & n69559 ;
  assign n69560 = ~n12230 ;
  assign n12359 = n69560 & n12358 ;
  assign n12360 = n12237 | n12359 ;
  assign n12362 = n12357 | n12360 ;
  assign n69561 = ~n12237 ;
  assign n12363 = n69561 & n12362 ;
  assign n69562 = ~n12227 ;
  assign n12364 = x74 & n69562 ;
  assign n69563 = ~n12222 ;
  assign n12365 = n69563 & n12364 ;
  assign n12366 = n12229 | n12365 ;
  assign n12367 = n12363 | n12366 ;
  assign n69564 = ~n12229 ;
  assign n12368 = n69564 & n12367 ;
  assign n69565 = ~n12219 ;
  assign n12369 = x75 & n69565 ;
  assign n69566 = ~n12214 ;
  assign n12370 = n69566 & n12369 ;
  assign n12371 = n12221 | n12370 ;
  assign n12373 = n12368 | n12371 ;
  assign n69567 = ~n12221 ;
  assign n12374 = n69567 & n12373 ;
  assign n69568 = ~n12211 ;
  assign n12375 = x76 & n69568 ;
  assign n69569 = ~n12206 ;
  assign n12376 = n69569 & n12375 ;
  assign n12377 = n12213 | n12376 ;
  assign n12378 = n12374 | n12377 ;
  assign n69570 = ~n12213 ;
  assign n12379 = n69570 & n12378 ;
  assign n69571 = ~n12203 ;
  assign n12380 = x77 & n69571 ;
  assign n69572 = ~n12198 ;
  assign n12381 = n69572 & n12380 ;
  assign n12382 = n12205 | n12381 ;
  assign n12384 = n12379 | n12382 ;
  assign n69573 = ~n12205 ;
  assign n12385 = n69573 & n12384 ;
  assign n69574 = ~n12195 ;
  assign n12386 = x78 & n69574 ;
  assign n69575 = ~n12190 ;
  assign n12387 = n69575 & n12386 ;
  assign n12388 = n12197 | n12387 ;
  assign n12389 = n12385 | n12388 ;
  assign n69576 = ~n12197 ;
  assign n12390 = n69576 & n12389 ;
  assign n69577 = ~n12187 ;
  assign n12391 = x79 & n69577 ;
  assign n69578 = ~n12182 ;
  assign n12392 = n69578 & n12391 ;
  assign n12393 = n12189 | n12392 ;
  assign n12395 = n12390 | n12393 ;
  assign n69579 = ~n12189 ;
  assign n12396 = n69579 & n12395 ;
  assign n69580 = ~n12179 ;
  assign n12397 = x80 & n69580 ;
  assign n69581 = ~n12174 ;
  assign n12398 = n69581 & n12397 ;
  assign n12399 = n12181 | n12398 ;
  assign n12400 = n12396 | n12399 ;
  assign n69582 = ~n12181 ;
  assign n12401 = n69582 & n12400 ;
  assign n69583 = ~n12171 ;
  assign n12402 = x81 & n69583 ;
  assign n69584 = ~n12166 ;
  assign n12403 = n69584 & n12402 ;
  assign n12404 = n12173 | n12403 ;
  assign n12406 = n12401 | n12404 ;
  assign n69585 = ~n12173 ;
  assign n12407 = n69585 & n12406 ;
  assign n69586 = ~n12163 ;
  assign n12408 = x82 & n69586 ;
  assign n69587 = ~n12158 ;
  assign n12409 = n69587 & n12408 ;
  assign n12410 = n12165 | n12409 ;
  assign n12411 = n12407 | n12410 ;
  assign n69588 = ~n12165 ;
  assign n12412 = n69588 & n12411 ;
  assign n69589 = ~n12155 ;
  assign n12413 = x83 & n69589 ;
  assign n69590 = ~n12150 ;
  assign n12414 = n69590 & n12413 ;
  assign n12415 = n12157 | n12414 ;
  assign n12417 = n12412 | n12415 ;
  assign n69591 = ~n12157 ;
  assign n12418 = n69591 & n12417 ;
  assign n69592 = ~n12147 ;
  assign n12419 = x84 & n69592 ;
  assign n69593 = ~n12142 ;
  assign n12420 = n69593 & n12419 ;
  assign n12421 = n12149 | n12420 ;
  assign n12422 = n12418 | n12421 ;
  assign n69594 = ~n12149 ;
  assign n12423 = n69594 & n12422 ;
  assign n69595 = ~n12139 ;
  assign n12424 = x85 & n69595 ;
  assign n69596 = ~n12134 ;
  assign n12425 = n69596 & n12424 ;
  assign n12426 = n12141 | n12425 ;
  assign n12428 = n12423 | n12426 ;
  assign n69597 = ~n12141 ;
  assign n12429 = n69597 & n12428 ;
  assign n69598 = ~n12131 ;
  assign n12430 = x86 & n69598 ;
  assign n69599 = ~n12126 ;
  assign n12431 = n69599 & n12430 ;
  assign n12432 = n12133 | n12431 ;
  assign n12433 = n12429 | n12432 ;
  assign n69600 = ~n12133 ;
  assign n12434 = n69600 & n12433 ;
  assign n69601 = ~n12123 ;
  assign n12435 = x87 & n69601 ;
  assign n69602 = ~n12118 ;
  assign n12436 = n69602 & n12435 ;
  assign n12437 = n12125 | n12436 ;
  assign n12439 = n12434 | n12437 ;
  assign n69603 = ~n12125 ;
  assign n12440 = n69603 & n12439 ;
  assign n69604 = ~n12115 ;
  assign n12441 = x88 & n69604 ;
  assign n69605 = ~n12110 ;
  assign n12442 = n69605 & n12441 ;
  assign n12443 = n12117 | n12442 ;
  assign n12444 = n12440 | n12443 ;
  assign n69606 = ~n12117 ;
  assign n12445 = n69606 & n12444 ;
  assign n69607 = ~n12107 ;
  assign n12446 = x89 & n69607 ;
  assign n69608 = ~n12102 ;
  assign n12447 = n69608 & n12446 ;
  assign n12448 = n12109 | n12447 ;
  assign n12450 = n12445 | n12448 ;
  assign n69609 = ~n12109 ;
  assign n12451 = n69609 & n12450 ;
  assign n69610 = ~n12099 ;
  assign n12452 = x90 & n69610 ;
  assign n69611 = ~n12094 ;
  assign n12453 = n69611 & n12452 ;
  assign n12454 = n12101 | n12453 ;
  assign n12455 = n12451 | n12454 ;
  assign n69612 = ~n12101 ;
  assign n12456 = n69612 & n12455 ;
  assign n69613 = ~n12091 ;
  assign n12457 = x91 & n69613 ;
  assign n69614 = ~n12086 ;
  assign n12458 = n69614 & n12457 ;
  assign n12459 = n12093 | n12458 ;
  assign n12461 = n12456 | n12459 ;
  assign n69615 = ~n12093 ;
  assign n12462 = n69615 & n12461 ;
  assign n69616 = ~n12083 ;
  assign n12463 = x92 & n69616 ;
  assign n69617 = ~n12078 ;
  assign n12464 = n69617 & n12463 ;
  assign n12465 = n12085 | n12464 ;
  assign n12466 = n12462 | n12465 ;
  assign n69618 = ~n12085 ;
  assign n12467 = n69618 & n12466 ;
  assign n69619 = ~n12075 ;
  assign n12468 = x93 & n69619 ;
  assign n69620 = ~n12070 ;
  assign n12469 = n69620 & n12468 ;
  assign n12470 = n12077 | n12469 ;
  assign n12472 = n12467 | n12470 ;
  assign n69621 = ~n12077 ;
  assign n12473 = n69621 & n12472 ;
  assign n69622 = ~n12067 ;
  assign n12474 = x94 & n69622 ;
  assign n69623 = ~n12062 ;
  assign n12475 = n69623 & n12474 ;
  assign n12476 = n12069 | n12475 ;
  assign n12477 = n12473 | n12476 ;
  assign n69624 = ~n12069 ;
  assign n12478 = n69624 & n12477 ;
  assign n69625 = ~n12059 ;
  assign n12479 = x95 & n69625 ;
  assign n69626 = ~n12054 ;
  assign n12480 = n69626 & n12479 ;
  assign n12481 = n12061 | n12480 ;
  assign n12483 = n12478 | n12481 ;
  assign n69627 = ~n12061 ;
  assign n12484 = n69627 & n12483 ;
  assign n69628 = ~n12051 ;
  assign n12485 = x96 & n69628 ;
  assign n69629 = ~n12046 ;
  assign n12486 = n69629 & n12485 ;
  assign n12487 = n12053 | n12486 ;
  assign n12488 = n12484 | n12487 ;
  assign n69630 = ~n12053 ;
  assign n12489 = n69630 & n12488 ;
  assign n69631 = ~n12043 ;
  assign n12490 = x97 & n69631 ;
  assign n69632 = ~n12038 ;
  assign n12491 = n69632 & n12490 ;
  assign n12492 = n12045 | n12491 ;
  assign n12494 = n12489 | n12492 ;
  assign n69633 = ~n12045 ;
  assign n12495 = n69633 & n12494 ;
  assign n69634 = ~n12035 ;
  assign n12496 = x98 & n69634 ;
  assign n69635 = ~n12030 ;
  assign n12497 = n69635 & n12496 ;
  assign n12498 = n12037 | n12497 ;
  assign n12499 = n12495 | n12498 ;
  assign n69636 = ~n12037 ;
  assign n12500 = n69636 & n12499 ;
  assign n69637 = ~n12027 ;
  assign n12501 = x99 & n69637 ;
  assign n69638 = ~n12022 ;
  assign n12502 = n69638 & n12501 ;
  assign n12503 = n12029 | n12502 ;
  assign n12505 = n12500 | n12503 ;
  assign n69639 = ~n12029 ;
  assign n12506 = n69639 & n12505 ;
  assign n69640 = ~n12019 ;
  assign n12507 = x100 & n69640 ;
  assign n69641 = ~n12014 ;
  assign n12508 = n69641 & n12507 ;
  assign n12509 = n12021 | n12508 ;
  assign n12510 = n12506 | n12509 ;
  assign n69642 = ~n12021 ;
  assign n12511 = n69642 & n12510 ;
  assign n69643 = ~n12011 ;
  assign n12512 = x101 & n69643 ;
  assign n69644 = ~n11933 ;
  assign n12513 = n69644 & n12512 ;
  assign n12514 = n12013 | n12513 ;
  assign n12516 = n12511 | n12514 ;
  assign n69645 = ~n12013 ;
  assign n12517 = n69645 & n12516 ;
  assign n12524 = n69528 & n12523 ;
  assign n155 = ~n11930 ;
  assign n12525 = n155 & n12521 ;
  assign n12526 = n11405 & n11930 ;
  assign n69647 = ~n12526 ;
  assign n12527 = x102 & n69647 ;
  assign n69648 = ~n12525 ;
  assign n12528 = n69648 & n12527 ;
  assign n12529 = n281 | n292 ;
  assign n12530 = n467 | n12529 ;
  assign n12531 = n465 | n12530 ;
  assign n12532 = n12528 | n12531 ;
  assign n12533 = n12524 | n12532 ;
  assign n12535 = n12517 | n12533 ;
  assign n69649 = ~n12534 ;
  assign n12536 = n69649 & n12535 ;
  assign n69650 = ~n12511 ;
  assign n12515 = n69650 & n12514 ;
  assign n12539 = n12302 | n12313 ;
  assign n12540 = x65 & n12539 ;
  assign n69651 = ~n12540 ;
  assign n12541 = n12317 & n69651 ;
  assign n12542 = n12319 | n12541 ;
  assign n12543 = n69537 & n12542 ;
  assign n12545 = n12324 | n12543 ;
  assign n12546 = n69540 & n12545 ;
  assign n12547 = n12289 | n12329 ;
  assign n12549 = n12546 | n12547 ;
  assign n12550 = n69543 & n12549 ;
  assign n12552 = n12334 | n12550 ;
  assign n12553 = n69546 & n12552 ;
  assign n12555 = n12339 | n12553 ;
  assign n12556 = n69549 & n12555 ;
  assign n12557 = n12344 | n12556 ;
  assign n12559 = n69552 & n12557 ;
  assign n12560 = n12349 | n12559 ;
  assign n12561 = n69555 & n12560 ;
  assign n12562 = n12355 | n12561 ;
  assign n12564 = n69558 & n12562 ;
  assign n12565 = n12360 | n12564 ;
  assign n12566 = n69561 & n12565 ;
  assign n12567 = n12366 | n12566 ;
  assign n12569 = n69564 & n12567 ;
  assign n12570 = n12371 | n12569 ;
  assign n12571 = n69567 & n12570 ;
  assign n12572 = n12377 | n12571 ;
  assign n12574 = n69570 & n12572 ;
  assign n12575 = n12382 | n12574 ;
  assign n12576 = n69573 & n12575 ;
  assign n12577 = n12388 | n12576 ;
  assign n12579 = n69576 & n12577 ;
  assign n12580 = n12393 | n12579 ;
  assign n12581 = n69579 & n12580 ;
  assign n12582 = n12399 | n12581 ;
  assign n12584 = n69582 & n12582 ;
  assign n12585 = n12404 | n12584 ;
  assign n12586 = n69585 & n12585 ;
  assign n12587 = n12410 | n12586 ;
  assign n12589 = n69588 & n12587 ;
  assign n12590 = n12415 | n12589 ;
  assign n12591 = n69591 & n12590 ;
  assign n12592 = n12421 | n12591 ;
  assign n12594 = n69594 & n12592 ;
  assign n12595 = n12426 | n12594 ;
  assign n12596 = n69597 & n12595 ;
  assign n12597 = n12432 | n12596 ;
  assign n12599 = n69600 & n12597 ;
  assign n12600 = n12437 | n12599 ;
  assign n12601 = n69603 & n12600 ;
  assign n12602 = n12443 | n12601 ;
  assign n12604 = n69606 & n12602 ;
  assign n12605 = n12448 | n12604 ;
  assign n12606 = n69609 & n12605 ;
  assign n12607 = n12454 | n12606 ;
  assign n12609 = n69612 & n12607 ;
  assign n12610 = n12459 | n12609 ;
  assign n12611 = n69615 & n12610 ;
  assign n12612 = n12465 | n12611 ;
  assign n12614 = n69618 & n12612 ;
  assign n12615 = n12470 | n12614 ;
  assign n12616 = n69621 & n12615 ;
  assign n12617 = n12476 | n12616 ;
  assign n12619 = n69624 & n12617 ;
  assign n12620 = n12481 | n12619 ;
  assign n12621 = n69627 & n12620 ;
  assign n12622 = n12487 | n12621 ;
  assign n12624 = n69630 & n12622 ;
  assign n12625 = n12492 | n12624 ;
  assign n12626 = n69633 & n12625 ;
  assign n12627 = n12498 | n12626 ;
  assign n12629 = n69636 & n12627 ;
  assign n12630 = n12503 | n12629 ;
  assign n12631 = n69639 & n12630 ;
  assign n12632 = n12509 | n12631 ;
  assign n12649 = n12021 | n12514 ;
  assign n69652 = ~n12649 ;
  assign n12650 = n12632 & n69652 ;
  assign n12651 = n12515 | n12650 ;
  assign n154 = ~n12536 ;
  assign n12652 = n154 & n12651 ;
  assign n12634 = n69642 & n12632 ;
  assign n12635 = n12514 | n12634 ;
  assign n12636 = n69645 & n12635 ;
  assign n12637 = n12533 | n12636 ;
  assign n12653 = n12012 & n69649 ;
  assign n12654 = n12637 & n12653 ;
  assign n12655 = n12652 | n12654 ;
  assign n12638 = n12013 | n12528 ;
  assign n12639 = n12524 | n12638 ;
  assign n69654 = ~n12639 ;
  assign n12640 = n12516 & n69654 ;
  assign n12641 = n12524 | n12528 ;
  assign n69655 = ~n12636 ;
  assign n12642 = n69655 & n12641 ;
  assign n12643 = n12640 | n12642 ;
  assign n12644 = n154 & n12643 ;
  assign n12645 = n11929 & n12523 ;
  assign n12646 = n12637 & n12645 ;
  assign n12647 = n12644 | n12646 ;
  assign n69656 = ~x103 ;
  assign n12648 = n69656 & n12647 ;
  assign n69657 = ~n12646 ;
  assign n13178 = x103 & n69657 ;
  assign n69658 = ~n12644 ;
  assign n13179 = n69658 & n13178 ;
  assign n13180 = n12648 | n13179 ;
  assign n12656 = n69528 & n12655 ;
  assign n69659 = ~n12631 ;
  assign n12633 = n12509 & n69659 ;
  assign n12657 = n12029 | n12509 ;
  assign n69660 = ~n12657 ;
  assign n12658 = n12505 & n69660 ;
  assign n12659 = n12633 | n12658 ;
  assign n12660 = n154 & n12659 ;
  assign n12661 = n12020 & n69649 ;
  assign n12662 = n12637 & n12661 ;
  assign n12663 = n12660 | n12662 ;
  assign n12664 = n69261 & n12663 ;
  assign n69661 = ~n12662 ;
  assign n13166 = x101 & n69661 ;
  assign n69662 = ~n12660 ;
  assign n13167 = n69662 & n13166 ;
  assign n13168 = n12664 | n13167 ;
  assign n69663 = ~n12500 ;
  assign n12504 = n69663 & n12503 ;
  assign n12665 = n12037 | n12503 ;
  assign n69664 = ~n12665 ;
  assign n12666 = n12627 & n69664 ;
  assign n12667 = n12504 | n12666 ;
  assign n12668 = n154 & n12667 ;
  assign n12669 = n12028 & n69649 ;
  assign n12670 = n12637 & n12669 ;
  assign n12671 = n12668 | n12670 ;
  assign n12672 = n69075 & n12671 ;
  assign n69665 = ~n12626 ;
  assign n12628 = n12498 & n69665 ;
  assign n12673 = n12045 | n12498 ;
  assign n69666 = ~n12673 ;
  assign n12674 = n12494 & n69666 ;
  assign n12675 = n12628 | n12674 ;
  assign n12676 = n154 & n12675 ;
  assign n12677 = n12036 & n69649 ;
  assign n12678 = n12637 & n12677 ;
  assign n12679 = n12676 | n12678 ;
  assign n12680 = n68993 & n12679 ;
  assign n69667 = ~n12678 ;
  assign n13154 = x99 & n69667 ;
  assign n69668 = ~n12676 ;
  assign n13155 = n69668 & n13154 ;
  assign n13156 = n12680 | n13155 ;
  assign n69669 = ~n12489 ;
  assign n12493 = n69669 & n12492 ;
  assign n12681 = n12053 | n12492 ;
  assign n69670 = ~n12681 ;
  assign n12682 = n12622 & n69670 ;
  assign n12683 = n12493 | n12682 ;
  assign n12684 = n154 & n12683 ;
  assign n12685 = n12044 & n69649 ;
  assign n12686 = n12637 & n12685 ;
  assign n12687 = n12684 | n12686 ;
  assign n12688 = n68716 & n12687 ;
  assign n69671 = ~n12621 ;
  assign n12623 = n12487 & n69671 ;
  assign n12689 = n12061 | n12487 ;
  assign n69672 = ~n12689 ;
  assign n12690 = n12483 & n69672 ;
  assign n12691 = n12623 | n12690 ;
  assign n12692 = n154 & n12691 ;
  assign n12693 = n12052 & n69649 ;
  assign n12694 = n12637 & n12693 ;
  assign n12695 = n12692 | n12694 ;
  assign n12696 = n68545 & n12695 ;
  assign n69673 = ~n12694 ;
  assign n13142 = x97 & n69673 ;
  assign n69674 = ~n12692 ;
  assign n13143 = n69674 & n13142 ;
  assign n13144 = n12696 | n13143 ;
  assign n69675 = ~n12478 ;
  assign n12482 = n69675 & n12481 ;
  assign n12697 = n12069 | n12481 ;
  assign n69676 = ~n12697 ;
  assign n12698 = n12617 & n69676 ;
  assign n12699 = n12482 | n12698 ;
  assign n12700 = n154 & n12699 ;
  assign n12701 = n12060 & n69649 ;
  assign n12702 = n12637 & n12701 ;
  assign n12703 = n12700 | n12702 ;
  assign n12704 = n68438 & n12703 ;
  assign n69677 = ~n12616 ;
  assign n12618 = n12476 & n69677 ;
  assign n12705 = n12077 | n12476 ;
  assign n69678 = ~n12705 ;
  assign n12706 = n12472 & n69678 ;
  assign n12707 = n12618 | n12706 ;
  assign n12708 = n154 & n12707 ;
  assign n12709 = n12068 & n69649 ;
  assign n12710 = n12637 & n12709 ;
  assign n12711 = n12708 | n12710 ;
  assign n12712 = n68214 & n12711 ;
  assign n69679 = ~n12710 ;
  assign n13130 = x95 & n69679 ;
  assign n69680 = ~n12708 ;
  assign n13131 = n69680 & n13130 ;
  assign n13132 = n12712 | n13131 ;
  assign n69681 = ~n12467 ;
  assign n12471 = n69681 & n12470 ;
  assign n12713 = n12085 | n12470 ;
  assign n69682 = ~n12713 ;
  assign n12714 = n12612 & n69682 ;
  assign n12715 = n12471 | n12714 ;
  assign n12716 = n154 & n12715 ;
  assign n12717 = n12076 & n69649 ;
  assign n12718 = n12637 & n12717 ;
  assign n12719 = n12716 | n12718 ;
  assign n12720 = n68058 & n12719 ;
  assign n69683 = ~n12611 ;
  assign n12613 = n12465 & n69683 ;
  assign n12721 = n12093 | n12465 ;
  assign n69684 = ~n12721 ;
  assign n12722 = n12461 & n69684 ;
  assign n12723 = n12613 | n12722 ;
  assign n12724 = n154 & n12723 ;
  assign n12725 = n12084 & n69649 ;
  assign n12726 = n12637 & n12725 ;
  assign n12727 = n12724 | n12726 ;
  assign n12728 = n67986 & n12727 ;
  assign n69685 = ~n12726 ;
  assign n13118 = x93 & n69685 ;
  assign n69686 = ~n12724 ;
  assign n13119 = n69686 & n13118 ;
  assign n13120 = n12728 | n13119 ;
  assign n69687 = ~n12456 ;
  assign n12460 = n69687 & n12459 ;
  assign n12729 = n12101 | n12459 ;
  assign n69688 = ~n12729 ;
  assign n12730 = n12607 & n69688 ;
  assign n12731 = n12460 | n12730 ;
  assign n12732 = n154 & n12731 ;
  assign n12733 = n12092 & n69649 ;
  assign n12734 = n12637 & n12733 ;
  assign n12735 = n12732 | n12734 ;
  assign n12736 = n67763 & n12735 ;
  assign n69689 = ~n12606 ;
  assign n12608 = n12454 & n69689 ;
  assign n12737 = n12109 | n12454 ;
  assign n69690 = ~n12737 ;
  assign n12738 = n12450 & n69690 ;
  assign n12739 = n12608 | n12738 ;
  assign n12740 = n154 & n12739 ;
  assign n12741 = n12100 & n69649 ;
  assign n12742 = n12637 & n12741 ;
  assign n12743 = n12740 | n12742 ;
  assign n12744 = n67622 & n12743 ;
  assign n69691 = ~n12742 ;
  assign n13106 = x91 & n69691 ;
  assign n69692 = ~n12740 ;
  assign n13107 = n69692 & n13106 ;
  assign n13108 = n12744 | n13107 ;
  assign n69693 = ~n12445 ;
  assign n12449 = n69693 & n12448 ;
  assign n12745 = n12117 | n12448 ;
  assign n69694 = ~n12745 ;
  assign n12746 = n12602 & n69694 ;
  assign n12747 = n12449 | n12746 ;
  assign n12748 = n154 & n12747 ;
  assign n12749 = n12108 & n69649 ;
  assign n12750 = n12637 & n12749 ;
  assign n12751 = n12748 | n12750 ;
  assign n12752 = n67531 & n12751 ;
  assign n69695 = ~n12601 ;
  assign n12603 = n12443 & n69695 ;
  assign n12753 = n12125 | n12443 ;
  assign n69696 = ~n12753 ;
  assign n12754 = n12439 & n69696 ;
  assign n12755 = n12603 | n12754 ;
  assign n12756 = n154 & n12755 ;
  assign n12757 = n12116 & n69649 ;
  assign n12758 = n12637 & n12757 ;
  assign n12759 = n12756 | n12758 ;
  assign n12760 = n67348 & n12759 ;
  assign n69697 = ~n12758 ;
  assign n13094 = x89 & n69697 ;
  assign n69698 = ~n12756 ;
  assign n13095 = n69698 & n13094 ;
  assign n13096 = n12760 | n13095 ;
  assign n69699 = ~n12434 ;
  assign n12438 = n69699 & n12437 ;
  assign n12761 = n12133 | n12437 ;
  assign n69700 = ~n12761 ;
  assign n12762 = n12597 & n69700 ;
  assign n12763 = n12438 | n12762 ;
  assign n12764 = n154 & n12763 ;
  assign n12765 = n12124 & n69649 ;
  assign n12766 = n12637 & n12765 ;
  assign n12767 = n12764 | n12766 ;
  assign n12768 = n67222 & n12767 ;
  assign n69701 = ~n12596 ;
  assign n12598 = n12432 & n69701 ;
  assign n12769 = n12141 | n12432 ;
  assign n69702 = ~n12769 ;
  assign n12770 = n12428 & n69702 ;
  assign n12771 = n12598 | n12770 ;
  assign n12772 = n154 & n12771 ;
  assign n12773 = n12132 & n69649 ;
  assign n12774 = n12637 & n12773 ;
  assign n12775 = n12772 | n12774 ;
  assign n12776 = n67164 & n12775 ;
  assign n69703 = ~n12774 ;
  assign n13082 = x87 & n69703 ;
  assign n69704 = ~n12772 ;
  assign n13083 = n69704 & n13082 ;
  assign n13084 = n12776 | n13083 ;
  assign n69705 = ~n12423 ;
  assign n12427 = n69705 & n12426 ;
  assign n12777 = n12149 | n12426 ;
  assign n69706 = ~n12777 ;
  assign n12778 = n12592 & n69706 ;
  assign n12779 = n12427 | n12778 ;
  assign n12780 = n154 & n12779 ;
  assign n12781 = n12140 & n69649 ;
  assign n12782 = n12637 & n12781 ;
  assign n12783 = n12780 | n12782 ;
  assign n12784 = n66979 & n12783 ;
  assign n69707 = ~n12591 ;
  assign n12593 = n12421 & n69707 ;
  assign n12785 = n12157 | n12421 ;
  assign n69708 = ~n12785 ;
  assign n12786 = n12417 & n69708 ;
  assign n12787 = n12593 | n12786 ;
  assign n12788 = n154 & n12787 ;
  assign n12789 = n12148 & n69649 ;
  assign n12790 = n12637 & n12789 ;
  assign n12791 = n12788 | n12790 ;
  assign n12792 = n66868 & n12791 ;
  assign n69709 = ~n12790 ;
  assign n13070 = x85 & n69709 ;
  assign n69710 = ~n12788 ;
  assign n13071 = n69710 & n13070 ;
  assign n13072 = n12792 | n13071 ;
  assign n69711 = ~n12412 ;
  assign n12416 = n69711 & n12415 ;
  assign n12793 = n12165 | n12415 ;
  assign n69712 = ~n12793 ;
  assign n12794 = n12587 & n69712 ;
  assign n12795 = n12416 | n12794 ;
  assign n12796 = n154 & n12795 ;
  assign n12797 = n12156 & n69649 ;
  assign n12798 = n12637 & n12797 ;
  assign n12799 = n12796 | n12798 ;
  assign n12800 = n66797 & n12799 ;
  assign n69713 = ~n12586 ;
  assign n12588 = n12410 & n69713 ;
  assign n12801 = n12173 | n12410 ;
  assign n69714 = ~n12801 ;
  assign n12802 = n12406 & n69714 ;
  assign n12803 = n12588 | n12802 ;
  assign n12804 = n154 & n12803 ;
  assign n12805 = n12164 & n69649 ;
  assign n12806 = n12637 & n12805 ;
  assign n12807 = n12804 | n12806 ;
  assign n12808 = n66654 & n12807 ;
  assign n69715 = ~n12806 ;
  assign n13058 = x83 & n69715 ;
  assign n69716 = ~n12804 ;
  assign n13059 = n69716 & n13058 ;
  assign n13060 = n12808 | n13059 ;
  assign n69717 = ~n12401 ;
  assign n12405 = n69717 & n12404 ;
  assign n12809 = n12181 | n12404 ;
  assign n69718 = ~n12809 ;
  assign n12810 = n12582 & n69718 ;
  assign n12811 = n12405 | n12810 ;
  assign n12812 = n154 & n12811 ;
  assign n12813 = n12172 & n69649 ;
  assign n12814 = n12637 & n12813 ;
  assign n12815 = n12812 | n12814 ;
  assign n12816 = n66560 & n12815 ;
  assign n69719 = ~n12581 ;
  assign n12583 = n12399 & n69719 ;
  assign n12817 = n12189 | n12399 ;
  assign n69720 = ~n12817 ;
  assign n12818 = n12395 & n69720 ;
  assign n12819 = n12583 | n12818 ;
  assign n12820 = n154 & n12819 ;
  assign n12821 = n12180 & n69649 ;
  assign n12822 = n12637 & n12821 ;
  assign n12823 = n12820 | n12822 ;
  assign n12824 = n66505 & n12823 ;
  assign n69721 = ~n12822 ;
  assign n13046 = x81 & n69721 ;
  assign n69722 = ~n12820 ;
  assign n13047 = n69722 & n13046 ;
  assign n13048 = n12824 | n13047 ;
  assign n69723 = ~n12390 ;
  assign n12394 = n69723 & n12393 ;
  assign n12825 = n12197 | n12393 ;
  assign n69724 = ~n12825 ;
  assign n12826 = n12577 & n69724 ;
  assign n12827 = n12394 | n12826 ;
  assign n12828 = n154 & n12827 ;
  assign n12829 = n12188 & n69649 ;
  assign n12830 = n12637 & n12829 ;
  assign n12831 = n12828 | n12830 ;
  assign n12832 = n66379 & n12831 ;
  assign n69725 = ~n12576 ;
  assign n12578 = n12388 & n69725 ;
  assign n12833 = n12205 | n12388 ;
  assign n69726 = ~n12833 ;
  assign n12834 = n12384 & n69726 ;
  assign n12835 = n12578 | n12834 ;
  assign n12836 = n154 & n12835 ;
  assign n12837 = n12196 & n69649 ;
  assign n12838 = n12637 & n12837 ;
  assign n12839 = n12836 | n12838 ;
  assign n12840 = n66299 & n12839 ;
  assign n69727 = ~n12838 ;
  assign n13034 = x79 & n69727 ;
  assign n69728 = ~n12836 ;
  assign n13035 = n69728 & n13034 ;
  assign n13036 = n12840 | n13035 ;
  assign n69729 = ~n12379 ;
  assign n12383 = n69729 & n12382 ;
  assign n12841 = n12213 | n12382 ;
  assign n69730 = ~n12841 ;
  assign n12842 = n12572 & n69730 ;
  assign n12843 = n12383 | n12842 ;
  assign n12844 = n154 & n12843 ;
  assign n12845 = n12204 & n69649 ;
  assign n12846 = n12637 & n12845 ;
  assign n12847 = n12844 | n12846 ;
  assign n12848 = n66244 & n12847 ;
  assign n69731 = ~n12571 ;
  assign n12573 = n12377 & n69731 ;
  assign n12849 = n12221 | n12377 ;
  assign n69732 = ~n12849 ;
  assign n12850 = n12373 & n69732 ;
  assign n12851 = n12573 | n12850 ;
  assign n12852 = n154 & n12851 ;
  assign n12853 = n12212 & n69649 ;
  assign n12854 = n12637 & n12853 ;
  assign n12855 = n12852 | n12854 ;
  assign n12856 = n66145 & n12855 ;
  assign n69733 = ~n12854 ;
  assign n13022 = x77 & n69733 ;
  assign n69734 = ~n12852 ;
  assign n13023 = n69734 & n13022 ;
  assign n13024 = n12856 | n13023 ;
  assign n69735 = ~n12368 ;
  assign n12372 = n69735 & n12371 ;
  assign n12857 = n12229 | n12371 ;
  assign n69736 = ~n12857 ;
  assign n12858 = n12567 & n69736 ;
  assign n12859 = n12372 | n12858 ;
  assign n12860 = n154 & n12859 ;
  assign n12861 = n12220 & n69649 ;
  assign n12862 = n12637 & n12861 ;
  assign n12863 = n12860 | n12862 ;
  assign n12864 = n66081 & n12863 ;
  assign n69737 = ~n12566 ;
  assign n12568 = n12366 & n69737 ;
  assign n12865 = n12237 | n12366 ;
  assign n69738 = ~n12865 ;
  assign n12866 = n12362 & n69738 ;
  assign n12867 = n12568 | n12866 ;
  assign n12868 = n154 & n12867 ;
  assign n12869 = n12228 & n69649 ;
  assign n12870 = n12637 & n12869 ;
  assign n12871 = n12868 | n12870 ;
  assign n12872 = n66043 & n12871 ;
  assign n69739 = ~n12870 ;
  assign n13010 = x75 & n69739 ;
  assign n69740 = ~n12868 ;
  assign n13011 = n69740 & n13010 ;
  assign n13012 = n12872 | n13011 ;
  assign n69741 = ~n12357 ;
  assign n12361 = n69741 & n12360 ;
  assign n12873 = n12245 | n12360 ;
  assign n69742 = ~n12873 ;
  assign n12874 = n12562 & n69742 ;
  assign n12875 = n12361 | n12874 ;
  assign n12876 = n154 & n12875 ;
  assign n12877 = n12236 & n69649 ;
  assign n12878 = n12637 & n12877 ;
  assign n12879 = n12876 | n12878 ;
  assign n12880 = n65960 & n12879 ;
  assign n69743 = ~n12561 ;
  assign n12563 = n12355 & n69743 ;
  assign n12881 = n12253 | n12355 ;
  assign n69744 = ~n12881 ;
  assign n12882 = n12351 & n69744 ;
  assign n12883 = n12563 | n12882 ;
  assign n12884 = n154 & n12883 ;
  assign n12885 = n12244 & n69649 ;
  assign n12886 = n12637 & n12885 ;
  assign n12887 = n12884 | n12886 ;
  assign n12888 = n65909 & n12887 ;
  assign n69745 = ~n12886 ;
  assign n12998 = x73 & n69745 ;
  assign n69746 = ~n12884 ;
  assign n12999 = n69746 & n12998 ;
  assign n13000 = n12888 | n12999 ;
  assign n69747 = ~n12346 ;
  assign n12350 = n69747 & n12349 ;
  assign n12889 = n12262 | n12349 ;
  assign n69748 = ~n12889 ;
  assign n12890 = n12557 & n69748 ;
  assign n12891 = n12350 | n12890 ;
  assign n12892 = n154 & n12891 ;
  assign n12893 = n12252 & n69649 ;
  assign n12894 = n12637 & n12893 ;
  assign n12895 = n12892 | n12894 ;
  assign n12896 = n65877 & n12895 ;
  assign n69749 = ~n12556 ;
  assign n12558 = n12344 & n69749 ;
  assign n12897 = n12271 | n12344 ;
  assign n69750 = ~n12897 ;
  assign n12898 = n12340 & n69750 ;
  assign n12899 = n12558 | n12898 ;
  assign n12900 = n154 & n12899 ;
  assign n12901 = n12261 & n69649 ;
  assign n12902 = n12637 & n12901 ;
  assign n12903 = n12900 | n12902 ;
  assign n12904 = n65820 & n12903 ;
  assign n69751 = ~n12902 ;
  assign n12986 = x71 & n69751 ;
  assign n69752 = ~n12900 ;
  assign n12987 = n69752 & n12986 ;
  assign n12988 = n12904 | n12987 ;
  assign n69753 = ~n12336 ;
  assign n12554 = n69753 & n12339 ;
  assign n12905 = n12280 | n12339 ;
  assign n69754 = ~n12905 ;
  assign n12906 = n12552 & n69754 ;
  assign n12907 = n12554 | n12906 ;
  assign n12908 = n154 & n12907 ;
  assign n12909 = n12270 & n69649 ;
  assign n12910 = n12637 & n12909 ;
  assign n12911 = n12908 | n12910 ;
  assign n12912 = n65791 & n12911 ;
  assign n69755 = ~n12550 ;
  assign n12551 = n12334 & n69755 ;
  assign n12913 = n12327 | n12547 ;
  assign n12914 = n12289 | n12334 ;
  assign n69756 = ~n12914 ;
  assign n12915 = n12913 & n69756 ;
  assign n12916 = n12551 | n12915 ;
  assign n12917 = n154 & n12916 ;
  assign n12918 = n12279 & n69649 ;
  assign n12919 = n12637 & n12918 ;
  assign n12920 = n12917 | n12919 ;
  assign n12921 = n65772 & n12920 ;
  assign n69757 = ~n12919 ;
  assign n12975 = x69 & n69757 ;
  assign n69758 = ~n12917 ;
  assign n12976 = n69758 & n12975 ;
  assign n12977 = n12921 | n12976 ;
  assign n69759 = ~n12327 ;
  assign n12548 = n69759 & n12547 ;
  assign n12922 = n12295 | n12547 ;
  assign n69760 = ~n12922 ;
  assign n12923 = n12326 & n69760 ;
  assign n12924 = n12548 | n12923 ;
  assign n12925 = n154 & n12924 ;
  assign n12926 = n12288 & n69649 ;
  assign n12927 = n12637 & n12926 ;
  assign n12928 = n12925 | n12927 ;
  assign n12929 = n65746 & n12928 ;
  assign n69761 = ~n12543 ;
  assign n12544 = n12325 & n69761 ;
  assign n12930 = n12321 | n12325 ;
  assign n69762 = ~n12930 ;
  assign n12931 = n12320 & n69762 ;
  assign n12932 = n12544 | n12931 ;
  assign n12933 = n154 & n12932 ;
  assign n12934 = n12294 & n69649 ;
  assign n12935 = n12637 & n12934 ;
  assign n12936 = n12933 | n12935 ;
  assign n12937 = n65721 & n12936 ;
  assign n69763 = ~n12935 ;
  assign n12965 = x67 & n69763 ;
  assign n69764 = ~n12933 ;
  assign n12966 = n69764 & n12965 ;
  assign n12967 = n12937 | n12966 ;
  assign n12938 = n12317 & n12319 ;
  assign n12939 = n69535 & n12938 ;
  assign n69765 = ~n12939 ;
  assign n12940 = n12542 & n69765 ;
  assign n12941 = n154 & n12940 ;
  assign n12942 = n12314 & n69649 ;
  assign n12943 = n12637 & n12942 ;
  assign n12944 = n12941 | n12943 ;
  assign n12945 = n65686 & n12944 ;
  assign n69766 = ~x24 ;
  assign n12955 = n69766 & x64 ;
  assign n12538 = n12319 & n154 ;
  assign n12946 = n69649 & n12637 ;
  assign n69767 = ~n12946 ;
  assign n12947 = x64 & n69767 ;
  assign n69768 = ~n12947 ;
  assign n12948 = x25 & n69768 ;
  assign n12949 = n12538 | n12948 ;
  assign n12950 = x65 & n12949 ;
  assign n12537 = x64 & n154 ;
  assign n69769 = ~n12537 ;
  assign n12951 = x25 & n69769 ;
  assign n12952 = n12319 & n69767 ;
  assign n12953 = x65 | n12952 ;
  assign n12954 = n12951 | n12953 ;
  assign n69770 = ~n12950 ;
  assign n12956 = n69770 & n12954 ;
  assign n12957 = n12955 | n12956 ;
  assign n12958 = n12538 | n12951 ;
  assign n12959 = n65670 & n12958 ;
  assign n69771 = ~n12959 ;
  assign n12960 = n12957 & n69771 ;
  assign n69772 = ~n12943 ;
  assign n12961 = x66 & n69772 ;
  assign n69773 = ~n12941 ;
  assign n12962 = n69773 & n12961 ;
  assign n12963 = n12945 | n12962 ;
  assign n12964 = n12960 | n12963 ;
  assign n69774 = ~n12945 ;
  assign n12968 = n69774 & n12964 ;
  assign n12969 = n12967 | n12968 ;
  assign n69775 = ~n12937 ;
  assign n12970 = n69775 & n12969 ;
  assign n69776 = ~n12927 ;
  assign n12971 = x68 & n69776 ;
  assign n69777 = ~n12925 ;
  assign n12972 = n69777 & n12971 ;
  assign n12973 = n12929 | n12972 ;
  assign n12974 = n12970 | n12973 ;
  assign n69778 = ~n12929 ;
  assign n12978 = n69778 & n12974 ;
  assign n12979 = n12977 | n12978 ;
  assign n69779 = ~n12921 ;
  assign n12980 = n69779 & n12979 ;
  assign n69780 = ~n12910 ;
  assign n12981 = x70 & n69780 ;
  assign n69781 = ~n12908 ;
  assign n12982 = n69781 & n12981 ;
  assign n12983 = n12912 | n12982 ;
  assign n12985 = n12980 | n12983 ;
  assign n69782 = ~n12912 ;
  assign n12990 = n69782 & n12985 ;
  assign n12991 = n12988 | n12990 ;
  assign n69783 = ~n12904 ;
  assign n12992 = n69783 & n12991 ;
  assign n69784 = ~n12894 ;
  assign n12993 = x72 & n69784 ;
  assign n69785 = ~n12892 ;
  assign n12994 = n69785 & n12993 ;
  assign n12995 = n12896 | n12994 ;
  assign n12997 = n12992 | n12995 ;
  assign n69786 = ~n12896 ;
  assign n13002 = n69786 & n12997 ;
  assign n13003 = n13000 | n13002 ;
  assign n69787 = ~n12888 ;
  assign n13004 = n69787 & n13003 ;
  assign n69788 = ~n12878 ;
  assign n13005 = x74 & n69788 ;
  assign n69789 = ~n12876 ;
  assign n13006 = n69789 & n13005 ;
  assign n13007 = n12880 | n13006 ;
  assign n13009 = n13004 | n13007 ;
  assign n69790 = ~n12880 ;
  assign n13014 = n69790 & n13009 ;
  assign n13015 = n13012 | n13014 ;
  assign n69791 = ~n12872 ;
  assign n13016 = n69791 & n13015 ;
  assign n69792 = ~n12862 ;
  assign n13017 = x76 & n69792 ;
  assign n69793 = ~n12860 ;
  assign n13018 = n69793 & n13017 ;
  assign n13019 = n12864 | n13018 ;
  assign n13021 = n13016 | n13019 ;
  assign n69794 = ~n12864 ;
  assign n13026 = n69794 & n13021 ;
  assign n13027 = n13024 | n13026 ;
  assign n69795 = ~n12856 ;
  assign n13028 = n69795 & n13027 ;
  assign n69796 = ~n12846 ;
  assign n13029 = x78 & n69796 ;
  assign n69797 = ~n12844 ;
  assign n13030 = n69797 & n13029 ;
  assign n13031 = n12848 | n13030 ;
  assign n13033 = n13028 | n13031 ;
  assign n69798 = ~n12848 ;
  assign n13038 = n69798 & n13033 ;
  assign n13039 = n13036 | n13038 ;
  assign n69799 = ~n12840 ;
  assign n13040 = n69799 & n13039 ;
  assign n69800 = ~n12830 ;
  assign n13041 = x80 & n69800 ;
  assign n69801 = ~n12828 ;
  assign n13042 = n69801 & n13041 ;
  assign n13043 = n12832 | n13042 ;
  assign n13045 = n13040 | n13043 ;
  assign n69802 = ~n12832 ;
  assign n13050 = n69802 & n13045 ;
  assign n13051 = n13048 | n13050 ;
  assign n69803 = ~n12824 ;
  assign n13052 = n69803 & n13051 ;
  assign n69804 = ~n12814 ;
  assign n13053 = x82 & n69804 ;
  assign n69805 = ~n12812 ;
  assign n13054 = n69805 & n13053 ;
  assign n13055 = n12816 | n13054 ;
  assign n13057 = n13052 | n13055 ;
  assign n69806 = ~n12816 ;
  assign n13062 = n69806 & n13057 ;
  assign n13063 = n13060 | n13062 ;
  assign n69807 = ~n12808 ;
  assign n13064 = n69807 & n13063 ;
  assign n69808 = ~n12798 ;
  assign n13065 = x84 & n69808 ;
  assign n69809 = ~n12796 ;
  assign n13066 = n69809 & n13065 ;
  assign n13067 = n12800 | n13066 ;
  assign n13069 = n13064 | n13067 ;
  assign n69810 = ~n12800 ;
  assign n13074 = n69810 & n13069 ;
  assign n13075 = n13072 | n13074 ;
  assign n69811 = ~n12792 ;
  assign n13076 = n69811 & n13075 ;
  assign n69812 = ~n12782 ;
  assign n13077 = x86 & n69812 ;
  assign n69813 = ~n12780 ;
  assign n13078 = n69813 & n13077 ;
  assign n13079 = n12784 | n13078 ;
  assign n13081 = n13076 | n13079 ;
  assign n69814 = ~n12784 ;
  assign n13086 = n69814 & n13081 ;
  assign n13087 = n13084 | n13086 ;
  assign n69815 = ~n12776 ;
  assign n13088 = n69815 & n13087 ;
  assign n69816 = ~n12766 ;
  assign n13089 = x88 & n69816 ;
  assign n69817 = ~n12764 ;
  assign n13090 = n69817 & n13089 ;
  assign n13091 = n12768 | n13090 ;
  assign n13093 = n13088 | n13091 ;
  assign n69818 = ~n12768 ;
  assign n13098 = n69818 & n13093 ;
  assign n13099 = n13096 | n13098 ;
  assign n69819 = ~n12760 ;
  assign n13100 = n69819 & n13099 ;
  assign n69820 = ~n12750 ;
  assign n13101 = x90 & n69820 ;
  assign n69821 = ~n12748 ;
  assign n13102 = n69821 & n13101 ;
  assign n13103 = n12752 | n13102 ;
  assign n13105 = n13100 | n13103 ;
  assign n69822 = ~n12752 ;
  assign n13110 = n69822 & n13105 ;
  assign n13111 = n13108 | n13110 ;
  assign n69823 = ~n12744 ;
  assign n13112 = n69823 & n13111 ;
  assign n69824 = ~n12734 ;
  assign n13113 = x92 & n69824 ;
  assign n69825 = ~n12732 ;
  assign n13114 = n69825 & n13113 ;
  assign n13115 = n12736 | n13114 ;
  assign n13117 = n13112 | n13115 ;
  assign n69826 = ~n12736 ;
  assign n13122 = n69826 & n13117 ;
  assign n13123 = n13120 | n13122 ;
  assign n69827 = ~n12728 ;
  assign n13124 = n69827 & n13123 ;
  assign n69828 = ~n12718 ;
  assign n13125 = x94 & n69828 ;
  assign n69829 = ~n12716 ;
  assign n13126 = n69829 & n13125 ;
  assign n13127 = n12720 | n13126 ;
  assign n13129 = n13124 | n13127 ;
  assign n69830 = ~n12720 ;
  assign n13134 = n69830 & n13129 ;
  assign n13135 = n13132 | n13134 ;
  assign n69831 = ~n12712 ;
  assign n13136 = n69831 & n13135 ;
  assign n69832 = ~n12702 ;
  assign n13137 = x96 & n69832 ;
  assign n69833 = ~n12700 ;
  assign n13138 = n69833 & n13137 ;
  assign n13139 = n12704 | n13138 ;
  assign n13141 = n13136 | n13139 ;
  assign n69834 = ~n12704 ;
  assign n13146 = n69834 & n13141 ;
  assign n13147 = n13144 | n13146 ;
  assign n69835 = ~n12696 ;
  assign n13148 = n69835 & n13147 ;
  assign n69836 = ~n12686 ;
  assign n13149 = x98 & n69836 ;
  assign n69837 = ~n12684 ;
  assign n13150 = n69837 & n13149 ;
  assign n13151 = n12688 | n13150 ;
  assign n13153 = n13148 | n13151 ;
  assign n69838 = ~n12688 ;
  assign n13158 = n69838 & n13153 ;
  assign n13159 = n13156 | n13158 ;
  assign n69839 = ~n12680 ;
  assign n13160 = n69839 & n13159 ;
  assign n69840 = ~n12670 ;
  assign n13161 = x100 & n69840 ;
  assign n69841 = ~n12668 ;
  assign n13162 = n69841 & n13161 ;
  assign n13163 = n12672 | n13162 ;
  assign n13165 = n13160 | n13163 ;
  assign n69842 = ~n12672 ;
  assign n13170 = n69842 & n13165 ;
  assign n13171 = n13168 | n13170 ;
  assign n69843 = ~n12664 ;
  assign n13172 = n69843 & n13171 ;
  assign n69844 = ~n12654 ;
  assign n13173 = x102 & n69844 ;
  assign n69845 = ~n12652 ;
  assign n13174 = n69845 & n13173 ;
  assign n13175 = n12656 | n13174 ;
  assign n13177 = n13172 | n13175 ;
  assign n69846 = ~n12656 ;
  assign n13181 = n69846 & n13177 ;
  assign n13182 = n13180 | n13181 ;
  assign n69847 = ~n12648 ;
  assign n13183 = n69847 & n13182 ;
  assign n13184 = n66858 | n67093 ;
  assign n13185 = n13183 | n13184 ;
  assign n13276 = n12655 & n13185 ;
  assign n13176 = n12664 | n13175 ;
  assign n13189 = x65 & n12958 ;
  assign n69848 = ~n13189 ;
  assign n13190 = n12954 & n69848 ;
  assign n13192 = n12955 | n13190 ;
  assign n13194 = n69771 & n13192 ;
  assign n13195 = n12963 | n13194 ;
  assign n13196 = n69774 & n13195 ;
  assign n13197 = n12967 | n13196 ;
  assign n13198 = n69775 & n13197 ;
  assign n13199 = n12973 | n13198 ;
  assign n13200 = n69778 & n13199 ;
  assign n13201 = n12977 | n13200 ;
  assign n13202 = n69779 & n13201 ;
  assign n13203 = n12983 | n13202 ;
  assign n13204 = n69782 & n13203 ;
  assign n13205 = n12988 | n13204 ;
  assign n13206 = n69783 & n13205 ;
  assign n13207 = n12995 | n13206 ;
  assign n13208 = n69786 & n13207 ;
  assign n13209 = n13000 | n13208 ;
  assign n13210 = n69787 & n13209 ;
  assign n13211 = n13007 | n13210 ;
  assign n13212 = n69790 & n13211 ;
  assign n13213 = n13012 | n13212 ;
  assign n13214 = n69791 & n13213 ;
  assign n13215 = n13019 | n13214 ;
  assign n13216 = n69794 & n13215 ;
  assign n13217 = n13024 | n13216 ;
  assign n13218 = n69795 & n13217 ;
  assign n13219 = n13031 | n13218 ;
  assign n13220 = n69798 & n13219 ;
  assign n13221 = n13036 | n13220 ;
  assign n13222 = n69799 & n13221 ;
  assign n13223 = n13043 | n13222 ;
  assign n13224 = n69802 & n13223 ;
  assign n13225 = n13048 | n13224 ;
  assign n13226 = n69803 & n13225 ;
  assign n13227 = n13055 | n13226 ;
  assign n13228 = n69806 & n13227 ;
  assign n13229 = n13060 | n13228 ;
  assign n13230 = n69807 & n13229 ;
  assign n13231 = n13067 | n13230 ;
  assign n13232 = n69810 & n13231 ;
  assign n13233 = n13072 | n13232 ;
  assign n13234 = n69811 & n13233 ;
  assign n13235 = n13079 | n13234 ;
  assign n13236 = n69814 & n13235 ;
  assign n13237 = n13084 | n13236 ;
  assign n13238 = n69815 & n13237 ;
  assign n13239 = n13091 | n13238 ;
  assign n13240 = n69818 & n13239 ;
  assign n13241 = n13096 | n13240 ;
  assign n13242 = n69819 & n13241 ;
  assign n13243 = n13103 | n13242 ;
  assign n13244 = n69822 & n13243 ;
  assign n13245 = n13108 | n13244 ;
  assign n13246 = n69823 & n13245 ;
  assign n13247 = n13115 | n13246 ;
  assign n13248 = n69826 & n13247 ;
  assign n13249 = n13120 | n13248 ;
  assign n13250 = n69827 & n13249 ;
  assign n13251 = n13127 | n13250 ;
  assign n13252 = n69830 & n13251 ;
  assign n13253 = n13132 | n13252 ;
  assign n13254 = n69831 & n13253 ;
  assign n13255 = n13139 | n13254 ;
  assign n13256 = n69834 & n13255 ;
  assign n13257 = n13144 | n13256 ;
  assign n13258 = n69835 & n13257 ;
  assign n13259 = n13151 | n13258 ;
  assign n13260 = n69838 & n13259 ;
  assign n13261 = n13156 | n13260 ;
  assign n13262 = n69839 & n13261 ;
  assign n13263 = n13163 | n13262 ;
  assign n13264 = n69842 & n13263 ;
  assign n13265 = n13168 | n13264 ;
  assign n69849 = ~n13176 ;
  assign n13277 = n69849 & n13265 ;
  assign n13266 = n69843 & n13265 ;
  assign n69850 = ~n13266 ;
  assign n13278 = n13175 & n69850 ;
  assign n13279 = n13277 | n13278 ;
  assign n69851 = ~n13184 ;
  assign n13280 = n69851 & n13279 ;
  assign n69852 = ~n13183 ;
  assign n13281 = n69852 & n13280 ;
  assign n13282 = n13276 | n13281 ;
  assign n69853 = ~n12647 ;
  assign n13186 = n69853 & n13185 ;
  assign n69854 = ~n13181 ;
  assign n13269 = n13180 & n69854 ;
  assign n13267 = n13175 | n13266 ;
  assign n13270 = n12656 | n13180 ;
  assign n69855 = ~n13270 ;
  assign n13271 = n13267 & n69855 ;
  assign n13272 = n13269 | n13271 ;
  assign n13273 = n13185 | n13272 ;
  assign n69856 = ~n13186 ;
  assign n13274 = n69856 & n13273 ;
  assign n69857 = ~x104 ;
  assign n13275 = n69857 & n13274 ;
  assign n13283 = n69656 & n13282 ;
  assign n13284 = n12663 & n13185 ;
  assign n13169 = n12672 | n13168 ;
  assign n69858 = ~n13169 ;
  assign n13285 = n13165 & n69858 ;
  assign n69859 = ~n13170 ;
  assign n13286 = n13168 & n69859 ;
  assign n13287 = n13285 | n13286 ;
  assign n13288 = n69851 & n13287 ;
  assign n13289 = n69852 & n13288 ;
  assign n13290 = n13284 | n13289 ;
  assign n13291 = n69528 & n13290 ;
  assign n13292 = n12671 & n13185 ;
  assign n13164 = n12680 | n13163 ;
  assign n69860 = ~n13164 ;
  assign n13293 = n69860 & n13261 ;
  assign n69861 = ~n13262 ;
  assign n13294 = n13163 & n69861 ;
  assign n13295 = n13293 | n13294 ;
  assign n13296 = n69851 & n13295 ;
  assign n13297 = n69852 & n13296 ;
  assign n13298 = n13292 | n13297 ;
  assign n13299 = n69261 & n13298 ;
  assign n13300 = n12679 & n13185 ;
  assign n13157 = n12688 | n13156 ;
  assign n69862 = ~n13157 ;
  assign n13301 = n13153 & n69862 ;
  assign n69863 = ~n13158 ;
  assign n13302 = n13156 & n69863 ;
  assign n13303 = n13301 | n13302 ;
  assign n13304 = n69851 & n13303 ;
  assign n13305 = n69852 & n13304 ;
  assign n13306 = n13300 | n13305 ;
  assign n13307 = n69075 & n13306 ;
  assign n13308 = n12687 & n13185 ;
  assign n13152 = n12696 | n13151 ;
  assign n69864 = ~n13152 ;
  assign n13309 = n69864 & n13257 ;
  assign n69865 = ~n13258 ;
  assign n13310 = n13151 & n69865 ;
  assign n13311 = n13309 | n13310 ;
  assign n13312 = n69851 & n13311 ;
  assign n13313 = n69852 & n13312 ;
  assign n13314 = n13308 | n13313 ;
  assign n13315 = n68993 & n13314 ;
  assign n13316 = n12695 & n13185 ;
  assign n13145 = n12704 | n13144 ;
  assign n69866 = ~n13145 ;
  assign n13317 = n13141 & n69866 ;
  assign n69867 = ~n13146 ;
  assign n13318 = n13144 & n69867 ;
  assign n13319 = n13317 | n13318 ;
  assign n13320 = n69851 & n13319 ;
  assign n13321 = n69852 & n13320 ;
  assign n13322 = n13316 | n13321 ;
  assign n13323 = n68716 & n13322 ;
  assign n13324 = n12703 & n13185 ;
  assign n13140 = n12712 | n13139 ;
  assign n69868 = ~n13140 ;
  assign n13325 = n69868 & n13253 ;
  assign n69869 = ~n13254 ;
  assign n13326 = n13139 & n69869 ;
  assign n13327 = n13325 | n13326 ;
  assign n13328 = n69851 & n13327 ;
  assign n13329 = n69852 & n13328 ;
  assign n13330 = n13324 | n13329 ;
  assign n13331 = n68545 & n13330 ;
  assign n13332 = n12711 & n13185 ;
  assign n13133 = n12720 | n13132 ;
  assign n69870 = ~n13133 ;
  assign n13333 = n13129 & n69870 ;
  assign n69871 = ~n13134 ;
  assign n13334 = n13132 & n69871 ;
  assign n13335 = n13333 | n13334 ;
  assign n13336 = n69851 & n13335 ;
  assign n13337 = n69852 & n13336 ;
  assign n13338 = n13332 | n13337 ;
  assign n13339 = n68438 & n13338 ;
  assign n13340 = n12719 & n13185 ;
  assign n13128 = n12728 | n13127 ;
  assign n69872 = ~n13128 ;
  assign n13341 = n69872 & n13249 ;
  assign n69873 = ~n13250 ;
  assign n13342 = n13127 & n69873 ;
  assign n13343 = n13341 | n13342 ;
  assign n13344 = n69851 & n13343 ;
  assign n13345 = n69852 & n13344 ;
  assign n13346 = n13340 | n13345 ;
  assign n13347 = n68214 & n13346 ;
  assign n13348 = n12727 & n13185 ;
  assign n13121 = n12736 | n13120 ;
  assign n69874 = ~n13121 ;
  assign n13349 = n13117 & n69874 ;
  assign n69875 = ~n13122 ;
  assign n13350 = n13120 & n69875 ;
  assign n13351 = n13349 | n13350 ;
  assign n13352 = n69851 & n13351 ;
  assign n13353 = n69852 & n13352 ;
  assign n13354 = n13348 | n13353 ;
  assign n13355 = n68058 & n13354 ;
  assign n13356 = n12735 & n13185 ;
  assign n13116 = n12744 | n13115 ;
  assign n69876 = ~n13116 ;
  assign n13357 = n69876 & n13245 ;
  assign n69877 = ~n13246 ;
  assign n13358 = n13115 & n69877 ;
  assign n13359 = n13357 | n13358 ;
  assign n13360 = n69851 & n13359 ;
  assign n13361 = n69852 & n13360 ;
  assign n13362 = n13356 | n13361 ;
  assign n13363 = n67986 & n13362 ;
  assign n13364 = n12743 & n13185 ;
  assign n13109 = n12752 | n13108 ;
  assign n69878 = ~n13109 ;
  assign n13365 = n13105 & n69878 ;
  assign n69879 = ~n13110 ;
  assign n13366 = n13108 & n69879 ;
  assign n13367 = n13365 | n13366 ;
  assign n13368 = n69851 & n13367 ;
  assign n13369 = n69852 & n13368 ;
  assign n13370 = n13364 | n13369 ;
  assign n13371 = n67763 & n13370 ;
  assign n13372 = n12751 & n13185 ;
  assign n13104 = n12760 | n13103 ;
  assign n69880 = ~n13104 ;
  assign n13373 = n69880 & n13241 ;
  assign n69881 = ~n13242 ;
  assign n13374 = n13103 & n69881 ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = n69851 & n13375 ;
  assign n13377 = n69852 & n13376 ;
  assign n13378 = n13372 | n13377 ;
  assign n13379 = n67622 & n13378 ;
  assign n13380 = n12759 & n13185 ;
  assign n13097 = n12768 | n13096 ;
  assign n69882 = ~n13097 ;
  assign n13381 = n13093 & n69882 ;
  assign n69883 = ~n13098 ;
  assign n13382 = n13096 & n69883 ;
  assign n13383 = n13381 | n13382 ;
  assign n13384 = n69851 & n13383 ;
  assign n13385 = n69852 & n13384 ;
  assign n13386 = n13380 | n13385 ;
  assign n13387 = n67531 & n13386 ;
  assign n13388 = n12767 & n13185 ;
  assign n13092 = n12776 | n13091 ;
  assign n69884 = ~n13092 ;
  assign n13389 = n69884 & n13237 ;
  assign n69885 = ~n13238 ;
  assign n13390 = n13091 & n69885 ;
  assign n13391 = n13389 | n13390 ;
  assign n13392 = n69851 & n13391 ;
  assign n13393 = n69852 & n13392 ;
  assign n13394 = n13388 | n13393 ;
  assign n13395 = n67348 & n13394 ;
  assign n13396 = n12775 & n13185 ;
  assign n13085 = n12784 | n13084 ;
  assign n69886 = ~n13085 ;
  assign n13397 = n13081 & n69886 ;
  assign n69887 = ~n13086 ;
  assign n13398 = n13084 & n69887 ;
  assign n13399 = n13397 | n13398 ;
  assign n13400 = n69851 & n13399 ;
  assign n13401 = n69852 & n13400 ;
  assign n13402 = n13396 | n13401 ;
  assign n13403 = n67222 & n13402 ;
  assign n13404 = n12783 & n13185 ;
  assign n13080 = n12792 | n13079 ;
  assign n69888 = ~n13080 ;
  assign n13405 = n69888 & n13233 ;
  assign n69889 = ~n13234 ;
  assign n13406 = n13079 & n69889 ;
  assign n13407 = n13405 | n13406 ;
  assign n13408 = n69851 & n13407 ;
  assign n13409 = n69852 & n13408 ;
  assign n13410 = n13404 | n13409 ;
  assign n13411 = n67164 & n13410 ;
  assign n13412 = n12791 & n13185 ;
  assign n13073 = n12800 | n13072 ;
  assign n69890 = ~n13073 ;
  assign n13413 = n13069 & n69890 ;
  assign n69891 = ~n13074 ;
  assign n13414 = n13072 & n69891 ;
  assign n13415 = n13413 | n13414 ;
  assign n13416 = n69851 & n13415 ;
  assign n13417 = n69852 & n13416 ;
  assign n13418 = n13412 | n13417 ;
  assign n13419 = n66979 & n13418 ;
  assign n13420 = n12799 & n13185 ;
  assign n13068 = n12808 | n13067 ;
  assign n69892 = ~n13068 ;
  assign n13421 = n69892 & n13229 ;
  assign n69893 = ~n13230 ;
  assign n13422 = n13067 & n69893 ;
  assign n13423 = n13421 | n13422 ;
  assign n13424 = n69851 & n13423 ;
  assign n13425 = n69852 & n13424 ;
  assign n13426 = n13420 | n13425 ;
  assign n13427 = n66868 & n13426 ;
  assign n13428 = n12807 & n13185 ;
  assign n13061 = n12816 | n13060 ;
  assign n69894 = ~n13061 ;
  assign n13429 = n13057 & n69894 ;
  assign n69895 = ~n13062 ;
  assign n13430 = n13060 & n69895 ;
  assign n13431 = n13429 | n13430 ;
  assign n13432 = n69851 & n13431 ;
  assign n13433 = n69852 & n13432 ;
  assign n13434 = n13428 | n13433 ;
  assign n13435 = n66797 & n13434 ;
  assign n13436 = n12815 & n13185 ;
  assign n13056 = n12824 | n13055 ;
  assign n69896 = ~n13056 ;
  assign n13437 = n69896 & n13225 ;
  assign n69897 = ~n13226 ;
  assign n13438 = n13055 & n69897 ;
  assign n13439 = n13437 | n13438 ;
  assign n13440 = n69851 & n13439 ;
  assign n13441 = n69852 & n13440 ;
  assign n13442 = n13436 | n13441 ;
  assign n13443 = n66654 & n13442 ;
  assign n13444 = n12823 & n13185 ;
  assign n13049 = n12832 | n13048 ;
  assign n69898 = ~n13049 ;
  assign n13445 = n13045 & n69898 ;
  assign n69899 = ~n13050 ;
  assign n13446 = n13048 & n69899 ;
  assign n13447 = n13445 | n13446 ;
  assign n13448 = n69851 & n13447 ;
  assign n13449 = n69852 & n13448 ;
  assign n13450 = n13444 | n13449 ;
  assign n13451 = n66560 & n13450 ;
  assign n13452 = n12831 & n13185 ;
  assign n13044 = n12840 | n13043 ;
  assign n69900 = ~n13044 ;
  assign n13453 = n69900 & n13221 ;
  assign n69901 = ~n13222 ;
  assign n13454 = n13043 & n69901 ;
  assign n13455 = n13453 | n13454 ;
  assign n13456 = n69851 & n13455 ;
  assign n13457 = n69852 & n13456 ;
  assign n13458 = n13452 | n13457 ;
  assign n13459 = n66505 & n13458 ;
  assign n13460 = n12839 & n13185 ;
  assign n13037 = n12848 | n13036 ;
  assign n69902 = ~n13037 ;
  assign n13461 = n13033 & n69902 ;
  assign n69903 = ~n13038 ;
  assign n13462 = n13036 & n69903 ;
  assign n13463 = n13461 | n13462 ;
  assign n13464 = n69851 & n13463 ;
  assign n13465 = n69852 & n13464 ;
  assign n13466 = n13460 | n13465 ;
  assign n13467 = n66379 & n13466 ;
  assign n13468 = n12847 & n13185 ;
  assign n13032 = n12856 | n13031 ;
  assign n69904 = ~n13032 ;
  assign n13469 = n69904 & n13217 ;
  assign n69905 = ~n13218 ;
  assign n13470 = n13031 & n69905 ;
  assign n13471 = n13469 | n13470 ;
  assign n13472 = n69851 & n13471 ;
  assign n13473 = n69852 & n13472 ;
  assign n13474 = n13468 | n13473 ;
  assign n13475 = n66299 & n13474 ;
  assign n13476 = n12855 & n13185 ;
  assign n13025 = n12864 | n13024 ;
  assign n69906 = ~n13025 ;
  assign n13477 = n13021 & n69906 ;
  assign n69907 = ~n13026 ;
  assign n13478 = n13024 & n69907 ;
  assign n13479 = n13477 | n13478 ;
  assign n13480 = n69851 & n13479 ;
  assign n13481 = n69852 & n13480 ;
  assign n13482 = n13476 | n13481 ;
  assign n13483 = n66244 & n13482 ;
  assign n13484 = n12863 & n13185 ;
  assign n13020 = n12872 | n13019 ;
  assign n69908 = ~n13020 ;
  assign n13485 = n69908 & n13213 ;
  assign n69909 = ~n13214 ;
  assign n13486 = n13019 & n69909 ;
  assign n13487 = n13485 | n13486 ;
  assign n13488 = n69851 & n13487 ;
  assign n13489 = n69852 & n13488 ;
  assign n13490 = n13484 | n13489 ;
  assign n13491 = n66145 & n13490 ;
  assign n13492 = n12871 & n13185 ;
  assign n13013 = n12880 | n13012 ;
  assign n69910 = ~n13013 ;
  assign n13493 = n13009 & n69910 ;
  assign n69911 = ~n13014 ;
  assign n13494 = n13012 & n69911 ;
  assign n13495 = n13493 | n13494 ;
  assign n13496 = n69851 & n13495 ;
  assign n13497 = n69852 & n13496 ;
  assign n13498 = n13492 | n13497 ;
  assign n13499 = n66081 & n13498 ;
  assign n13500 = n12879 & n13185 ;
  assign n13008 = n12888 | n13007 ;
  assign n69912 = ~n13008 ;
  assign n13501 = n69912 & n13209 ;
  assign n69913 = ~n13210 ;
  assign n13502 = n13007 & n69913 ;
  assign n13503 = n13501 | n13502 ;
  assign n13504 = n69851 & n13503 ;
  assign n13505 = n69852 & n13504 ;
  assign n13506 = n13500 | n13505 ;
  assign n13507 = n66043 & n13506 ;
  assign n13508 = n12887 & n13185 ;
  assign n13001 = n12896 | n13000 ;
  assign n69914 = ~n13001 ;
  assign n13509 = n12997 & n69914 ;
  assign n69915 = ~n13002 ;
  assign n13510 = n13000 & n69915 ;
  assign n13511 = n13509 | n13510 ;
  assign n13512 = n69851 & n13511 ;
  assign n13513 = n69852 & n13512 ;
  assign n13514 = n13508 | n13513 ;
  assign n13515 = n65960 & n13514 ;
  assign n13516 = n12895 & n13185 ;
  assign n12996 = n12904 | n12995 ;
  assign n69916 = ~n12996 ;
  assign n13517 = n69916 & n13205 ;
  assign n69917 = ~n13206 ;
  assign n13518 = n12995 & n69917 ;
  assign n13519 = n13517 | n13518 ;
  assign n13520 = n69851 & n13519 ;
  assign n13521 = n69852 & n13520 ;
  assign n13522 = n13516 | n13521 ;
  assign n13523 = n65909 & n13522 ;
  assign n13524 = n12903 & n13185 ;
  assign n12989 = n12912 | n12988 ;
  assign n69918 = ~n12989 ;
  assign n13525 = n12985 & n69918 ;
  assign n69919 = ~n12990 ;
  assign n13526 = n12988 & n69919 ;
  assign n13527 = n13525 | n13526 ;
  assign n13528 = n69851 & n13527 ;
  assign n13529 = n69852 & n13528 ;
  assign n13530 = n13524 | n13529 ;
  assign n13531 = n65877 & n13530 ;
  assign n13532 = n12911 & n13185 ;
  assign n12984 = n12921 | n12983 ;
  assign n69920 = ~n12984 ;
  assign n13533 = n69920 & n13201 ;
  assign n69921 = ~n13202 ;
  assign n13534 = n12983 & n69921 ;
  assign n13535 = n13533 | n13534 ;
  assign n13536 = n69851 & n13535 ;
  assign n13537 = n69852 & n13536 ;
  assign n13538 = n13532 | n13537 ;
  assign n13539 = n65820 & n13538 ;
  assign n13540 = n12920 & n13185 ;
  assign n13188 = n12929 | n12977 ;
  assign n69922 = ~n13188 ;
  assign n13541 = n12974 & n69922 ;
  assign n69923 = ~n12978 ;
  assign n13542 = n12977 & n69923 ;
  assign n13543 = n13541 | n13542 ;
  assign n13544 = n69851 & n13543 ;
  assign n13545 = n69852 & n13544 ;
  assign n13546 = n13540 | n13545 ;
  assign n13547 = n65791 & n13546 ;
  assign n13548 = n12928 & n13185 ;
  assign n13549 = n12937 | n12973 ;
  assign n69924 = ~n13549 ;
  assign n13550 = n13197 & n69924 ;
  assign n69925 = ~n13198 ;
  assign n13551 = n12973 & n69925 ;
  assign n13552 = n13550 | n13551 ;
  assign n13553 = n69851 & n13552 ;
  assign n13554 = n69852 & n13553 ;
  assign n13555 = n13548 | n13554 ;
  assign n13556 = n65772 & n13555 ;
  assign n13557 = n12936 & n13185 ;
  assign n13558 = n12945 | n12967 ;
  assign n69926 = ~n13558 ;
  assign n13559 = n13195 & n69926 ;
  assign n69927 = ~n12968 ;
  assign n13560 = n12967 & n69927 ;
  assign n13561 = n13559 | n13560 ;
  assign n13562 = n69851 & n13561 ;
  assign n13563 = n69852 & n13562 ;
  assign n13564 = n13557 | n13563 ;
  assign n13565 = n65746 & n13564 ;
  assign n13566 = n12944 & n13185 ;
  assign n13193 = n12959 | n12963 ;
  assign n69928 = ~n13193 ;
  assign n13567 = n12957 & n69928 ;
  assign n69929 = ~n13194 ;
  assign n13568 = n12963 & n69929 ;
  assign n13569 = n13567 | n13568 ;
  assign n13570 = n69851 & n13569 ;
  assign n13571 = n69852 & n13570 ;
  assign n13572 = n13566 | n13571 ;
  assign n13573 = n65721 & n13572 ;
  assign n13187 = n12958 & n13185 ;
  assign n13191 = n12954 & n12955 ;
  assign n13574 = n69770 & n13191 ;
  assign n13575 = n13184 | n13574 ;
  assign n69930 = ~n13575 ;
  assign n13576 = n12957 & n69930 ;
  assign n13577 = n69852 & n13576 ;
  assign n13578 = n13187 | n13577 ;
  assign n13579 = n65686 & n13578 ;
  assign n13586 = n69371 & n12955 ;
  assign n13587 = n69372 & n13586 ;
  assign n13588 = n67021 & n13587 ;
  assign n13589 = n69852 & n13588 ;
  assign n13580 = x64 & n69857 ;
  assign n13581 = n69530 & n13580 ;
  assign n13582 = n69531 & n13581 ;
  assign n13583 = n67026 & n13582 ;
  assign n13268 = n69846 & n13267 ;
  assign n13597 = n13180 | n13268 ;
  assign n13598 = n69847 & n13597 ;
  assign n69931 = ~n13598 ;
  assign n13599 = n13583 & n69931 ;
  assign n69932 = ~n13599 ;
  assign n13600 = x24 & n69932 ;
  assign n13601 = n13589 | n13600 ;
  assign n13602 = n65670 & n13601 ;
  assign n13584 = n69852 & n13583 ;
  assign n69933 = ~n13584 ;
  assign n13585 = x24 & n69933 ;
  assign n13590 = n13585 | n13589 ;
  assign n13591 = x65 & n13590 ;
  assign n13593 = x65 | n13589 ;
  assign n13594 = n13585 | n13593 ;
  assign n69934 = ~n13591 ;
  assign n13595 = n69934 & n13594 ;
  assign n69935 = ~x23 ;
  assign n13596 = n69935 & x64 ;
  assign n13603 = n13595 | n13596 ;
  assign n69936 = ~n13602 ;
  assign n13604 = n69936 & n13603 ;
  assign n69937 = ~n13577 ;
  assign n13605 = x66 & n69937 ;
  assign n69938 = ~n13187 ;
  assign n13606 = n69938 & n13605 ;
  assign n13607 = n13579 | n13606 ;
  assign n13608 = n13604 | n13607 ;
  assign n69939 = ~n13579 ;
  assign n13609 = n69939 & n13608 ;
  assign n69940 = ~n13571 ;
  assign n13610 = x67 & n69940 ;
  assign n69941 = ~n13566 ;
  assign n13611 = n69941 & n13610 ;
  assign n13612 = n13573 | n13611 ;
  assign n13613 = n13609 | n13612 ;
  assign n69942 = ~n13573 ;
  assign n13614 = n69942 & n13613 ;
  assign n69943 = ~n13563 ;
  assign n13615 = x68 & n69943 ;
  assign n69944 = ~n13557 ;
  assign n13616 = n69944 & n13615 ;
  assign n13617 = n13565 | n13616 ;
  assign n13618 = n13614 | n13617 ;
  assign n69945 = ~n13565 ;
  assign n13619 = n69945 & n13618 ;
  assign n69946 = ~n13554 ;
  assign n13620 = x69 & n69946 ;
  assign n69947 = ~n13548 ;
  assign n13621 = n69947 & n13620 ;
  assign n13622 = n13556 | n13621 ;
  assign n13623 = n13619 | n13622 ;
  assign n69948 = ~n13556 ;
  assign n13624 = n69948 & n13623 ;
  assign n69949 = ~n13545 ;
  assign n13625 = x70 & n69949 ;
  assign n69950 = ~n13540 ;
  assign n13626 = n69950 & n13625 ;
  assign n13627 = n13547 | n13626 ;
  assign n13629 = n13624 | n13627 ;
  assign n69951 = ~n13547 ;
  assign n13630 = n69951 & n13629 ;
  assign n69952 = ~n13537 ;
  assign n13631 = x71 & n69952 ;
  assign n69953 = ~n13532 ;
  assign n13632 = n69953 & n13631 ;
  assign n13633 = n13539 | n13632 ;
  assign n13634 = n13630 | n13633 ;
  assign n69954 = ~n13539 ;
  assign n13635 = n69954 & n13634 ;
  assign n69955 = ~n13529 ;
  assign n13636 = x72 & n69955 ;
  assign n69956 = ~n13524 ;
  assign n13637 = n69956 & n13636 ;
  assign n13638 = n13531 | n13637 ;
  assign n13640 = n13635 | n13638 ;
  assign n69957 = ~n13531 ;
  assign n13641 = n69957 & n13640 ;
  assign n69958 = ~n13521 ;
  assign n13642 = x73 & n69958 ;
  assign n69959 = ~n13516 ;
  assign n13643 = n69959 & n13642 ;
  assign n13644 = n13523 | n13643 ;
  assign n13645 = n13641 | n13644 ;
  assign n69960 = ~n13523 ;
  assign n13646 = n69960 & n13645 ;
  assign n69961 = ~n13513 ;
  assign n13647 = x74 & n69961 ;
  assign n69962 = ~n13508 ;
  assign n13648 = n69962 & n13647 ;
  assign n13649 = n13515 | n13648 ;
  assign n13651 = n13646 | n13649 ;
  assign n69963 = ~n13515 ;
  assign n13652 = n69963 & n13651 ;
  assign n69964 = ~n13505 ;
  assign n13653 = x75 & n69964 ;
  assign n69965 = ~n13500 ;
  assign n13654 = n69965 & n13653 ;
  assign n13655 = n13507 | n13654 ;
  assign n13656 = n13652 | n13655 ;
  assign n69966 = ~n13507 ;
  assign n13657 = n69966 & n13656 ;
  assign n69967 = ~n13497 ;
  assign n13658 = x76 & n69967 ;
  assign n69968 = ~n13492 ;
  assign n13659 = n69968 & n13658 ;
  assign n13660 = n13499 | n13659 ;
  assign n13662 = n13657 | n13660 ;
  assign n69969 = ~n13499 ;
  assign n13663 = n69969 & n13662 ;
  assign n69970 = ~n13489 ;
  assign n13664 = x77 & n69970 ;
  assign n69971 = ~n13484 ;
  assign n13665 = n69971 & n13664 ;
  assign n13666 = n13491 | n13665 ;
  assign n13667 = n13663 | n13666 ;
  assign n69972 = ~n13491 ;
  assign n13668 = n69972 & n13667 ;
  assign n69973 = ~n13481 ;
  assign n13669 = x78 & n69973 ;
  assign n69974 = ~n13476 ;
  assign n13670 = n69974 & n13669 ;
  assign n13671 = n13483 | n13670 ;
  assign n13673 = n13668 | n13671 ;
  assign n69975 = ~n13483 ;
  assign n13674 = n69975 & n13673 ;
  assign n69976 = ~n13473 ;
  assign n13675 = x79 & n69976 ;
  assign n69977 = ~n13468 ;
  assign n13676 = n69977 & n13675 ;
  assign n13677 = n13475 | n13676 ;
  assign n13678 = n13674 | n13677 ;
  assign n69978 = ~n13475 ;
  assign n13679 = n69978 & n13678 ;
  assign n69979 = ~n13465 ;
  assign n13680 = x80 & n69979 ;
  assign n69980 = ~n13460 ;
  assign n13681 = n69980 & n13680 ;
  assign n13682 = n13467 | n13681 ;
  assign n13684 = n13679 | n13682 ;
  assign n69981 = ~n13467 ;
  assign n13685 = n69981 & n13684 ;
  assign n69982 = ~n13457 ;
  assign n13686 = x81 & n69982 ;
  assign n69983 = ~n13452 ;
  assign n13687 = n69983 & n13686 ;
  assign n13688 = n13459 | n13687 ;
  assign n13689 = n13685 | n13688 ;
  assign n69984 = ~n13459 ;
  assign n13690 = n69984 & n13689 ;
  assign n69985 = ~n13449 ;
  assign n13691 = x82 & n69985 ;
  assign n69986 = ~n13444 ;
  assign n13692 = n69986 & n13691 ;
  assign n13693 = n13451 | n13692 ;
  assign n13695 = n13690 | n13693 ;
  assign n69987 = ~n13451 ;
  assign n13696 = n69987 & n13695 ;
  assign n69988 = ~n13441 ;
  assign n13697 = x83 & n69988 ;
  assign n69989 = ~n13436 ;
  assign n13698 = n69989 & n13697 ;
  assign n13699 = n13443 | n13698 ;
  assign n13700 = n13696 | n13699 ;
  assign n69990 = ~n13443 ;
  assign n13701 = n69990 & n13700 ;
  assign n69991 = ~n13433 ;
  assign n13702 = x84 & n69991 ;
  assign n69992 = ~n13428 ;
  assign n13703 = n69992 & n13702 ;
  assign n13704 = n13435 | n13703 ;
  assign n13706 = n13701 | n13704 ;
  assign n69993 = ~n13435 ;
  assign n13707 = n69993 & n13706 ;
  assign n69994 = ~n13425 ;
  assign n13708 = x85 & n69994 ;
  assign n69995 = ~n13420 ;
  assign n13709 = n69995 & n13708 ;
  assign n13710 = n13427 | n13709 ;
  assign n13711 = n13707 | n13710 ;
  assign n69996 = ~n13427 ;
  assign n13712 = n69996 & n13711 ;
  assign n69997 = ~n13417 ;
  assign n13713 = x86 & n69997 ;
  assign n69998 = ~n13412 ;
  assign n13714 = n69998 & n13713 ;
  assign n13715 = n13419 | n13714 ;
  assign n13717 = n13712 | n13715 ;
  assign n69999 = ~n13419 ;
  assign n13718 = n69999 & n13717 ;
  assign n70000 = ~n13409 ;
  assign n13719 = x87 & n70000 ;
  assign n70001 = ~n13404 ;
  assign n13720 = n70001 & n13719 ;
  assign n13721 = n13411 | n13720 ;
  assign n13722 = n13718 | n13721 ;
  assign n70002 = ~n13411 ;
  assign n13723 = n70002 & n13722 ;
  assign n70003 = ~n13401 ;
  assign n13724 = x88 & n70003 ;
  assign n70004 = ~n13396 ;
  assign n13725 = n70004 & n13724 ;
  assign n13726 = n13403 | n13725 ;
  assign n13728 = n13723 | n13726 ;
  assign n70005 = ~n13403 ;
  assign n13729 = n70005 & n13728 ;
  assign n70006 = ~n13393 ;
  assign n13730 = x89 & n70006 ;
  assign n70007 = ~n13388 ;
  assign n13731 = n70007 & n13730 ;
  assign n13732 = n13395 | n13731 ;
  assign n13733 = n13729 | n13732 ;
  assign n70008 = ~n13395 ;
  assign n13734 = n70008 & n13733 ;
  assign n70009 = ~n13385 ;
  assign n13735 = x90 & n70009 ;
  assign n70010 = ~n13380 ;
  assign n13736 = n70010 & n13735 ;
  assign n13737 = n13387 | n13736 ;
  assign n13739 = n13734 | n13737 ;
  assign n70011 = ~n13387 ;
  assign n13740 = n70011 & n13739 ;
  assign n70012 = ~n13377 ;
  assign n13741 = x91 & n70012 ;
  assign n70013 = ~n13372 ;
  assign n13742 = n70013 & n13741 ;
  assign n13743 = n13379 | n13742 ;
  assign n13744 = n13740 | n13743 ;
  assign n70014 = ~n13379 ;
  assign n13745 = n70014 & n13744 ;
  assign n70015 = ~n13369 ;
  assign n13746 = x92 & n70015 ;
  assign n70016 = ~n13364 ;
  assign n13747 = n70016 & n13746 ;
  assign n13748 = n13371 | n13747 ;
  assign n13750 = n13745 | n13748 ;
  assign n70017 = ~n13371 ;
  assign n13751 = n70017 & n13750 ;
  assign n70018 = ~n13361 ;
  assign n13752 = x93 & n70018 ;
  assign n70019 = ~n13356 ;
  assign n13753 = n70019 & n13752 ;
  assign n13754 = n13363 | n13753 ;
  assign n13755 = n13751 | n13754 ;
  assign n70020 = ~n13363 ;
  assign n13756 = n70020 & n13755 ;
  assign n70021 = ~n13353 ;
  assign n13757 = x94 & n70021 ;
  assign n70022 = ~n13348 ;
  assign n13758 = n70022 & n13757 ;
  assign n13759 = n13355 | n13758 ;
  assign n13761 = n13756 | n13759 ;
  assign n70023 = ~n13355 ;
  assign n13762 = n70023 & n13761 ;
  assign n70024 = ~n13345 ;
  assign n13763 = x95 & n70024 ;
  assign n70025 = ~n13340 ;
  assign n13764 = n70025 & n13763 ;
  assign n13765 = n13347 | n13764 ;
  assign n13766 = n13762 | n13765 ;
  assign n70026 = ~n13347 ;
  assign n13767 = n70026 & n13766 ;
  assign n70027 = ~n13337 ;
  assign n13768 = x96 & n70027 ;
  assign n70028 = ~n13332 ;
  assign n13769 = n70028 & n13768 ;
  assign n13770 = n13339 | n13769 ;
  assign n13772 = n13767 | n13770 ;
  assign n70029 = ~n13339 ;
  assign n13773 = n70029 & n13772 ;
  assign n70030 = ~n13329 ;
  assign n13774 = x97 & n70030 ;
  assign n70031 = ~n13324 ;
  assign n13775 = n70031 & n13774 ;
  assign n13776 = n13331 | n13775 ;
  assign n13777 = n13773 | n13776 ;
  assign n70032 = ~n13331 ;
  assign n13778 = n70032 & n13777 ;
  assign n70033 = ~n13321 ;
  assign n13779 = x98 & n70033 ;
  assign n70034 = ~n13316 ;
  assign n13780 = n70034 & n13779 ;
  assign n13781 = n13323 | n13780 ;
  assign n13783 = n13778 | n13781 ;
  assign n70035 = ~n13323 ;
  assign n13784 = n70035 & n13783 ;
  assign n70036 = ~n13313 ;
  assign n13785 = x99 & n70036 ;
  assign n70037 = ~n13308 ;
  assign n13786 = n70037 & n13785 ;
  assign n13787 = n13315 | n13786 ;
  assign n13788 = n13784 | n13787 ;
  assign n70038 = ~n13315 ;
  assign n13789 = n70038 & n13788 ;
  assign n70039 = ~n13305 ;
  assign n13790 = x100 & n70039 ;
  assign n70040 = ~n13300 ;
  assign n13791 = n70040 & n13790 ;
  assign n13792 = n13307 | n13791 ;
  assign n13794 = n13789 | n13792 ;
  assign n70041 = ~n13307 ;
  assign n13795 = n70041 & n13794 ;
  assign n70042 = ~n13297 ;
  assign n13796 = x101 & n70042 ;
  assign n70043 = ~n13292 ;
  assign n13797 = n70043 & n13796 ;
  assign n13798 = n13299 | n13797 ;
  assign n13799 = n13795 | n13798 ;
  assign n70044 = ~n13299 ;
  assign n13800 = n70044 & n13799 ;
  assign n70045 = ~n13289 ;
  assign n13801 = x102 & n70045 ;
  assign n70046 = ~n13284 ;
  assign n13802 = n70046 & n13801 ;
  assign n13803 = n13291 | n13802 ;
  assign n13805 = n13800 | n13803 ;
  assign n70047 = ~n13291 ;
  assign n13806 = n70047 & n13805 ;
  assign n70048 = ~n13281 ;
  assign n13807 = x103 & n70048 ;
  assign n70049 = ~n13276 ;
  assign n13808 = n70049 & n13807 ;
  assign n13809 = n13283 | n13808 ;
  assign n13810 = n13806 | n13809 ;
  assign n70050 = ~n13283 ;
  assign n13811 = n70050 & n13810 ;
  assign n153 = ~n13185 ;
  assign n13812 = n153 & n13272 ;
  assign n13813 = n12647 & n13185 ;
  assign n70052 = ~n13813 ;
  assign n13814 = x104 & n70052 ;
  assign n70053 = ~n13812 ;
  assign n13815 = n70053 & n13814 ;
  assign n13816 = n13275 | n13815 ;
  assign n13818 = n13811 | n13816 ;
  assign n70054 = ~n13275 ;
  assign n13819 = n70054 & n13818 ;
  assign n13820 = n279 | n293 ;
  assign n13821 = n13819 | n13820 ;
  assign n13822 = n13282 & n13821 ;
  assign n13592 = n65670 & n13590 ;
  assign n13823 = x65 & n13601 ;
  assign n70055 = ~n13823 ;
  assign n13824 = n13594 & n70055 ;
  assign n13825 = n13596 | n13824 ;
  assign n70056 = ~n13592 ;
  assign n13826 = n70056 & n13825 ;
  assign n13827 = n13607 | n13826 ;
  assign n13828 = n69939 & n13827 ;
  assign n13829 = n13611 | n13828 ;
  assign n13831 = n69942 & n13829 ;
  assign n13833 = n13617 | n13831 ;
  assign n13834 = n69945 & n13833 ;
  assign n13836 = n13622 | n13834 ;
  assign n13837 = n69948 & n13836 ;
  assign n13838 = n13627 | n13837 ;
  assign n13839 = n69951 & n13838 ;
  assign n13840 = n13633 | n13839 ;
  assign n13842 = n69954 & n13840 ;
  assign n13843 = n13638 | n13842 ;
  assign n13844 = n69957 & n13843 ;
  assign n13845 = n13644 | n13844 ;
  assign n13847 = n69960 & n13845 ;
  assign n13848 = n13649 | n13847 ;
  assign n13849 = n69963 & n13848 ;
  assign n13850 = n13655 | n13849 ;
  assign n13852 = n69966 & n13850 ;
  assign n13853 = n13660 | n13852 ;
  assign n13854 = n69969 & n13853 ;
  assign n13855 = n13666 | n13854 ;
  assign n13857 = n69972 & n13855 ;
  assign n13858 = n13671 | n13857 ;
  assign n13859 = n69975 & n13858 ;
  assign n13860 = n13677 | n13859 ;
  assign n13862 = n69978 & n13860 ;
  assign n13863 = n13682 | n13862 ;
  assign n13864 = n69981 & n13863 ;
  assign n13865 = n13688 | n13864 ;
  assign n13867 = n69984 & n13865 ;
  assign n13868 = n13693 | n13867 ;
  assign n13869 = n69987 & n13868 ;
  assign n13870 = n13699 | n13869 ;
  assign n13872 = n69990 & n13870 ;
  assign n13873 = n13704 | n13872 ;
  assign n13874 = n69993 & n13873 ;
  assign n13875 = n13710 | n13874 ;
  assign n13877 = n69996 & n13875 ;
  assign n13878 = n13715 | n13877 ;
  assign n13879 = n69999 & n13878 ;
  assign n13880 = n13721 | n13879 ;
  assign n13882 = n70002 & n13880 ;
  assign n13883 = n13726 | n13882 ;
  assign n13884 = n70005 & n13883 ;
  assign n13885 = n13732 | n13884 ;
  assign n13887 = n70008 & n13885 ;
  assign n13888 = n13737 | n13887 ;
  assign n13889 = n70011 & n13888 ;
  assign n13890 = n13743 | n13889 ;
  assign n13892 = n70014 & n13890 ;
  assign n13893 = n13748 | n13892 ;
  assign n13894 = n70017 & n13893 ;
  assign n13895 = n13754 | n13894 ;
  assign n13897 = n70020 & n13895 ;
  assign n13898 = n13759 | n13897 ;
  assign n13899 = n70023 & n13898 ;
  assign n13900 = n13765 | n13899 ;
  assign n13902 = n70026 & n13900 ;
  assign n13903 = n13770 | n13902 ;
  assign n13904 = n70029 & n13903 ;
  assign n13905 = n13776 | n13904 ;
  assign n13907 = n70032 & n13905 ;
  assign n13908 = n13781 | n13907 ;
  assign n13909 = n70035 & n13908 ;
  assign n13910 = n13787 | n13909 ;
  assign n13912 = n70038 & n13910 ;
  assign n13913 = n13792 | n13912 ;
  assign n13914 = n70041 & n13913 ;
  assign n13915 = n13798 | n13914 ;
  assign n13917 = n70044 & n13915 ;
  assign n13918 = n13803 | n13917 ;
  assign n13919 = n70047 & n13918 ;
  assign n70057 = ~n13919 ;
  assign n13920 = n13809 & n70057 ;
  assign n13922 = n13291 | n13809 ;
  assign n70058 = ~n13922 ;
  assign n13923 = n13805 & n70058 ;
  assign n13924 = n13920 | n13923 ;
  assign n70059 = ~n13820 ;
  assign n13925 = n70059 & n13924 ;
  assign n70060 = ~n13819 ;
  assign n13926 = n70060 & n13925 ;
  assign n13927 = n13822 | n13926 ;
  assign n13928 = n69857 & n13927 ;
  assign n70061 = ~n13926 ;
  assign n14454 = x104 & n70061 ;
  assign n70062 = ~n13822 ;
  assign n14455 = n70062 & n14454 ;
  assign n14456 = n13928 | n14455 ;
  assign n13929 = n13290 & n13821 ;
  assign n70063 = ~n13800 ;
  assign n13804 = n70063 & n13803 ;
  assign n13930 = n13299 | n13803 ;
  assign n70064 = ~n13930 ;
  assign n13931 = n13915 & n70064 ;
  assign n13932 = n13804 | n13931 ;
  assign n13933 = n70059 & n13932 ;
  assign n13934 = n70060 & n13933 ;
  assign n13935 = n13929 | n13934 ;
  assign n13936 = n69656 & n13935 ;
  assign n13937 = n13298 & n13821 ;
  assign n70065 = ~n13914 ;
  assign n13916 = n13798 & n70065 ;
  assign n13938 = n13307 | n13798 ;
  assign n70066 = ~n13938 ;
  assign n13939 = n13794 & n70066 ;
  assign n13940 = n13916 | n13939 ;
  assign n13941 = n70059 & n13940 ;
  assign n13942 = n70060 & n13941 ;
  assign n13943 = n13937 | n13942 ;
  assign n13944 = n69528 & n13943 ;
  assign n70067 = ~n13942 ;
  assign n14443 = x102 & n70067 ;
  assign n70068 = ~n13937 ;
  assign n14444 = n70068 & n14443 ;
  assign n14445 = n13944 | n14444 ;
  assign n13945 = n13306 & n13821 ;
  assign n70069 = ~n13789 ;
  assign n13793 = n70069 & n13792 ;
  assign n13946 = n13315 | n13792 ;
  assign n70070 = ~n13946 ;
  assign n13947 = n13910 & n70070 ;
  assign n13948 = n13793 | n13947 ;
  assign n13949 = n70059 & n13948 ;
  assign n13950 = n70060 & n13949 ;
  assign n13951 = n13945 | n13950 ;
  assign n13952 = n69261 & n13951 ;
  assign n13953 = n13314 & n13821 ;
  assign n70071 = ~n13909 ;
  assign n13911 = n13787 & n70071 ;
  assign n13954 = n13323 | n13787 ;
  assign n70072 = ~n13954 ;
  assign n13955 = n13783 & n70072 ;
  assign n13956 = n13911 | n13955 ;
  assign n13957 = n70059 & n13956 ;
  assign n13958 = n70060 & n13957 ;
  assign n13959 = n13953 | n13958 ;
  assign n13960 = n69075 & n13959 ;
  assign n70073 = ~n13958 ;
  assign n14433 = x100 & n70073 ;
  assign n70074 = ~n13953 ;
  assign n14434 = n70074 & n14433 ;
  assign n14435 = n13960 | n14434 ;
  assign n13961 = n13322 & n13821 ;
  assign n70075 = ~n13778 ;
  assign n13782 = n70075 & n13781 ;
  assign n13962 = n13331 | n13781 ;
  assign n70076 = ~n13962 ;
  assign n13963 = n13905 & n70076 ;
  assign n13964 = n13782 | n13963 ;
  assign n13965 = n70059 & n13964 ;
  assign n13966 = n70060 & n13965 ;
  assign n13967 = n13961 | n13966 ;
  assign n13968 = n68993 & n13967 ;
  assign n13969 = n13330 & n13821 ;
  assign n70077 = ~n13904 ;
  assign n13906 = n13776 & n70077 ;
  assign n13970 = n13339 | n13776 ;
  assign n70078 = ~n13970 ;
  assign n13971 = n13772 & n70078 ;
  assign n13972 = n13906 | n13971 ;
  assign n13973 = n70059 & n13972 ;
  assign n13974 = n70060 & n13973 ;
  assign n13975 = n13969 | n13974 ;
  assign n13976 = n68716 & n13975 ;
  assign n70079 = ~n13974 ;
  assign n14423 = x98 & n70079 ;
  assign n70080 = ~n13969 ;
  assign n14424 = n70080 & n14423 ;
  assign n14425 = n13976 | n14424 ;
  assign n13977 = n13338 & n13821 ;
  assign n70081 = ~n13767 ;
  assign n13771 = n70081 & n13770 ;
  assign n13978 = n13347 | n13770 ;
  assign n70082 = ~n13978 ;
  assign n13979 = n13900 & n70082 ;
  assign n13980 = n13771 | n13979 ;
  assign n13981 = n70059 & n13980 ;
  assign n13982 = n70060 & n13981 ;
  assign n13983 = n13977 | n13982 ;
  assign n13984 = n68545 & n13983 ;
  assign n13985 = n13346 & n13821 ;
  assign n70083 = ~n13899 ;
  assign n13901 = n13765 & n70083 ;
  assign n13986 = n13355 | n13765 ;
  assign n70084 = ~n13986 ;
  assign n13987 = n13761 & n70084 ;
  assign n13988 = n13901 | n13987 ;
  assign n13989 = n70059 & n13988 ;
  assign n13990 = n70060 & n13989 ;
  assign n13991 = n13985 | n13990 ;
  assign n13992 = n68438 & n13991 ;
  assign n70085 = ~n13990 ;
  assign n14413 = x96 & n70085 ;
  assign n70086 = ~n13985 ;
  assign n14414 = n70086 & n14413 ;
  assign n14415 = n13992 | n14414 ;
  assign n13993 = n13354 & n13821 ;
  assign n70087 = ~n13756 ;
  assign n13760 = n70087 & n13759 ;
  assign n13994 = n13363 | n13759 ;
  assign n70088 = ~n13994 ;
  assign n13995 = n13895 & n70088 ;
  assign n13996 = n13760 | n13995 ;
  assign n13997 = n70059 & n13996 ;
  assign n13998 = n70060 & n13997 ;
  assign n13999 = n13993 | n13998 ;
  assign n14000 = n68214 & n13999 ;
  assign n14001 = n13362 & n13821 ;
  assign n70089 = ~n13894 ;
  assign n13896 = n13754 & n70089 ;
  assign n14002 = n13371 | n13754 ;
  assign n70090 = ~n14002 ;
  assign n14003 = n13750 & n70090 ;
  assign n14004 = n13896 | n14003 ;
  assign n14005 = n70059 & n14004 ;
  assign n14006 = n70060 & n14005 ;
  assign n14007 = n14001 | n14006 ;
  assign n14008 = n68058 & n14007 ;
  assign n70091 = ~n14006 ;
  assign n14403 = x94 & n70091 ;
  assign n70092 = ~n14001 ;
  assign n14404 = n70092 & n14403 ;
  assign n14405 = n14008 | n14404 ;
  assign n14009 = n13370 & n13821 ;
  assign n70093 = ~n13745 ;
  assign n13749 = n70093 & n13748 ;
  assign n14010 = n13379 | n13748 ;
  assign n70094 = ~n14010 ;
  assign n14011 = n13890 & n70094 ;
  assign n14012 = n13749 | n14011 ;
  assign n14013 = n70059 & n14012 ;
  assign n14014 = n70060 & n14013 ;
  assign n14015 = n14009 | n14014 ;
  assign n14016 = n67986 & n14015 ;
  assign n14017 = n13378 & n13821 ;
  assign n70095 = ~n13889 ;
  assign n13891 = n13743 & n70095 ;
  assign n14018 = n13387 | n13743 ;
  assign n70096 = ~n14018 ;
  assign n14019 = n13739 & n70096 ;
  assign n14020 = n13891 | n14019 ;
  assign n14021 = n70059 & n14020 ;
  assign n14022 = n70060 & n14021 ;
  assign n14023 = n14017 | n14022 ;
  assign n14024 = n67763 & n14023 ;
  assign n70097 = ~n14022 ;
  assign n14393 = x92 & n70097 ;
  assign n70098 = ~n14017 ;
  assign n14394 = n70098 & n14393 ;
  assign n14395 = n14024 | n14394 ;
  assign n14025 = n13386 & n13821 ;
  assign n70099 = ~n13734 ;
  assign n13738 = n70099 & n13737 ;
  assign n14026 = n13395 | n13737 ;
  assign n70100 = ~n14026 ;
  assign n14027 = n13885 & n70100 ;
  assign n14028 = n13738 | n14027 ;
  assign n14029 = n70059 & n14028 ;
  assign n14030 = n70060 & n14029 ;
  assign n14031 = n14025 | n14030 ;
  assign n14032 = n67622 & n14031 ;
  assign n14033 = n13394 & n13821 ;
  assign n70101 = ~n13884 ;
  assign n13886 = n13732 & n70101 ;
  assign n14034 = n13403 | n13732 ;
  assign n70102 = ~n14034 ;
  assign n14035 = n13728 & n70102 ;
  assign n14036 = n13886 | n14035 ;
  assign n14037 = n70059 & n14036 ;
  assign n14038 = n70060 & n14037 ;
  assign n14039 = n14033 | n14038 ;
  assign n14040 = n67531 & n14039 ;
  assign n70103 = ~n14038 ;
  assign n14383 = x90 & n70103 ;
  assign n70104 = ~n14033 ;
  assign n14384 = n70104 & n14383 ;
  assign n14385 = n14040 | n14384 ;
  assign n14041 = n13402 & n13821 ;
  assign n70105 = ~n13723 ;
  assign n13727 = n70105 & n13726 ;
  assign n14042 = n13411 | n13726 ;
  assign n70106 = ~n14042 ;
  assign n14043 = n13880 & n70106 ;
  assign n14044 = n13727 | n14043 ;
  assign n14045 = n70059 & n14044 ;
  assign n14046 = n70060 & n14045 ;
  assign n14047 = n14041 | n14046 ;
  assign n14048 = n67348 & n14047 ;
  assign n14049 = n13410 & n13821 ;
  assign n70107 = ~n13879 ;
  assign n13881 = n13721 & n70107 ;
  assign n14050 = n13419 | n13721 ;
  assign n70108 = ~n14050 ;
  assign n14051 = n13717 & n70108 ;
  assign n14052 = n13881 | n14051 ;
  assign n14053 = n70059 & n14052 ;
  assign n14054 = n70060 & n14053 ;
  assign n14055 = n14049 | n14054 ;
  assign n14056 = n67222 & n14055 ;
  assign n70109 = ~n14054 ;
  assign n14373 = x88 & n70109 ;
  assign n70110 = ~n14049 ;
  assign n14374 = n70110 & n14373 ;
  assign n14375 = n14056 | n14374 ;
  assign n14057 = n13418 & n13821 ;
  assign n70111 = ~n13712 ;
  assign n13716 = n70111 & n13715 ;
  assign n14058 = n13427 | n13715 ;
  assign n70112 = ~n14058 ;
  assign n14059 = n13875 & n70112 ;
  assign n14060 = n13716 | n14059 ;
  assign n14061 = n70059 & n14060 ;
  assign n14062 = n70060 & n14061 ;
  assign n14063 = n14057 | n14062 ;
  assign n14064 = n67164 & n14063 ;
  assign n14065 = n13426 & n13821 ;
  assign n70113 = ~n13874 ;
  assign n13876 = n13710 & n70113 ;
  assign n14066 = n13435 | n13710 ;
  assign n70114 = ~n14066 ;
  assign n14067 = n13706 & n70114 ;
  assign n14068 = n13876 | n14067 ;
  assign n14069 = n70059 & n14068 ;
  assign n14070 = n70060 & n14069 ;
  assign n14071 = n14065 | n14070 ;
  assign n14072 = n66979 & n14071 ;
  assign n70115 = ~n14070 ;
  assign n14362 = x86 & n70115 ;
  assign n70116 = ~n14065 ;
  assign n14363 = n70116 & n14362 ;
  assign n14364 = n14072 | n14363 ;
  assign n14073 = n13434 & n13821 ;
  assign n70117 = ~n13701 ;
  assign n13705 = n70117 & n13704 ;
  assign n14074 = n13443 | n13704 ;
  assign n70118 = ~n14074 ;
  assign n14075 = n13870 & n70118 ;
  assign n14076 = n13705 | n14075 ;
  assign n14077 = n70059 & n14076 ;
  assign n14078 = n70060 & n14077 ;
  assign n14079 = n14073 | n14078 ;
  assign n14080 = n66868 & n14079 ;
  assign n14081 = n13442 & n13821 ;
  assign n70119 = ~n13869 ;
  assign n13871 = n13699 & n70119 ;
  assign n14082 = n13451 | n13699 ;
  assign n70120 = ~n14082 ;
  assign n14083 = n13695 & n70120 ;
  assign n14084 = n13871 | n14083 ;
  assign n14085 = n70059 & n14084 ;
  assign n14086 = n70060 & n14085 ;
  assign n14087 = n14081 | n14086 ;
  assign n14088 = n66797 & n14087 ;
  assign n70121 = ~n14086 ;
  assign n14352 = x84 & n70121 ;
  assign n70122 = ~n14081 ;
  assign n14353 = n70122 & n14352 ;
  assign n14354 = n14088 | n14353 ;
  assign n14089 = n13450 & n13821 ;
  assign n70123 = ~n13690 ;
  assign n13694 = n70123 & n13693 ;
  assign n14090 = n13459 | n13693 ;
  assign n70124 = ~n14090 ;
  assign n14091 = n13865 & n70124 ;
  assign n14092 = n13694 | n14091 ;
  assign n14093 = n70059 & n14092 ;
  assign n14094 = n70060 & n14093 ;
  assign n14095 = n14089 | n14094 ;
  assign n14096 = n66654 & n14095 ;
  assign n14097 = n13458 & n13821 ;
  assign n70125 = ~n13864 ;
  assign n13866 = n13688 & n70125 ;
  assign n14098 = n13467 | n13688 ;
  assign n70126 = ~n14098 ;
  assign n14099 = n13684 & n70126 ;
  assign n14100 = n13866 | n14099 ;
  assign n14101 = n70059 & n14100 ;
  assign n14102 = n70060 & n14101 ;
  assign n14103 = n14097 | n14102 ;
  assign n14104 = n66560 & n14103 ;
  assign n70127 = ~n14102 ;
  assign n14342 = x82 & n70127 ;
  assign n70128 = ~n14097 ;
  assign n14343 = n70128 & n14342 ;
  assign n14344 = n14104 | n14343 ;
  assign n14105 = n13466 & n13821 ;
  assign n70129 = ~n13679 ;
  assign n13683 = n70129 & n13682 ;
  assign n14106 = n13475 | n13682 ;
  assign n70130 = ~n14106 ;
  assign n14107 = n13860 & n70130 ;
  assign n14108 = n13683 | n14107 ;
  assign n14109 = n70059 & n14108 ;
  assign n14110 = n70060 & n14109 ;
  assign n14111 = n14105 | n14110 ;
  assign n14112 = n66505 & n14111 ;
  assign n14113 = n13474 & n13821 ;
  assign n70131 = ~n13859 ;
  assign n13861 = n13677 & n70131 ;
  assign n14114 = n13483 | n13677 ;
  assign n70132 = ~n14114 ;
  assign n14115 = n13673 & n70132 ;
  assign n14116 = n13861 | n14115 ;
  assign n14117 = n70059 & n14116 ;
  assign n14118 = n70060 & n14117 ;
  assign n14119 = n14113 | n14118 ;
  assign n14120 = n66379 & n14119 ;
  assign n70133 = ~n14118 ;
  assign n14331 = x80 & n70133 ;
  assign n70134 = ~n14113 ;
  assign n14332 = n70134 & n14331 ;
  assign n14333 = n14120 | n14332 ;
  assign n14121 = n13482 & n13821 ;
  assign n70135 = ~n13668 ;
  assign n13672 = n70135 & n13671 ;
  assign n14122 = n13491 | n13671 ;
  assign n70136 = ~n14122 ;
  assign n14123 = n13855 & n70136 ;
  assign n14124 = n13672 | n14123 ;
  assign n14125 = n70059 & n14124 ;
  assign n14126 = n70060 & n14125 ;
  assign n14127 = n14121 | n14126 ;
  assign n14128 = n66299 & n14127 ;
  assign n14129 = n13490 & n13821 ;
  assign n70137 = ~n13854 ;
  assign n13856 = n13666 & n70137 ;
  assign n14130 = n13499 | n13666 ;
  assign n70138 = ~n14130 ;
  assign n14131 = n13662 & n70138 ;
  assign n14132 = n13856 | n14131 ;
  assign n14133 = n70059 & n14132 ;
  assign n14134 = n70060 & n14133 ;
  assign n14135 = n14129 | n14134 ;
  assign n14136 = n66244 & n14135 ;
  assign n70139 = ~n14134 ;
  assign n14321 = x78 & n70139 ;
  assign n70140 = ~n14129 ;
  assign n14322 = n70140 & n14321 ;
  assign n14323 = n14136 | n14322 ;
  assign n14137 = n13498 & n13821 ;
  assign n70141 = ~n13657 ;
  assign n13661 = n70141 & n13660 ;
  assign n14138 = n13507 | n13660 ;
  assign n70142 = ~n14138 ;
  assign n14139 = n13850 & n70142 ;
  assign n14140 = n13661 | n14139 ;
  assign n14141 = n70059 & n14140 ;
  assign n14142 = n70060 & n14141 ;
  assign n14143 = n14137 | n14142 ;
  assign n14144 = n66145 & n14143 ;
  assign n14145 = n13506 & n13821 ;
  assign n70143 = ~n13849 ;
  assign n13851 = n13655 & n70143 ;
  assign n14146 = n13515 | n13655 ;
  assign n70144 = ~n14146 ;
  assign n14147 = n13651 & n70144 ;
  assign n14148 = n13851 | n14147 ;
  assign n14149 = n70059 & n14148 ;
  assign n14150 = n70060 & n14149 ;
  assign n14151 = n14145 | n14150 ;
  assign n14152 = n66081 & n14151 ;
  assign n70145 = ~n14150 ;
  assign n14310 = x76 & n70145 ;
  assign n70146 = ~n14145 ;
  assign n14311 = n70146 & n14310 ;
  assign n14312 = n14152 | n14311 ;
  assign n14153 = n13514 & n13821 ;
  assign n70147 = ~n13646 ;
  assign n13650 = n70147 & n13649 ;
  assign n14154 = n13523 | n13649 ;
  assign n70148 = ~n14154 ;
  assign n14155 = n13845 & n70148 ;
  assign n14156 = n13650 | n14155 ;
  assign n14157 = n70059 & n14156 ;
  assign n14158 = n70060 & n14157 ;
  assign n14159 = n14153 | n14158 ;
  assign n14160 = n66043 & n14159 ;
  assign n14161 = n13522 & n13821 ;
  assign n70149 = ~n13844 ;
  assign n13846 = n13644 & n70149 ;
  assign n14162 = n13531 | n13644 ;
  assign n70150 = ~n14162 ;
  assign n14163 = n13640 & n70150 ;
  assign n14164 = n13846 | n14163 ;
  assign n14165 = n70059 & n14164 ;
  assign n14166 = n70060 & n14165 ;
  assign n14167 = n14161 | n14166 ;
  assign n14168 = n65960 & n14167 ;
  assign n70151 = ~n14166 ;
  assign n14299 = x74 & n70151 ;
  assign n70152 = ~n14161 ;
  assign n14300 = n70152 & n14299 ;
  assign n14301 = n14168 | n14300 ;
  assign n14169 = n13530 & n13821 ;
  assign n70153 = ~n13635 ;
  assign n13639 = n70153 & n13638 ;
  assign n14170 = n13539 | n13638 ;
  assign n70154 = ~n14170 ;
  assign n14171 = n13840 & n70154 ;
  assign n14172 = n13639 | n14171 ;
  assign n14173 = n70059 & n14172 ;
  assign n14174 = n70060 & n14173 ;
  assign n14175 = n14169 | n14174 ;
  assign n14176 = n65909 & n14175 ;
  assign n14177 = n13538 & n13821 ;
  assign n70155 = ~n13839 ;
  assign n13841 = n13633 & n70155 ;
  assign n14178 = n13547 | n13633 ;
  assign n70156 = ~n14178 ;
  assign n14179 = n13629 & n70156 ;
  assign n14180 = n13841 | n14179 ;
  assign n14181 = n70059 & n14180 ;
  assign n14182 = n70060 & n14181 ;
  assign n14183 = n14177 | n14182 ;
  assign n14184 = n65877 & n14183 ;
  assign n70157 = ~n14182 ;
  assign n14288 = x72 & n70157 ;
  assign n70158 = ~n14177 ;
  assign n14289 = n70158 & n14288 ;
  assign n14290 = n14184 | n14289 ;
  assign n14185 = n13546 & n13821 ;
  assign n70159 = ~n13624 ;
  assign n13628 = n70159 & n13627 ;
  assign n14186 = n13556 | n13627 ;
  assign n70160 = ~n14186 ;
  assign n14187 = n13836 & n70160 ;
  assign n14188 = n13628 | n14187 ;
  assign n14189 = n70059 & n14188 ;
  assign n14190 = n70060 & n14189 ;
  assign n14191 = n14185 | n14190 ;
  assign n14192 = n65820 & n14191 ;
  assign n14193 = n13555 & n13821 ;
  assign n70161 = ~n13834 ;
  assign n13835 = n13622 & n70161 ;
  assign n14194 = n13565 | n13622 ;
  assign n70162 = ~n14194 ;
  assign n14195 = n13833 & n70162 ;
  assign n14196 = n13835 | n14195 ;
  assign n14197 = n70059 & n14196 ;
  assign n14198 = n70060 & n14197 ;
  assign n14199 = n14193 | n14198 ;
  assign n14200 = n65791 & n14199 ;
  assign n70163 = ~n14198 ;
  assign n14278 = x70 & n70163 ;
  assign n70164 = ~n14193 ;
  assign n14279 = n70164 & n14278 ;
  assign n14280 = n14200 | n14279 ;
  assign n14201 = n13564 & n13821 ;
  assign n70165 = ~n13614 ;
  assign n13832 = n70165 & n13617 ;
  assign n14202 = n13612 | n13828 ;
  assign n14203 = n13573 | n13617 ;
  assign n70166 = ~n14203 ;
  assign n14204 = n14202 & n70166 ;
  assign n14205 = n13832 | n14204 ;
  assign n14206 = n70059 & n14205 ;
  assign n14207 = n70060 & n14206 ;
  assign n14208 = n14201 | n14207 ;
  assign n14209 = n65772 & n14208 ;
  assign n14210 = n13572 & n13821 ;
  assign n70167 = ~n13828 ;
  assign n13830 = n13612 & n70167 ;
  assign n14211 = n13579 | n13612 ;
  assign n70168 = ~n14211 ;
  assign n14212 = n13827 & n70168 ;
  assign n14213 = n13830 | n14212 ;
  assign n14214 = n70059 & n14213 ;
  assign n14215 = n70060 & n14214 ;
  assign n14216 = n14210 | n14215 ;
  assign n14217 = n65746 & n14216 ;
  assign n70169 = ~n14215 ;
  assign n14268 = x68 & n70169 ;
  assign n70170 = ~n14210 ;
  assign n14269 = n70170 & n14268 ;
  assign n14270 = n14217 | n14269 ;
  assign n14218 = n13578 & n13821 ;
  assign n14219 = n13602 | n13607 ;
  assign n70171 = ~n14219 ;
  assign n14220 = n13825 & n70171 ;
  assign n70172 = ~n13604 ;
  assign n14221 = n70172 & n13607 ;
  assign n14222 = n14220 | n14221 ;
  assign n14223 = n70059 & n14222 ;
  assign n14224 = n70060 & n14223 ;
  assign n14225 = n14218 | n14224 ;
  assign n14227 = n65721 & n14225 ;
  assign n13921 = n13809 | n13919 ;
  assign n14228 = n70050 & n13921 ;
  assign n14229 = n13816 | n14228 ;
  assign n14230 = n70054 & n14229 ;
  assign n14231 = n13820 | n14230 ;
  assign n14232 = n13601 & n14231 ;
  assign n14233 = n13594 & n13596 ;
  assign n14234 = n70055 & n14233 ;
  assign n14235 = n13820 | n14234 ;
  assign n70173 = ~n14235 ;
  assign n14236 = n13825 & n70173 ;
  assign n14237 = n70060 & n14236 ;
  assign n14238 = n14232 | n14237 ;
  assign n14239 = n65686 & n14238 ;
  assign n14258 = n13590 & n13821 ;
  assign n70174 = ~n14237 ;
  assign n14259 = x66 & n70174 ;
  assign n70175 = ~n14258 ;
  assign n14260 = n70175 & n14259 ;
  assign n14261 = n14239 | n14260 ;
  assign n70176 = ~x105 ;
  assign n14240 = x64 & n70176 ;
  assign n70177 = ~n65444 ;
  assign n14241 = n70177 & n14240 ;
  assign n70178 = ~n65527 ;
  assign n14242 = n70178 & n14241 ;
  assign n14243 = n66510 & n14242 ;
  assign n70179 = ~n14230 ;
  assign n14244 = n70179 & n14243 ;
  assign n70180 = ~n14244 ;
  assign n14245 = x23 & n70180 ;
  assign n14246 = n69530 & n13596 ;
  assign n14247 = n69531 & n14246 ;
  assign n14248 = n67026 & n14247 ;
  assign n14249 = n70060 & n14248 ;
  assign n14250 = n14245 | n14249 ;
  assign n14251 = x65 & n14250 ;
  assign n14252 = x65 | n14249 ;
  assign n14253 = n14245 | n14252 ;
  assign n70181 = ~n14251 ;
  assign n14254 = n70181 & n14253 ;
  assign n70182 = ~x22 ;
  assign n14255 = n70182 & x64 ;
  assign n14256 = n14254 | n14255 ;
  assign n14257 = n65670 & n14250 ;
  assign n70183 = ~n14257 ;
  assign n14262 = n14256 & n70183 ;
  assign n14263 = n14261 | n14262 ;
  assign n70184 = ~n14239 ;
  assign n14264 = n70184 & n14263 ;
  assign n70185 = ~n14224 ;
  assign n14226 = x67 & n70185 ;
  assign n70186 = ~n14218 ;
  assign n14265 = n70186 & n14226 ;
  assign n14266 = n14227 | n14265 ;
  assign n14267 = n14264 | n14266 ;
  assign n70187 = ~n14227 ;
  assign n14271 = n70187 & n14267 ;
  assign n14272 = n14270 | n14271 ;
  assign n70188 = ~n14217 ;
  assign n14273 = n70188 & n14272 ;
  assign n70189 = ~n14207 ;
  assign n14274 = x69 & n70189 ;
  assign n70190 = ~n14201 ;
  assign n14275 = n70190 & n14274 ;
  assign n14276 = n14209 | n14275 ;
  assign n14277 = n14273 | n14276 ;
  assign n70191 = ~n14209 ;
  assign n14281 = n70191 & n14277 ;
  assign n14282 = n14280 | n14281 ;
  assign n70192 = ~n14200 ;
  assign n14283 = n70192 & n14282 ;
  assign n70193 = ~n14190 ;
  assign n14284 = x71 & n70193 ;
  assign n70194 = ~n14185 ;
  assign n14285 = n70194 & n14284 ;
  assign n14286 = n14192 | n14285 ;
  assign n14287 = n14283 | n14286 ;
  assign n70195 = ~n14192 ;
  assign n14291 = n70195 & n14287 ;
  assign n14292 = n14290 | n14291 ;
  assign n70196 = ~n14184 ;
  assign n14293 = n70196 & n14292 ;
  assign n70197 = ~n14174 ;
  assign n14294 = x73 & n70197 ;
  assign n70198 = ~n14169 ;
  assign n14295 = n70198 & n14294 ;
  assign n14296 = n14176 | n14295 ;
  assign n14298 = n14293 | n14296 ;
  assign n70199 = ~n14176 ;
  assign n14302 = n70199 & n14298 ;
  assign n14303 = n14301 | n14302 ;
  assign n70200 = ~n14168 ;
  assign n14304 = n70200 & n14303 ;
  assign n70201 = ~n14158 ;
  assign n14305 = x75 & n70201 ;
  assign n70202 = ~n14153 ;
  assign n14306 = n70202 & n14305 ;
  assign n14307 = n14160 | n14306 ;
  assign n14309 = n14304 | n14307 ;
  assign n70203 = ~n14160 ;
  assign n14313 = n70203 & n14309 ;
  assign n14314 = n14312 | n14313 ;
  assign n70204 = ~n14152 ;
  assign n14315 = n70204 & n14314 ;
  assign n70205 = ~n14142 ;
  assign n14316 = x77 & n70205 ;
  assign n70206 = ~n14137 ;
  assign n14317 = n70206 & n14316 ;
  assign n14318 = n14144 | n14317 ;
  assign n14320 = n14315 | n14318 ;
  assign n70207 = ~n14144 ;
  assign n14324 = n70207 & n14320 ;
  assign n14325 = n14323 | n14324 ;
  assign n70208 = ~n14136 ;
  assign n14326 = n70208 & n14325 ;
  assign n70209 = ~n14126 ;
  assign n14327 = x79 & n70209 ;
  assign n70210 = ~n14121 ;
  assign n14328 = n70210 & n14327 ;
  assign n14329 = n14128 | n14328 ;
  assign n14330 = n14326 | n14329 ;
  assign n70211 = ~n14128 ;
  assign n14335 = n70211 & n14330 ;
  assign n14336 = n14333 | n14335 ;
  assign n70212 = ~n14120 ;
  assign n14337 = n70212 & n14336 ;
  assign n70213 = ~n14110 ;
  assign n14338 = x81 & n70213 ;
  assign n70214 = ~n14105 ;
  assign n14339 = n70214 & n14338 ;
  assign n14340 = n14112 | n14339 ;
  assign n14341 = n14337 | n14340 ;
  assign n70215 = ~n14112 ;
  assign n14345 = n70215 & n14341 ;
  assign n14346 = n14344 | n14345 ;
  assign n70216 = ~n14104 ;
  assign n14347 = n70216 & n14346 ;
  assign n70217 = ~n14094 ;
  assign n14348 = x83 & n70217 ;
  assign n70218 = ~n14089 ;
  assign n14349 = n70218 & n14348 ;
  assign n14350 = n14096 | n14349 ;
  assign n14351 = n14347 | n14350 ;
  assign n70219 = ~n14096 ;
  assign n14355 = n70219 & n14351 ;
  assign n14356 = n14354 | n14355 ;
  assign n70220 = ~n14088 ;
  assign n14357 = n70220 & n14356 ;
  assign n70221 = ~n14078 ;
  assign n14358 = x85 & n70221 ;
  assign n70222 = ~n14073 ;
  assign n14359 = n70222 & n14358 ;
  assign n14360 = n14080 | n14359 ;
  assign n14361 = n14357 | n14360 ;
  assign n70223 = ~n14080 ;
  assign n14365 = n70223 & n14361 ;
  assign n14366 = n14364 | n14365 ;
  assign n70224 = ~n14072 ;
  assign n14367 = n70224 & n14366 ;
  assign n70225 = ~n14062 ;
  assign n14368 = x87 & n70225 ;
  assign n70226 = ~n14057 ;
  assign n14369 = n70226 & n14368 ;
  assign n14370 = n14064 | n14369 ;
  assign n14372 = n14367 | n14370 ;
  assign n70227 = ~n14064 ;
  assign n14376 = n70227 & n14372 ;
  assign n14377 = n14375 | n14376 ;
  assign n70228 = ~n14056 ;
  assign n14378 = n70228 & n14377 ;
  assign n70229 = ~n14046 ;
  assign n14379 = x89 & n70229 ;
  assign n70230 = ~n14041 ;
  assign n14380 = n70230 & n14379 ;
  assign n14381 = n14048 | n14380 ;
  assign n14382 = n14378 | n14381 ;
  assign n70231 = ~n14048 ;
  assign n14386 = n70231 & n14382 ;
  assign n14387 = n14385 | n14386 ;
  assign n70232 = ~n14040 ;
  assign n14388 = n70232 & n14387 ;
  assign n70233 = ~n14030 ;
  assign n14389 = x91 & n70233 ;
  assign n70234 = ~n14025 ;
  assign n14390 = n70234 & n14389 ;
  assign n14391 = n14032 | n14390 ;
  assign n14392 = n14388 | n14391 ;
  assign n70235 = ~n14032 ;
  assign n14396 = n70235 & n14392 ;
  assign n14397 = n14395 | n14396 ;
  assign n70236 = ~n14024 ;
  assign n14398 = n70236 & n14397 ;
  assign n70237 = ~n14014 ;
  assign n14399 = x93 & n70237 ;
  assign n70238 = ~n14009 ;
  assign n14400 = n70238 & n14399 ;
  assign n14401 = n14016 | n14400 ;
  assign n14402 = n14398 | n14401 ;
  assign n70239 = ~n14016 ;
  assign n14406 = n70239 & n14402 ;
  assign n14407 = n14405 | n14406 ;
  assign n70240 = ~n14008 ;
  assign n14408 = n70240 & n14407 ;
  assign n70241 = ~n13998 ;
  assign n14409 = x95 & n70241 ;
  assign n70242 = ~n13993 ;
  assign n14410 = n70242 & n14409 ;
  assign n14411 = n14000 | n14410 ;
  assign n14412 = n14408 | n14411 ;
  assign n70243 = ~n14000 ;
  assign n14416 = n70243 & n14412 ;
  assign n14417 = n14415 | n14416 ;
  assign n70244 = ~n13992 ;
  assign n14418 = n70244 & n14417 ;
  assign n70245 = ~n13982 ;
  assign n14419 = x97 & n70245 ;
  assign n70246 = ~n13977 ;
  assign n14420 = n70246 & n14419 ;
  assign n14421 = n13984 | n14420 ;
  assign n14422 = n14418 | n14421 ;
  assign n70247 = ~n13984 ;
  assign n14426 = n70247 & n14422 ;
  assign n14427 = n14425 | n14426 ;
  assign n70248 = ~n13976 ;
  assign n14428 = n70248 & n14427 ;
  assign n70249 = ~n13966 ;
  assign n14429 = x99 & n70249 ;
  assign n70250 = ~n13961 ;
  assign n14430 = n70250 & n14429 ;
  assign n14431 = n13968 | n14430 ;
  assign n14432 = n14428 | n14431 ;
  assign n70251 = ~n13968 ;
  assign n14436 = n70251 & n14432 ;
  assign n14437 = n14435 | n14436 ;
  assign n70252 = ~n13960 ;
  assign n14438 = n70252 & n14437 ;
  assign n70253 = ~n13950 ;
  assign n14439 = x101 & n70253 ;
  assign n70254 = ~n13945 ;
  assign n14440 = n70254 & n14439 ;
  assign n14441 = n13952 | n14440 ;
  assign n14442 = n14438 | n14441 ;
  assign n70255 = ~n13952 ;
  assign n14447 = n70255 & n14442 ;
  assign n14448 = n14445 | n14447 ;
  assign n70256 = ~n13944 ;
  assign n14449 = n70256 & n14448 ;
  assign n70257 = ~n13934 ;
  assign n14450 = x103 & n70257 ;
  assign n70258 = ~n13929 ;
  assign n14451 = n70258 & n14450 ;
  assign n14452 = n13936 | n14451 ;
  assign n14453 = n14449 | n14452 ;
  assign n70259 = ~n13936 ;
  assign n14457 = n70259 & n14453 ;
  assign n14458 = n14456 | n14457 ;
  assign n70260 = ~n13928 ;
  assign n14459 = n70260 & n14458 ;
  assign n70261 = ~n13811 ;
  assign n13817 = n70261 & n13816 ;
  assign n14460 = n13283 | n13816 ;
  assign n70262 = ~n14460 ;
  assign n14461 = n13921 & n70262 ;
  assign n14462 = n13817 | n14461 ;
  assign n14463 = n13821 | n14462 ;
  assign n70263 = ~n13274 ;
  assign n14464 = n70263 & n13821 ;
  assign n70264 = ~n14464 ;
  assign n14465 = n14463 & n70264 ;
  assign n14466 = n70176 & n14465 ;
  assign n152 = ~n13821 ;
  assign n14467 = n152 & n14462 ;
  assign n14468 = n13274 & n13821 ;
  assign n70266 = ~n14468 ;
  assign n14469 = x105 & n70266 ;
  assign n70267 = ~n14467 ;
  assign n14470 = n70267 & n14469 ;
  assign n14471 = n65444 | n65527 ;
  assign n14472 = n66858 | n14471 ;
  assign n14473 = n14470 | n14472 ;
  assign n14474 = n14466 | n14473 ;
  assign n14475 = n14459 | n14474 ;
  assign n14476 = n70059 & n14465 ;
  assign n70268 = ~n14476 ;
  assign n14477 = n14475 & n70268 ;
  assign n70269 = ~n14457 ;
  assign n14573 = n14456 & n70269 ;
  assign n14490 = n70060 & n14243 ;
  assign n70270 = ~n14490 ;
  assign n14491 = x23 & n70270 ;
  assign n14492 = n14249 | n14491 ;
  assign n14493 = x65 & n14492 ;
  assign n70271 = ~n14493 ;
  assign n14494 = n14253 & n70271 ;
  assign n14495 = n14255 | n14494 ;
  assign n14496 = n70183 & n14495 ;
  assign n14497 = n14261 | n14496 ;
  assign n14498 = n70184 & n14497 ;
  assign n14499 = n14266 | n14498 ;
  assign n14500 = n70187 & n14499 ;
  assign n14501 = n14270 | n14500 ;
  assign n14502 = n70188 & n14501 ;
  assign n14503 = n14276 | n14502 ;
  assign n14504 = n70191 & n14503 ;
  assign n14505 = n14280 | n14504 ;
  assign n14506 = n70192 & n14505 ;
  assign n14507 = n14286 | n14506 ;
  assign n14508 = n70195 & n14507 ;
  assign n14509 = n14290 | n14508 ;
  assign n14510 = n70196 & n14509 ;
  assign n14511 = n14296 | n14510 ;
  assign n14512 = n70199 & n14511 ;
  assign n14513 = n14301 | n14512 ;
  assign n14514 = n70200 & n14513 ;
  assign n14515 = n14307 | n14514 ;
  assign n14516 = n70203 & n14515 ;
  assign n14517 = n14312 | n14516 ;
  assign n14518 = n70204 & n14517 ;
  assign n14519 = n14318 | n14518 ;
  assign n14520 = n70207 & n14519 ;
  assign n14521 = n14323 | n14520 ;
  assign n14522 = n70208 & n14521 ;
  assign n14523 = n14329 | n14522 ;
  assign n14524 = n70211 & n14523 ;
  assign n14525 = n14333 | n14524 ;
  assign n14526 = n70212 & n14525 ;
  assign n14527 = n14340 | n14526 ;
  assign n14528 = n70215 & n14527 ;
  assign n14529 = n14344 | n14528 ;
  assign n14530 = n70216 & n14529 ;
  assign n14531 = n14350 | n14530 ;
  assign n14532 = n70219 & n14531 ;
  assign n14533 = n14354 | n14532 ;
  assign n14534 = n70220 & n14533 ;
  assign n14535 = n14360 | n14534 ;
  assign n14536 = n70223 & n14535 ;
  assign n14537 = n14364 | n14536 ;
  assign n14538 = n70224 & n14537 ;
  assign n14539 = n14370 | n14538 ;
  assign n14540 = n70227 & n14539 ;
  assign n14541 = n14375 | n14540 ;
  assign n14542 = n70228 & n14541 ;
  assign n14543 = n14381 | n14542 ;
  assign n14544 = n70231 & n14543 ;
  assign n14545 = n14385 | n14544 ;
  assign n14546 = n70232 & n14545 ;
  assign n14547 = n14391 | n14546 ;
  assign n14548 = n70235 & n14547 ;
  assign n14549 = n14395 | n14548 ;
  assign n14550 = n70236 & n14549 ;
  assign n14551 = n14401 | n14550 ;
  assign n14552 = n70239 & n14551 ;
  assign n14553 = n14405 | n14552 ;
  assign n14554 = n70240 & n14553 ;
  assign n14555 = n14411 | n14554 ;
  assign n14556 = n70243 & n14555 ;
  assign n14557 = n14415 | n14556 ;
  assign n14558 = n70244 & n14557 ;
  assign n14559 = n14421 | n14558 ;
  assign n14560 = n70247 & n14559 ;
  assign n14561 = n14425 | n14560 ;
  assign n14562 = n70248 & n14561 ;
  assign n14563 = n14431 | n14562 ;
  assign n14564 = n70251 & n14563 ;
  assign n14565 = n14435 | n14564 ;
  assign n14566 = n70252 & n14565 ;
  assign n14567 = n14441 | n14566 ;
  assign n14568 = n70255 & n14567 ;
  assign n14569 = n14445 | n14568 ;
  assign n14570 = n70256 & n14569 ;
  assign n14571 = n14452 | n14570 ;
  assign n14574 = n13936 | n14456 ;
  assign n70272 = ~n14574 ;
  assign n14575 = n14571 & n70272 ;
  assign n14576 = n14573 | n14575 ;
  assign n151 = ~n14477 ;
  assign n14577 = n151 & n14576 ;
  assign n14578 = n13927 & n70268 ;
  assign n14579 = n14475 & n14578 ;
  assign n14580 = n14577 | n14579 ;
  assign n14479 = n13928 | n14470 ;
  assign n14480 = n14466 | n14479 ;
  assign n70274 = ~n14480 ;
  assign n14481 = n14458 & n70274 ;
  assign n14482 = n14466 | n14470 ;
  assign n70275 = ~n14459 ;
  assign n14483 = n70275 & n14482 ;
  assign n14484 = n14481 | n14483 ;
  assign n14485 = n151 & n14484 ;
  assign n14486 = n13820 & n14465 ;
  assign n14487 = n14475 & n14486 ;
  assign n14488 = n14485 | n14487 ;
  assign n70276 = ~x106 ;
  assign n14489 = n70276 & n14488 ;
  assign n14581 = n70176 & n14580 ;
  assign n70277 = ~n14570 ;
  assign n14582 = n14452 & n70277 ;
  assign n14583 = n13944 | n14452 ;
  assign n70278 = ~n14583 ;
  assign n14584 = n14448 & n70278 ;
  assign n14585 = n14582 | n14584 ;
  assign n14586 = n151 & n14585 ;
  assign n14587 = n13935 & n70268 ;
  assign n14588 = n14475 & n14587 ;
  assign n14589 = n14586 | n14588 ;
  assign n14590 = n69857 & n14589 ;
  assign n70279 = ~n14447 ;
  assign n14591 = n14445 & n70279 ;
  assign n14446 = n13952 | n14445 ;
  assign n70280 = ~n14446 ;
  assign n14592 = n14442 & n70280 ;
  assign n14593 = n14591 | n14592 ;
  assign n14594 = n151 & n14593 ;
  assign n14595 = n13943 & n70268 ;
  assign n14596 = n14475 & n14595 ;
  assign n14597 = n14594 | n14596 ;
  assign n14598 = n69656 & n14597 ;
  assign n70281 = ~n14566 ;
  assign n14599 = n14441 & n70281 ;
  assign n14600 = n13960 | n14441 ;
  assign n70282 = ~n14600 ;
  assign n14601 = n14437 & n70282 ;
  assign n14602 = n14599 | n14601 ;
  assign n14603 = n151 & n14602 ;
  assign n14604 = n13951 & n70268 ;
  assign n14605 = n14475 & n14604 ;
  assign n14606 = n14603 | n14605 ;
  assign n14607 = n69528 & n14606 ;
  assign n70283 = ~n14436 ;
  assign n14608 = n14435 & n70283 ;
  assign n14609 = n13968 | n14435 ;
  assign n70284 = ~n14609 ;
  assign n14610 = n14563 & n70284 ;
  assign n14611 = n14608 | n14610 ;
  assign n14612 = n151 & n14611 ;
  assign n14613 = n13959 & n70268 ;
  assign n14614 = n14475 & n14613 ;
  assign n14615 = n14612 | n14614 ;
  assign n14616 = n69261 & n14615 ;
  assign n70285 = ~n14562 ;
  assign n14617 = n14431 & n70285 ;
  assign n14618 = n13976 | n14431 ;
  assign n70286 = ~n14618 ;
  assign n14619 = n14427 & n70286 ;
  assign n14620 = n14617 | n14619 ;
  assign n14621 = n151 & n14620 ;
  assign n14622 = n13967 & n70268 ;
  assign n14623 = n14475 & n14622 ;
  assign n14624 = n14621 | n14623 ;
  assign n14625 = n69075 & n14624 ;
  assign n70287 = ~n14426 ;
  assign n14626 = n14425 & n70287 ;
  assign n14627 = n13984 | n14425 ;
  assign n70288 = ~n14627 ;
  assign n14628 = n14559 & n70288 ;
  assign n14629 = n14626 | n14628 ;
  assign n14630 = n151 & n14629 ;
  assign n14631 = n13975 & n70268 ;
  assign n14632 = n14475 & n14631 ;
  assign n14633 = n14630 | n14632 ;
  assign n14634 = n68993 & n14633 ;
  assign n70289 = ~n14558 ;
  assign n14635 = n14421 & n70289 ;
  assign n14636 = n13992 | n14421 ;
  assign n70290 = ~n14636 ;
  assign n14637 = n14417 & n70290 ;
  assign n14638 = n14635 | n14637 ;
  assign n14639 = n151 & n14638 ;
  assign n14640 = n13983 & n70268 ;
  assign n14641 = n14475 & n14640 ;
  assign n14642 = n14639 | n14641 ;
  assign n14643 = n68716 & n14642 ;
  assign n70291 = ~n14416 ;
  assign n14644 = n14415 & n70291 ;
  assign n14645 = n14000 | n14415 ;
  assign n70292 = ~n14645 ;
  assign n14646 = n14555 & n70292 ;
  assign n14647 = n14644 | n14646 ;
  assign n14648 = n151 & n14647 ;
  assign n14649 = n13991 & n70268 ;
  assign n14650 = n14475 & n14649 ;
  assign n14651 = n14648 | n14650 ;
  assign n14652 = n68545 & n14651 ;
  assign n70293 = ~n14554 ;
  assign n14653 = n14411 & n70293 ;
  assign n14654 = n14008 | n14411 ;
  assign n70294 = ~n14654 ;
  assign n14655 = n14407 & n70294 ;
  assign n14656 = n14653 | n14655 ;
  assign n14657 = n151 & n14656 ;
  assign n14658 = n13999 & n70268 ;
  assign n14659 = n14475 & n14658 ;
  assign n14660 = n14657 | n14659 ;
  assign n14661 = n68438 & n14660 ;
  assign n70295 = ~n14406 ;
  assign n14662 = n14405 & n70295 ;
  assign n14663 = n14016 | n14405 ;
  assign n70296 = ~n14663 ;
  assign n14664 = n14551 & n70296 ;
  assign n14665 = n14662 | n14664 ;
  assign n14666 = n151 & n14665 ;
  assign n14667 = n14007 & n70268 ;
  assign n14668 = n14475 & n14667 ;
  assign n14669 = n14666 | n14668 ;
  assign n14670 = n68214 & n14669 ;
  assign n70297 = ~n14550 ;
  assign n14671 = n14401 & n70297 ;
  assign n14672 = n14024 | n14401 ;
  assign n70298 = ~n14672 ;
  assign n14673 = n14397 & n70298 ;
  assign n14674 = n14671 | n14673 ;
  assign n14675 = n151 & n14674 ;
  assign n14676 = n14015 & n70268 ;
  assign n14677 = n14475 & n14676 ;
  assign n14678 = n14675 | n14677 ;
  assign n14679 = n68058 & n14678 ;
  assign n70299 = ~n14396 ;
  assign n14680 = n14395 & n70299 ;
  assign n14681 = n14032 | n14395 ;
  assign n70300 = ~n14681 ;
  assign n14682 = n14547 & n70300 ;
  assign n14683 = n14680 | n14682 ;
  assign n14684 = n151 & n14683 ;
  assign n14685 = n14023 & n70268 ;
  assign n14686 = n14475 & n14685 ;
  assign n14687 = n14684 | n14686 ;
  assign n14688 = n67986 & n14687 ;
  assign n70301 = ~n14546 ;
  assign n14689 = n14391 & n70301 ;
  assign n14690 = n14040 | n14391 ;
  assign n70302 = ~n14690 ;
  assign n14691 = n14387 & n70302 ;
  assign n14692 = n14689 | n14691 ;
  assign n14693 = n151 & n14692 ;
  assign n14694 = n14031 & n70268 ;
  assign n14695 = n14475 & n14694 ;
  assign n14696 = n14693 | n14695 ;
  assign n14697 = n67763 & n14696 ;
  assign n70303 = ~n14386 ;
  assign n14698 = n14385 & n70303 ;
  assign n14699 = n14048 | n14385 ;
  assign n70304 = ~n14699 ;
  assign n14700 = n14543 & n70304 ;
  assign n14701 = n14698 | n14700 ;
  assign n14702 = n151 & n14701 ;
  assign n14703 = n14039 & n70268 ;
  assign n14704 = n14475 & n14703 ;
  assign n14705 = n14702 | n14704 ;
  assign n14706 = n67622 & n14705 ;
  assign n70305 = ~n14542 ;
  assign n14707 = n14381 & n70305 ;
  assign n14708 = n14056 | n14381 ;
  assign n70306 = ~n14708 ;
  assign n14709 = n14377 & n70306 ;
  assign n14710 = n14707 | n14709 ;
  assign n14711 = n151 & n14710 ;
  assign n14712 = n14047 & n70268 ;
  assign n14713 = n14475 & n14712 ;
  assign n14714 = n14711 | n14713 ;
  assign n14715 = n67531 & n14714 ;
  assign n70307 = ~n14376 ;
  assign n14716 = n14375 & n70307 ;
  assign n14717 = n14064 | n14375 ;
  assign n70308 = ~n14717 ;
  assign n14718 = n14539 & n70308 ;
  assign n14719 = n14716 | n14718 ;
  assign n14720 = n151 & n14719 ;
  assign n14721 = n14055 & n70268 ;
  assign n14722 = n14475 & n14721 ;
  assign n14723 = n14720 | n14722 ;
  assign n14724 = n67348 & n14723 ;
  assign n70309 = ~n14538 ;
  assign n14725 = n14370 & n70309 ;
  assign n14371 = n14072 | n14370 ;
  assign n70310 = ~n14371 ;
  assign n14726 = n70310 & n14537 ;
  assign n14727 = n14725 | n14726 ;
  assign n14728 = n151 & n14727 ;
  assign n14729 = n14063 & n70268 ;
  assign n14730 = n14475 & n14729 ;
  assign n14731 = n14728 | n14730 ;
  assign n14732 = n67222 & n14731 ;
  assign n70311 = ~n14365 ;
  assign n14733 = n14364 & n70311 ;
  assign n14734 = n14080 | n14364 ;
  assign n70312 = ~n14734 ;
  assign n14735 = n14535 & n70312 ;
  assign n14736 = n14733 | n14735 ;
  assign n14737 = n151 & n14736 ;
  assign n14738 = n14071 & n70268 ;
  assign n14739 = n14475 & n14738 ;
  assign n14740 = n14737 | n14739 ;
  assign n14741 = n67164 & n14740 ;
  assign n70313 = ~n14534 ;
  assign n14742 = n14360 & n70313 ;
  assign n14743 = n14088 | n14360 ;
  assign n70314 = ~n14743 ;
  assign n14744 = n14356 & n70314 ;
  assign n14745 = n14742 | n14744 ;
  assign n14746 = n151 & n14745 ;
  assign n14747 = n14079 & n70268 ;
  assign n14748 = n14475 & n14747 ;
  assign n14749 = n14746 | n14748 ;
  assign n14750 = n66979 & n14749 ;
  assign n70315 = ~n14355 ;
  assign n14751 = n14354 & n70315 ;
  assign n14752 = n14096 | n14354 ;
  assign n70316 = ~n14752 ;
  assign n14753 = n14531 & n70316 ;
  assign n14754 = n14751 | n14753 ;
  assign n14755 = n151 & n14754 ;
  assign n14756 = n14087 & n70268 ;
  assign n14757 = n14475 & n14756 ;
  assign n14758 = n14755 | n14757 ;
  assign n14759 = n66868 & n14758 ;
  assign n70317 = ~n14530 ;
  assign n14760 = n14350 & n70317 ;
  assign n14761 = n14104 | n14350 ;
  assign n70318 = ~n14761 ;
  assign n14762 = n14346 & n70318 ;
  assign n14763 = n14760 | n14762 ;
  assign n14764 = n151 & n14763 ;
  assign n14765 = n14095 & n70268 ;
  assign n14766 = n14475 & n14765 ;
  assign n14767 = n14764 | n14766 ;
  assign n14768 = n66797 & n14767 ;
  assign n70319 = ~n14345 ;
  assign n14769 = n14344 & n70319 ;
  assign n14770 = n14112 | n14344 ;
  assign n70320 = ~n14770 ;
  assign n14771 = n14527 & n70320 ;
  assign n14772 = n14769 | n14771 ;
  assign n14773 = n151 & n14772 ;
  assign n14774 = n14103 & n70268 ;
  assign n14775 = n14475 & n14774 ;
  assign n14776 = n14773 | n14775 ;
  assign n14777 = n66654 & n14776 ;
  assign n70321 = ~n14526 ;
  assign n14778 = n14340 & n70321 ;
  assign n14779 = n14120 | n14340 ;
  assign n70322 = ~n14779 ;
  assign n14780 = n14336 & n70322 ;
  assign n14781 = n14778 | n14780 ;
  assign n14782 = n151 & n14781 ;
  assign n14783 = n14111 & n70268 ;
  assign n14784 = n14475 & n14783 ;
  assign n14785 = n14782 | n14784 ;
  assign n14786 = n66560 & n14785 ;
  assign n70323 = ~n14335 ;
  assign n14787 = n14333 & n70323 ;
  assign n14334 = n14128 | n14333 ;
  assign n70324 = ~n14334 ;
  assign n14788 = n14330 & n70324 ;
  assign n14789 = n14787 | n14788 ;
  assign n14790 = n151 & n14789 ;
  assign n14791 = n14119 & n70268 ;
  assign n14792 = n14475 & n14791 ;
  assign n14793 = n14790 | n14792 ;
  assign n14794 = n66505 & n14793 ;
  assign n70325 = ~n14522 ;
  assign n14795 = n14329 & n70325 ;
  assign n14796 = n14136 | n14329 ;
  assign n70326 = ~n14796 ;
  assign n14797 = n14325 & n70326 ;
  assign n14798 = n14795 | n14797 ;
  assign n14799 = n151 & n14798 ;
  assign n14800 = n14127 & n70268 ;
  assign n14801 = n14475 & n14800 ;
  assign n14802 = n14799 | n14801 ;
  assign n14803 = n66379 & n14802 ;
  assign n70327 = ~n14324 ;
  assign n14804 = n14323 & n70327 ;
  assign n14805 = n14144 | n14323 ;
  assign n70328 = ~n14805 ;
  assign n14806 = n14519 & n70328 ;
  assign n14807 = n14804 | n14806 ;
  assign n14808 = n151 & n14807 ;
  assign n14809 = n14135 & n70268 ;
  assign n14810 = n14475 & n14809 ;
  assign n14811 = n14808 | n14810 ;
  assign n14812 = n66299 & n14811 ;
  assign n70329 = ~n14518 ;
  assign n14813 = n14318 & n70329 ;
  assign n14319 = n14152 | n14318 ;
  assign n70330 = ~n14319 ;
  assign n14814 = n70330 & n14517 ;
  assign n14815 = n14813 | n14814 ;
  assign n14816 = n151 & n14815 ;
  assign n14817 = n14143 & n70268 ;
  assign n14818 = n14475 & n14817 ;
  assign n14819 = n14816 | n14818 ;
  assign n14820 = n66244 & n14819 ;
  assign n70331 = ~n14313 ;
  assign n14821 = n14312 & n70331 ;
  assign n14822 = n14160 | n14312 ;
  assign n70332 = ~n14822 ;
  assign n14823 = n14515 & n70332 ;
  assign n14824 = n14821 | n14823 ;
  assign n14825 = n151 & n14824 ;
  assign n14826 = n14151 & n70268 ;
  assign n14827 = n14475 & n14826 ;
  assign n14828 = n14825 | n14827 ;
  assign n14829 = n66145 & n14828 ;
  assign n70333 = ~n14514 ;
  assign n14830 = n14307 & n70333 ;
  assign n14308 = n14168 | n14307 ;
  assign n70334 = ~n14308 ;
  assign n14831 = n70334 & n14513 ;
  assign n14832 = n14830 | n14831 ;
  assign n14833 = n151 & n14832 ;
  assign n14834 = n14159 & n70268 ;
  assign n14835 = n14475 & n14834 ;
  assign n14836 = n14833 | n14835 ;
  assign n14837 = n66081 & n14836 ;
  assign n70335 = ~n14302 ;
  assign n14838 = n14301 & n70335 ;
  assign n14839 = n14176 | n14301 ;
  assign n70336 = ~n14839 ;
  assign n14840 = n14511 & n70336 ;
  assign n14841 = n14838 | n14840 ;
  assign n14842 = n151 & n14841 ;
  assign n14843 = n14167 & n70268 ;
  assign n14844 = n14475 & n14843 ;
  assign n14845 = n14842 | n14844 ;
  assign n14846 = n66043 & n14845 ;
  assign n70337 = ~n14510 ;
  assign n14847 = n14296 & n70337 ;
  assign n14297 = n14184 | n14296 ;
  assign n70338 = ~n14297 ;
  assign n14848 = n70338 & n14509 ;
  assign n14849 = n14847 | n14848 ;
  assign n14850 = n151 & n14849 ;
  assign n14851 = n14175 & n70268 ;
  assign n14852 = n14475 & n14851 ;
  assign n14853 = n14850 | n14852 ;
  assign n14854 = n65960 & n14853 ;
  assign n70339 = ~n14291 ;
  assign n14855 = n14290 & n70339 ;
  assign n14856 = n14192 | n14290 ;
  assign n70340 = ~n14856 ;
  assign n14857 = n14507 & n70340 ;
  assign n14858 = n14855 | n14857 ;
  assign n14859 = n151 & n14858 ;
  assign n14860 = n14183 & n70268 ;
  assign n14861 = n14475 & n14860 ;
  assign n14862 = n14859 | n14861 ;
  assign n14863 = n65909 & n14862 ;
  assign n70341 = ~n14506 ;
  assign n14864 = n14286 & n70341 ;
  assign n14865 = n14200 | n14286 ;
  assign n70342 = ~n14865 ;
  assign n14866 = n14282 & n70342 ;
  assign n14867 = n14864 | n14866 ;
  assign n14868 = n151 & n14867 ;
  assign n14869 = n14191 & n70268 ;
  assign n14870 = n14475 & n14869 ;
  assign n14871 = n14868 | n14870 ;
  assign n14872 = n65877 & n14871 ;
  assign n70343 = ~n14281 ;
  assign n14873 = n14280 & n70343 ;
  assign n14874 = n14209 | n14280 ;
  assign n70344 = ~n14874 ;
  assign n14875 = n14503 & n70344 ;
  assign n14876 = n14873 | n14875 ;
  assign n14877 = n151 & n14876 ;
  assign n14878 = n14199 & n70268 ;
  assign n14879 = n14475 & n14878 ;
  assign n14880 = n14877 | n14879 ;
  assign n14881 = n65820 & n14880 ;
  assign n70345 = ~n14502 ;
  assign n14882 = n14276 & n70345 ;
  assign n14883 = n14217 | n14276 ;
  assign n70346 = ~n14883 ;
  assign n14884 = n14272 & n70346 ;
  assign n14885 = n14882 | n14884 ;
  assign n14886 = n151 & n14885 ;
  assign n14887 = n14208 & n70268 ;
  assign n14888 = n14475 & n14887 ;
  assign n14889 = n14886 | n14888 ;
  assign n14890 = n65791 & n14889 ;
  assign n70347 = ~n14271 ;
  assign n14891 = n14270 & n70347 ;
  assign n14892 = n14227 | n14270 ;
  assign n70348 = ~n14892 ;
  assign n14893 = n14499 & n70348 ;
  assign n14894 = n14891 | n14893 ;
  assign n14895 = n151 & n14894 ;
  assign n14896 = n14216 & n70268 ;
  assign n14897 = n14475 & n14896 ;
  assign n14898 = n14895 | n14897 ;
  assign n14899 = n65772 & n14898 ;
  assign n70349 = ~n14498 ;
  assign n14901 = n14266 & n70349 ;
  assign n14900 = n14239 | n14266 ;
  assign n70350 = ~n14900 ;
  assign n14902 = n14497 & n70350 ;
  assign n14903 = n14901 | n14902 ;
  assign n14904 = n151 & n14903 ;
  assign n14905 = n14225 & n70268 ;
  assign n14906 = n14475 & n14905 ;
  assign n14907 = n14904 | n14906 ;
  assign n14908 = n65746 & n14907 ;
  assign n70351 = ~n14262 ;
  assign n14910 = n14261 & n70351 ;
  assign n14909 = n14257 | n14261 ;
  assign n70352 = ~n14909 ;
  assign n14911 = n14256 & n70352 ;
  assign n14912 = n14910 | n14911 ;
  assign n14913 = n151 & n14912 ;
  assign n14914 = n14238 & n70268 ;
  assign n14915 = n14475 & n14914 ;
  assign n14916 = n14913 | n14915 ;
  assign n14917 = n65721 & n14916 ;
  assign n14918 = n14253 & n14255 ;
  assign n14919 = n70181 & n14918 ;
  assign n70353 = ~n14919 ;
  assign n14920 = n14256 & n70353 ;
  assign n14921 = n151 & n14920 ;
  assign n14922 = n14250 & n70268 ;
  assign n14923 = n14475 & n14922 ;
  assign n14924 = n14921 | n14923 ;
  assign n14925 = n65686 & n14924 ;
  assign n14478 = n14255 & n151 ;
  assign n14926 = x64 & n151 ;
  assign n70354 = ~n14926 ;
  assign n14927 = x22 & n70354 ;
  assign n14928 = n14478 | n14927 ;
  assign n14941 = n65670 & n14928 ;
  assign n14572 = n70259 & n14571 ;
  assign n14929 = n14456 | n14572 ;
  assign n14930 = n70260 & n14929 ;
  assign n14931 = n14474 | n14930 ;
  assign n14932 = n70268 & n14931 ;
  assign n70355 = ~n14932 ;
  assign n14933 = x64 & n70355 ;
  assign n70356 = ~n14933 ;
  assign n14934 = x22 & n70356 ;
  assign n14935 = n14478 | n14934 ;
  assign n14936 = x65 & n14935 ;
  assign n14937 = x65 | n14478 ;
  assign n14938 = n14934 | n14937 ;
  assign n70357 = ~n14936 ;
  assign n14939 = n70357 & n14938 ;
  assign n70358 = ~x21 ;
  assign n14940 = n70358 & x64 ;
  assign n14942 = n14939 | n14940 ;
  assign n70359 = ~n14941 ;
  assign n14943 = n70359 & n14942 ;
  assign n70360 = ~n14923 ;
  assign n14944 = x66 & n70360 ;
  assign n70361 = ~n14921 ;
  assign n14945 = n70361 & n14944 ;
  assign n14946 = n14925 | n14945 ;
  assign n14947 = n14943 | n14946 ;
  assign n70362 = ~n14925 ;
  assign n14948 = n70362 & n14947 ;
  assign n70363 = ~n14915 ;
  assign n14949 = x67 & n70363 ;
  assign n70364 = ~n14913 ;
  assign n14950 = n70364 & n14949 ;
  assign n14951 = n14917 | n14950 ;
  assign n14952 = n14948 | n14951 ;
  assign n70365 = ~n14917 ;
  assign n14953 = n70365 & n14952 ;
  assign n70366 = ~n14906 ;
  assign n14954 = x68 & n70366 ;
  assign n70367 = ~n14904 ;
  assign n14955 = n70367 & n14954 ;
  assign n14956 = n14908 | n14955 ;
  assign n14957 = n14953 | n14956 ;
  assign n70368 = ~n14908 ;
  assign n14958 = n70368 & n14957 ;
  assign n70369 = ~n14897 ;
  assign n14959 = x69 & n70369 ;
  assign n70370 = ~n14895 ;
  assign n14960 = n70370 & n14959 ;
  assign n14961 = n14899 | n14960 ;
  assign n14962 = n14958 | n14961 ;
  assign n70371 = ~n14899 ;
  assign n14963 = n70371 & n14962 ;
  assign n70372 = ~n14888 ;
  assign n14964 = x70 & n70372 ;
  assign n70373 = ~n14886 ;
  assign n14965 = n70373 & n14964 ;
  assign n14966 = n14963 | n14965 ;
  assign n70374 = ~n14890 ;
  assign n14967 = n70374 & n14966 ;
  assign n70375 = ~n14879 ;
  assign n14968 = x71 & n70375 ;
  assign n70376 = ~n14877 ;
  assign n14969 = n70376 & n14968 ;
  assign n14970 = n14881 | n14969 ;
  assign n14971 = n14967 | n14970 ;
  assign n70377 = ~n14881 ;
  assign n14972 = n70377 & n14971 ;
  assign n70378 = ~n14870 ;
  assign n14973 = x72 & n70378 ;
  assign n70379 = ~n14868 ;
  assign n14974 = n70379 & n14973 ;
  assign n14975 = n14872 | n14974 ;
  assign n14977 = n14972 | n14975 ;
  assign n70380 = ~n14872 ;
  assign n14978 = n70380 & n14977 ;
  assign n70381 = ~n14861 ;
  assign n14979 = x73 & n70381 ;
  assign n70382 = ~n14859 ;
  assign n14980 = n70382 & n14979 ;
  assign n14981 = n14863 | n14980 ;
  assign n14982 = n14978 | n14981 ;
  assign n70383 = ~n14863 ;
  assign n14983 = n70383 & n14982 ;
  assign n70384 = ~n14852 ;
  assign n14984 = x74 & n70384 ;
  assign n70385 = ~n14850 ;
  assign n14985 = n70385 & n14984 ;
  assign n14986 = n14854 | n14985 ;
  assign n14988 = n14983 | n14986 ;
  assign n70386 = ~n14854 ;
  assign n14989 = n70386 & n14988 ;
  assign n70387 = ~n14844 ;
  assign n14990 = x75 & n70387 ;
  assign n70388 = ~n14842 ;
  assign n14991 = n70388 & n14990 ;
  assign n14992 = n14846 | n14991 ;
  assign n14993 = n14989 | n14992 ;
  assign n70389 = ~n14846 ;
  assign n14994 = n70389 & n14993 ;
  assign n70390 = ~n14835 ;
  assign n14995 = x76 & n70390 ;
  assign n70391 = ~n14833 ;
  assign n14996 = n70391 & n14995 ;
  assign n14997 = n14837 | n14996 ;
  assign n14999 = n14994 | n14997 ;
  assign n70392 = ~n14837 ;
  assign n15000 = n70392 & n14999 ;
  assign n70393 = ~n14827 ;
  assign n15001 = x77 & n70393 ;
  assign n70394 = ~n14825 ;
  assign n15002 = n70394 & n15001 ;
  assign n15003 = n14829 | n15002 ;
  assign n15004 = n15000 | n15003 ;
  assign n70395 = ~n14829 ;
  assign n15005 = n70395 & n15004 ;
  assign n70396 = ~n14818 ;
  assign n15006 = x78 & n70396 ;
  assign n70397 = ~n14816 ;
  assign n15007 = n70397 & n15006 ;
  assign n15008 = n14820 | n15007 ;
  assign n15010 = n15005 | n15008 ;
  assign n70398 = ~n14820 ;
  assign n15011 = n70398 & n15010 ;
  assign n70399 = ~n14810 ;
  assign n15012 = x79 & n70399 ;
  assign n70400 = ~n14808 ;
  assign n15013 = n70400 & n15012 ;
  assign n15014 = n14812 | n15013 ;
  assign n15015 = n15011 | n15014 ;
  assign n70401 = ~n14812 ;
  assign n15016 = n70401 & n15015 ;
  assign n70402 = ~n14801 ;
  assign n15017 = x80 & n70402 ;
  assign n70403 = ~n14799 ;
  assign n15018 = n70403 & n15017 ;
  assign n15019 = n14803 | n15018 ;
  assign n15021 = n15016 | n15019 ;
  assign n70404 = ~n14803 ;
  assign n15022 = n70404 & n15021 ;
  assign n70405 = ~n14792 ;
  assign n15023 = x81 & n70405 ;
  assign n70406 = ~n14790 ;
  assign n15024 = n70406 & n15023 ;
  assign n15025 = n14794 | n15024 ;
  assign n15026 = n15022 | n15025 ;
  assign n70407 = ~n14794 ;
  assign n15027 = n70407 & n15026 ;
  assign n70408 = ~n14784 ;
  assign n15028 = x82 & n70408 ;
  assign n70409 = ~n14782 ;
  assign n15029 = n70409 & n15028 ;
  assign n15030 = n14786 | n15029 ;
  assign n15032 = n15027 | n15030 ;
  assign n70410 = ~n14786 ;
  assign n15033 = n70410 & n15032 ;
  assign n70411 = ~n14775 ;
  assign n15034 = x83 & n70411 ;
  assign n70412 = ~n14773 ;
  assign n15035 = n70412 & n15034 ;
  assign n15036 = n14777 | n15035 ;
  assign n15037 = n15033 | n15036 ;
  assign n70413 = ~n14777 ;
  assign n15038 = n70413 & n15037 ;
  assign n70414 = ~n14766 ;
  assign n15039 = x84 & n70414 ;
  assign n70415 = ~n14764 ;
  assign n15040 = n70415 & n15039 ;
  assign n15041 = n14768 | n15040 ;
  assign n15043 = n15038 | n15041 ;
  assign n70416 = ~n14768 ;
  assign n15044 = n70416 & n15043 ;
  assign n70417 = ~n14757 ;
  assign n15045 = x85 & n70417 ;
  assign n70418 = ~n14755 ;
  assign n15046 = n70418 & n15045 ;
  assign n15047 = n14759 | n15046 ;
  assign n15048 = n15044 | n15047 ;
  assign n70419 = ~n14759 ;
  assign n15049 = n70419 & n15048 ;
  assign n70420 = ~n14748 ;
  assign n15050 = x86 & n70420 ;
  assign n70421 = ~n14746 ;
  assign n15051 = n70421 & n15050 ;
  assign n15052 = n14750 | n15051 ;
  assign n15054 = n15049 | n15052 ;
  assign n70422 = ~n14750 ;
  assign n15055 = n70422 & n15054 ;
  assign n70423 = ~n14739 ;
  assign n15056 = x87 & n70423 ;
  assign n70424 = ~n14737 ;
  assign n15057 = n70424 & n15056 ;
  assign n15058 = n14741 | n15057 ;
  assign n15059 = n15055 | n15058 ;
  assign n70425 = ~n14741 ;
  assign n15060 = n70425 & n15059 ;
  assign n70426 = ~n14730 ;
  assign n15061 = x88 & n70426 ;
  assign n70427 = ~n14728 ;
  assign n15062 = n70427 & n15061 ;
  assign n15063 = n14732 | n15062 ;
  assign n15065 = n15060 | n15063 ;
  assign n70428 = ~n14732 ;
  assign n15066 = n70428 & n15065 ;
  assign n70429 = ~n14722 ;
  assign n15067 = x89 & n70429 ;
  assign n70430 = ~n14720 ;
  assign n15068 = n70430 & n15067 ;
  assign n15069 = n14724 | n15068 ;
  assign n15070 = n15066 | n15069 ;
  assign n70431 = ~n14724 ;
  assign n15071 = n70431 & n15070 ;
  assign n70432 = ~n14713 ;
  assign n15072 = x90 & n70432 ;
  assign n70433 = ~n14711 ;
  assign n15073 = n70433 & n15072 ;
  assign n15074 = n14715 | n15073 ;
  assign n15076 = n15071 | n15074 ;
  assign n70434 = ~n14715 ;
  assign n15077 = n70434 & n15076 ;
  assign n70435 = ~n14704 ;
  assign n15078 = x91 & n70435 ;
  assign n70436 = ~n14702 ;
  assign n15079 = n70436 & n15078 ;
  assign n15080 = n14706 | n15079 ;
  assign n15081 = n15077 | n15080 ;
  assign n70437 = ~n14706 ;
  assign n15082 = n70437 & n15081 ;
  assign n70438 = ~n14695 ;
  assign n15083 = x92 & n70438 ;
  assign n70439 = ~n14693 ;
  assign n15084 = n70439 & n15083 ;
  assign n15085 = n14697 | n15084 ;
  assign n15087 = n15082 | n15085 ;
  assign n70440 = ~n14697 ;
  assign n15088 = n70440 & n15087 ;
  assign n70441 = ~n14686 ;
  assign n15089 = x93 & n70441 ;
  assign n70442 = ~n14684 ;
  assign n15090 = n70442 & n15089 ;
  assign n15091 = n14688 | n15090 ;
  assign n15092 = n15088 | n15091 ;
  assign n70443 = ~n14688 ;
  assign n15093 = n70443 & n15092 ;
  assign n70444 = ~n14677 ;
  assign n15094 = x94 & n70444 ;
  assign n70445 = ~n14675 ;
  assign n15095 = n70445 & n15094 ;
  assign n15096 = n14679 | n15095 ;
  assign n15098 = n15093 | n15096 ;
  assign n70446 = ~n14679 ;
  assign n15099 = n70446 & n15098 ;
  assign n70447 = ~n14668 ;
  assign n15100 = x95 & n70447 ;
  assign n70448 = ~n14666 ;
  assign n15101 = n70448 & n15100 ;
  assign n15102 = n14670 | n15101 ;
  assign n15103 = n15099 | n15102 ;
  assign n70449 = ~n14670 ;
  assign n15104 = n70449 & n15103 ;
  assign n70450 = ~n14659 ;
  assign n15105 = x96 & n70450 ;
  assign n70451 = ~n14657 ;
  assign n15106 = n70451 & n15105 ;
  assign n15107 = n14661 | n15106 ;
  assign n15109 = n15104 | n15107 ;
  assign n70452 = ~n14661 ;
  assign n15110 = n70452 & n15109 ;
  assign n70453 = ~n14650 ;
  assign n15111 = x97 & n70453 ;
  assign n70454 = ~n14648 ;
  assign n15112 = n70454 & n15111 ;
  assign n15113 = n14652 | n15112 ;
  assign n15114 = n15110 | n15113 ;
  assign n70455 = ~n14652 ;
  assign n15115 = n70455 & n15114 ;
  assign n70456 = ~n14641 ;
  assign n15116 = x98 & n70456 ;
  assign n70457 = ~n14639 ;
  assign n15117 = n70457 & n15116 ;
  assign n15118 = n14643 | n15117 ;
  assign n15120 = n15115 | n15118 ;
  assign n70458 = ~n14643 ;
  assign n15121 = n70458 & n15120 ;
  assign n70459 = ~n14632 ;
  assign n15122 = x99 & n70459 ;
  assign n70460 = ~n14630 ;
  assign n15123 = n70460 & n15122 ;
  assign n15124 = n14634 | n15123 ;
  assign n15125 = n15121 | n15124 ;
  assign n70461 = ~n14634 ;
  assign n15126 = n70461 & n15125 ;
  assign n70462 = ~n14623 ;
  assign n15127 = x100 & n70462 ;
  assign n70463 = ~n14621 ;
  assign n15128 = n70463 & n15127 ;
  assign n15129 = n14625 | n15128 ;
  assign n15131 = n15126 | n15129 ;
  assign n70464 = ~n14625 ;
  assign n15132 = n70464 & n15131 ;
  assign n70465 = ~n14614 ;
  assign n15133 = x101 & n70465 ;
  assign n70466 = ~n14612 ;
  assign n15134 = n70466 & n15133 ;
  assign n15135 = n14616 | n15134 ;
  assign n15136 = n15132 | n15135 ;
  assign n70467 = ~n14616 ;
  assign n15137 = n70467 & n15136 ;
  assign n70468 = ~n14605 ;
  assign n15138 = x102 & n70468 ;
  assign n70469 = ~n14603 ;
  assign n15139 = n70469 & n15138 ;
  assign n15140 = n14607 | n15139 ;
  assign n15142 = n15137 | n15140 ;
  assign n70470 = ~n14607 ;
  assign n15143 = n70470 & n15142 ;
  assign n70471 = ~n14596 ;
  assign n15144 = x103 & n70471 ;
  assign n70472 = ~n14594 ;
  assign n15145 = n70472 & n15144 ;
  assign n15146 = n14598 | n15145 ;
  assign n15147 = n15143 | n15146 ;
  assign n70473 = ~n14598 ;
  assign n15148 = n70473 & n15147 ;
  assign n70474 = ~n14588 ;
  assign n15149 = x104 & n70474 ;
  assign n70475 = ~n14586 ;
  assign n15150 = n70475 & n15149 ;
  assign n15151 = n14590 | n15150 ;
  assign n15153 = n15148 | n15151 ;
  assign n70476 = ~n14590 ;
  assign n15154 = n70476 & n15153 ;
  assign n70477 = ~n14579 ;
  assign n15155 = x105 & n70477 ;
  assign n70478 = ~n14577 ;
  assign n15156 = n70478 & n15155 ;
  assign n15157 = n14581 | n15156 ;
  assign n15158 = n15154 | n15157 ;
  assign n70479 = ~n14581 ;
  assign n15159 = n70479 & n15158 ;
  assign n70480 = ~n14487 ;
  assign n15160 = x106 & n70480 ;
  assign n70481 = ~n14485 ;
  assign n15161 = n70481 & n15160 ;
  assign n15162 = n14489 | n15161 ;
  assign n15164 = n15159 | n15162 ;
  assign n70482 = ~n14489 ;
  assign n15165 = n70482 & n15164 ;
  assign n15166 = n289 | n291 ;
  assign n15167 = n279 | n15166 ;
  assign n15168 = n15165 | n15167 ;
  assign n15169 = n14580 & n15168 ;
  assign n15170 = x65 & n14928 ;
  assign n70483 = ~n15170 ;
  assign n15171 = n14938 & n70483 ;
  assign n15172 = n14940 | n15171 ;
  assign n15173 = n70359 & n15172 ;
  assign n15174 = n14946 | n15173 ;
  assign n15175 = n70362 & n15174 ;
  assign n15177 = n14951 | n15175 ;
  assign n15178 = n70365 & n15177 ;
  assign n15180 = n14956 | n15178 ;
  assign n15181 = n70368 & n15180 ;
  assign n15182 = n14960 | n15181 ;
  assign n15184 = n70371 & n15182 ;
  assign n15185 = n14890 | n14965 ;
  assign n15187 = n15184 | n15185 ;
  assign n15188 = n70374 & n15187 ;
  assign n15189 = n14970 | n15188 ;
  assign n15191 = n70377 & n15189 ;
  assign n15192 = n14975 | n15191 ;
  assign n15193 = n70380 & n15192 ;
  assign n15194 = n14981 | n15193 ;
  assign n15196 = n70383 & n15194 ;
  assign n15197 = n14986 | n15196 ;
  assign n15198 = n70386 & n15197 ;
  assign n15199 = n14992 | n15198 ;
  assign n15201 = n70389 & n15199 ;
  assign n15202 = n14997 | n15201 ;
  assign n15203 = n70392 & n15202 ;
  assign n15204 = n15003 | n15203 ;
  assign n15206 = n70395 & n15204 ;
  assign n15207 = n15008 | n15206 ;
  assign n15208 = n70398 & n15207 ;
  assign n15209 = n15014 | n15208 ;
  assign n15211 = n70401 & n15209 ;
  assign n15212 = n15019 | n15211 ;
  assign n15213 = n70404 & n15212 ;
  assign n15214 = n15025 | n15213 ;
  assign n15216 = n70407 & n15214 ;
  assign n15217 = n15030 | n15216 ;
  assign n15218 = n70410 & n15217 ;
  assign n15219 = n15036 | n15218 ;
  assign n15221 = n70413 & n15219 ;
  assign n15222 = n15041 | n15221 ;
  assign n15223 = n70416 & n15222 ;
  assign n15224 = n15047 | n15223 ;
  assign n15226 = n70419 & n15224 ;
  assign n15227 = n15052 | n15226 ;
  assign n15228 = n70422 & n15227 ;
  assign n15229 = n15058 | n15228 ;
  assign n15231 = n70425 & n15229 ;
  assign n15232 = n15063 | n15231 ;
  assign n15233 = n70428 & n15232 ;
  assign n15234 = n15069 | n15233 ;
  assign n15236 = n70431 & n15234 ;
  assign n15237 = n15074 | n15236 ;
  assign n15238 = n70434 & n15237 ;
  assign n15239 = n15080 | n15238 ;
  assign n15241 = n70437 & n15239 ;
  assign n15242 = n15085 | n15241 ;
  assign n15243 = n70440 & n15242 ;
  assign n15244 = n15091 | n15243 ;
  assign n15246 = n70443 & n15244 ;
  assign n15247 = n15096 | n15246 ;
  assign n15248 = n70446 & n15247 ;
  assign n15249 = n15102 | n15248 ;
  assign n15251 = n70449 & n15249 ;
  assign n15252 = n15107 | n15251 ;
  assign n15253 = n70452 & n15252 ;
  assign n15254 = n15113 | n15253 ;
  assign n15256 = n70455 & n15254 ;
  assign n15257 = n15118 | n15256 ;
  assign n15258 = n70458 & n15257 ;
  assign n15259 = n15124 | n15258 ;
  assign n15261 = n70461 & n15259 ;
  assign n15262 = n15129 | n15261 ;
  assign n15263 = n70464 & n15262 ;
  assign n15264 = n15135 | n15263 ;
  assign n15266 = n70467 & n15264 ;
  assign n15267 = n15140 | n15266 ;
  assign n15268 = n70470 & n15267 ;
  assign n15269 = n15146 | n15268 ;
  assign n15271 = n70473 & n15269 ;
  assign n15272 = n15151 | n15271 ;
  assign n15273 = n70476 & n15272 ;
  assign n70484 = ~n15273 ;
  assign n15274 = n15157 & n70484 ;
  assign n15276 = n14590 | n15157 ;
  assign n70485 = ~n15276 ;
  assign n15277 = n15153 & n70485 ;
  assign n15278 = n15274 | n15277 ;
  assign n70486 = ~n15167 ;
  assign n15279 = n70486 & n15278 ;
  assign n70487 = ~n15165 ;
  assign n15280 = n70487 & n15279 ;
  assign n15281 = n15169 | n15280 ;
  assign n15282 = n70276 & n15281 ;
  assign n70488 = ~n15280 ;
  assign n15838 = x106 & n70488 ;
  assign n70489 = ~n15169 ;
  assign n15839 = n70489 & n15838 ;
  assign n15840 = n15282 | n15839 ;
  assign n15283 = n14589 & n15168 ;
  assign n70490 = ~n15148 ;
  assign n15152 = n70490 & n15151 ;
  assign n15284 = n14598 | n15151 ;
  assign n70491 = ~n15284 ;
  assign n15285 = n15269 & n70491 ;
  assign n15286 = n15152 | n15285 ;
  assign n15287 = n70486 & n15286 ;
  assign n15288 = n70487 & n15287 ;
  assign n15289 = n15283 | n15288 ;
  assign n15290 = n70176 & n15289 ;
  assign n15291 = n14597 & n15168 ;
  assign n70492 = ~n15268 ;
  assign n15270 = n15146 & n70492 ;
  assign n15292 = n14607 | n15146 ;
  assign n70493 = ~n15292 ;
  assign n15293 = n15142 & n70493 ;
  assign n15294 = n15270 | n15293 ;
  assign n15295 = n70486 & n15294 ;
  assign n15296 = n70487 & n15295 ;
  assign n15297 = n15291 | n15296 ;
  assign n15298 = n69857 & n15297 ;
  assign n70494 = ~n15296 ;
  assign n15826 = x104 & n70494 ;
  assign n70495 = ~n15291 ;
  assign n15827 = n70495 & n15826 ;
  assign n15828 = n15298 | n15827 ;
  assign n15299 = n14606 & n15168 ;
  assign n70496 = ~n15137 ;
  assign n15141 = n70496 & n15140 ;
  assign n15300 = n14616 | n15140 ;
  assign n70497 = ~n15300 ;
  assign n15301 = n15264 & n70497 ;
  assign n15302 = n15141 | n15301 ;
  assign n15303 = n70486 & n15302 ;
  assign n15304 = n70487 & n15303 ;
  assign n15305 = n15299 | n15304 ;
  assign n15306 = n69656 & n15305 ;
  assign n15307 = n14615 & n15168 ;
  assign n70498 = ~n15263 ;
  assign n15265 = n15135 & n70498 ;
  assign n15308 = n14625 | n15135 ;
  assign n70499 = ~n15308 ;
  assign n15309 = n15131 & n70499 ;
  assign n15310 = n15265 | n15309 ;
  assign n15311 = n70486 & n15310 ;
  assign n15312 = n70487 & n15311 ;
  assign n15313 = n15307 | n15312 ;
  assign n15314 = n69528 & n15313 ;
  assign n70500 = ~n15312 ;
  assign n15816 = x102 & n70500 ;
  assign n70501 = ~n15307 ;
  assign n15817 = n70501 & n15816 ;
  assign n15818 = n15314 | n15817 ;
  assign n15315 = n14624 & n15168 ;
  assign n70502 = ~n15126 ;
  assign n15130 = n70502 & n15129 ;
  assign n15316 = n14634 | n15129 ;
  assign n70503 = ~n15316 ;
  assign n15317 = n15259 & n70503 ;
  assign n15318 = n15130 | n15317 ;
  assign n15319 = n70486 & n15318 ;
  assign n15320 = n70487 & n15319 ;
  assign n15321 = n15315 | n15320 ;
  assign n15322 = n69261 & n15321 ;
  assign n15323 = n14633 & n15168 ;
  assign n70504 = ~n15258 ;
  assign n15260 = n15124 & n70504 ;
  assign n15324 = n14643 | n15124 ;
  assign n70505 = ~n15324 ;
  assign n15325 = n15120 & n70505 ;
  assign n15326 = n15260 | n15325 ;
  assign n15327 = n70486 & n15326 ;
  assign n15328 = n70487 & n15327 ;
  assign n15329 = n15323 | n15328 ;
  assign n15330 = n69075 & n15329 ;
  assign n70506 = ~n15328 ;
  assign n15805 = x100 & n70506 ;
  assign n70507 = ~n15323 ;
  assign n15806 = n70507 & n15805 ;
  assign n15807 = n15330 | n15806 ;
  assign n15331 = n14642 & n15168 ;
  assign n70508 = ~n15115 ;
  assign n15119 = n70508 & n15118 ;
  assign n15332 = n14652 | n15118 ;
  assign n70509 = ~n15332 ;
  assign n15333 = n15254 & n70509 ;
  assign n15334 = n15119 | n15333 ;
  assign n15335 = n70486 & n15334 ;
  assign n15336 = n70487 & n15335 ;
  assign n15337 = n15331 | n15336 ;
  assign n15338 = n68993 & n15337 ;
  assign n15339 = n14651 & n15168 ;
  assign n70510 = ~n15253 ;
  assign n15255 = n15113 & n70510 ;
  assign n15340 = n14661 | n15113 ;
  assign n70511 = ~n15340 ;
  assign n15341 = n15109 & n70511 ;
  assign n15342 = n15255 | n15341 ;
  assign n15343 = n70486 & n15342 ;
  assign n15344 = n70487 & n15343 ;
  assign n15345 = n15339 | n15344 ;
  assign n15346 = n68716 & n15345 ;
  assign n70512 = ~n15344 ;
  assign n15794 = x98 & n70512 ;
  assign n70513 = ~n15339 ;
  assign n15795 = n70513 & n15794 ;
  assign n15796 = n15346 | n15795 ;
  assign n15347 = n14660 & n15168 ;
  assign n70514 = ~n15104 ;
  assign n15108 = n70514 & n15107 ;
  assign n15348 = n14670 | n15107 ;
  assign n70515 = ~n15348 ;
  assign n15349 = n15249 & n70515 ;
  assign n15350 = n15108 | n15349 ;
  assign n15351 = n70486 & n15350 ;
  assign n15352 = n70487 & n15351 ;
  assign n15353 = n15347 | n15352 ;
  assign n15354 = n68545 & n15353 ;
  assign n15355 = n14669 & n15168 ;
  assign n70516 = ~n15248 ;
  assign n15250 = n15102 & n70516 ;
  assign n15356 = n14679 | n15102 ;
  assign n70517 = ~n15356 ;
  assign n15357 = n15098 & n70517 ;
  assign n15358 = n15250 | n15357 ;
  assign n15359 = n70486 & n15358 ;
  assign n15360 = n70487 & n15359 ;
  assign n15361 = n15355 | n15360 ;
  assign n15362 = n68438 & n15361 ;
  assign n70518 = ~n15360 ;
  assign n15784 = x96 & n70518 ;
  assign n70519 = ~n15355 ;
  assign n15785 = n70519 & n15784 ;
  assign n15786 = n15362 | n15785 ;
  assign n15363 = n14678 & n15168 ;
  assign n70520 = ~n15093 ;
  assign n15097 = n70520 & n15096 ;
  assign n15364 = n14688 | n15096 ;
  assign n70521 = ~n15364 ;
  assign n15365 = n15244 & n70521 ;
  assign n15366 = n15097 | n15365 ;
  assign n15367 = n70486 & n15366 ;
  assign n15368 = n70487 & n15367 ;
  assign n15369 = n15363 | n15368 ;
  assign n15370 = n68214 & n15369 ;
  assign n15371 = n14687 & n15168 ;
  assign n70522 = ~n15243 ;
  assign n15245 = n15091 & n70522 ;
  assign n15372 = n14697 | n15091 ;
  assign n70523 = ~n15372 ;
  assign n15373 = n15087 & n70523 ;
  assign n15374 = n15245 | n15373 ;
  assign n15375 = n70486 & n15374 ;
  assign n15376 = n70487 & n15375 ;
  assign n15377 = n15371 | n15376 ;
  assign n15378 = n68058 & n15377 ;
  assign n70524 = ~n15376 ;
  assign n15774 = x94 & n70524 ;
  assign n70525 = ~n15371 ;
  assign n15775 = n70525 & n15774 ;
  assign n15776 = n15378 | n15775 ;
  assign n15379 = n14696 & n15168 ;
  assign n70526 = ~n15082 ;
  assign n15086 = n70526 & n15085 ;
  assign n15380 = n14706 | n15085 ;
  assign n70527 = ~n15380 ;
  assign n15381 = n15239 & n70527 ;
  assign n15382 = n15086 | n15381 ;
  assign n15383 = n70486 & n15382 ;
  assign n15384 = n70487 & n15383 ;
  assign n15385 = n15379 | n15384 ;
  assign n15386 = n67986 & n15385 ;
  assign n15387 = n14705 & n15168 ;
  assign n70528 = ~n15238 ;
  assign n15240 = n15080 & n70528 ;
  assign n15388 = n14715 | n15080 ;
  assign n70529 = ~n15388 ;
  assign n15389 = n15076 & n70529 ;
  assign n15390 = n15240 | n15389 ;
  assign n15391 = n70486 & n15390 ;
  assign n15392 = n70487 & n15391 ;
  assign n15393 = n15387 | n15392 ;
  assign n15394 = n67763 & n15393 ;
  assign n70530 = ~n15392 ;
  assign n15763 = x92 & n70530 ;
  assign n70531 = ~n15387 ;
  assign n15764 = n70531 & n15763 ;
  assign n15765 = n15394 | n15764 ;
  assign n15395 = n14714 & n15168 ;
  assign n70532 = ~n15071 ;
  assign n15075 = n70532 & n15074 ;
  assign n15396 = n14724 | n15074 ;
  assign n70533 = ~n15396 ;
  assign n15397 = n15234 & n70533 ;
  assign n15398 = n15075 | n15397 ;
  assign n15399 = n70486 & n15398 ;
  assign n15400 = n70487 & n15399 ;
  assign n15401 = n15395 | n15400 ;
  assign n15402 = n67622 & n15401 ;
  assign n15403 = n14723 & n15168 ;
  assign n70534 = ~n15233 ;
  assign n15235 = n15069 & n70534 ;
  assign n15404 = n14732 | n15069 ;
  assign n70535 = ~n15404 ;
  assign n15405 = n15065 & n70535 ;
  assign n15406 = n15235 | n15405 ;
  assign n15407 = n70486 & n15406 ;
  assign n15408 = n70487 & n15407 ;
  assign n15409 = n15403 | n15408 ;
  assign n15410 = n67531 & n15409 ;
  assign n70536 = ~n15408 ;
  assign n15752 = x90 & n70536 ;
  assign n70537 = ~n15403 ;
  assign n15753 = n70537 & n15752 ;
  assign n15754 = n15410 | n15753 ;
  assign n15411 = n14731 & n15168 ;
  assign n70538 = ~n15060 ;
  assign n15064 = n70538 & n15063 ;
  assign n15412 = n14741 | n15063 ;
  assign n70539 = ~n15412 ;
  assign n15413 = n15229 & n70539 ;
  assign n15414 = n15064 | n15413 ;
  assign n15415 = n70486 & n15414 ;
  assign n15416 = n70487 & n15415 ;
  assign n15417 = n15411 | n15416 ;
  assign n15418 = n67348 & n15417 ;
  assign n15419 = n14740 & n15168 ;
  assign n70540 = ~n15228 ;
  assign n15230 = n15058 & n70540 ;
  assign n15420 = n14750 | n15058 ;
  assign n70541 = ~n15420 ;
  assign n15421 = n15054 & n70541 ;
  assign n15422 = n15230 | n15421 ;
  assign n15423 = n70486 & n15422 ;
  assign n15424 = n70487 & n15423 ;
  assign n15425 = n15419 | n15424 ;
  assign n15426 = n67222 & n15425 ;
  assign n70542 = ~n15424 ;
  assign n15741 = x88 & n70542 ;
  assign n70543 = ~n15419 ;
  assign n15742 = n70543 & n15741 ;
  assign n15743 = n15426 | n15742 ;
  assign n15427 = n14749 & n15168 ;
  assign n70544 = ~n15049 ;
  assign n15053 = n70544 & n15052 ;
  assign n15428 = n14759 | n15052 ;
  assign n70545 = ~n15428 ;
  assign n15429 = n15224 & n70545 ;
  assign n15430 = n15053 | n15429 ;
  assign n15431 = n70486 & n15430 ;
  assign n15432 = n70487 & n15431 ;
  assign n15433 = n15427 | n15432 ;
  assign n15434 = n67164 & n15433 ;
  assign n15435 = n14758 & n15168 ;
  assign n70546 = ~n15223 ;
  assign n15225 = n15047 & n70546 ;
  assign n15436 = n14768 | n15047 ;
  assign n70547 = ~n15436 ;
  assign n15437 = n15043 & n70547 ;
  assign n15438 = n15225 | n15437 ;
  assign n15439 = n70486 & n15438 ;
  assign n15440 = n70487 & n15439 ;
  assign n15441 = n15435 | n15440 ;
  assign n15442 = n66979 & n15441 ;
  assign n70548 = ~n15440 ;
  assign n15731 = x86 & n70548 ;
  assign n70549 = ~n15435 ;
  assign n15732 = n70549 & n15731 ;
  assign n15733 = n15442 | n15732 ;
  assign n15443 = n14767 & n15168 ;
  assign n70550 = ~n15038 ;
  assign n15042 = n70550 & n15041 ;
  assign n15444 = n14777 | n15041 ;
  assign n70551 = ~n15444 ;
  assign n15445 = n15219 & n70551 ;
  assign n15446 = n15042 | n15445 ;
  assign n15447 = n70486 & n15446 ;
  assign n15448 = n70487 & n15447 ;
  assign n15449 = n15443 | n15448 ;
  assign n15450 = n66868 & n15449 ;
  assign n15451 = n14776 & n15168 ;
  assign n70552 = ~n15218 ;
  assign n15220 = n15036 & n70552 ;
  assign n15452 = n14786 | n15036 ;
  assign n70553 = ~n15452 ;
  assign n15453 = n15032 & n70553 ;
  assign n15454 = n15220 | n15453 ;
  assign n15455 = n70486 & n15454 ;
  assign n15456 = n70487 & n15455 ;
  assign n15457 = n15451 | n15456 ;
  assign n15458 = n66797 & n15457 ;
  assign n70554 = ~n15456 ;
  assign n15720 = x84 & n70554 ;
  assign n70555 = ~n15451 ;
  assign n15721 = n70555 & n15720 ;
  assign n15722 = n15458 | n15721 ;
  assign n15459 = n14785 & n15168 ;
  assign n70556 = ~n15027 ;
  assign n15031 = n70556 & n15030 ;
  assign n15460 = n14794 | n15030 ;
  assign n70557 = ~n15460 ;
  assign n15461 = n15214 & n70557 ;
  assign n15462 = n15031 | n15461 ;
  assign n15463 = n70486 & n15462 ;
  assign n15464 = n70487 & n15463 ;
  assign n15465 = n15459 | n15464 ;
  assign n15466 = n66654 & n15465 ;
  assign n15467 = n14793 & n15168 ;
  assign n70558 = ~n15213 ;
  assign n15215 = n15025 & n70558 ;
  assign n15468 = n14803 | n15025 ;
  assign n70559 = ~n15468 ;
  assign n15469 = n15021 & n70559 ;
  assign n15470 = n15215 | n15469 ;
  assign n15471 = n70486 & n15470 ;
  assign n15472 = n70487 & n15471 ;
  assign n15473 = n15467 | n15472 ;
  assign n15474 = n66560 & n15473 ;
  assign n70560 = ~n15472 ;
  assign n15709 = x82 & n70560 ;
  assign n70561 = ~n15467 ;
  assign n15710 = n70561 & n15709 ;
  assign n15711 = n15474 | n15710 ;
  assign n15475 = n14802 & n15168 ;
  assign n70562 = ~n15016 ;
  assign n15020 = n70562 & n15019 ;
  assign n15476 = n14812 | n15019 ;
  assign n70563 = ~n15476 ;
  assign n15477 = n15209 & n70563 ;
  assign n15478 = n15020 | n15477 ;
  assign n15479 = n70486 & n15478 ;
  assign n15480 = n70487 & n15479 ;
  assign n15481 = n15475 | n15480 ;
  assign n15482 = n66505 & n15481 ;
  assign n15483 = n14811 & n15168 ;
  assign n70564 = ~n15208 ;
  assign n15210 = n15014 & n70564 ;
  assign n15484 = n14820 | n15014 ;
  assign n70565 = ~n15484 ;
  assign n15485 = n15010 & n70565 ;
  assign n15486 = n15210 | n15485 ;
  assign n15487 = n70486 & n15486 ;
  assign n15488 = n70487 & n15487 ;
  assign n15489 = n15483 | n15488 ;
  assign n15490 = n66379 & n15489 ;
  assign n70566 = ~n15488 ;
  assign n15697 = x80 & n70566 ;
  assign n70567 = ~n15483 ;
  assign n15698 = n70567 & n15697 ;
  assign n15699 = n15490 | n15698 ;
  assign n15491 = n14819 & n15168 ;
  assign n70568 = ~n15005 ;
  assign n15009 = n70568 & n15008 ;
  assign n15492 = n14829 | n15008 ;
  assign n70569 = ~n15492 ;
  assign n15493 = n15204 & n70569 ;
  assign n15494 = n15009 | n15493 ;
  assign n15495 = n70486 & n15494 ;
  assign n15496 = n70487 & n15495 ;
  assign n15497 = n15491 | n15496 ;
  assign n15498 = n66299 & n15497 ;
  assign n15499 = n14828 & n15168 ;
  assign n70570 = ~n15203 ;
  assign n15205 = n15003 & n70570 ;
  assign n15500 = n14837 | n15003 ;
  assign n70571 = ~n15500 ;
  assign n15501 = n14999 & n70571 ;
  assign n15502 = n15205 | n15501 ;
  assign n15503 = n70486 & n15502 ;
  assign n15504 = n70487 & n15503 ;
  assign n15505 = n15499 | n15504 ;
  assign n15506 = n66244 & n15505 ;
  assign n70572 = ~n15504 ;
  assign n15687 = x78 & n70572 ;
  assign n70573 = ~n15499 ;
  assign n15688 = n70573 & n15687 ;
  assign n15689 = n15506 | n15688 ;
  assign n15507 = n14836 & n15168 ;
  assign n70574 = ~n14994 ;
  assign n14998 = n70574 & n14997 ;
  assign n15508 = n14846 | n14997 ;
  assign n70575 = ~n15508 ;
  assign n15509 = n15199 & n70575 ;
  assign n15510 = n14998 | n15509 ;
  assign n15511 = n70486 & n15510 ;
  assign n15512 = n70487 & n15511 ;
  assign n15513 = n15507 | n15512 ;
  assign n15514 = n66145 & n15513 ;
  assign n15515 = n14845 & n15168 ;
  assign n70576 = ~n15198 ;
  assign n15200 = n14992 & n70576 ;
  assign n15516 = n14854 | n14992 ;
  assign n70577 = ~n15516 ;
  assign n15517 = n14988 & n70577 ;
  assign n15518 = n15200 | n15517 ;
  assign n15519 = n70486 & n15518 ;
  assign n15520 = n70487 & n15519 ;
  assign n15521 = n15515 | n15520 ;
  assign n15522 = n66081 & n15521 ;
  assign n70578 = ~n15520 ;
  assign n15677 = x76 & n70578 ;
  assign n70579 = ~n15515 ;
  assign n15678 = n70579 & n15677 ;
  assign n15679 = n15522 | n15678 ;
  assign n15523 = n14853 & n15168 ;
  assign n70580 = ~n14983 ;
  assign n14987 = n70580 & n14986 ;
  assign n15524 = n14863 | n14986 ;
  assign n70581 = ~n15524 ;
  assign n15525 = n15194 & n70581 ;
  assign n15526 = n14987 | n15525 ;
  assign n15527 = n70486 & n15526 ;
  assign n15528 = n70487 & n15527 ;
  assign n15529 = n15523 | n15528 ;
  assign n15530 = n66043 & n15529 ;
  assign n15531 = n14862 & n15168 ;
  assign n70582 = ~n15193 ;
  assign n15195 = n14981 & n70582 ;
  assign n15532 = n14872 | n14981 ;
  assign n70583 = ~n15532 ;
  assign n15533 = n14977 & n70583 ;
  assign n15534 = n15195 | n15533 ;
  assign n15535 = n70486 & n15534 ;
  assign n15536 = n70487 & n15535 ;
  assign n15537 = n15531 | n15536 ;
  assign n15538 = n65960 & n15537 ;
  assign n70584 = ~n15536 ;
  assign n15666 = x74 & n70584 ;
  assign n70585 = ~n15531 ;
  assign n15667 = n70585 & n15666 ;
  assign n15668 = n15538 | n15667 ;
  assign n15539 = n14871 & n15168 ;
  assign n70586 = ~n14972 ;
  assign n14976 = n70586 & n14975 ;
  assign n15540 = n14881 | n14975 ;
  assign n70587 = ~n15540 ;
  assign n15541 = n15189 & n70587 ;
  assign n15542 = n14976 | n15541 ;
  assign n15543 = n70486 & n15542 ;
  assign n15544 = n70487 & n15543 ;
  assign n15545 = n15539 | n15544 ;
  assign n15546 = n65909 & n15545 ;
  assign n15547 = n14880 & n15168 ;
  assign n70588 = ~n15188 ;
  assign n15190 = n14970 & n70588 ;
  assign n15548 = n14963 | n15185 ;
  assign n15549 = n14890 | n14970 ;
  assign n70589 = ~n15549 ;
  assign n15550 = n15548 & n70589 ;
  assign n15551 = n15190 | n15550 ;
  assign n15552 = n70486 & n15551 ;
  assign n15553 = n70487 & n15552 ;
  assign n15554 = n15547 | n15553 ;
  assign n15555 = n65877 & n15554 ;
  assign n70590 = ~n15553 ;
  assign n15656 = x72 & n70590 ;
  assign n70591 = ~n15547 ;
  assign n15657 = n70591 & n15656 ;
  assign n15658 = n15555 | n15657 ;
  assign n15556 = n14889 & n15168 ;
  assign n70592 = ~n14963 ;
  assign n15186 = n70592 & n15185 ;
  assign n15557 = n14961 | n15181 ;
  assign n15558 = n14899 | n15185 ;
  assign n70593 = ~n15558 ;
  assign n15559 = n15557 & n70593 ;
  assign n15560 = n15186 | n15559 ;
  assign n15561 = n70486 & n15560 ;
  assign n15562 = n70487 & n15561 ;
  assign n15563 = n15556 | n15562 ;
  assign n15564 = n65820 & n15563 ;
  assign n15565 = n14898 & n15168 ;
  assign n70594 = ~n15181 ;
  assign n15183 = n14961 & n70594 ;
  assign n15566 = n14908 | n14961 ;
  assign n70595 = ~n15566 ;
  assign n15567 = n14957 & n70595 ;
  assign n15568 = n15183 | n15567 ;
  assign n15569 = n70486 & n15568 ;
  assign n15570 = n70487 & n15569 ;
  assign n15571 = n15565 | n15570 ;
  assign n15572 = n65791 & n15571 ;
  assign n70596 = ~n15570 ;
  assign n15646 = x70 & n70596 ;
  assign n70597 = ~n15565 ;
  assign n15647 = n70597 & n15646 ;
  assign n15648 = n15572 | n15647 ;
  assign n15573 = n14907 & n15168 ;
  assign n70598 = ~n14953 ;
  assign n15179 = n70598 & n14956 ;
  assign n15574 = n14917 | n14956 ;
  assign n70599 = ~n15574 ;
  assign n15575 = n15177 & n70599 ;
  assign n15576 = n15179 | n15575 ;
  assign n15577 = n70486 & n15576 ;
  assign n15578 = n70487 & n15577 ;
  assign n15579 = n15573 | n15578 ;
  assign n15580 = n65772 & n15579 ;
  assign n15581 = n14916 & n15168 ;
  assign n70600 = ~n15175 ;
  assign n15176 = n14951 & n70600 ;
  assign n15582 = n14925 | n14951 ;
  assign n70601 = ~n15582 ;
  assign n15583 = n15174 & n70601 ;
  assign n15584 = n15176 | n15583 ;
  assign n15585 = n70486 & n15584 ;
  assign n15586 = n70487 & n15585 ;
  assign n15587 = n15581 | n15586 ;
  assign n15588 = n65746 & n15587 ;
  assign n70602 = ~n15586 ;
  assign n15636 = x68 & n70602 ;
  assign n70603 = ~n15581 ;
  assign n15637 = n70603 & n15636 ;
  assign n15638 = n15588 | n15637 ;
  assign n15589 = n14924 & n15168 ;
  assign n15590 = n14941 | n14946 ;
  assign n70604 = ~n15590 ;
  assign n15591 = n15172 & n70604 ;
  assign n70605 = ~n14943 ;
  assign n15592 = n70605 & n14946 ;
  assign n15593 = n15591 | n15592 ;
  assign n15594 = n70486 & n15593 ;
  assign n15595 = n70487 & n15594 ;
  assign n15596 = n15589 | n15595 ;
  assign n15597 = n65721 & n15596 ;
  assign n15598 = n14935 & n15168 ;
  assign n15599 = n14938 & n14940 ;
  assign n15600 = n70483 & n15599 ;
  assign n15601 = n15167 | n15600 ;
  assign n70606 = ~n15601 ;
  assign n15602 = n15172 & n70606 ;
  assign n15603 = n70487 & n15602 ;
  assign n15604 = n15598 | n15603 ;
  assign n15605 = n65686 & n15604 ;
  assign n70607 = ~n15603 ;
  assign n15626 = x66 & n70607 ;
  assign n70608 = ~n15598 ;
  assign n15627 = n70608 & n15626 ;
  assign n15628 = n15605 | n15627 ;
  assign n15275 = n15157 | n15273 ;
  assign n15606 = n70479 & n15275 ;
  assign n15607 = n15162 | n15606 ;
  assign n15608 = n70482 & n15607 ;
  assign n70609 = ~x107 ;
  assign n15609 = x64 & n70609 ;
  assign n15610 = n70178 & n15609 ;
  assign n15611 = n66510 & n15610 ;
  assign n70610 = ~n15608 ;
  assign n15612 = n70610 & n15611 ;
  assign n70611 = ~n15612 ;
  assign n15613 = x21 & n70611 ;
  assign n70612 = ~n291 ;
  assign n15614 = n70612 & n14940 ;
  assign n70613 = ~n289 ;
  assign n15615 = n70613 & n15614 ;
  assign n15616 = n66715 & n15615 ;
  assign n15617 = n70487 & n15616 ;
  assign n15618 = n15613 | n15617 ;
  assign n15619 = x65 & n15618 ;
  assign n15620 = x65 | n15617 ;
  assign n15621 = n15613 | n15620 ;
  assign n70614 = ~n15619 ;
  assign n15622 = n70614 & n15621 ;
  assign n70615 = ~x20 ;
  assign n15623 = n70615 & x64 ;
  assign n15624 = n15622 | n15623 ;
  assign n15625 = n65670 & n15618 ;
  assign n70616 = ~n15625 ;
  assign n15629 = n15624 & n70616 ;
  assign n15630 = n15628 | n15629 ;
  assign n70617 = ~n15605 ;
  assign n15631 = n70617 & n15630 ;
  assign n70618 = ~n15595 ;
  assign n15632 = x67 & n70618 ;
  assign n70619 = ~n15589 ;
  assign n15633 = n70619 & n15632 ;
  assign n15634 = n15597 | n15633 ;
  assign n15635 = n15631 | n15634 ;
  assign n70620 = ~n15597 ;
  assign n15639 = n70620 & n15635 ;
  assign n15640 = n15638 | n15639 ;
  assign n70621 = ~n15588 ;
  assign n15641 = n70621 & n15640 ;
  assign n70622 = ~n15578 ;
  assign n15642 = x69 & n70622 ;
  assign n70623 = ~n15573 ;
  assign n15643 = n70623 & n15642 ;
  assign n15644 = n15580 | n15643 ;
  assign n15645 = n15641 | n15644 ;
  assign n70624 = ~n15580 ;
  assign n15649 = n70624 & n15645 ;
  assign n15650 = n15648 | n15649 ;
  assign n70625 = ~n15572 ;
  assign n15651 = n70625 & n15650 ;
  assign n70626 = ~n15562 ;
  assign n15652 = x71 & n70626 ;
  assign n70627 = ~n15556 ;
  assign n15653 = n70627 & n15652 ;
  assign n15654 = n15564 | n15653 ;
  assign n15655 = n15651 | n15654 ;
  assign n70628 = ~n15564 ;
  assign n15659 = n70628 & n15655 ;
  assign n15660 = n15658 | n15659 ;
  assign n70629 = ~n15555 ;
  assign n15661 = n70629 & n15660 ;
  assign n70630 = ~n15544 ;
  assign n15662 = x73 & n70630 ;
  assign n70631 = ~n15539 ;
  assign n15663 = n70631 & n15662 ;
  assign n15664 = n15546 | n15663 ;
  assign n15665 = n15661 | n15664 ;
  assign n70632 = ~n15546 ;
  assign n15670 = n70632 & n15665 ;
  assign n15671 = n15668 | n15670 ;
  assign n70633 = ~n15538 ;
  assign n15672 = n70633 & n15671 ;
  assign n70634 = ~n15528 ;
  assign n15673 = x75 & n70634 ;
  assign n70635 = ~n15523 ;
  assign n15674 = n70635 & n15673 ;
  assign n15675 = n15530 | n15674 ;
  assign n15676 = n15672 | n15675 ;
  assign n70636 = ~n15530 ;
  assign n15680 = n70636 & n15676 ;
  assign n15681 = n15679 | n15680 ;
  assign n70637 = ~n15522 ;
  assign n15682 = n70637 & n15681 ;
  assign n70638 = ~n15512 ;
  assign n15683 = x77 & n70638 ;
  assign n70639 = ~n15507 ;
  assign n15684 = n70639 & n15683 ;
  assign n15685 = n15514 | n15684 ;
  assign n15686 = n15682 | n15685 ;
  assign n70640 = ~n15514 ;
  assign n15690 = n70640 & n15686 ;
  assign n15691 = n15689 | n15690 ;
  assign n70641 = ~n15506 ;
  assign n15692 = n70641 & n15691 ;
  assign n70642 = ~n15496 ;
  assign n15693 = x79 & n70642 ;
  assign n70643 = ~n15491 ;
  assign n15694 = n70643 & n15693 ;
  assign n15695 = n15498 | n15694 ;
  assign n15696 = n15692 | n15695 ;
  assign n70644 = ~n15498 ;
  assign n15701 = n70644 & n15696 ;
  assign n15702 = n15699 | n15701 ;
  assign n70645 = ~n15490 ;
  assign n15703 = n70645 & n15702 ;
  assign n70646 = ~n15480 ;
  assign n15704 = x81 & n70646 ;
  assign n70647 = ~n15475 ;
  assign n15705 = n70647 & n15704 ;
  assign n15706 = n15482 | n15705 ;
  assign n15708 = n15703 | n15706 ;
  assign n70648 = ~n15482 ;
  assign n15713 = n70648 & n15708 ;
  assign n15714 = n15711 | n15713 ;
  assign n70649 = ~n15474 ;
  assign n15715 = n70649 & n15714 ;
  assign n70650 = ~n15464 ;
  assign n15716 = x83 & n70650 ;
  assign n70651 = ~n15459 ;
  assign n15717 = n70651 & n15716 ;
  assign n15718 = n15466 | n15717 ;
  assign n15719 = n15715 | n15718 ;
  assign n70652 = ~n15466 ;
  assign n15723 = n70652 & n15719 ;
  assign n15724 = n15722 | n15723 ;
  assign n70653 = ~n15458 ;
  assign n15725 = n70653 & n15724 ;
  assign n70654 = ~n15448 ;
  assign n15726 = x85 & n70654 ;
  assign n70655 = ~n15443 ;
  assign n15727 = n70655 & n15726 ;
  assign n15728 = n15450 | n15727 ;
  assign n15730 = n15725 | n15728 ;
  assign n70656 = ~n15450 ;
  assign n15734 = n70656 & n15730 ;
  assign n15735 = n15733 | n15734 ;
  assign n70657 = ~n15442 ;
  assign n15736 = n70657 & n15735 ;
  assign n70658 = ~n15432 ;
  assign n15737 = x87 & n70658 ;
  assign n70659 = ~n15427 ;
  assign n15738 = n70659 & n15737 ;
  assign n15739 = n15434 | n15738 ;
  assign n15740 = n15736 | n15739 ;
  assign n70660 = ~n15434 ;
  assign n15744 = n70660 & n15740 ;
  assign n15745 = n15743 | n15744 ;
  assign n70661 = ~n15426 ;
  assign n15746 = n70661 & n15745 ;
  assign n70662 = ~n15416 ;
  assign n15747 = x89 & n70662 ;
  assign n70663 = ~n15411 ;
  assign n15748 = n70663 & n15747 ;
  assign n15749 = n15418 | n15748 ;
  assign n15751 = n15746 | n15749 ;
  assign n70664 = ~n15418 ;
  assign n15755 = n70664 & n15751 ;
  assign n15756 = n15754 | n15755 ;
  assign n70665 = ~n15410 ;
  assign n15757 = n70665 & n15756 ;
  assign n70666 = ~n15400 ;
  assign n15758 = x91 & n70666 ;
  assign n70667 = ~n15395 ;
  assign n15759 = n70667 & n15758 ;
  assign n15760 = n15402 | n15759 ;
  assign n15762 = n15757 | n15760 ;
  assign n70668 = ~n15402 ;
  assign n15767 = n70668 & n15762 ;
  assign n15768 = n15765 | n15767 ;
  assign n70669 = ~n15394 ;
  assign n15769 = n70669 & n15768 ;
  assign n70670 = ~n15384 ;
  assign n15770 = x93 & n70670 ;
  assign n70671 = ~n15379 ;
  assign n15771 = n70671 & n15770 ;
  assign n15772 = n15386 | n15771 ;
  assign n15773 = n15769 | n15772 ;
  assign n70672 = ~n15386 ;
  assign n15777 = n70672 & n15773 ;
  assign n15778 = n15776 | n15777 ;
  assign n70673 = ~n15378 ;
  assign n15779 = n70673 & n15778 ;
  assign n70674 = ~n15368 ;
  assign n15780 = x95 & n70674 ;
  assign n70675 = ~n15363 ;
  assign n15781 = n70675 & n15780 ;
  assign n15782 = n15370 | n15781 ;
  assign n15783 = n15779 | n15782 ;
  assign n70676 = ~n15370 ;
  assign n15787 = n70676 & n15783 ;
  assign n15788 = n15786 | n15787 ;
  assign n70677 = ~n15362 ;
  assign n15789 = n70677 & n15788 ;
  assign n70678 = ~n15352 ;
  assign n15790 = x97 & n70678 ;
  assign n70679 = ~n15347 ;
  assign n15791 = n70679 & n15790 ;
  assign n15792 = n15354 | n15791 ;
  assign n15793 = n15789 | n15792 ;
  assign n70680 = ~n15354 ;
  assign n15798 = n70680 & n15793 ;
  assign n15799 = n15796 | n15798 ;
  assign n70681 = ~n15346 ;
  assign n15800 = n70681 & n15799 ;
  assign n70682 = ~n15336 ;
  assign n15801 = x99 & n70682 ;
  assign n70683 = ~n15331 ;
  assign n15802 = n70683 & n15801 ;
  assign n15803 = n15338 | n15802 ;
  assign n15804 = n15800 | n15803 ;
  assign n70684 = ~n15338 ;
  assign n15809 = n70684 & n15804 ;
  assign n15810 = n15807 | n15809 ;
  assign n70685 = ~n15330 ;
  assign n15811 = n70685 & n15810 ;
  assign n70686 = ~n15320 ;
  assign n15812 = x101 & n70686 ;
  assign n70687 = ~n15315 ;
  assign n15813 = n70687 & n15812 ;
  assign n15814 = n15322 | n15813 ;
  assign n15815 = n15811 | n15814 ;
  assign n70688 = ~n15322 ;
  assign n15819 = n70688 & n15815 ;
  assign n15820 = n15818 | n15819 ;
  assign n70689 = ~n15314 ;
  assign n15821 = n70689 & n15820 ;
  assign n70690 = ~n15304 ;
  assign n15822 = x103 & n70690 ;
  assign n70691 = ~n15299 ;
  assign n15823 = n70691 & n15822 ;
  assign n15824 = n15306 | n15823 ;
  assign n15825 = n15821 | n15824 ;
  assign n70692 = ~n15306 ;
  assign n15830 = n70692 & n15825 ;
  assign n15831 = n15828 | n15830 ;
  assign n70693 = ~n15298 ;
  assign n15832 = n70693 & n15831 ;
  assign n70694 = ~n15288 ;
  assign n15833 = x105 & n70694 ;
  assign n70695 = ~n15283 ;
  assign n15834 = n70695 & n15833 ;
  assign n15835 = n15290 | n15834 ;
  assign n15837 = n15832 | n15835 ;
  assign n70696 = ~n15290 ;
  assign n15842 = n70696 & n15837 ;
  assign n15843 = n15840 | n15842 ;
  assign n70697 = ~n15282 ;
  assign n15844 = n70697 & n15843 ;
  assign n70698 = ~n15159 ;
  assign n15163 = n70698 & n15162 ;
  assign n15845 = n14581 | n15162 ;
  assign n70699 = ~n15845 ;
  assign n15846 = n15275 & n70699 ;
  assign n15847 = n15163 | n15846 ;
  assign n15848 = n15168 | n15847 ;
  assign n70700 = ~n14488 ;
  assign n15849 = n70700 & n15168 ;
  assign n70701 = ~n15849 ;
  assign n15850 = n15848 & n70701 ;
  assign n15851 = n70609 & n15850 ;
  assign n150 = ~n15168 ;
  assign n15852 = n150 & n15847 ;
  assign n15853 = n14488 & n15168 ;
  assign n70703 = ~n15853 ;
  assign n15854 = x107 & n70703 ;
  assign n70704 = ~n15852 ;
  assign n15855 = n70704 & n15854 ;
  assign n15857 = n15855 | n15856 ;
  assign n15858 = n15851 | n15857 ;
  assign n15859 = n15844 | n15858 ;
  assign n15860 = n70486 & n15850 ;
  assign n70705 = ~n15860 ;
  assign n15861 = n15859 & n70705 ;
  assign n16561 = n15282 | n15855 ;
  assign n16562 = n15851 | n16561 ;
  assign n70706 = ~n16562 ;
  assign n16563 = n15843 & n70706 ;
  assign n15871 = n70487 & n15611 ;
  assign n70707 = ~n15871 ;
  assign n15872 = x21 & n70707 ;
  assign n15873 = n15617 | n15872 ;
  assign n15874 = x65 & n15873 ;
  assign n70708 = ~n15874 ;
  assign n15875 = n15621 & n70708 ;
  assign n15876 = n15623 | n15875 ;
  assign n15877 = n70616 & n15876 ;
  assign n15878 = n15628 | n15877 ;
  assign n15879 = n70617 & n15878 ;
  assign n15880 = n15634 | n15879 ;
  assign n15881 = n70620 & n15880 ;
  assign n15882 = n15638 | n15881 ;
  assign n15883 = n70621 & n15882 ;
  assign n15884 = n15644 | n15883 ;
  assign n15885 = n70624 & n15884 ;
  assign n15886 = n15648 | n15885 ;
  assign n15887 = n70625 & n15886 ;
  assign n15888 = n15654 | n15887 ;
  assign n15889 = n70628 & n15888 ;
  assign n15890 = n15658 | n15889 ;
  assign n15891 = n70629 & n15890 ;
  assign n15892 = n15664 | n15891 ;
  assign n15893 = n70632 & n15892 ;
  assign n15894 = n15668 | n15893 ;
  assign n15895 = n70633 & n15894 ;
  assign n15896 = n15675 | n15895 ;
  assign n15897 = n70636 & n15896 ;
  assign n15898 = n15679 | n15897 ;
  assign n15899 = n70637 & n15898 ;
  assign n15900 = n15685 | n15899 ;
  assign n15901 = n70640 & n15900 ;
  assign n15902 = n15689 | n15901 ;
  assign n15903 = n70641 & n15902 ;
  assign n15904 = n15695 | n15903 ;
  assign n15905 = n70644 & n15904 ;
  assign n15906 = n15699 | n15905 ;
  assign n15907 = n70645 & n15906 ;
  assign n15908 = n15706 | n15907 ;
  assign n15909 = n70648 & n15908 ;
  assign n15910 = n15711 | n15909 ;
  assign n15911 = n70649 & n15910 ;
  assign n15912 = n15718 | n15911 ;
  assign n15913 = n70652 & n15912 ;
  assign n15914 = n15722 | n15913 ;
  assign n15915 = n70653 & n15914 ;
  assign n15916 = n15728 | n15915 ;
  assign n15917 = n70656 & n15916 ;
  assign n15918 = n15733 | n15917 ;
  assign n15919 = n70657 & n15918 ;
  assign n15920 = n15739 | n15919 ;
  assign n15921 = n70660 & n15920 ;
  assign n15922 = n15743 | n15921 ;
  assign n15923 = n70661 & n15922 ;
  assign n15924 = n15749 | n15923 ;
  assign n15925 = n70664 & n15924 ;
  assign n15926 = n15754 | n15925 ;
  assign n15927 = n70665 & n15926 ;
  assign n15928 = n15760 | n15927 ;
  assign n15929 = n70668 & n15928 ;
  assign n15930 = n15765 | n15929 ;
  assign n15931 = n70669 & n15930 ;
  assign n15932 = n15772 | n15931 ;
  assign n15933 = n70672 & n15932 ;
  assign n15934 = n15776 | n15933 ;
  assign n15935 = n70673 & n15934 ;
  assign n15936 = n15782 | n15935 ;
  assign n15937 = n70676 & n15936 ;
  assign n15938 = n15786 | n15937 ;
  assign n15939 = n70677 & n15938 ;
  assign n15940 = n15792 | n15939 ;
  assign n15941 = n70680 & n15940 ;
  assign n15942 = n15796 | n15941 ;
  assign n15943 = n70681 & n15942 ;
  assign n15944 = n15803 | n15943 ;
  assign n15945 = n70684 & n15944 ;
  assign n15946 = n15807 | n15945 ;
  assign n15947 = n70685 & n15946 ;
  assign n15948 = n15814 | n15947 ;
  assign n15949 = n70688 & n15948 ;
  assign n15950 = n15818 | n15949 ;
  assign n15951 = n70689 & n15950 ;
  assign n15952 = n15824 | n15951 ;
  assign n15953 = n70692 & n15952 ;
  assign n15954 = n15828 | n15953 ;
  assign n15955 = n70693 & n15954 ;
  assign n16312 = n15835 | n15955 ;
  assign n16313 = n70696 & n16312 ;
  assign n16314 = n15840 | n16313 ;
  assign n16315 = n70697 & n16314 ;
  assign n16564 = n15851 | n15855 ;
  assign n70709 = ~n16315 ;
  assign n16565 = n70709 & n16564 ;
  assign n16566 = n16563 | n16565 ;
  assign n149 = ~n15861 ;
  assign n16567 = n149 & n16566 ;
  assign n16568 = n15167 & n15850 ;
  assign n16569 = n15859 & n16568 ;
  assign n16570 = n16567 | n16569 ;
  assign n70711 = ~n15856 ;
  assign n16577 = n70711 & n16570 ;
  assign n70712 = ~n15842 ;
  assign n15863 = n15840 & n70712 ;
  assign n15841 = n15290 | n15840 ;
  assign n70713 = ~n15841 ;
  assign n15864 = n15837 & n70713 ;
  assign n15865 = n15863 | n15864 ;
  assign n15866 = n149 & n15865 ;
  assign n15867 = n15281 & n70705 ;
  assign n15868 = n15859 & n15867 ;
  assign n15869 = n15866 | n15868 ;
  assign n15870 = n70609 & n15869 ;
  assign n70714 = ~n15955 ;
  assign n15956 = n15835 & n70714 ;
  assign n15836 = n15298 | n15835 ;
  assign n70715 = ~n15836 ;
  assign n15957 = n70715 & n15954 ;
  assign n15958 = n15956 | n15957 ;
  assign n15959 = n149 & n15958 ;
  assign n15960 = n15289 & n70705 ;
  assign n15961 = n15859 & n15960 ;
  assign n15962 = n15959 | n15961 ;
  assign n15963 = n70276 & n15962 ;
  assign n70716 = ~n15830 ;
  assign n15964 = n15828 & n70716 ;
  assign n15829 = n15306 | n15828 ;
  assign n70717 = ~n15829 ;
  assign n15965 = n15825 & n70717 ;
  assign n15966 = n15964 | n15965 ;
  assign n15967 = n149 & n15966 ;
  assign n15968 = n15297 & n70705 ;
  assign n15969 = n15859 & n15968 ;
  assign n15970 = n15967 | n15969 ;
  assign n15971 = n70176 & n15970 ;
  assign n70718 = ~n15951 ;
  assign n15972 = n15824 & n70718 ;
  assign n15973 = n15314 | n15824 ;
  assign n70719 = ~n15973 ;
  assign n15974 = n15820 & n70719 ;
  assign n15975 = n15972 | n15974 ;
  assign n15976 = n149 & n15975 ;
  assign n15977 = n15305 & n70705 ;
  assign n15978 = n15859 & n15977 ;
  assign n15979 = n15976 | n15978 ;
  assign n15980 = n69857 & n15979 ;
  assign n70720 = ~n15819 ;
  assign n15981 = n15818 & n70720 ;
  assign n15982 = n15322 | n15818 ;
  assign n70721 = ~n15982 ;
  assign n15983 = n15948 & n70721 ;
  assign n15984 = n15981 | n15983 ;
  assign n15985 = n149 & n15984 ;
  assign n15986 = n15313 & n70705 ;
  assign n15987 = n15859 & n15986 ;
  assign n15988 = n15985 | n15987 ;
  assign n15989 = n69656 & n15988 ;
  assign n70722 = ~n15947 ;
  assign n15990 = n15814 & n70722 ;
  assign n15991 = n15330 | n15814 ;
  assign n70723 = ~n15991 ;
  assign n15992 = n15810 & n70723 ;
  assign n15993 = n15990 | n15992 ;
  assign n15994 = n149 & n15993 ;
  assign n15995 = n15321 & n70705 ;
  assign n15996 = n15859 & n15995 ;
  assign n15997 = n15994 | n15996 ;
  assign n15998 = n69528 & n15997 ;
  assign n70724 = ~n15809 ;
  assign n15999 = n15807 & n70724 ;
  assign n15808 = n15338 | n15807 ;
  assign n70725 = ~n15808 ;
  assign n16000 = n15804 & n70725 ;
  assign n16001 = n15999 | n16000 ;
  assign n16002 = n149 & n16001 ;
  assign n16003 = n15329 & n70705 ;
  assign n16004 = n15859 & n16003 ;
  assign n16005 = n16002 | n16004 ;
  assign n16006 = n69261 & n16005 ;
  assign n70726 = ~n15943 ;
  assign n16007 = n15803 & n70726 ;
  assign n16008 = n15346 | n15803 ;
  assign n70727 = ~n16008 ;
  assign n16009 = n15799 & n70727 ;
  assign n16010 = n16007 | n16009 ;
  assign n16011 = n149 & n16010 ;
  assign n16012 = n15337 & n70705 ;
  assign n16013 = n15859 & n16012 ;
  assign n16014 = n16011 | n16013 ;
  assign n16015 = n69075 & n16014 ;
  assign n70728 = ~n15798 ;
  assign n16016 = n15796 & n70728 ;
  assign n15797 = n15354 | n15796 ;
  assign n70729 = ~n15797 ;
  assign n16017 = n15793 & n70729 ;
  assign n16018 = n16016 | n16017 ;
  assign n16019 = n149 & n16018 ;
  assign n16020 = n15345 & n70705 ;
  assign n16021 = n15859 & n16020 ;
  assign n16022 = n16019 | n16021 ;
  assign n16023 = n68993 & n16022 ;
  assign n70730 = ~n15939 ;
  assign n16024 = n15792 & n70730 ;
  assign n16025 = n15362 | n15792 ;
  assign n70731 = ~n16025 ;
  assign n16026 = n15788 & n70731 ;
  assign n16027 = n16024 | n16026 ;
  assign n16028 = n149 & n16027 ;
  assign n16029 = n15353 & n70705 ;
  assign n16030 = n15859 & n16029 ;
  assign n16031 = n16028 | n16030 ;
  assign n16032 = n68716 & n16031 ;
  assign n70732 = ~n15787 ;
  assign n16033 = n15786 & n70732 ;
  assign n16034 = n15370 | n15786 ;
  assign n70733 = ~n16034 ;
  assign n16035 = n15936 & n70733 ;
  assign n16036 = n16033 | n16035 ;
  assign n16037 = n149 & n16036 ;
  assign n16038 = n15361 & n70705 ;
  assign n16039 = n15859 & n16038 ;
  assign n16040 = n16037 | n16039 ;
  assign n16041 = n68545 & n16040 ;
  assign n70734 = ~n15935 ;
  assign n16042 = n15782 & n70734 ;
  assign n16043 = n15378 | n15782 ;
  assign n70735 = ~n16043 ;
  assign n16044 = n15778 & n70735 ;
  assign n16045 = n16042 | n16044 ;
  assign n16046 = n149 & n16045 ;
  assign n16047 = n15369 & n70705 ;
  assign n16048 = n15859 & n16047 ;
  assign n16049 = n16046 | n16048 ;
  assign n16050 = n68438 & n16049 ;
  assign n70736 = ~n15777 ;
  assign n16051 = n15776 & n70736 ;
  assign n16052 = n15386 | n15776 ;
  assign n70737 = ~n16052 ;
  assign n16053 = n15932 & n70737 ;
  assign n16054 = n16051 | n16053 ;
  assign n16055 = n149 & n16054 ;
  assign n16056 = n15377 & n70705 ;
  assign n16057 = n15859 & n16056 ;
  assign n16058 = n16055 | n16057 ;
  assign n16059 = n68214 & n16058 ;
  assign n70738 = ~n15931 ;
  assign n16060 = n15772 & n70738 ;
  assign n16061 = n15394 | n15772 ;
  assign n70739 = ~n16061 ;
  assign n16062 = n15768 & n70739 ;
  assign n16063 = n16060 | n16062 ;
  assign n16064 = n149 & n16063 ;
  assign n16065 = n15385 & n70705 ;
  assign n16066 = n15859 & n16065 ;
  assign n16067 = n16064 | n16066 ;
  assign n16068 = n68058 & n16067 ;
  assign n70740 = ~n15767 ;
  assign n16069 = n15765 & n70740 ;
  assign n15766 = n15402 | n15765 ;
  assign n70741 = ~n15766 ;
  assign n16070 = n15762 & n70741 ;
  assign n16071 = n16069 | n16070 ;
  assign n16072 = n149 & n16071 ;
  assign n16073 = n15393 & n70705 ;
  assign n16074 = n15859 & n16073 ;
  assign n16075 = n16072 | n16074 ;
  assign n16076 = n67986 & n16075 ;
  assign n70742 = ~n15927 ;
  assign n16077 = n15760 & n70742 ;
  assign n15761 = n15410 | n15760 ;
  assign n70743 = ~n15761 ;
  assign n16078 = n70743 & n15926 ;
  assign n16079 = n16077 | n16078 ;
  assign n16080 = n149 & n16079 ;
  assign n16081 = n15401 & n70705 ;
  assign n16082 = n15859 & n16081 ;
  assign n16083 = n16080 | n16082 ;
  assign n16084 = n67763 & n16083 ;
  assign n70744 = ~n15755 ;
  assign n16085 = n15754 & n70744 ;
  assign n16086 = n15418 | n15754 ;
  assign n70745 = ~n16086 ;
  assign n16087 = n15924 & n70745 ;
  assign n16088 = n16085 | n16087 ;
  assign n16089 = n149 & n16088 ;
  assign n16090 = n15409 & n70705 ;
  assign n16091 = n15859 & n16090 ;
  assign n16092 = n16089 | n16091 ;
  assign n16093 = n67622 & n16092 ;
  assign n70746 = ~n15923 ;
  assign n16094 = n15749 & n70746 ;
  assign n15750 = n15426 | n15749 ;
  assign n70747 = ~n15750 ;
  assign n16095 = n70747 & n15922 ;
  assign n16096 = n16094 | n16095 ;
  assign n16097 = n149 & n16096 ;
  assign n16098 = n15417 & n70705 ;
  assign n16099 = n15859 & n16098 ;
  assign n16100 = n16097 | n16099 ;
  assign n16101 = n67531 & n16100 ;
  assign n70748 = ~n15744 ;
  assign n16102 = n15743 & n70748 ;
  assign n16103 = n15434 | n15743 ;
  assign n70749 = ~n16103 ;
  assign n16104 = n15920 & n70749 ;
  assign n16105 = n16102 | n16104 ;
  assign n16106 = n149 & n16105 ;
  assign n16107 = n15425 & n70705 ;
  assign n16108 = n15859 & n16107 ;
  assign n16109 = n16106 | n16108 ;
  assign n16110 = n67348 & n16109 ;
  assign n70750 = ~n15919 ;
  assign n16111 = n15739 & n70750 ;
  assign n16112 = n15442 | n15739 ;
  assign n70751 = ~n16112 ;
  assign n16113 = n15735 & n70751 ;
  assign n16114 = n16111 | n16113 ;
  assign n16115 = n149 & n16114 ;
  assign n16116 = n15433 & n70705 ;
  assign n16117 = n15859 & n16116 ;
  assign n16118 = n16115 | n16117 ;
  assign n16119 = n67222 & n16118 ;
  assign n70752 = ~n15734 ;
  assign n16120 = n15733 & n70752 ;
  assign n16121 = n15450 | n15733 ;
  assign n70753 = ~n16121 ;
  assign n16122 = n15916 & n70753 ;
  assign n16123 = n16120 | n16122 ;
  assign n16124 = n149 & n16123 ;
  assign n16125 = n15441 & n70705 ;
  assign n16126 = n15859 & n16125 ;
  assign n16127 = n16124 | n16126 ;
  assign n16128 = n67164 & n16127 ;
  assign n70754 = ~n15915 ;
  assign n16129 = n15728 & n70754 ;
  assign n15729 = n15458 | n15728 ;
  assign n70755 = ~n15729 ;
  assign n16130 = n70755 & n15914 ;
  assign n16131 = n16129 | n16130 ;
  assign n16132 = n149 & n16131 ;
  assign n16133 = n15449 & n70705 ;
  assign n16134 = n15859 & n16133 ;
  assign n16135 = n16132 | n16134 ;
  assign n16136 = n66979 & n16135 ;
  assign n70756 = ~n15723 ;
  assign n16137 = n15722 & n70756 ;
  assign n16138 = n15466 | n15722 ;
  assign n70757 = ~n16138 ;
  assign n16139 = n15912 & n70757 ;
  assign n16140 = n16137 | n16139 ;
  assign n16141 = n149 & n16140 ;
  assign n16142 = n15457 & n70705 ;
  assign n16143 = n15859 & n16142 ;
  assign n16144 = n16141 | n16143 ;
  assign n16145 = n66868 & n16144 ;
  assign n70758 = ~n15911 ;
  assign n16146 = n15718 & n70758 ;
  assign n16147 = n15474 | n15718 ;
  assign n70759 = ~n16147 ;
  assign n16148 = n15714 & n70759 ;
  assign n16149 = n16146 | n16148 ;
  assign n16150 = n149 & n16149 ;
  assign n16151 = n15465 & n70705 ;
  assign n16152 = n15859 & n16151 ;
  assign n16153 = n16150 | n16152 ;
  assign n16154 = n66797 & n16153 ;
  assign n70760 = ~n15713 ;
  assign n16155 = n15711 & n70760 ;
  assign n15712 = n15482 | n15711 ;
  assign n70761 = ~n15712 ;
  assign n16156 = n15708 & n70761 ;
  assign n16157 = n16155 | n16156 ;
  assign n16158 = n149 & n16157 ;
  assign n16159 = n15473 & n70705 ;
  assign n16160 = n15859 & n16159 ;
  assign n16161 = n16158 | n16160 ;
  assign n16162 = n66654 & n16161 ;
  assign n70762 = ~n15907 ;
  assign n16163 = n15706 & n70762 ;
  assign n15707 = n15490 | n15706 ;
  assign n70763 = ~n15707 ;
  assign n16164 = n70763 & n15906 ;
  assign n16165 = n16163 | n16164 ;
  assign n16166 = n149 & n16165 ;
  assign n16167 = n15481 & n70705 ;
  assign n16168 = n15859 & n16167 ;
  assign n16169 = n16166 | n16168 ;
  assign n16170 = n66560 & n16169 ;
  assign n70764 = ~n15701 ;
  assign n16171 = n15699 & n70764 ;
  assign n15700 = n15498 | n15699 ;
  assign n70765 = ~n15700 ;
  assign n16172 = n15696 & n70765 ;
  assign n16173 = n16171 | n16172 ;
  assign n16174 = n149 & n16173 ;
  assign n16175 = n15489 & n70705 ;
  assign n16176 = n15859 & n16175 ;
  assign n16177 = n16174 | n16176 ;
  assign n16178 = n66505 & n16177 ;
  assign n70766 = ~n15903 ;
  assign n16179 = n15695 & n70766 ;
  assign n16180 = n15506 | n15695 ;
  assign n70767 = ~n16180 ;
  assign n16181 = n15691 & n70767 ;
  assign n16182 = n16179 | n16181 ;
  assign n16183 = n149 & n16182 ;
  assign n16184 = n15497 & n70705 ;
  assign n16185 = n15859 & n16184 ;
  assign n16186 = n16183 | n16185 ;
  assign n16187 = n66379 & n16186 ;
  assign n70768 = ~n15690 ;
  assign n16188 = n15689 & n70768 ;
  assign n16189 = n15514 | n15689 ;
  assign n70769 = ~n16189 ;
  assign n16190 = n15900 & n70769 ;
  assign n16191 = n16188 | n16190 ;
  assign n16192 = n149 & n16191 ;
  assign n16193 = n15505 & n70705 ;
  assign n16194 = n15859 & n16193 ;
  assign n16195 = n16192 | n16194 ;
  assign n16196 = n66299 & n16195 ;
  assign n70770 = ~n15899 ;
  assign n16197 = n15685 & n70770 ;
  assign n16198 = n15522 | n15685 ;
  assign n70771 = ~n16198 ;
  assign n16199 = n15681 & n70771 ;
  assign n16200 = n16197 | n16199 ;
  assign n16201 = n149 & n16200 ;
  assign n16202 = n15513 & n70705 ;
  assign n16203 = n15859 & n16202 ;
  assign n16204 = n16201 | n16203 ;
  assign n16205 = n66244 & n16204 ;
  assign n70772 = ~n15680 ;
  assign n16206 = n15679 & n70772 ;
  assign n16207 = n15530 | n15679 ;
  assign n70773 = ~n16207 ;
  assign n16208 = n15896 & n70773 ;
  assign n16209 = n16206 | n16208 ;
  assign n16210 = n149 & n16209 ;
  assign n16211 = n15521 & n70705 ;
  assign n16212 = n15859 & n16211 ;
  assign n16213 = n16210 | n16212 ;
  assign n16214 = n66145 & n16213 ;
  assign n70774 = ~n15895 ;
  assign n16215 = n15675 & n70774 ;
  assign n16216 = n15538 | n15675 ;
  assign n70775 = ~n16216 ;
  assign n16217 = n15671 & n70775 ;
  assign n16218 = n16215 | n16217 ;
  assign n16219 = n149 & n16218 ;
  assign n16220 = n15529 & n70705 ;
  assign n16221 = n15859 & n16220 ;
  assign n16222 = n16219 | n16221 ;
  assign n16223 = n66081 & n16222 ;
  assign n70776 = ~n15670 ;
  assign n16224 = n15668 & n70776 ;
  assign n15669 = n15546 | n15668 ;
  assign n70777 = ~n15669 ;
  assign n16225 = n15665 & n70777 ;
  assign n16226 = n16224 | n16225 ;
  assign n16227 = n149 & n16226 ;
  assign n16228 = n15537 & n70705 ;
  assign n16229 = n15859 & n16228 ;
  assign n16230 = n16227 | n16229 ;
  assign n16231 = n66043 & n16230 ;
  assign n70778 = ~n15891 ;
  assign n16232 = n15664 & n70778 ;
  assign n16233 = n15555 | n15664 ;
  assign n70779 = ~n16233 ;
  assign n16234 = n15660 & n70779 ;
  assign n16235 = n16232 | n16234 ;
  assign n16236 = n149 & n16235 ;
  assign n16237 = n15545 & n70705 ;
  assign n16238 = n15859 & n16237 ;
  assign n16239 = n16236 | n16238 ;
  assign n16240 = n65960 & n16239 ;
  assign n70780 = ~n15659 ;
  assign n16241 = n15658 & n70780 ;
  assign n16242 = n15564 | n15658 ;
  assign n70781 = ~n16242 ;
  assign n16243 = n15888 & n70781 ;
  assign n16244 = n16241 | n16243 ;
  assign n16245 = n149 & n16244 ;
  assign n16246 = n15554 & n70705 ;
  assign n16247 = n15859 & n16246 ;
  assign n16248 = n16245 | n16247 ;
  assign n16249 = n65909 & n16248 ;
  assign n70782 = ~n15887 ;
  assign n16250 = n15654 & n70782 ;
  assign n16251 = n15572 | n15654 ;
  assign n70783 = ~n16251 ;
  assign n16252 = n15650 & n70783 ;
  assign n16253 = n16250 | n16252 ;
  assign n16254 = n149 & n16253 ;
  assign n16255 = n15563 & n70705 ;
  assign n16256 = n15859 & n16255 ;
  assign n16257 = n16254 | n16256 ;
  assign n16258 = n65877 & n16257 ;
  assign n70784 = ~n15649 ;
  assign n16259 = n15648 & n70784 ;
  assign n16260 = n15580 | n15648 ;
  assign n70785 = ~n16260 ;
  assign n16261 = n15884 & n70785 ;
  assign n16262 = n16259 | n16261 ;
  assign n16263 = n149 & n16262 ;
  assign n16264 = n15571 & n70705 ;
  assign n16265 = n15859 & n16264 ;
  assign n16266 = n16263 | n16265 ;
  assign n16267 = n65820 & n16266 ;
  assign n70786 = ~n15883 ;
  assign n16268 = n15644 & n70786 ;
  assign n16269 = n15588 | n15644 ;
  assign n70787 = ~n16269 ;
  assign n16270 = n15640 & n70787 ;
  assign n16271 = n16268 | n16270 ;
  assign n16272 = n149 & n16271 ;
  assign n16273 = n15579 & n70705 ;
  assign n16274 = n15859 & n16273 ;
  assign n16275 = n16272 | n16274 ;
  assign n16276 = n65791 & n16275 ;
  assign n70788 = ~n15639 ;
  assign n16278 = n15638 & n70788 ;
  assign n16277 = n15597 | n15638 ;
  assign n70789 = ~n16277 ;
  assign n16279 = n15635 & n70789 ;
  assign n16280 = n16278 | n16279 ;
  assign n16281 = n149 & n16280 ;
  assign n16282 = n15587 & n70705 ;
  assign n16283 = n15859 & n16282 ;
  assign n16284 = n16281 | n16283 ;
  assign n16285 = n65772 & n16284 ;
  assign n70790 = ~n15879 ;
  assign n16287 = n15634 & n70790 ;
  assign n16286 = n15605 | n15634 ;
  assign n70791 = ~n16286 ;
  assign n16288 = n15878 & n70791 ;
  assign n16289 = n16287 | n16288 ;
  assign n16290 = n149 & n16289 ;
  assign n16291 = n15596 & n70705 ;
  assign n16292 = n15859 & n16291 ;
  assign n16293 = n16290 | n16292 ;
  assign n16294 = n65746 & n16293 ;
  assign n70792 = ~n15629 ;
  assign n16296 = n15628 & n70792 ;
  assign n16295 = n15625 | n15628 ;
  assign n70793 = ~n16295 ;
  assign n16297 = n15624 & n70793 ;
  assign n16298 = n16296 | n16297 ;
  assign n16299 = n149 & n16298 ;
  assign n16300 = n15604 & n70705 ;
  assign n16301 = n15859 & n16300 ;
  assign n16302 = n16299 | n16301 ;
  assign n16303 = n65721 & n16302 ;
  assign n16304 = n15621 & n15623 ;
  assign n16305 = n70614 & n16304 ;
  assign n70794 = ~n16305 ;
  assign n16306 = n15624 & n70794 ;
  assign n16307 = n149 & n16306 ;
  assign n16308 = n15618 & n70705 ;
  assign n16309 = n15859 & n16308 ;
  assign n16310 = n16307 | n16309 ;
  assign n16311 = n65686 & n16310 ;
  assign n15862 = n15623 & n149 ;
  assign n16320 = x64 & n149 ;
  assign n70795 = ~n16320 ;
  assign n16321 = x20 & n70795 ;
  assign n16322 = n15862 | n16321 ;
  assign n16324 = x65 & n16322 ;
  assign n16316 = n15858 | n16315 ;
  assign n16317 = n70705 & n16316 ;
  assign n70796 = ~n16317 ;
  assign n16318 = x64 & n70796 ;
  assign n70797 = ~n16318 ;
  assign n16319 = x20 & n70797 ;
  assign n16323 = x65 | n15862 ;
  assign n16325 = n16319 | n16323 ;
  assign n70798 = ~n16324 ;
  assign n16326 = n70798 & n16325 ;
  assign n70799 = ~x19 ;
  assign n16327 = n70799 & x64 ;
  assign n16328 = n16326 | n16327 ;
  assign n16329 = n65670 & n16322 ;
  assign n70800 = ~n16329 ;
  assign n16330 = n16328 & n70800 ;
  assign n70801 = ~n16309 ;
  assign n16331 = x66 & n70801 ;
  assign n70802 = ~n16307 ;
  assign n16332 = n70802 & n16331 ;
  assign n16333 = n16311 | n16332 ;
  assign n16334 = n16330 | n16333 ;
  assign n70803 = ~n16311 ;
  assign n16335 = n70803 & n16334 ;
  assign n70804 = ~n16301 ;
  assign n16336 = x67 & n70804 ;
  assign n70805 = ~n16299 ;
  assign n16337 = n70805 & n16336 ;
  assign n16338 = n16303 | n16337 ;
  assign n16339 = n16335 | n16338 ;
  assign n70806 = ~n16303 ;
  assign n16340 = n70806 & n16339 ;
  assign n70807 = ~n16292 ;
  assign n16341 = x68 & n70807 ;
  assign n70808 = ~n16290 ;
  assign n16342 = n70808 & n16341 ;
  assign n16343 = n16294 | n16342 ;
  assign n16344 = n16340 | n16343 ;
  assign n70809 = ~n16294 ;
  assign n16345 = n70809 & n16344 ;
  assign n70810 = ~n16283 ;
  assign n16346 = x69 & n70810 ;
  assign n70811 = ~n16281 ;
  assign n16347 = n70811 & n16346 ;
  assign n16348 = n16285 | n16347 ;
  assign n16350 = n16345 | n16348 ;
  assign n70812 = ~n16285 ;
  assign n16351 = n70812 & n16350 ;
  assign n70813 = ~n16274 ;
  assign n16352 = x70 & n70813 ;
  assign n70814 = ~n16272 ;
  assign n16353 = n70814 & n16352 ;
  assign n16354 = n16276 | n16353 ;
  assign n16355 = n16351 | n16354 ;
  assign n70815 = ~n16276 ;
  assign n16356 = n70815 & n16355 ;
  assign n70816 = ~n16265 ;
  assign n16357 = x71 & n70816 ;
  assign n70817 = ~n16263 ;
  assign n16358 = n70817 & n16357 ;
  assign n16359 = n16267 | n16358 ;
  assign n16361 = n16356 | n16359 ;
  assign n70818 = ~n16267 ;
  assign n16362 = n70818 & n16361 ;
  assign n70819 = ~n16256 ;
  assign n16363 = x72 & n70819 ;
  assign n70820 = ~n16254 ;
  assign n16364 = n70820 & n16363 ;
  assign n16365 = n16258 | n16364 ;
  assign n16366 = n16362 | n16365 ;
  assign n70821 = ~n16258 ;
  assign n16367 = n70821 & n16366 ;
  assign n70822 = ~n16247 ;
  assign n16368 = x73 & n70822 ;
  assign n70823 = ~n16245 ;
  assign n16369 = n70823 & n16368 ;
  assign n16370 = n16249 | n16369 ;
  assign n16372 = n16367 | n16370 ;
  assign n70824 = ~n16249 ;
  assign n16373 = n70824 & n16372 ;
  assign n70825 = ~n16238 ;
  assign n16374 = x74 & n70825 ;
  assign n70826 = ~n16236 ;
  assign n16375 = n70826 & n16374 ;
  assign n16376 = n16240 | n16375 ;
  assign n16377 = n16373 | n16376 ;
  assign n70827 = ~n16240 ;
  assign n16378 = n70827 & n16377 ;
  assign n70828 = ~n16229 ;
  assign n16379 = x75 & n70828 ;
  assign n70829 = ~n16227 ;
  assign n16380 = n70829 & n16379 ;
  assign n16381 = n16231 | n16380 ;
  assign n16383 = n16378 | n16381 ;
  assign n70830 = ~n16231 ;
  assign n16384 = n70830 & n16383 ;
  assign n70831 = ~n16221 ;
  assign n16385 = x76 & n70831 ;
  assign n70832 = ~n16219 ;
  assign n16386 = n70832 & n16385 ;
  assign n16387 = n16223 | n16386 ;
  assign n16388 = n16384 | n16387 ;
  assign n70833 = ~n16223 ;
  assign n16389 = n70833 & n16388 ;
  assign n70834 = ~n16212 ;
  assign n16390 = x77 & n70834 ;
  assign n70835 = ~n16210 ;
  assign n16391 = n70835 & n16390 ;
  assign n16392 = n16214 | n16391 ;
  assign n16394 = n16389 | n16392 ;
  assign n70836 = ~n16214 ;
  assign n16395 = n70836 & n16394 ;
  assign n70837 = ~n16203 ;
  assign n16396 = x78 & n70837 ;
  assign n70838 = ~n16201 ;
  assign n16397 = n70838 & n16396 ;
  assign n16398 = n16205 | n16397 ;
  assign n16399 = n16395 | n16398 ;
  assign n70839 = ~n16205 ;
  assign n16400 = n70839 & n16399 ;
  assign n70840 = ~n16194 ;
  assign n16401 = x79 & n70840 ;
  assign n70841 = ~n16192 ;
  assign n16402 = n70841 & n16401 ;
  assign n16403 = n16196 | n16402 ;
  assign n16405 = n16400 | n16403 ;
  assign n70842 = ~n16196 ;
  assign n16406 = n70842 & n16405 ;
  assign n70843 = ~n16185 ;
  assign n16407 = x80 & n70843 ;
  assign n70844 = ~n16183 ;
  assign n16408 = n70844 & n16407 ;
  assign n16409 = n16187 | n16408 ;
  assign n16410 = n16406 | n16409 ;
  assign n70845 = ~n16187 ;
  assign n16411 = n70845 & n16410 ;
  assign n70846 = ~n16176 ;
  assign n16412 = x81 & n70846 ;
  assign n70847 = ~n16174 ;
  assign n16413 = n70847 & n16412 ;
  assign n16414 = n16178 | n16413 ;
  assign n16416 = n16411 | n16414 ;
  assign n70848 = ~n16178 ;
  assign n16417 = n70848 & n16416 ;
  assign n70849 = ~n16168 ;
  assign n16418 = x82 & n70849 ;
  assign n70850 = ~n16166 ;
  assign n16419 = n70850 & n16418 ;
  assign n16420 = n16170 | n16419 ;
  assign n16421 = n16417 | n16420 ;
  assign n70851 = ~n16170 ;
  assign n16422 = n70851 & n16421 ;
  assign n70852 = ~n16160 ;
  assign n16423 = x83 & n70852 ;
  assign n70853 = ~n16158 ;
  assign n16424 = n70853 & n16423 ;
  assign n16425 = n16162 | n16424 ;
  assign n16427 = n16422 | n16425 ;
  assign n70854 = ~n16162 ;
  assign n16428 = n70854 & n16427 ;
  assign n70855 = ~n16152 ;
  assign n16429 = x84 & n70855 ;
  assign n70856 = ~n16150 ;
  assign n16430 = n70856 & n16429 ;
  assign n16431 = n16154 | n16430 ;
  assign n16432 = n16428 | n16431 ;
  assign n70857 = ~n16154 ;
  assign n16433 = n70857 & n16432 ;
  assign n70858 = ~n16143 ;
  assign n16434 = x85 & n70858 ;
  assign n70859 = ~n16141 ;
  assign n16435 = n70859 & n16434 ;
  assign n16436 = n16145 | n16435 ;
  assign n16438 = n16433 | n16436 ;
  assign n70860 = ~n16145 ;
  assign n16439 = n70860 & n16438 ;
  assign n70861 = ~n16134 ;
  assign n16440 = x86 & n70861 ;
  assign n70862 = ~n16132 ;
  assign n16441 = n70862 & n16440 ;
  assign n16442 = n16136 | n16441 ;
  assign n16443 = n16439 | n16442 ;
  assign n70863 = ~n16136 ;
  assign n16444 = n70863 & n16443 ;
  assign n70864 = ~n16126 ;
  assign n16445 = x87 & n70864 ;
  assign n70865 = ~n16124 ;
  assign n16446 = n70865 & n16445 ;
  assign n16447 = n16128 | n16446 ;
  assign n16449 = n16444 | n16447 ;
  assign n70866 = ~n16128 ;
  assign n16450 = n70866 & n16449 ;
  assign n70867 = ~n16117 ;
  assign n16451 = x88 & n70867 ;
  assign n70868 = ~n16115 ;
  assign n16452 = n70868 & n16451 ;
  assign n16453 = n16119 | n16452 ;
  assign n16454 = n16450 | n16453 ;
  assign n70869 = ~n16119 ;
  assign n16455 = n70869 & n16454 ;
  assign n70870 = ~n16108 ;
  assign n16456 = x89 & n70870 ;
  assign n70871 = ~n16106 ;
  assign n16457 = n70871 & n16456 ;
  assign n16458 = n16110 | n16457 ;
  assign n16460 = n16455 | n16458 ;
  assign n70872 = ~n16110 ;
  assign n16461 = n70872 & n16460 ;
  assign n70873 = ~n16099 ;
  assign n16462 = x90 & n70873 ;
  assign n70874 = ~n16097 ;
  assign n16463 = n70874 & n16462 ;
  assign n16464 = n16101 | n16463 ;
  assign n16465 = n16461 | n16464 ;
  assign n70875 = ~n16101 ;
  assign n16466 = n70875 & n16465 ;
  assign n70876 = ~n16091 ;
  assign n16467 = x91 & n70876 ;
  assign n70877 = ~n16089 ;
  assign n16468 = n70877 & n16467 ;
  assign n16469 = n16093 | n16468 ;
  assign n16471 = n16466 | n16469 ;
  assign n70878 = ~n16093 ;
  assign n16472 = n70878 & n16471 ;
  assign n70879 = ~n16082 ;
  assign n16473 = x92 & n70879 ;
  assign n70880 = ~n16080 ;
  assign n16474 = n70880 & n16473 ;
  assign n16475 = n16084 | n16474 ;
  assign n16476 = n16472 | n16475 ;
  assign n70881 = ~n16084 ;
  assign n16477 = n70881 & n16476 ;
  assign n70882 = ~n16074 ;
  assign n16478 = x93 & n70882 ;
  assign n70883 = ~n16072 ;
  assign n16479 = n70883 & n16478 ;
  assign n16480 = n16076 | n16479 ;
  assign n16482 = n16477 | n16480 ;
  assign n70884 = ~n16076 ;
  assign n16483 = n70884 & n16482 ;
  assign n70885 = ~n16066 ;
  assign n16484 = x94 & n70885 ;
  assign n70886 = ~n16064 ;
  assign n16485 = n70886 & n16484 ;
  assign n16486 = n16068 | n16485 ;
  assign n16487 = n16483 | n16486 ;
  assign n70887 = ~n16068 ;
  assign n16488 = n70887 & n16487 ;
  assign n70888 = ~n16057 ;
  assign n16489 = x95 & n70888 ;
  assign n70889 = ~n16055 ;
  assign n16490 = n70889 & n16489 ;
  assign n16491 = n16059 | n16490 ;
  assign n16493 = n16488 | n16491 ;
  assign n70890 = ~n16059 ;
  assign n16494 = n70890 & n16493 ;
  assign n70891 = ~n16048 ;
  assign n16495 = x96 & n70891 ;
  assign n70892 = ~n16046 ;
  assign n16496 = n70892 & n16495 ;
  assign n16497 = n16050 | n16496 ;
  assign n16498 = n16494 | n16497 ;
  assign n70893 = ~n16050 ;
  assign n16499 = n70893 & n16498 ;
  assign n70894 = ~n16039 ;
  assign n16500 = x97 & n70894 ;
  assign n70895 = ~n16037 ;
  assign n16501 = n70895 & n16500 ;
  assign n16502 = n16041 | n16501 ;
  assign n16504 = n16499 | n16502 ;
  assign n70896 = ~n16041 ;
  assign n16505 = n70896 & n16504 ;
  assign n70897 = ~n16030 ;
  assign n16506 = x98 & n70897 ;
  assign n70898 = ~n16028 ;
  assign n16507 = n70898 & n16506 ;
  assign n16508 = n16032 | n16507 ;
  assign n16509 = n16505 | n16508 ;
  assign n70899 = ~n16032 ;
  assign n16510 = n70899 & n16509 ;
  assign n70900 = ~n16021 ;
  assign n16511 = x99 & n70900 ;
  assign n70901 = ~n16019 ;
  assign n16512 = n70901 & n16511 ;
  assign n16513 = n16023 | n16512 ;
  assign n16515 = n16510 | n16513 ;
  assign n70902 = ~n16023 ;
  assign n16516 = n70902 & n16515 ;
  assign n70903 = ~n16013 ;
  assign n16517 = x100 & n70903 ;
  assign n70904 = ~n16011 ;
  assign n16518 = n70904 & n16517 ;
  assign n16519 = n16015 | n16518 ;
  assign n16520 = n16516 | n16519 ;
  assign n70905 = ~n16015 ;
  assign n16521 = n70905 & n16520 ;
  assign n70906 = ~n16004 ;
  assign n16522 = x101 & n70906 ;
  assign n70907 = ~n16002 ;
  assign n16523 = n70907 & n16522 ;
  assign n16524 = n16006 | n16523 ;
  assign n16526 = n16521 | n16524 ;
  assign n70908 = ~n16006 ;
  assign n16527 = n70908 & n16526 ;
  assign n70909 = ~n15996 ;
  assign n16528 = x102 & n70909 ;
  assign n70910 = ~n15994 ;
  assign n16529 = n70910 & n16528 ;
  assign n16530 = n15998 | n16529 ;
  assign n16531 = n16527 | n16530 ;
  assign n70911 = ~n15998 ;
  assign n16532 = n70911 & n16531 ;
  assign n70912 = ~n15987 ;
  assign n16533 = x103 & n70912 ;
  assign n70913 = ~n15985 ;
  assign n16534 = n70913 & n16533 ;
  assign n16535 = n15989 | n16534 ;
  assign n16537 = n16532 | n16535 ;
  assign n70914 = ~n15989 ;
  assign n16538 = n70914 & n16537 ;
  assign n70915 = ~n15978 ;
  assign n16539 = x104 & n70915 ;
  assign n70916 = ~n15976 ;
  assign n16540 = n70916 & n16539 ;
  assign n16541 = n15980 | n16540 ;
  assign n16542 = n16538 | n16541 ;
  assign n70917 = ~n15980 ;
  assign n16543 = n70917 & n16542 ;
  assign n70918 = ~n15969 ;
  assign n16544 = x105 & n70918 ;
  assign n70919 = ~n15967 ;
  assign n16545 = n70919 & n16544 ;
  assign n16546 = n15971 | n16545 ;
  assign n16548 = n16543 | n16546 ;
  assign n70920 = ~n15971 ;
  assign n16549 = n70920 & n16548 ;
  assign n70921 = ~n15961 ;
  assign n16550 = x106 & n70921 ;
  assign n70922 = ~n15959 ;
  assign n16551 = n70922 & n16550 ;
  assign n16552 = n15963 | n16551 ;
  assign n16553 = n16549 | n16552 ;
  assign n70923 = ~n15963 ;
  assign n16554 = n70923 & n16553 ;
  assign n70924 = ~n15868 ;
  assign n16555 = x107 & n70924 ;
  assign n70925 = ~n15866 ;
  assign n16556 = n70925 & n16555 ;
  assign n16557 = n15870 | n16556 ;
  assign n16559 = n16554 | n16557 ;
  assign n70926 = ~n15870 ;
  assign n16560 = n70926 & n16559 ;
  assign n70927 = ~x108 ;
  assign n16571 = n70927 & n16570 ;
  assign n70928 = ~n16569 ;
  assign n16572 = x108 & n70928 ;
  assign n70929 = ~n16567 ;
  assign n16573 = n70929 & n16572 ;
  assign n16574 = n465 | n467 ;
  assign n16575 = n16573 | n16574 ;
  assign n16576 = n16571 | n16575 ;
  assign n16578 = n16560 | n16576 ;
  assign n70930 = ~n16577 ;
  assign n16579 = n70930 & n16578 ;
  assign n16693 = n15870 | n16573 ;
  assign n16694 = n16571 | n16693 ;
  assign n70931 = ~n16694 ;
  assign n16695 = n16559 & n70931 ;
  assign n16582 = n15862 | n16319 ;
  assign n16583 = x65 & n16582 ;
  assign n70932 = ~n16583 ;
  assign n16584 = n16325 & n70932 ;
  assign n16585 = n16327 | n16584 ;
  assign n16586 = n70800 & n16585 ;
  assign n16587 = n16333 | n16586 ;
  assign n16588 = n70803 & n16587 ;
  assign n16590 = n16338 | n16588 ;
  assign n16591 = n70806 & n16590 ;
  assign n16593 = n16343 | n16591 ;
  assign n16594 = n70809 & n16593 ;
  assign n16595 = n16348 | n16594 ;
  assign n16596 = n70812 & n16595 ;
  assign n16597 = n16354 | n16596 ;
  assign n16599 = n70815 & n16597 ;
  assign n16600 = n16359 | n16599 ;
  assign n16601 = n70818 & n16600 ;
  assign n16602 = n16365 | n16601 ;
  assign n16604 = n70821 & n16602 ;
  assign n16605 = n16370 | n16604 ;
  assign n16606 = n70824 & n16605 ;
  assign n16607 = n16376 | n16606 ;
  assign n16609 = n70827 & n16607 ;
  assign n16610 = n16381 | n16609 ;
  assign n16611 = n70830 & n16610 ;
  assign n16612 = n16387 | n16611 ;
  assign n16614 = n70833 & n16612 ;
  assign n16615 = n16392 | n16614 ;
  assign n16616 = n70836 & n16615 ;
  assign n16617 = n16398 | n16616 ;
  assign n16619 = n70839 & n16617 ;
  assign n16620 = n16403 | n16619 ;
  assign n16621 = n70842 & n16620 ;
  assign n16622 = n16409 | n16621 ;
  assign n16624 = n70845 & n16622 ;
  assign n16625 = n16414 | n16624 ;
  assign n16626 = n70848 & n16625 ;
  assign n16627 = n16420 | n16626 ;
  assign n16629 = n70851 & n16627 ;
  assign n16630 = n16425 | n16629 ;
  assign n16631 = n70854 & n16630 ;
  assign n16632 = n16431 | n16631 ;
  assign n16634 = n70857 & n16632 ;
  assign n16635 = n16436 | n16634 ;
  assign n16636 = n70860 & n16635 ;
  assign n16637 = n16442 | n16636 ;
  assign n16639 = n70863 & n16637 ;
  assign n16640 = n16447 | n16639 ;
  assign n16641 = n70866 & n16640 ;
  assign n16642 = n16453 | n16641 ;
  assign n16644 = n70869 & n16642 ;
  assign n16645 = n16458 | n16644 ;
  assign n16646 = n70872 & n16645 ;
  assign n16647 = n16464 | n16646 ;
  assign n16649 = n70875 & n16647 ;
  assign n16650 = n16469 | n16649 ;
  assign n16651 = n70878 & n16650 ;
  assign n16652 = n16475 | n16651 ;
  assign n16654 = n70881 & n16652 ;
  assign n16655 = n16480 | n16654 ;
  assign n16656 = n70884 & n16655 ;
  assign n16657 = n16486 | n16656 ;
  assign n16659 = n70887 & n16657 ;
  assign n16660 = n16491 | n16659 ;
  assign n16661 = n70890 & n16660 ;
  assign n16662 = n16497 | n16661 ;
  assign n16664 = n70893 & n16662 ;
  assign n16665 = n16502 | n16664 ;
  assign n16666 = n70896 & n16665 ;
  assign n16667 = n16508 | n16666 ;
  assign n16669 = n70899 & n16667 ;
  assign n16670 = n16513 | n16669 ;
  assign n16671 = n70902 & n16670 ;
  assign n16672 = n16519 | n16671 ;
  assign n16674 = n70905 & n16672 ;
  assign n16675 = n16524 | n16674 ;
  assign n16676 = n70908 & n16675 ;
  assign n16677 = n16530 | n16676 ;
  assign n16679 = n70911 & n16677 ;
  assign n16680 = n16535 | n16679 ;
  assign n16681 = n70914 & n16680 ;
  assign n16682 = n16541 | n16681 ;
  assign n16684 = n70917 & n16682 ;
  assign n16685 = n16546 | n16684 ;
  assign n16686 = n70920 & n16685 ;
  assign n16687 = n16552 | n16686 ;
  assign n16689 = n70923 & n16687 ;
  assign n16690 = n16557 | n16689 ;
  assign n16691 = n70926 & n16690 ;
  assign n16696 = n16571 | n16573 ;
  assign n70933 = ~n16691 ;
  assign n16697 = n70933 & n16696 ;
  assign n16698 = n16695 | n16697 ;
  assign n148 = ~n16579 ;
  assign n16699 = n148 & n16698 ;
  assign n16692 = n16576 | n16691 ;
  assign n16700 = n15856 & n16570 ;
  assign n16701 = n16692 & n16700 ;
  assign n16702 = n16699 | n16701 ;
  assign n70935 = ~x109 ;
  assign n16703 = n70935 & n16702 ;
  assign n70936 = ~n16701 ;
  assign n17317 = x109 & n70936 ;
  assign n70937 = ~n16699 ;
  assign n17318 = n70937 & n17317 ;
  assign n17319 = n16703 | n17318 ;
  assign n70938 = ~n16554 ;
  assign n16558 = n70938 & n16557 ;
  assign n16704 = n15963 | n16557 ;
  assign n70939 = ~n16704 ;
  assign n16705 = n16687 & n70939 ;
  assign n16706 = n16558 | n16705 ;
  assign n16707 = n148 & n16706 ;
  assign n16708 = n15869 & n70930 ;
  assign n16709 = n16692 & n16708 ;
  assign n16710 = n16707 | n16709 ;
  assign n16711 = n70927 & n16710 ;
  assign n70940 = ~n16686 ;
  assign n16688 = n16552 & n70940 ;
  assign n16712 = n15971 | n16552 ;
  assign n70941 = ~n16712 ;
  assign n16713 = n16548 & n70941 ;
  assign n16714 = n16688 | n16713 ;
  assign n16715 = n148 & n16714 ;
  assign n16716 = n15962 & n70930 ;
  assign n16717 = n16692 & n16716 ;
  assign n16718 = n16715 | n16717 ;
  assign n16719 = n70609 & n16718 ;
  assign n70942 = ~n16717 ;
  assign n17305 = x107 & n70942 ;
  assign n70943 = ~n16715 ;
  assign n17306 = n70943 & n17305 ;
  assign n17307 = n16719 | n17306 ;
  assign n70944 = ~n16543 ;
  assign n16547 = n70944 & n16546 ;
  assign n16720 = n15980 | n16546 ;
  assign n70945 = ~n16720 ;
  assign n16721 = n16682 & n70945 ;
  assign n16722 = n16547 | n16721 ;
  assign n16723 = n148 & n16722 ;
  assign n16724 = n15970 & n70930 ;
  assign n16725 = n16692 & n16724 ;
  assign n16726 = n16723 | n16725 ;
  assign n16727 = n70276 & n16726 ;
  assign n70946 = ~n16681 ;
  assign n16683 = n16541 & n70946 ;
  assign n16728 = n15989 | n16541 ;
  assign n70947 = ~n16728 ;
  assign n16729 = n16537 & n70947 ;
  assign n16730 = n16683 | n16729 ;
  assign n16731 = n148 & n16730 ;
  assign n16732 = n15979 & n70930 ;
  assign n16733 = n16692 & n16732 ;
  assign n16734 = n16731 | n16733 ;
  assign n16735 = n70176 & n16734 ;
  assign n70948 = ~n16733 ;
  assign n17293 = x105 & n70948 ;
  assign n70949 = ~n16731 ;
  assign n17294 = n70949 & n17293 ;
  assign n17295 = n16735 | n17294 ;
  assign n70950 = ~n16532 ;
  assign n16536 = n70950 & n16535 ;
  assign n16736 = n15998 | n16535 ;
  assign n70951 = ~n16736 ;
  assign n16737 = n16677 & n70951 ;
  assign n16738 = n16536 | n16737 ;
  assign n16739 = n148 & n16738 ;
  assign n16740 = n15988 & n70930 ;
  assign n16741 = n16692 & n16740 ;
  assign n16742 = n16739 | n16741 ;
  assign n16743 = n69857 & n16742 ;
  assign n70952 = ~n16676 ;
  assign n16678 = n16530 & n70952 ;
  assign n16744 = n16006 | n16530 ;
  assign n70953 = ~n16744 ;
  assign n16745 = n16526 & n70953 ;
  assign n16746 = n16678 | n16745 ;
  assign n16747 = n148 & n16746 ;
  assign n16748 = n15997 & n70930 ;
  assign n16749 = n16692 & n16748 ;
  assign n16750 = n16747 | n16749 ;
  assign n16751 = n69656 & n16750 ;
  assign n70954 = ~n16749 ;
  assign n17281 = x103 & n70954 ;
  assign n70955 = ~n16747 ;
  assign n17282 = n70955 & n17281 ;
  assign n17283 = n16751 | n17282 ;
  assign n70956 = ~n16521 ;
  assign n16525 = n70956 & n16524 ;
  assign n16752 = n16015 | n16524 ;
  assign n70957 = ~n16752 ;
  assign n16753 = n16672 & n70957 ;
  assign n16754 = n16525 | n16753 ;
  assign n16755 = n148 & n16754 ;
  assign n16756 = n16005 & n70930 ;
  assign n16757 = n16692 & n16756 ;
  assign n16758 = n16755 | n16757 ;
  assign n16759 = n69528 & n16758 ;
  assign n70958 = ~n16671 ;
  assign n16673 = n16519 & n70958 ;
  assign n16760 = n16023 | n16519 ;
  assign n70959 = ~n16760 ;
  assign n16761 = n16515 & n70959 ;
  assign n16762 = n16673 | n16761 ;
  assign n16763 = n148 & n16762 ;
  assign n16764 = n16014 & n70930 ;
  assign n16765 = n16692 & n16764 ;
  assign n16766 = n16763 | n16765 ;
  assign n16767 = n69261 & n16766 ;
  assign n70960 = ~n16765 ;
  assign n17269 = x101 & n70960 ;
  assign n70961 = ~n16763 ;
  assign n17270 = n70961 & n17269 ;
  assign n17271 = n16767 | n17270 ;
  assign n70962 = ~n16510 ;
  assign n16514 = n70962 & n16513 ;
  assign n16768 = n16032 | n16513 ;
  assign n70963 = ~n16768 ;
  assign n16769 = n16667 & n70963 ;
  assign n16770 = n16514 | n16769 ;
  assign n16771 = n148 & n16770 ;
  assign n16772 = n16022 & n70930 ;
  assign n16773 = n16692 & n16772 ;
  assign n16774 = n16771 | n16773 ;
  assign n16775 = n69075 & n16774 ;
  assign n70964 = ~n16666 ;
  assign n16668 = n16508 & n70964 ;
  assign n16776 = n16041 | n16508 ;
  assign n70965 = ~n16776 ;
  assign n16777 = n16504 & n70965 ;
  assign n16778 = n16668 | n16777 ;
  assign n16779 = n148 & n16778 ;
  assign n16780 = n16031 & n70930 ;
  assign n16781 = n16692 & n16780 ;
  assign n16782 = n16779 | n16781 ;
  assign n16783 = n68993 & n16782 ;
  assign n70966 = ~n16781 ;
  assign n17257 = x99 & n70966 ;
  assign n70967 = ~n16779 ;
  assign n17258 = n70967 & n17257 ;
  assign n17259 = n16783 | n17258 ;
  assign n70968 = ~n16499 ;
  assign n16503 = n70968 & n16502 ;
  assign n16784 = n16050 | n16502 ;
  assign n70969 = ~n16784 ;
  assign n16785 = n16662 & n70969 ;
  assign n16786 = n16503 | n16785 ;
  assign n16787 = n148 & n16786 ;
  assign n16788 = n16040 & n70930 ;
  assign n16789 = n16692 & n16788 ;
  assign n16790 = n16787 | n16789 ;
  assign n16791 = n68716 & n16790 ;
  assign n70970 = ~n16661 ;
  assign n16663 = n16497 & n70970 ;
  assign n16792 = n16059 | n16497 ;
  assign n70971 = ~n16792 ;
  assign n16793 = n16493 & n70971 ;
  assign n16794 = n16663 | n16793 ;
  assign n16795 = n148 & n16794 ;
  assign n16796 = n16049 & n70930 ;
  assign n16797 = n16692 & n16796 ;
  assign n16798 = n16795 | n16797 ;
  assign n16799 = n68545 & n16798 ;
  assign n70972 = ~n16797 ;
  assign n17245 = x97 & n70972 ;
  assign n70973 = ~n16795 ;
  assign n17246 = n70973 & n17245 ;
  assign n17247 = n16799 | n17246 ;
  assign n70974 = ~n16488 ;
  assign n16492 = n70974 & n16491 ;
  assign n16800 = n16068 | n16491 ;
  assign n70975 = ~n16800 ;
  assign n16801 = n16657 & n70975 ;
  assign n16802 = n16492 | n16801 ;
  assign n16803 = n148 & n16802 ;
  assign n16804 = n16058 & n70930 ;
  assign n16805 = n16692 & n16804 ;
  assign n16806 = n16803 | n16805 ;
  assign n16807 = n68438 & n16806 ;
  assign n70976 = ~n16656 ;
  assign n16658 = n16486 & n70976 ;
  assign n16808 = n16076 | n16486 ;
  assign n70977 = ~n16808 ;
  assign n16809 = n16482 & n70977 ;
  assign n16810 = n16658 | n16809 ;
  assign n16811 = n148 & n16810 ;
  assign n16812 = n16067 & n70930 ;
  assign n16813 = n16692 & n16812 ;
  assign n16814 = n16811 | n16813 ;
  assign n16815 = n68214 & n16814 ;
  assign n70978 = ~n16813 ;
  assign n17233 = x95 & n70978 ;
  assign n70979 = ~n16811 ;
  assign n17234 = n70979 & n17233 ;
  assign n17235 = n16815 | n17234 ;
  assign n70980 = ~n16477 ;
  assign n16481 = n70980 & n16480 ;
  assign n16816 = n16084 | n16480 ;
  assign n70981 = ~n16816 ;
  assign n16817 = n16652 & n70981 ;
  assign n16818 = n16481 | n16817 ;
  assign n16819 = n148 & n16818 ;
  assign n16820 = n16075 & n70930 ;
  assign n16821 = n16692 & n16820 ;
  assign n16822 = n16819 | n16821 ;
  assign n16823 = n68058 & n16822 ;
  assign n70982 = ~n16651 ;
  assign n16653 = n16475 & n70982 ;
  assign n16824 = n16093 | n16475 ;
  assign n70983 = ~n16824 ;
  assign n16825 = n16471 & n70983 ;
  assign n16826 = n16653 | n16825 ;
  assign n16827 = n148 & n16826 ;
  assign n16828 = n16083 & n70930 ;
  assign n16829 = n16692 & n16828 ;
  assign n16830 = n16827 | n16829 ;
  assign n16831 = n67986 & n16830 ;
  assign n70984 = ~n16829 ;
  assign n17221 = x93 & n70984 ;
  assign n70985 = ~n16827 ;
  assign n17222 = n70985 & n17221 ;
  assign n17223 = n16831 | n17222 ;
  assign n70986 = ~n16466 ;
  assign n16470 = n70986 & n16469 ;
  assign n16832 = n16101 | n16469 ;
  assign n70987 = ~n16832 ;
  assign n16833 = n16647 & n70987 ;
  assign n16834 = n16470 | n16833 ;
  assign n16835 = n148 & n16834 ;
  assign n16836 = n16092 & n70930 ;
  assign n16837 = n16692 & n16836 ;
  assign n16838 = n16835 | n16837 ;
  assign n16839 = n67763 & n16838 ;
  assign n70988 = ~n16646 ;
  assign n16648 = n16464 & n70988 ;
  assign n16840 = n16110 | n16464 ;
  assign n70989 = ~n16840 ;
  assign n16841 = n16460 & n70989 ;
  assign n16842 = n16648 | n16841 ;
  assign n16843 = n148 & n16842 ;
  assign n16844 = n16100 & n70930 ;
  assign n16845 = n16692 & n16844 ;
  assign n16846 = n16843 | n16845 ;
  assign n16847 = n67622 & n16846 ;
  assign n70990 = ~n16845 ;
  assign n17209 = x91 & n70990 ;
  assign n70991 = ~n16843 ;
  assign n17210 = n70991 & n17209 ;
  assign n17211 = n16847 | n17210 ;
  assign n70992 = ~n16455 ;
  assign n16459 = n70992 & n16458 ;
  assign n16848 = n16119 | n16458 ;
  assign n70993 = ~n16848 ;
  assign n16849 = n16642 & n70993 ;
  assign n16850 = n16459 | n16849 ;
  assign n16851 = n148 & n16850 ;
  assign n16852 = n16109 & n70930 ;
  assign n16853 = n16692 & n16852 ;
  assign n16854 = n16851 | n16853 ;
  assign n16855 = n67531 & n16854 ;
  assign n70994 = ~n16641 ;
  assign n16643 = n16453 & n70994 ;
  assign n16856 = n16128 | n16453 ;
  assign n70995 = ~n16856 ;
  assign n16857 = n16449 & n70995 ;
  assign n16858 = n16643 | n16857 ;
  assign n16859 = n148 & n16858 ;
  assign n16860 = n16118 & n70930 ;
  assign n16861 = n16692 & n16860 ;
  assign n16862 = n16859 | n16861 ;
  assign n16863 = n67348 & n16862 ;
  assign n70996 = ~n16861 ;
  assign n17197 = x89 & n70996 ;
  assign n70997 = ~n16859 ;
  assign n17198 = n70997 & n17197 ;
  assign n17199 = n16863 | n17198 ;
  assign n70998 = ~n16444 ;
  assign n16448 = n70998 & n16447 ;
  assign n16864 = n16136 | n16447 ;
  assign n70999 = ~n16864 ;
  assign n16865 = n16637 & n70999 ;
  assign n16866 = n16448 | n16865 ;
  assign n16867 = n148 & n16866 ;
  assign n16868 = n16127 & n70930 ;
  assign n16869 = n16692 & n16868 ;
  assign n16870 = n16867 | n16869 ;
  assign n16871 = n67222 & n16870 ;
  assign n71000 = ~n16636 ;
  assign n16638 = n16442 & n71000 ;
  assign n16872 = n16145 | n16442 ;
  assign n71001 = ~n16872 ;
  assign n16873 = n16438 & n71001 ;
  assign n16874 = n16638 | n16873 ;
  assign n16875 = n148 & n16874 ;
  assign n16876 = n16135 & n70930 ;
  assign n16877 = n16692 & n16876 ;
  assign n16878 = n16875 | n16877 ;
  assign n16879 = n67164 & n16878 ;
  assign n71002 = ~n16877 ;
  assign n17185 = x87 & n71002 ;
  assign n71003 = ~n16875 ;
  assign n17186 = n71003 & n17185 ;
  assign n17187 = n16879 | n17186 ;
  assign n71004 = ~n16433 ;
  assign n16437 = n71004 & n16436 ;
  assign n16880 = n16154 | n16436 ;
  assign n71005 = ~n16880 ;
  assign n16881 = n16632 & n71005 ;
  assign n16882 = n16437 | n16881 ;
  assign n16883 = n148 & n16882 ;
  assign n16884 = n16144 & n70930 ;
  assign n16885 = n16692 & n16884 ;
  assign n16886 = n16883 | n16885 ;
  assign n16887 = n66979 & n16886 ;
  assign n71006 = ~n16631 ;
  assign n16633 = n16431 & n71006 ;
  assign n16888 = n16162 | n16431 ;
  assign n71007 = ~n16888 ;
  assign n16889 = n16427 & n71007 ;
  assign n16890 = n16633 | n16889 ;
  assign n16891 = n148 & n16890 ;
  assign n16892 = n16153 & n70930 ;
  assign n16893 = n16692 & n16892 ;
  assign n16894 = n16891 | n16893 ;
  assign n16895 = n66868 & n16894 ;
  assign n71008 = ~n16893 ;
  assign n17173 = x85 & n71008 ;
  assign n71009 = ~n16891 ;
  assign n17174 = n71009 & n17173 ;
  assign n17175 = n16895 | n17174 ;
  assign n71010 = ~n16422 ;
  assign n16426 = n71010 & n16425 ;
  assign n16896 = n16170 | n16425 ;
  assign n71011 = ~n16896 ;
  assign n16897 = n16627 & n71011 ;
  assign n16898 = n16426 | n16897 ;
  assign n16899 = n148 & n16898 ;
  assign n16900 = n16161 & n70930 ;
  assign n16901 = n16692 & n16900 ;
  assign n16902 = n16899 | n16901 ;
  assign n16903 = n66797 & n16902 ;
  assign n71012 = ~n16626 ;
  assign n16628 = n16420 & n71012 ;
  assign n16904 = n16178 | n16420 ;
  assign n71013 = ~n16904 ;
  assign n16905 = n16416 & n71013 ;
  assign n16906 = n16628 | n16905 ;
  assign n16907 = n148 & n16906 ;
  assign n16908 = n16169 & n70930 ;
  assign n16909 = n16692 & n16908 ;
  assign n16910 = n16907 | n16909 ;
  assign n16911 = n66654 & n16910 ;
  assign n71014 = ~n16909 ;
  assign n17161 = x83 & n71014 ;
  assign n71015 = ~n16907 ;
  assign n17162 = n71015 & n17161 ;
  assign n17163 = n16911 | n17162 ;
  assign n71016 = ~n16411 ;
  assign n16415 = n71016 & n16414 ;
  assign n16912 = n16187 | n16414 ;
  assign n71017 = ~n16912 ;
  assign n16913 = n16622 & n71017 ;
  assign n16914 = n16415 | n16913 ;
  assign n16915 = n148 & n16914 ;
  assign n16916 = n16177 & n70930 ;
  assign n16917 = n16692 & n16916 ;
  assign n16918 = n16915 | n16917 ;
  assign n16919 = n66560 & n16918 ;
  assign n71018 = ~n16621 ;
  assign n16623 = n16409 & n71018 ;
  assign n16920 = n16196 | n16409 ;
  assign n71019 = ~n16920 ;
  assign n16921 = n16405 & n71019 ;
  assign n16922 = n16623 | n16921 ;
  assign n16923 = n148 & n16922 ;
  assign n16924 = n16186 & n70930 ;
  assign n16925 = n16692 & n16924 ;
  assign n16926 = n16923 | n16925 ;
  assign n16927 = n66505 & n16926 ;
  assign n71020 = ~n16925 ;
  assign n17149 = x81 & n71020 ;
  assign n71021 = ~n16923 ;
  assign n17150 = n71021 & n17149 ;
  assign n17151 = n16927 | n17150 ;
  assign n71022 = ~n16400 ;
  assign n16404 = n71022 & n16403 ;
  assign n16928 = n16205 | n16403 ;
  assign n71023 = ~n16928 ;
  assign n16929 = n16617 & n71023 ;
  assign n16930 = n16404 | n16929 ;
  assign n16931 = n148 & n16930 ;
  assign n16932 = n16195 & n70930 ;
  assign n16933 = n16692 & n16932 ;
  assign n16934 = n16931 | n16933 ;
  assign n16935 = n66379 & n16934 ;
  assign n71024 = ~n16616 ;
  assign n16618 = n16398 & n71024 ;
  assign n16936 = n16214 | n16398 ;
  assign n71025 = ~n16936 ;
  assign n16937 = n16394 & n71025 ;
  assign n16938 = n16618 | n16937 ;
  assign n16939 = n148 & n16938 ;
  assign n16940 = n16204 & n70930 ;
  assign n16941 = n16692 & n16940 ;
  assign n16942 = n16939 | n16941 ;
  assign n16943 = n66299 & n16942 ;
  assign n71026 = ~n16941 ;
  assign n17137 = x79 & n71026 ;
  assign n71027 = ~n16939 ;
  assign n17138 = n71027 & n17137 ;
  assign n17139 = n16943 | n17138 ;
  assign n71028 = ~n16389 ;
  assign n16393 = n71028 & n16392 ;
  assign n16944 = n16223 | n16392 ;
  assign n71029 = ~n16944 ;
  assign n16945 = n16612 & n71029 ;
  assign n16946 = n16393 | n16945 ;
  assign n16947 = n148 & n16946 ;
  assign n16948 = n16213 & n70930 ;
  assign n16949 = n16692 & n16948 ;
  assign n16950 = n16947 | n16949 ;
  assign n16951 = n66244 & n16950 ;
  assign n71030 = ~n16611 ;
  assign n16613 = n16387 & n71030 ;
  assign n16952 = n16231 | n16387 ;
  assign n71031 = ~n16952 ;
  assign n16953 = n16383 & n71031 ;
  assign n16954 = n16613 | n16953 ;
  assign n16955 = n148 & n16954 ;
  assign n16956 = n16222 & n70930 ;
  assign n16957 = n16692 & n16956 ;
  assign n16958 = n16955 | n16957 ;
  assign n16959 = n66145 & n16958 ;
  assign n71032 = ~n16957 ;
  assign n17125 = x77 & n71032 ;
  assign n71033 = ~n16955 ;
  assign n17126 = n71033 & n17125 ;
  assign n17127 = n16959 | n17126 ;
  assign n71034 = ~n16378 ;
  assign n16382 = n71034 & n16381 ;
  assign n16960 = n16240 | n16381 ;
  assign n71035 = ~n16960 ;
  assign n16961 = n16607 & n71035 ;
  assign n16962 = n16382 | n16961 ;
  assign n16963 = n148 & n16962 ;
  assign n16964 = n16230 & n70930 ;
  assign n16965 = n16692 & n16964 ;
  assign n16966 = n16963 | n16965 ;
  assign n16967 = n66081 & n16966 ;
  assign n71036 = ~n16606 ;
  assign n16608 = n16376 & n71036 ;
  assign n16968 = n16249 | n16376 ;
  assign n71037 = ~n16968 ;
  assign n16969 = n16372 & n71037 ;
  assign n16970 = n16608 | n16969 ;
  assign n16971 = n148 & n16970 ;
  assign n16972 = n16239 & n70930 ;
  assign n16973 = n16692 & n16972 ;
  assign n16974 = n16971 | n16973 ;
  assign n16975 = n66043 & n16974 ;
  assign n71038 = ~n16973 ;
  assign n17113 = x75 & n71038 ;
  assign n71039 = ~n16971 ;
  assign n17114 = n71039 & n17113 ;
  assign n17115 = n16975 | n17114 ;
  assign n71040 = ~n16367 ;
  assign n16371 = n71040 & n16370 ;
  assign n16976 = n16258 | n16370 ;
  assign n71041 = ~n16976 ;
  assign n16977 = n16602 & n71041 ;
  assign n16978 = n16371 | n16977 ;
  assign n16979 = n148 & n16978 ;
  assign n16980 = n16248 & n70930 ;
  assign n16981 = n16692 & n16980 ;
  assign n16982 = n16979 | n16981 ;
  assign n16983 = n65960 & n16982 ;
  assign n71042 = ~n16601 ;
  assign n16603 = n16365 & n71042 ;
  assign n16984 = n16267 | n16365 ;
  assign n71043 = ~n16984 ;
  assign n16985 = n16361 & n71043 ;
  assign n16986 = n16603 | n16985 ;
  assign n16987 = n148 & n16986 ;
  assign n16988 = n16257 & n70930 ;
  assign n16989 = n16692 & n16988 ;
  assign n16990 = n16987 | n16989 ;
  assign n16991 = n65909 & n16990 ;
  assign n71044 = ~n16989 ;
  assign n17101 = x73 & n71044 ;
  assign n71045 = ~n16987 ;
  assign n17102 = n71045 & n17101 ;
  assign n17103 = n16991 | n17102 ;
  assign n71046 = ~n16356 ;
  assign n16360 = n71046 & n16359 ;
  assign n16992 = n16276 | n16359 ;
  assign n71047 = ~n16992 ;
  assign n16993 = n16597 & n71047 ;
  assign n16994 = n16360 | n16993 ;
  assign n16995 = n148 & n16994 ;
  assign n16996 = n16266 & n70930 ;
  assign n16997 = n16692 & n16996 ;
  assign n16998 = n16995 | n16997 ;
  assign n16999 = n65877 & n16998 ;
  assign n71048 = ~n16596 ;
  assign n16598 = n16354 & n71048 ;
  assign n17000 = n16285 | n16354 ;
  assign n71049 = ~n17000 ;
  assign n17001 = n16350 & n71049 ;
  assign n17002 = n16598 | n17001 ;
  assign n17003 = n148 & n17002 ;
  assign n17004 = n16275 & n70930 ;
  assign n17005 = n16692 & n17004 ;
  assign n17006 = n17003 | n17005 ;
  assign n17007 = n65820 & n17006 ;
  assign n71050 = ~n17005 ;
  assign n17089 = x71 & n71050 ;
  assign n71051 = ~n17003 ;
  assign n17090 = n71051 & n17089 ;
  assign n17091 = n17007 | n17090 ;
  assign n71052 = ~n16345 ;
  assign n16349 = n71052 & n16348 ;
  assign n17008 = n16294 | n16348 ;
  assign n71053 = ~n17008 ;
  assign n17009 = n16593 & n71053 ;
  assign n17010 = n16349 | n17009 ;
  assign n17011 = n148 & n17010 ;
  assign n17012 = n16284 & n70930 ;
  assign n17013 = n16692 & n17012 ;
  assign n17014 = n17011 | n17013 ;
  assign n17015 = n65791 & n17014 ;
  assign n71054 = ~n16591 ;
  assign n16592 = n16343 & n71054 ;
  assign n17016 = n16303 | n16343 ;
  assign n71055 = ~n17016 ;
  assign n17017 = n16339 & n71055 ;
  assign n17018 = n16592 | n17017 ;
  assign n17019 = n148 & n17018 ;
  assign n17020 = n16293 & n70930 ;
  assign n17021 = n16692 & n17020 ;
  assign n17022 = n17019 | n17021 ;
  assign n17023 = n65772 & n17022 ;
  assign n71056 = ~n17021 ;
  assign n17078 = x69 & n71056 ;
  assign n71057 = ~n17019 ;
  assign n17079 = n71057 & n17078 ;
  assign n17080 = n17023 | n17079 ;
  assign n71058 = ~n16335 ;
  assign n16589 = n71058 & n16338 ;
  assign n17024 = n16311 | n16338 ;
  assign n71059 = ~n17024 ;
  assign n17025 = n16334 & n71059 ;
  assign n17026 = n16589 | n17025 ;
  assign n17027 = n148 & n17026 ;
  assign n17028 = n16302 & n70930 ;
  assign n17029 = n16692 & n17028 ;
  assign n17030 = n17027 | n17029 ;
  assign n17031 = n65746 & n17030 ;
  assign n71060 = ~n16330 ;
  assign n17033 = n71060 & n16333 ;
  assign n17032 = n16329 | n16333 ;
  assign n71061 = ~n17032 ;
  assign n17034 = n16328 & n71061 ;
  assign n17035 = n17033 | n17034 ;
  assign n17036 = n148 & n17035 ;
  assign n17037 = n16310 & n70930 ;
  assign n17038 = n16692 & n17037 ;
  assign n17039 = n17036 | n17038 ;
  assign n17040 = n65721 & n17039 ;
  assign n71062 = ~n17038 ;
  assign n17068 = x67 & n71062 ;
  assign n71063 = ~n17036 ;
  assign n17069 = n71063 & n17068 ;
  assign n17070 = n17040 | n17069 ;
  assign n17041 = n16325 & n16327 ;
  assign n17042 = n70798 & n17041 ;
  assign n71064 = ~n17042 ;
  assign n17043 = n16585 & n71064 ;
  assign n17044 = n148 & n17043 ;
  assign n17045 = n16322 & n70930 ;
  assign n17046 = n16692 & n17045 ;
  assign n17047 = n17044 | n17046 ;
  assign n17048 = n65686 & n17047 ;
  assign n71065 = ~x18 ;
  assign n17058 = n71065 & x64 ;
  assign n16580 = n16327 & n148 ;
  assign n17049 = n70930 & n16692 ;
  assign n71066 = ~n17049 ;
  assign n17050 = x64 & n71066 ;
  assign n71067 = ~n17050 ;
  assign n17051 = x19 & n71067 ;
  assign n17052 = n16580 | n17051 ;
  assign n17053 = x65 & n17052 ;
  assign n16581 = x64 & n148 ;
  assign n71068 = ~n16581 ;
  assign n17054 = x19 & n71068 ;
  assign n17055 = n16327 & n71066 ;
  assign n17056 = x65 | n17055 ;
  assign n17057 = n17054 | n17056 ;
  assign n71069 = ~n17053 ;
  assign n17059 = n71069 & n17057 ;
  assign n17060 = n17058 | n17059 ;
  assign n17061 = n16580 | n17054 ;
  assign n17062 = n65670 & n17061 ;
  assign n71070 = ~n17062 ;
  assign n17063 = n17060 & n71070 ;
  assign n71071 = ~n17046 ;
  assign n17064 = x66 & n71071 ;
  assign n71072 = ~n17044 ;
  assign n17065 = n71072 & n17064 ;
  assign n17066 = n17048 | n17065 ;
  assign n17067 = n17063 | n17066 ;
  assign n71073 = ~n17048 ;
  assign n17071 = n71073 & n17067 ;
  assign n17072 = n17070 | n17071 ;
  assign n71074 = ~n17040 ;
  assign n17073 = n71074 & n17072 ;
  assign n71075 = ~n17029 ;
  assign n17074 = x68 & n71075 ;
  assign n71076 = ~n17027 ;
  assign n17075 = n71076 & n17074 ;
  assign n17076 = n17031 | n17075 ;
  assign n17077 = n17073 | n17076 ;
  assign n71077 = ~n17031 ;
  assign n17081 = n71077 & n17077 ;
  assign n17082 = n17080 | n17081 ;
  assign n71078 = ~n17023 ;
  assign n17083 = n71078 & n17082 ;
  assign n71079 = ~n17013 ;
  assign n17084 = x70 & n71079 ;
  assign n71080 = ~n17011 ;
  assign n17085 = n71080 & n17084 ;
  assign n17086 = n17015 | n17085 ;
  assign n17088 = n17083 | n17086 ;
  assign n71081 = ~n17015 ;
  assign n17093 = n71081 & n17088 ;
  assign n17094 = n17091 | n17093 ;
  assign n71082 = ~n17007 ;
  assign n17095 = n71082 & n17094 ;
  assign n71083 = ~n16997 ;
  assign n17096 = x72 & n71083 ;
  assign n71084 = ~n16995 ;
  assign n17097 = n71084 & n17096 ;
  assign n17098 = n16999 | n17097 ;
  assign n17100 = n17095 | n17098 ;
  assign n71085 = ~n16999 ;
  assign n17105 = n71085 & n17100 ;
  assign n17106 = n17103 | n17105 ;
  assign n71086 = ~n16991 ;
  assign n17107 = n71086 & n17106 ;
  assign n71087 = ~n16981 ;
  assign n17108 = x74 & n71087 ;
  assign n71088 = ~n16979 ;
  assign n17109 = n71088 & n17108 ;
  assign n17110 = n16983 | n17109 ;
  assign n17112 = n17107 | n17110 ;
  assign n71089 = ~n16983 ;
  assign n17117 = n71089 & n17112 ;
  assign n17118 = n17115 | n17117 ;
  assign n71090 = ~n16975 ;
  assign n17119 = n71090 & n17118 ;
  assign n71091 = ~n16965 ;
  assign n17120 = x76 & n71091 ;
  assign n71092 = ~n16963 ;
  assign n17121 = n71092 & n17120 ;
  assign n17122 = n16967 | n17121 ;
  assign n17124 = n17119 | n17122 ;
  assign n71093 = ~n16967 ;
  assign n17129 = n71093 & n17124 ;
  assign n17130 = n17127 | n17129 ;
  assign n71094 = ~n16959 ;
  assign n17131 = n71094 & n17130 ;
  assign n71095 = ~n16949 ;
  assign n17132 = x78 & n71095 ;
  assign n71096 = ~n16947 ;
  assign n17133 = n71096 & n17132 ;
  assign n17134 = n16951 | n17133 ;
  assign n17136 = n17131 | n17134 ;
  assign n71097 = ~n16951 ;
  assign n17141 = n71097 & n17136 ;
  assign n17142 = n17139 | n17141 ;
  assign n71098 = ~n16943 ;
  assign n17143 = n71098 & n17142 ;
  assign n71099 = ~n16933 ;
  assign n17144 = x80 & n71099 ;
  assign n71100 = ~n16931 ;
  assign n17145 = n71100 & n17144 ;
  assign n17146 = n16935 | n17145 ;
  assign n17148 = n17143 | n17146 ;
  assign n71101 = ~n16935 ;
  assign n17153 = n71101 & n17148 ;
  assign n17154 = n17151 | n17153 ;
  assign n71102 = ~n16927 ;
  assign n17155 = n71102 & n17154 ;
  assign n71103 = ~n16917 ;
  assign n17156 = x82 & n71103 ;
  assign n71104 = ~n16915 ;
  assign n17157 = n71104 & n17156 ;
  assign n17158 = n16919 | n17157 ;
  assign n17160 = n17155 | n17158 ;
  assign n71105 = ~n16919 ;
  assign n17165 = n71105 & n17160 ;
  assign n17166 = n17163 | n17165 ;
  assign n71106 = ~n16911 ;
  assign n17167 = n71106 & n17166 ;
  assign n71107 = ~n16901 ;
  assign n17168 = x84 & n71107 ;
  assign n71108 = ~n16899 ;
  assign n17169 = n71108 & n17168 ;
  assign n17170 = n16903 | n17169 ;
  assign n17172 = n17167 | n17170 ;
  assign n71109 = ~n16903 ;
  assign n17177 = n71109 & n17172 ;
  assign n17178 = n17175 | n17177 ;
  assign n71110 = ~n16895 ;
  assign n17179 = n71110 & n17178 ;
  assign n71111 = ~n16885 ;
  assign n17180 = x86 & n71111 ;
  assign n71112 = ~n16883 ;
  assign n17181 = n71112 & n17180 ;
  assign n17182 = n16887 | n17181 ;
  assign n17184 = n17179 | n17182 ;
  assign n71113 = ~n16887 ;
  assign n17189 = n71113 & n17184 ;
  assign n17190 = n17187 | n17189 ;
  assign n71114 = ~n16879 ;
  assign n17191 = n71114 & n17190 ;
  assign n71115 = ~n16869 ;
  assign n17192 = x88 & n71115 ;
  assign n71116 = ~n16867 ;
  assign n17193 = n71116 & n17192 ;
  assign n17194 = n16871 | n17193 ;
  assign n17196 = n17191 | n17194 ;
  assign n71117 = ~n16871 ;
  assign n17201 = n71117 & n17196 ;
  assign n17202 = n17199 | n17201 ;
  assign n71118 = ~n16863 ;
  assign n17203 = n71118 & n17202 ;
  assign n71119 = ~n16853 ;
  assign n17204 = x90 & n71119 ;
  assign n71120 = ~n16851 ;
  assign n17205 = n71120 & n17204 ;
  assign n17206 = n16855 | n17205 ;
  assign n17208 = n17203 | n17206 ;
  assign n71121 = ~n16855 ;
  assign n17213 = n71121 & n17208 ;
  assign n17214 = n17211 | n17213 ;
  assign n71122 = ~n16847 ;
  assign n17215 = n71122 & n17214 ;
  assign n71123 = ~n16837 ;
  assign n17216 = x92 & n71123 ;
  assign n71124 = ~n16835 ;
  assign n17217 = n71124 & n17216 ;
  assign n17218 = n16839 | n17217 ;
  assign n17220 = n17215 | n17218 ;
  assign n71125 = ~n16839 ;
  assign n17225 = n71125 & n17220 ;
  assign n17226 = n17223 | n17225 ;
  assign n71126 = ~n16831 ;
  assign n17227 = n71126 & n17226 ;
  assign n71127 = ~n16821 ;
  assign n17228 = x94 & n71127 ;
  assign n71128 = ~n16819 ;
  assign n17229 = n71128 & n17228 ;
  assign n17230 = n16823 | n17229 ;
  assign n17232 = n17227 | n17230 ;
  assign n71129 = ~n16823 ;
  assign n17237 = n71129 & n17232 ;
  assign n17238 = n17235 | n17237 ;
  assign n71130 = ~n16815 ;
  assign n17239 = n71130 & n17238 ;
  assign n71131 = ~n16805 ;
  assign n17240 = x96 & n71131 ;
  assign n71132 = ~n16803 ;
  assign n17241 = n71132 & n17240 ;
  assign n17242 = n16807 | n17241 ;
  assign n17244 = n17239 | n17242 ;
  assign n71133 = ~n16807 ;
  assign n17249 = n71133 & n17244 ;
  assign n17250 = n17247 | n17249 ;
  assign n71134 = ~n16799 ;
  assign n17251 = n71134 & n17250 ;
  assign n71135 = ~n16789 ;
  assign n17252 = x98 & n71135 ;
  assign n71136 = ~n16787 ;
  assign n17253 = n71136 & n17252 ;
  assign n17254 = n16791 | n17253 ;
  assign n17256 = n17251 | n17254 ;
  assign n71137 = ~n16791 ;
  assign n17261 = n71137 & n17256 ;
  assign n17262 = n17259 | n17261 ;
  assign n71138 = ~n16783 ;
  assign n17263 = n71138 & n17262 ;
  assign n71139 = ~n16773 ;
  assign n17264 = x100 & n71139 ;
  assign n71140 = ~n16771 ;
  assign n17265 = n71140 & n17264 ;
  assign n17266 = n16775 | n17265 ;
  assign n17268 = n17263 | n17266 ;
  assign n71141 = ~n16775 ;
  assign n17273 = n71141 & n17268 ;
  assign n17274 = n17271 | n17273 ;
  assign n71142 = ~n16767 ;
  assign n17275 = n71142 & n17274 ;
  assign n71143 = ~n16757 ;
  assign n17276 = x102 & n71143 ;
  assign n71144 = ~n16755 ;
  assign n17277 = n71144 & n17276 ;
  assign n17278 = n16759 | n17277 ;
  assign n17280 = n17275 | n17278 ;
  assign n71145 = ~n16759 ;
  assign n17285 = n71145 & n17280 ;
  assign n17286 = n17283 | n17285 ;
  assign n71146 = ~n16751 ;
  assign n17287 = n71146 & n17286 ;
  assign n71147 = ~n16741 ;
  assign n17288 = x104 & n71147 ;
  assign n71148 = ~n16739 ;
  assign n17289 = n71148 & n17288 ;
  assign n17290 = n16743 | n17289 ;
  assign n17292 = n17287 | n17290 ;
  assign n71149 = ~n16743 ;
  assign n17297 = n71149 & n17292 ;
  assign n17298 = n17295 | n17297 ;
  assign n71150 = ~n16735 ;
  assign n17299 = n71150 & n17298 ;
  assign n71151 = ~n16725 ;
  assign n17300 = x106 & n71151 ;
  assign n71152 = ~n16723 ;
  assign n17301 = n71152 & n17300 ;
  assign n17302 = n16727 | n17301 ;
  assign n17304 = n17299 | n17302 ;
  assign n71153 = ~n16727 ;
  assign n17309 = n71153 & n17304 ;
  assign n17310 = n17307 | n17309 ;
  assign n71154 = ~n16719 ;
  assign n17311 = n71154 & n17310 ;
  assign n71155 = ~n16709 ;
  assign n17312 = x108 & n71155 ;
  assign n71156 = ~n16707 ;
  assign n17313 = n71156 & n17312 ;
  assign n17314 = n16711 | n17313 ;
  assign n17316 = n17311 | n17314 ;
  assign n71157 = ~n16711 ;
  assign n17320 = n71157 & n17316 ;
  assign n17321 = n17319 | n17320 ;
  assign n71158 = ~n16703 ;
  assign n17322 = n71158 & n17321 ;
  assign n17325 = n17322 | n17324 ;
  assign n71159 = ~n16702 ;
  assign n17327 = n71159 & n17325 ;
  assign n71160 = ~n17320 ;
  assign n18035 = n17319 & n71160 ;
  assign n17330 = x65 & n17061 ;
  assign n71161 = ~n17330 ;
  assign n17331 = n17057 & n71161 ;
  assign n17333 = n17058 | n17331 ;
  assign n17335 = n71070 & n17333 ;
  assign n17336 = n17066 | n17335 ;
  assign n17337 = n71073 & n17336 ;
  assign n17338 = n17070 | n17337 ;
  assign n17339 = n71074 & n17338 ;
  assign n17340 = n17076 | n17339 ;
  assign n17341 = n71077 & n17340 ;
  assign n17342 = n17080 | n17341 ;
  assign n17343 = n71078 & n17342 ;
  assign n17344 = n17086 | n17343 ;
  assign n17345 = n71081 & n17344 ;
  assign n17346 = n17091 | n17345 ;
  assign n17347 = n71082 & n17346 ;
  assign n17348 = n17098 | n17347 ;
  assign n17349 = n71085 & n17348 ;
  assign n17350 = n17103 | n17349 ;
  assign n17351 = n71086 & n17350 ;
  assign n17352 = n17110 | n17351 ;
  assign n17353 = n71089 & n17352 ;
  assign n17354 = n17115 | n17353 ;
  assign n17355 = n71090 & n17354 ;
  assign n17356 = n17122 | n17355 ;
  assign n17357 = n71093 & n17356 ;
  assign n17358 = n17127 | n17357 ;
  assign n17359 = n71094 & n17358 ;
  assign n17360 = n17134 | n17359 ;
  assign n17361 = n71097 & n17360 ;
  assign n17362 = n17139 | n17361 ;
  assign n17363 = n71098 & n17362 ;
  assign n17364 = n17146 | n17363 ;
  assign n17365 = n71101 & n17364 ;
  assign n17366 = n17151 | n17365 ;
  assign n17367 = n71102 & n17366 ;
  assign n17368 = n17158 | n17367 ;
  assign n17369 = n71105 & n17368 ;
  assign n17370 = n17163 | n17369 ;
  assign n17371 = n71106 & n17370 ;
  assign n17372 = n17170 | n17371 ;
  assign n17373 = n71109 & n17372 ;
  assign n17374 = n17175 | n17373 ;
  assign n17375 = n71110 & n17374 ;
  assign n17376 = n17182 | n17375 ;
  assign n17377 = n71113 & n17376 ;
  assign n17378 = n17187 | n17377 ;
  assign n17379 = n71114 & n17378 ;
  assign n17380 = n17194 | n17379 ;
  assign n17381 = n71117 & n17380 ;
  assign n17382 = n17199 | n17381 ;
  assign n17383 = n71118 & n17382 ;
  assign n17384 = n17206 | n17383 ;
  assign n17385 = n71121 & n17384 ;
  assign n17386 = n17211 | n17385 ;
  assign n17387 = n71122 & n17386 ;
  assign n17388 = n17218 | n17387 ;
  assign n17389 = n71125 & n17388 ;
  assign n17390 = n17223 | n17389 ;
  assign n17391 = n71126 & n17390 ;
  assign n17392 = n17230 | n17391 ;
  assign n17393 = n71129 & n17392 ;
  assign n17394 = n17235 | n17393 ;
  assign n17395 = n71130 & n17394 ;
  assign n17396 = n17242 | n17395 ;
  assign n17397 = n71133 & n17396 ;
  assign n17398 = n17247 | n17397 ;
  assign n17399 = n71134 & n17398 ;
  assign n17400 = n17254 | n17399 ;
  assign n17401 = n71137 & n17400 ;
  assign n17402 = n17259 | n17401 ;
  assign n17403 = n71138 & n17402 ;
  assign n17404 = n17266 | n17403 ;
  assign n17405 = n71141 & n17404 ;
  assign n17406 = n17271 | n17405 ;
  assign n17407 = n71142 & n17406 ;
  assign n17408 = n17278 | n17407 ;
  assign n17409 = n71145 & n17408 ;
  assign n17410 = n17283 | n17409 ;
  assign n17411 = n71146 & n17410 ;
  assign n17412 = n17290 | n17411 ;
  assign n17413 = n71149 & n17412 ;
  assign n17414 = n17295 | n17413 ;
  assign n17415 = n71150 & n17414 ;
  assign n17416 = n17302 | n17415 ;
  assign n17417 = n71153 & n17416 ;
  assign n17418 = n17307 | n17417 ;
  assign n17420 = n71154 & n17418 ;
  assign n17777 = n17314 | n17420 ;
  assign n18036 = n16711 | n17319 ;
  assign n71162 = ~n18036 ;
  assign n18037 = n17777 & n71162 ;
  assign n18038 = n18035 | n18037 ;
  assign n18039 = n17325 | n18038 ;
  assign n71163 = ~n17327 ;
  assign n18040 = n71163 & n18039 ;
  assign n71164 = ~n17324 ;
  assign n18050 = n71164 & n18040 ;
  assign n17328 = n16710 & n17325 ;
  assign n17315 = n16719 | n17314 ;
  assign n71165 = ~n17315 ;
  assign n17419 = n71165 & n17418 ;
  assign n71166 = ~n17420 ;
  assign n17421 = n17314 & n71166 ;
  assign n17422 = n17419 | n17421 ;
  assign n17423 = n71164 & n17422 ;
  assign n71167 = ~n17322 ;
  assign n17424 = n71167 & n17423 ;
  assign n17425 = n17328 | n17424 ;
  assign n17426 = n70935 & n17425 ;
  assign n17427 = n16718 & n17325 ;
  assign n17308 = n16727 | n17307 ;
  assign n71168 = ~n17308 ;
  assign n17428 = n17304 & n71168 ;
  assign n71169 = ~n17309 ;
  assign n17429 = n17307 & n71169 ;
  assign n17430 = n17428 | n17429 ;
  assign n17431 = n71164 & n17430 ;
  assign n17432 = n71167 & n17431 ;
  assign n17433 = n17427 | n17432 ;
  assign n17434 = n70927 & n17433 ;
  assign n17435 = n16726 & n17325 ;
  assign n17303 = n16735 | n17302 ;
  assign n71170 = ~n17303 ;
  assign n17436 = n71170 & n17414 ;
  assign n71171 = ~n17415 ;
  assign n17437 = n17302 & n71171 ;
  assign n17438 = n17436 | n17437 ;
  assign n17439 = n71164 & n17438 ;
  assign n17440 = n71167 & n17439 ;
  assign n17441 = n17435 | n17440 ;
  assign n17442 = n70609 & n17441 ;
  assign n17443 = n16734 & n17325 ;
  assign n17296 = n16743 | n17295 ;
  assign n71172 = ~n17296 ;
  assign n17444 = n17292 & n71172 ;
  assign n71173 = ~n17297 ;
  assign n17445 = n17295 & n71173 ;
  assign n17446 = n17444 | n17445 ;
  assign n17447 = n71164 & n17446 ;
  assign n17448 = n71167 & n17447 ;
  assign n17449 = n17443 | n17448 ;
  assign n17450 = n70276 & n17449 ;
  assign n17451 = n16742 & n17325 ;
  assign n17291 = n16751 | n17290 ;
  assign n71174 = ~n17291 ;
  assign n17452 = n71174 & n17410 ;
  assign n71175 = ~n17411 ;
  assign n17453 = n17290 & n71175 ;
  assign n17454 = n17452 | n17453 ;
  assign n17455 = n71164 & n17454 ;
  assign n17456 = n71167 & n17455 ;
  assign n17457 = n17451 | n17456 ;
  assign n17458 = n70176 & n17457 ;
  assign n17459 = n16750 & n17325 ;
  assign n17284 = n16759 | n17283 ;
  assign n71176 = ~n17284 ;
  assign n17460 = n17280 & n71176 ;
  assign n71177 = ~n17285 ;
  assign n17461 = n17283 & n71177 ;
  assign n17462 = n17460 | n17461 ;
  assign n17463 = n71164 & n17462 ;
  assign n17464 = n71167 & n17463 ;
  assign n17465 = n17459 | n17464 ;
  assign n17466 = n69857 & n17465 ;
  assign n17467 = n16758 & n17325 ;
  assign n17279 = n16767 | n17278 ;
  assign n71178 = ~n17279 ;
  assign n17468 = n71178 & n17406 ;
  assign n71179 = ~n17407 ;
  assign n17469 = n17278 & n71179 ;
  assign n17470 = n17468 | n17469 ;
  assign n17471 = n71164 & n17470 ;
  assign n17472 = n71167 & n17471 ;
  assign n17473 = n17467 | n17472 ;
  assign n17474 = n69656 & n17473 ;
  assign n17475 = n16766 & n17325 ;
  assign n17272 = n16775 | n17271 ;
  assign n71180 = ~n17272 ;
  assign n17476 = n17268 & n71180 ;
  assign n71181 = ~n17273 ;
  assign n17477 = n17271 & n71181 ;
  assign n17478 = n17476 | n17477 ;
  assign n17479 = n71164 & n17478 ;
  assign n17480 = n71167 & n17479 ;
  assign n17481 = n17475 | n17480 ;
  assign n17482 = n69528 & n17481 ;
  assign n17483 = n16774 & n17325 ;
  assign n17267 = n16783 | n17266 ;
  assign n71182 = ~n17267 ;
  assign n17484 = n71182 & n17402 ;
  assign n71183 = ~n17403 ;
  assign n17485 = n17266 & n71183 ;
  assign n17486 = n17484 | n17485 ;
  assign n17487 = n71164 & n17486 ;
  assign n17488 = n71167 & n17487 ;
  assign n17489 = n17483 | n17488 ;
  assign n17490 = n69261 & n17489 ;
  assign n17491 = n16782 & n17325 ;
  assign n17260 = n16791 | n17259 ;
  assign n71184 = ~n17260 ;
  assign n17492 = n17256 & n71184 ;
  assign n71185 = ~n17261 ;
  assign n17493 = n17259 & n71185 ;
  assign n17494 = n17492 | n17493 ;
  assign n17495 = n71164 & n17494 ;
  assign n17496 = n71167 & n17495 ;
  assign n17497 = n17491 | n17496 ;
  assign n17498 = n69075 & n17497 ;
  assign n17499 = n16790 & n17325 ;
  assign n17255 = n16799 | n17254 ;
  assign n71186 = ~n17255 ;
  assign n17500 = n71186 & n17398 ;
  assign n71187 = ~n17399 ;
  assign n17501 = n17254 & n71187 ;
  assign n17502 = n17500 | n17501 ;
  assign n17503 = n71164 & n17502 ;
  assign n17504 = n71167 & n17503 ;
  assign n17505 = n17499 | n17504 ;
  assign n17506 = n68993 & n17505 ;
  assign n17507 = n16798 & n17325 ;
  assign n17248 = n16807 | n17247 ;
  assign n71188 = ~n17248 ;
  assign n17508 = n17244 & n71188 ;
  assign n71189 = ~n17249 ;
  assign n17509 = n17247 & n71189 ;
  assign n17510 = n17508 | n17509 ;
  assign n17511 = n71164 & n17510 ;
  assign n17512 = n71167 & n17511 ;
  assign n17513 = n17507 | n17512 ;
  assign n17514 = n68716 & n17513 ;
  assign n17515 = n16806 & n17325 ;
  assign n17243 = n16815 | n17242 ;
  assign n71190 = ~n17243 ;
  assign n17516 = n71190 & n17394 ;
  assign n71191 = ~n17395 ;
  assign n17517 = n17242 & n71191 ;
  assign n17518 = n17516 | n17517 ;
  assign n17519 = n71164 & n17518 ;
  assign n17520 = n71167 & n17519 ;
  assign n17521 = n17515 | n17520 ;
  assign n17522 = n68545 & n17521 ;
  assign n17523 = n16814 & n17325 ;
  assign n17236 = n16823 | n17235 ;
  assign n71192 = ~n17236 ;
  assign n17524 = n17232 & n71192 ;
  assign n71193 = ~n17237 ;
  assign n17525 = n17235 & n71193 ;
  assign n17526 = n17524 | n17525 ;
  assign n17527 = n71164 & n17526 ;
  assign n17528 = n71167 & n17527 ;
  assign n17529 = n17523 | n17528 ;
  assign n17530 = n68438 & n17529 ;
  assign n17531 = n16822 & n17325 ;
  assign n17231 = n16831 | n17230 ;
  assign n71194 = ~n17231 ;
  assign n17532 = n71194 & n17390 ;
  assign n71195 = ~n17391 ;
  assign n17533 = n17230 & n71195 ;
  assign n17534 = n17532 | n17533 ;
  assign n17535 = n71164 & n17534 ;
  assign n17536 = n71167 & n17535 ;
  assign n17537 = n17531 | n17536 ;
  assign n17538 = n68214 & n17537 ;
  assign n17539 = n16830 & n17325 ;
  assign n17224 = n16839 | n17223 ;
  assign n71196 = ~n17224 ;
  assign n17540 = n17220 & n71196 ;
  assign n71197 = ~n17225 ;
  assign n17541 = n17223 & n71197 ;
  assign n17542 = n17540 | n17541 ;
  assign n17543 = n71164 & n17542 ;
  assign n17544 = n71167 & n17543 ;
  assign n17545 = n17539 | n17544 ;
  assign n17546 = n68058 & n17545 ;
  assign n17547 = n16838 & n17325 ;
  assign n17219 = n16847 | n17218 ;
  assign n71198 = ~n17219 ;
  assign n17548 = n71198 & n17386 ;
  assign n71199 = ~n17387 ;
  assign n17549 = n17218 & n71199 ;
  assign n17550 = n17548 | n17549 ;
  assign n17551 = n71164 & n17550 ;
  assign n17552 = n71167 & n17551 ;
  assign n17553 = n17547 | n17552 ;
  assign n17554 = n67986 & n17553 ;
  assign n17555 = n16846 & n17325 ;
  assign n17212 = n16855 | n17211 ;
  assign n71200 = ~n17212 ;
  assign n17556 = n17208 & n71200 ;
  assign n71201 = ~n17213 ;
  assign n17557 = n17211 & n71201 ;
  assign n17558 = n17556 | n17557 ;
  assign n17559 = n71164 & n17558 ;
  assign n17560 = n71167 & n17559 ;
  assign n17561 = n17555 | n17560 ;
  assign n17562 = n67763 & n17561 ;
  assign n17563 = n16854 & n17325 ;
  assign n17207 = n16863 | n17206 ;
  assign n71202 = ~n17207 ;
  assign n17564 = n71202 & n17382 ;
  assign n71203 = ~n17383 ;
  assign n17565 = n17206 & n71203 ;
  assign n17566 = n17564 | n17565 ;
  assign n17567 = n71164 & n17566 ;
  assign n17568 = n71167 & n17567 ;
  assign n17569 = n17563 | n17568 ;
  assign n17570 = n67622 & n17569 ;
  assign n17571 = n16862 & n17325 ;
  assign n17200 = n16871 | n17199 ;
  assign n71204 = ~n17200 ;
  assign n17572 = n17196 & n71204 ;
  assign n71205 = ~n17201 ;
  assign n17573 = n17199 & n71205 ;
  assign n17574 = n17572 | n17573 ;
  assign n17575 = n71164 & n17574 ;
  assign n17576 = n71167 & n17575 ;
  assign n17577 = n17571 | n17576 ;
  assign n17578 = n67531 & n17577 ;
  assign n17579 = n16870 & n17325 ;
  assign n17195 = n16879 | n17194 ;
  assign n71206 = ~n17195 ;
  assign n17580 = n71206 & n17378 ;
  assign n71207 = ~n17379 ;
  assign n17581 = n17194 & n71207 ;
  assign n17582 = n17580 | n17581 ;
  assign n17583 = n71164 & n17582 ;
  assign n17584 = n71167 & n17583 ;
  assign n17585 = n17579 | n17584 ;
  assign n17586 = n67348 & n17585 ;
  assign n17587 = n16878 & n17325 ;
  assign n17188 = n16887 | n17187 ;
  assign n71208 = ~n17188 ;
  assign n17588 = n17184 & n71208 ;
  assign n71209 = ~n17189 ;
  assign n17589 = n17187 & n71209 ;
  assign n17590 = n17588 | n17589 ;
  assign n17591 = n71164 & n17590 ;
  assign n17592 = n71167 & n17591 ;
  assign n17593 = n17587 | n17592 ;
  assign n17594 = n67222 & n17593 ;
  assign n17595 = n16886 & n17325 ;
  assign n17183 = n16895 | n17182 ;
  assign n71210 = ~n17183 ;
  assign n17596 = n71210 & n17374 ;
  assign n71211 = ~n17375 ;
  assign n17597 = n17182 & n71211 ;
  assign n17598 = n17596 | n17597 ;
  assign n17599 = n71164 & n17598 ;
  assign n17600 = n71167 & n17599 ;
  assign n17601 = n17595 | n17600 ;
  assign n17602 = n67164 & n17601 ;
  assign n17603 = n16894 & n17325 ;
  assign n17176 = n16903 | n17175 ;
  assign n71212 = ~n17176 ;
  assign n17604 = n17172 & n71212 ;
  assign n71213 = ~n17177 ;
  assign n17605 = n17175 & n71213 ;
  assign n17606 = n17604 | n17605 ;
  assign n17607 = n71164 & n17606 ;
  assign n17608 = n71167 & n17607 ;
  assign n17609 = n17603 | n17608 ;
  assign n17610 = n66979 & n17609 ;
  assign n17611 = n16902 & n17325 ;
  assign n17171 = n16911 | n17170 ;
  assign n71214 = ~n17171 ;
  assign n17612 = n71214 & n17370 ;
  assign n71215 = ~n17371 ;
  assign n17613 = n17170 & n71215 ;
  assign n17614 = n17612 | n17613 ;
  assign n17615 = n71164 & n17614 ;
  assign n17616 = n71167 & n17615 ;
  assign n17617 = n17611 | n17616 ;
  assign n17618 = n66868 & n17617 ;
  assign n17619 = n16910 & n17325 ;
  assign n17164 = n16919 | n17163 ;
  assign n71216 = ~n17164 ;
  assign n17620 = n17160 & n71216 ;
  assign n71217 = ~n17165 ;
  assign n17621 = n17163 & n71217 ;
  assign n17622 = n17620 | n17621 ;
  assign n17623 = n71164 & n17622 ;
  assign n17624 = n71167 & n17623 ;
  assign n17625 = n17619 | n17624 ;
  assign n17626 = n66797 & n17625 ;
  assign n17627 = n16918 & n17325 ;
  assign n17159 = n16927 | n17158 ;
  assign n71218 = ~n17159 ;
  assign n17628 = n71218 & n17366 ;
  assign n71219 = ~n17367 ;
  assign n17629 = n17158 & n71219 ;
  assign n17630 = n17628 | n17629 ;
  assign n17631 = n71164 & n17630 ;
  assign n17632 = n71167 & n17631 ;
  assign n17633 = n17627 | n17632 ;
  assign n17634 = n66654 & n17633 ;
  assign n17635 = n16926 & n17325 ;
  assign n17152 = n16935 | n17151 ;
  assign n71220 = ~n17152 ;
  assign n17636 = n17148 & n71220 ;
  assign n71221 = ~n17153 ;
  assign n17637 = n17151 & n71221 ;
  assign n17638 = n17636 | n17637 ;
  assign n17639 = n71164 & n17638 ;
  assign n17640 = n71167 & n17639 ;
  assign n17641 = n17635 | n17640 ;
  assign n17642 = n66560 & n17641 ;
  assign n17643 = n16934 & n17325 ;
  assign n17147 = n16943 | n17146 ;
  assign n71222 = ~n17147 ;
  assign n17644 = n71222 & n17362 ;
  assign n71223 = ~n17363 ;
  assign n17645 = n17146 & n71223 ;
  assign n17646 = n17644 | n17645 ;
  assign n17647 = n71164 & n17646 ;
  assign n17648 = n71167 & n17647 ;
  assign n17649 = n17643 | n17648 ;
  assign n17650 = n66505 & n17649 ;
  assign n17651 = n16942 & n17325 ;
  assign n17140 = n16951 | n17139 ;
  assign n71224 = ~n17140 ;
  assign n17652 = n17136 & n71224 ;
  assign n71225 = ~n17141 ;
  assign n17653 = n17139 & n71225 ;
  assign n17654 = n17652 | n17653 ;
  assign n17655 = n71164 & n17654 ;
  assign n17656 = n71167 & n17655 ;
  assign n17657 = n17651 | n17656 ;
  assign n17658 = n66379 & n17657 ;
  assign n17659 = n16950 & n17325 ;
  assign n17135 = n16959 | n17134 ;
  assign n71226 = ~n17135 ;
  assign n17660 = n71226 & n17358 ;
  assign n71227 = ~n17359 ;
  assign n17661 = n17134 & n71227 ;
  assign n17662 = n17660 | n17661 ;
  assign n17663 = n71164 & n17662 ;
  assign n17664 = n71167 & n17663 ;
  assign n17665 = n17659 | n17664 ;
  assign n17666 = n66299 & n17665 ;
  assign n17667 = n16958 & n17325 ;
  assign n17128 = n16967 | n17127 ;
  assign n71228 = ~n17128 ;
  assign n17668 = n17124 & n71228 ;
  assign n71229 = ~n17129 ;
  assign n17669 = n17127 & n71229 ;
  assign n17670 = n17668 | n17669 ;
  assign n17671 = n71164 & n17670 ;
  assign n17672 = n71167 & n17671 ;
  assign n17673 = n17667 | n17672 ;
  assign n17674 = n66244 & n17673 ;
  assign n17675 = n16966 & n17325 ;
  assign n17123 = n16975 | n17122 ;
  assign n71230 = ~n17123 ;
  assign n17676 = n71230 & n17354 ;
  assign n71231 = ~n17355 ;
  assign n17677 = n17122 & n71231 ;
  assign n17678 = n17676 | n17677 ;
  assign n17679 = n71164 & n17678 ;
  assign n17680 = n71167 & n17679 ;
  assign n17681 = n17675 | n17680 ;
  assign n17682 = n66145 & n17681 ;
  assign n17683 = n16974 & n17325 ;
  assign n17116 = n16983 | n17115 ;
  assign n71232 = ~n17116 ;
  assign n17684 = n17112 & n71232 ;
  assign n71233 = ~n17117 ;
  assign n17685 = n17115 & n71233 ;
  assign n17686 = n17684 | n17685 ;
  assign n17687 = n71164 & n17686 ;
  assign n17688 = n71167 & n17687 ;
  assign n17689 = n17683 | n17688 ;
  assign n17690 = n66081 & n17689 ;
  assign n17691 = n16982 & n17325 ;
  assign n17111 = n16991 | n17110 ;
  assign n71234 = ~n17111 ;
  assign n17692 = n71234 & n17350 ;
  assign n71235 = ~n17351 ;
  assign n17693 = n17110 & n71235 ;
  assign n17694 = n17692 | n17693 ;
  assign n17695 = n71164 & n17694 ;
  assign n17696 = n71167 & n17695 ;
  assign n17697 = n17691 | n17696 ;
  assign n17698 = n66043 & n17697 ;
  assign n17699 = n16990 & n17325 ;
  assign n17104 = n16999 | n17103 ;
  assign n71236 = ~n17104 ;
  assign n17700 = n17100 & n71236 ;
  assign n71237 = ~n17105 ;
  assign n17701 = n17103 & n71237 ;
  assign n17702 = n17700 | n17701 ;
  assign n17703 = n71164 & n17702 ;
  assign n17704 = n71167 & n17703 ;
  assign n17705 = n17699 | n17704 ;
  assign n17706 = n65960 & n17705 ;
  assign n17707 = n16998 & n17325 ;
  assign n17099 = n17007 | n17098 ;
  assign n71238 = ~n17099 ;
  assign n17708 = n71238 & n17346 ;
  assign n71239 = ~n17347 ;
  assign n17709 = n17098 & n71239 ;
  assign n17710 = n17708 | n17709 ;
  assign n17711 = n71164 & n17710 ;
  assign n17712 = n71167 & n17711 ;
  assign n17713 = n17707 | n17712 ;
  assign n17714 = n65909 & n17713 ;
  assign n17715 = n17006 & n17325 ;
  assign n17092 = n17015 | n17091 ;
  assign n71240 = ~n17092 ;
  assign n17716 = n17088 & n71240 ;
  assign n71241 = ~n17093 ;
  assign n17717 = n17091 & n71241 ;
  assign n17718 = n17716 | n17717 ;
  assign n17719 = n71164 & n17718 ;
  assign n17720 = n71167 & n17719 ;
  assign n17721 = n17715 | n17720 ;
  assign n17722 = n65877 & n17721 ;
  assign n17723 = n17014 & n17325 ;
  assign n17087 = n17023 | n17086 ;
  assign n71242 = ~n17087 ;
  assign n17724 = n71242 & n17342 ;
  assign n71243 = ~n17343 ;
  assign n17725 = n17086 & n71243 ;
  assign n17726 = n17724 | n17725 ;
  assign n17727 = n71164 & n17726 ;
  assign n17728 = n71167 & n17727 ;
  assign n17729 = n17723 | n17728 ;
  assign n17730 = n65820 & n17729 ;
  assign n17731 = n17022 & n17325 ;
  assign n17329 = n17031 | n17080 ;
  assign n71244 = ~n17329 ;
  assign n17732 = n17077 & n71244 ;
  assign n71245 = ~n17081 ;
  assign n17733 = n17080 & n71245 ;
  assign n17734 = n17732 | n17733 ;
  assign n17735 = n71164 & n17734 ;
  assign n17736 = n71167 & n17735 ;
  assign n17737 = n17731 | n17736 ;
  assign n17738 = n65791 & n17737 ;
  assign n17739 = n17030 & n17325 ;
  assign n17740 = n17040 | n17076 ;
  assign n71246 = ~n17740 ;
  assign n17741 = n17338 & n71246 ;
  assign n71247 = ~n17339 ;
  assign n17742 = n17076 & n71247 ;
  assign n17743 = n17741 | n17742 ;
  assign n17744 = n71164 & n17743 ;
  assign n17745 = n71167 & n17744 ;
  assign n17746 = n17739 | n17745 ;
  assign n17747 = n65772 & n17746 ;
  assign n17748 = n17039 & n17325 ;
  assign n17749 = n17048 | n17070 ;
  assign n71248 = ~n17749 ;
  assign n17750 = n17336 & n71248 ;
  assign n71249 = ~n17071 ;
  assign n17751 = n17070 & n71249 ;
  assign n17752 = n17750 | n17751 ;
  assign n17753 = n71164 & n17752 ;
  assign n17754 = n71167 & n17753 ;
  assign n17755 = n17748 | n17754 ;
  assign n17756 = n65746 & n17755 ;
  assign n17757 = n17047 & n17325 ;
  assign n17334 = n17062 | n17066 ;
  assign n71250 = ~n17334 ;
  assign n17758 = n17060 & n71250 ;
  assign n71251 = ~n17335 ;
  assign n17759 = n17066 & n71251 ;
  assign n17760 = n17758 | n17759 ;
  assign n17761 = n71164 & n17760 ;
  assign n17762 = n71167 & n17761 ;
  assign n17763 = n17757 | n17762 ;
  assign n17764 = n65721 & n17763 ;
  assign n17326 = n17061 & n17325 ;
  assign n17332 = n17057 & n17058 ;
  assign n17765 = n71069 & n17332 ;
  assign n17766 = n17324 | n17765 ;
  assign n71252 = ~n17766 ;
  assign n17767 = n17060 & n71252 ;
  assign n17768 = n71167 & n17767 ;
  assign n17769 = n17326 | n17768 ;
  assign n17770 = n65686 & n17769 ;
  assign n71253 = ~x110 ;
  assign n17771 = x64 & n71253 ;
  assign n71254 = ~n288 ;
  assign n17772 = n71254 & n17771 ;
  assign n71255 = ~n271 ;
  assign n17773 = n71255 & n17772 ;
  assign n17774 = n67026 & n17773 ;
  assign n17778 = n71157 & n17777 ;
  assign n17779 = n17319 | n17778 ;
  assign n17780 = n71158 & n17779 ;
  assign n71256 = ~n17780 ;
  assign n17781 = n17774 & n71256 ;
  assign n71257 = ~n17781 ;
  assign n17782 = x18 & n71257 ;
  assign n71258 = ~n65519 ;
  assign n17783 = n71258 & n17058 ;
  assign n71259 = ~n65504 ;
  assign n17784 = n71259 & n17783 ;
  assign n17785 = n67021 & n17784 ;
  assign n17786 = n71167 & n17785 ;
  assign n17787 = n17782 | n17786 ;
  assign n17789 = x65 & n17787 ;
  assign n17775 = n71167 & n17774 ;
  assign n71260 = ~n17775 ;
  assign n17776 = x18 & n71260 ;
  assign n17788 = x65 | n17786 ;
  assign n17790 = n17776 | n17788 ;
  assign n71261 = ~n17789 ;
  assign n17791 = n71261 & n17790 ;
  assign n71262 = ~x17 ;
  assign n17792 = n71262 & x64 ;
  assign n17793 = n17791 | n17792 ;
  assign n17794 = n65670 & n17787 ;
  assign n71263 = ~n17794 ;
  assign n17795 = n17793 & n71263 ;
  assign n71264 = ~n17768 ;
  assign n17796 = x66 & n71264 ;
  assign n71265 = ~n17326 ;
  assign n17797 = n71265 & n17796 ;
  assign n17798 = n17770 | n17797 ;
  assign n17799 = n17795 | n17798 ;
  assign n71266 = ~n17770 ;
  assign n17800 = n71266 & n17799 ;
  assign n71267 = ~n17762 ;
  assign n17801 = x67 & n71267 ;
  assign n71268 = ~n17757 ;
  assign n17802 = n71268 & n17801 ;
  assign n17803 = n17800 | n17802 ;
  assign n71269 = ~n17764 ;
  assign n17804 = n71269 & n17803 ;
  assign n71270 = ~n17754 ;
  assign n17805 = x68 & n71270 ;
  assign n71271 = ~n17748 ;
  assign n17806 = n71271 & n17805 ;
  assign n17807 = n17756 | n17806 ;
  assign n17808 = n17804 | n17807 ;
  assign n71272 = ~n17756 ;
  assign n17809 = n71272 & n17808 ;
  assign n71273 = ~n17745 ;
  assign n17810 = x69 & n71273 ;
  assign n71274 = ~n17739 ;
  assign n17811 = n71274 & n17810 ;
  assign n17812 = n17747 | n17811 ;
  assign n17813 = n17809 | n17812 ;
  assign n71275 = ~n17747 ;
  assign n17814 = n71275 & n17813 ;
  assign n71276 = ~n17736 ;
  assign n17815 = x70 & n71276 ;
  assign n71277 = ~n17731 ;
  assign n17816 = n71277 & n17815 ;
  assign n17817 = n17738 | n17816 ;
  assign n17818 = n17814 | n17817 ;
  assign n71278 = ~n17738 ;
  assign n17819 = n71278 & n17818 ;
  assign n71279 = ~n17728 ;
  assign n17820 = x71 & n71279 ;
  assign n71280 = ~n17723 ;
  assign n17821 = n71280 & n17820 ;
  assign n17822 = n17730 | n17821 ;
  assign n17824 = n17819 | n17822 ;
  assign n71281 = ~n17730 ;
  assign n17825 = n71281 & n17824 ;
  assign n71282 = ~n17720 ;
  assign n17826 = x72 & n71282 ;
  assign n71283 = ~n17715 ;
  assign n17827 = n71283 & n17826 ;
  assign n17828 = n17722 | n17827 ;
  assign n17829 = n17825 | n17828 ;
  assign n71284 = ~n17722 ;
  assign n17830 = n71284 & n17829 ;
  assign n71285 = ~n17712 ;
  assign n17831 = x73 & n71285 ;
  assign n71286 = ~n17707 ;
  assign n17832 = n71286 & n17831 ;
  assign n17833 = n17714 | n17832 ;
  assign n17835 = n17830 | n17833 ;
  assign n71287 = ~n17714 ;
  assign n17836 = n71287 & n17835 ;
  assign n71288 = ~n17704 ;
  assign n17837 = x74 & n71288 ;
  assign n71289 = ~n17699 ;
  assign n17838 = n71289 & n17837 ;
  assign n17839 = n17706 | n17838 ;
  assign n17840 = n17836 | n17839 ;
  assign n71290 = ~n17706 ;
  assign n17841 = n71290 & n17840 ;
  assign n71291 = ~n17696 ;
  assign n17842 = x75 & n71291 ;
  assign n71292 = ~n17691 ;
  assign n17843 = n71292 & n17842 ;
  assign n17844 = n17698 | n17843 ;
  assign n17846 = n17841 | n17844 ;
  assign n71293 = ~n17698 ;
  assign n17847 = n71293 & n17846 ;
  assign n71294 = ~n17688 ;
  assign n17848 = x76 & n71294 ;
  assign n71295 = ~n17683 ;
  assign n17849 = n71295 & n17848 ;
  assign n17850 = n17690 | n17849 ;
  assign n17851 = n17847 | n17850 ;
  assign n71296 = ~n17690 ;
  assign n17852 = n71296 & n17851 ;
  assign n71297 = ~n17680 ;
  assign n17853 = x77 & n71297 ;
  assign n71298 = ~n17675 ;
  assign n17854 = n71298 & n17853 ;
  assign n17855 = n17682 | n17854 ;
  assign n17857 = n17852 | n17855 ;
  assign n71299 = ~n17682 ;
  assign n17858 = n71299 & n17857 ;
  assign n71300 = ~n17672 ;
  assign n17859 = x78 & n71300 ;
  assign n71301 = ~n17667 ;
  assign n17860 = n71301 & n17859 ;
  assign n17861 = n17674 | n17860 ;
  assign n17862 = n17858 | n17861 ;
  assign n71302 = ~n17674 ;
  assign n17863 = n71302 & n17862 ;
  assign n71303 = ~n17664 ;
  assign n17864 = x79 & n71303 ;
  assign n71304 = ~n17659 ;
  assign n17865 = n71304 & n17864 ;
  assign n17866 = n17666 | n17865 ;
  assign n17868 = n17863 | n17866 ;
  assign n71305 = ~n17666 ;
  assign n17869 = n71305 & n17868 ;
  assign n71306 = ~n17656 ;
  assign n17870 = x80 & n71306 ;
  assign n71307 = ~n17651 ;
  assign n17871 = n71307 & n17870 ;
  assign n17872 = n17658 | n17871 ;
  assign n17873 = n17869 | n17872 ;
  assign n71308 = ~n17658 ;
  assign n17874 = n71308 & n17873 ;
  assign n71309 = ~n17648 ;
  assign n17875 = x81 & n71309 ;
  assign n71310 = ~n17643 ;
  assign n17876 = n71310 & n17875 ;
  assign n17877 = n17650 | n17876 ;
  assign n17879 = n17874 | n17877 ;
  assign n71311 = ~n17650 ;
  assign n17880 = n71311 & n17879 ;
  assign n71312 = ~n17640 ;
  assign n17881 = x82 & n71312 ;
  assign n71313 = ~n17635 ;
  assign n17882 = n71313 & n17881 ;
  assign n17883 = n17642 | n17882 ;
  assign n17884 = n17880 | n17883 ;
  assign n71314 = ~n17642 ;
  assign n17885 = n71314 & n17884 ;
  assign n71315 = ~n17632 ;
  assign n17886 = x83 & n71315 ;
  assign n71316 = ~n17627 ;
  assign n17887 = n71316 & n17886 ;
  assign n17888 = n17634 | n17887 ;
  assign n17890 = n17885 | n17888 ;
  assign n71317 = ~n17634 ;
  assign n17891 = n71317 & n17890 ;
  assign n71318 = ~n17624 ;
  assign n17892 = x84 & n71318 ;
  assign n71319 = ~n17619 ;
  assign n17893 = n71319 & n17892 ;
  assign n17894 = n17626 | n17893 ;
  assign n17895 = n17891 | n17894 ;
  assign n71320 = ~n17626 ;
  assign n17896 = n71320 & n17895 ;
  assign n71321 = ~n17616 ;
  assign n17897 = x85 & n71321 ;
  assign n71322 = ~n17611 ;
  assign n17898 = n71322 & n17897 ;
  assign n17899 = n17618 | n17898 ;
  assign n17901 = n17896 | n17899 ;
  assign n71323 = ~n17618 ;
  assign n17902 = n71323 & n17901 ;
  assign n71324 = ~n17608 ;
  assign n17903 = x86 & n71324 ;
  assign n71325 = ~n17603 ;
  assign n17904 = n71325 & n17903 ;
  assign n17905 = n17610 | n17904 ;
  assign n17906 = n17902 | n17905 ;
  assign n71326 = ~n17610 ;
  assign n17907 = n71326 & n17906 ;
  assign n71327 = ~n17600 ;
  assign n17908 = x87 & n71327 ;
  assign n71328 = ~n17595 ;
  assign n17909 = n71328 & n17908 ;
  assign n17910 = n17602 | n17909 ;
  assign n17912 = n17907 | n17910 ;
  assign n71329 = ~n17602 ;
  assign n17913 = n71329 & n17912 ;
  assign n71330 = ~n17592 ;
  assign n17914 = x88 & n71330 ;
  assign n71331 = ~n17587 ;
  assign n17915 = n71331 & n17914 ;
  assign n17916 = n17594 | n17915 ;
  assign n17917 = n17913 | n17916 ;
  assign n71332 = ~n17594 ;
  assign n17918 = n71332 & n17917 ;
  assign n71333 = ~n17584 ;
  assign n17919 = x89 & n71333 ;
  assign n71334 = ~n17579 ;
  assign n17920 = n71334 & n17919 ;
  assign n17921 = n17586 | n17920 ;
  assign n17923 = n17918 | n17921 ;
  assign n71335 = ~n17586 ;
  assign n17924 = n71335 & n17923 ;
  assign n71336 = ~n17576 ;
  assign n17925 = x90 & n71336 ;
  assign n71337 = ~n17571 ;
  assign n17926 = n71337 & n17925 ;
  assign n17927 = n17578 | n17926 ;
  assign n17928 = n17924 | n17927 ;
  assign n71338 = ~n17578 ;
  assign n17929 = n71338 & n17928 ;
  assign n71339 = ~n17568 ;
  assign n17930 = x91 & n71339 ;
  assign n71340 = ~n17563 ;
  assign n17931 = n71340 & n17930 ;
  assign n17932 = n17570 | n17931 ;
  assign n17934 = n17929 | n17932 ;
  assign n71341 = ~n17570 ;
  assign n17935 = n71341 & n17934 ;
  assign n71342 = ~n17560 ;
  assign n17936 = x92 & n71342 ;
  assign n71343 = ~n17555 ;
  assign n17937 = n71343 & n17936 ;
  assign n17938 = n17562 | n17937 ;
  assign n17939 = n17935 | n17938 ;
  assign n71344 = ~n17562 ;
  assign n17940 = n71344 & n17939 ;
  assign n71345 = ~n17552 ;
  assign n17941 = x93 & n71345 ;
  assign n71346 = ~n17547 ;
  assign n17942 = n71346 & n17941 ;
  assign n17943 = n17554 | n17942 ;
  assign n17945 = n17940 | n17943 ;
  assign n71347 = ~n17554 ;
  assign n17946 = n71347 & n17945 ;
  assign n71348 = ~n17544 ;
  assign n17947 = x94 & n71348 ;
  assign n71349 = ~n17539 ;
  assign n17948 = n71349 & n17947 ;
  assign n17949 = n17546 | n17948 ;
  assign n17950 = n17946 | n17949 ;
  assign n71350 = ~n17546 ;
  assign n17951 = n71350 & n17950 ;
  assign n71351 = ~n17536 ;
  assign n17952 = x95 & n71351 ;
  assign n71352 = ~n17531 ;
  assign n17953 = n71352 & n17952 ;
  assign n17954 = n17538 | n17953 ;
  assign n17956 = n17951 | n17954 ;
  assign n71353 = ~n17538 ;
  assign n17957 = n71353 & n17956 ;
  assign n71354 = ~n17528 ;
  assign n17958 = x96 & n71354 ;
  assign n71355 = ~n17523 ;
  assign n17959 = n71355 & n17958 ;
  assign n17960 = n17530 | n17959 ;
  assign n17961 = n17957 | n17960 ;
  assign n71356 = ~n17530 ;
  assign n17962 = n71356 & n17961 ;
  assign n71357 = ~n17520 ;
  assign n17963 = x97 & n71357 ;
  assign n71358 = ~n17515 ;
  assign n17964 = n71358 & n17963 ;
  assign n17965 = n17522 | n17964 ;
  assign n17967 = n17962 | n17965 ;
  assign n71359 = ~n17522 ;
  assign n17968 = n71359 & n17967 ;
  assign n71360 = ~n17512 ;
  assign n17969 = x98 & n71360 ;
  assign n71361 = ~n17507 ;
  assign n17970 = n71361 & n17969 ;
  assign n17971 = n17514 | n17970 ;
  assign n17972 = n17968 | n17971 ;
  assign n71362 = ~n17514 ;
  assign n17973 = n71362 & n17972 ;
  assign n71363 = ~n17504 ;
  assign n17974 = x99 & n71363 ;
  assign n71364 = ~n17499 ;
  assign n17975 = n71364 & n17974 ;
  assign n17976 = n17506 | n17975 ;
  assign n17978 = n17973 | n17976 ;
  assign n71365 = ~n17506 ;
  assign n17979 = n71365 & n17978 ;
  assign n71366 = ~n17496 ;
  assign n17980 = x100 & n71366 ;
  assign n71367 = ~n17491 ;
  assign n17981 = n71367 & n17980 ;
  assign n17982 = n17498 | n17981 ;
  assign n17983 = n17979 | n17982 ;
  assign n71368 = ~n17498 ;
  assign n17984 = n71368 & n17983 ;
  assign n71369 = ~n17488 ;
  assign n17985 = x101 & n71369 ;
  assign n71370 = ~n17483 ;
  assign n17986 = n71370 & n17985 ;
  assign n17987 = n17490 | n17986 ;
  assign n17989 = n17984 | n17987 ;
  assign n71371 = ~n17490 ;
  assign n17990 = n71371 & n17989 ;
  assign n71372 = ~n17480 ;
  assign n17991 = x102 & n71372 ;
  assign n71373 = ~n17475 ;
  assign n17992 = n71373 & n17991 ;
  assign n17993 = n17482 | n17992 ;
  assign n17994 = n17990 | n17993 ;
  assign n71374 = ~n17482 ;
  assign n17995 = n71374 & n17994 ;
  assign n71375 = ~n17472 ;
  assign n17996 = x103 & n71375 ;
  assign n71376 = ~n17467 ;
  assign n17997 = n71376 & n17996 ;
  assign n17998 = n17474 | n17997 ;
  assign n18000 = n17995 | n17998 ;
  assign n71377 = ~n17474 ;
  assign n18001 = n71377 & n18000 ;
  assign n71378 = ~n17464 ;
  assign n18002 = x104 & n71378 ;
  assign n71379 = ~n17459 ;
  assign n18003 = n71379 & n18002 ;
  assign n18004 = n17466 | n18003 ;
  assign n18005 = n18001 | n18004 ;
  assign n71380 = ~n17466 ;
  assign n18006 = n71380 & n18005 ;
  assign n71381 = ~n17456 ;
  assign n18007 = x105 & n71381 ;
  assign n71382 = ~n17451 ;
  assign n18008 = n71382 & n18007 ;
  assign n18009 = n17458 | n18008 ;
  assign n18011 = n18006 | n18009 ;
  assign n71383 = ~n17458 ;
  assign n18012 = n71383 & n18011 ;
  assign n71384 = ~n17448 ;
  assign n18013 = x106 & n71384 ;
  assign n71385 = ~n17443 ;
  assign n18014 = n71385 & n18013 ;
  assign n18015 = n17450 | n18014 ;
  assign n18016 = n18012 | n18015 ;
  assign n71386 = ~n17450 ;
  assign n18017 = n71386 & n18016 ;
  assign n71387 = ~n17440 ;
  assign n18018 = x107 & n71387 ;
  assign n71388 = ~n17435 ;
  assign n18019 = n71388 & n18018 ;
  assign n18020 = n17442 | n18019 ;
  assign n18022 = n18017 | n18020 ;
  assign n71389 = ~n17442 ;
  assign n18023 = n71389 & n18022 ;
  assign n71390 = ~n17432 ;
  assign n18024 = x108 & n71390 ;
  assign n71391 = ~n17427 ;
  assign n18025 = n71391 & n18024 ;
  assign n18026 = n17434 | n18025 ;
  assign n18027 = n18023 | n18026 ;
  assign n71392 = ~n17434 ;
  assign n18028 = n71392 & n18027 ;
  assign n71393 = ~n17424 ;
  assign n18029 = x109 & n71393 ;
  assign n71394 = ~n17328 ;
  assign n18030 = n71394 & n18029 ;
  assign n18031 = n17426 | n18030 ;
  assign n18033 = n18028 | n18031 ;
  assign n71395 = ~n17426 ;
  assign n18034 = n71395 & n18033 ;
  assign n18041 = n71253 & n18040 ;
  assign n147 = ~n17325 ;
  assign n18042 = n147 & n18038 ;
  assign n18043 = n16702 & n17325 ;
  assign n71397 = ~n18043 ;
  assign n18044 = x110 & n71397 ;
  assign n71398 = ~n18042 ;
  assign n18045 = n71398 & n18044 ;
  assign n18046 = n271 | n288 ;
  assign n18047 = n465 | n18046 ;
  assign n18048 = n18045 | n18047 ;
  assign n18049 = n18041 | n18048 ;
  assign n18051 = n18034 | n18049 ;
  assign n71399 = ~n18050 ;
  assign n18052 = n71399 & n18051 ;
  assign n71400 = ~n18028 ;
  assign n18032 = n71400 & n18031 ;
  assign n18055 = n17776 | n17786 ;
  assign n18056 = x65 & n18055 ;
  assign n71401 = ~n18056 ;
  assign n18057 = n17790 & n71401 ;
  assign n18058 = n17792 | n18057 ;
  assign n18059 = n71263 & n18058 ;
  assign n18061 = n17797 | n18059 ;
  assign n18062 = n71266 & n18061 ;
  assign n18063 = n17764 | n17802 ;
  assign n18065 = n18062 | n18063 ;
  assign n18066 = n71269 & n18065 ;
  assign n18068 = n17807 | n18066 ;
  assign n18069 = n71272 & n18068 ;
  assign n18071 = n17812 | n18069 ;
  assign n18072 = n71275 & n18071 ;
  assign n18073 = n17817 | n18072 ;
  assign n18075 = n71278 & n18073 ;
  assign n18076 = n17822 | n18075 ;
  assign n18077 = n71281 & n18076 ;
  assign n18078 = n17828 | n18077 ;
  assign n18080 = n71284 & n18078 ;
  assign n18081 = n17833 | n18080 ;
  assign n18082 = n71287 & n18081 ;
  assign n18083 = n17839 | n18082 ;
  assign n18085 = n71290 & n18083 ;
  assign n18086 = n17844 | n18085 ;
  assign n18087 = n71293 & n18086 ;
  assign n18088 = n17850 | n18087 ;
  assign n18090 = n71296 & n18088 ;
  assign n18091 = n17855 | n18090 ;
  assign n18092 = n71299 & n18091 ;
  assign n18093 = n17861 | n18092 ;
  assign n18095 = n71302 & n18093 ;
  assign n18096 = n17866 | n18095 ;
  assign n18097 = n71305 & n18096 ;
  assign n18098 = n17872 | n18097 ;
  assign n18100 = n71308 & n18098 ;
  assign n18101 = n17877 | n18100 ;
  assign n18102 = n71311 & n18101 ;
  assign n18103 = n17883 | n18102 ;
  assign n18105 = n71314 & n18103 ;
  assign n18106 = n17888 | n18105 ;
  assign n18107 = n71317 & n18106 ;
  assign n18108 = n17894 | n18107 ;
  assign n18110 = n71320 & n18108 ;
  assign n18111 = n17899 | n18110 ;
  assign n18112 = n71323 & n18111 ;
  assign n18113 = n17905 | n18112 ;
  assign n18115 = n71326 & n18113 ;
  assign n18116 = n17910 | n18115 ;
  assign n18117 = n71329 & n18116 ;
  assign n18118 = n17916 | n18117 ;
  assign n18120 = n71332 & n18118 ;
  assign n18121 = n17921 | n18120 ;
  assign n18122 = n71335 & n18121 ;
  assign n18123 = n17927 | n18122 ;
  assign n18125 = n71338 & n18123 ;
  assign n18126 = n17932 | n18125 ;
  assign n18127 = n71341 & n18126 ;
  assign n18128 = n17938 | n18127 ;
  assign n18130 = n71344 & n18128 ;
  assign n18131 = n17943 | n18130 ;
  assign n18132 = n71347 & n18131 ;
  assign n18133 = n17949 | n18132 ;
  assign n18135 = n71350 & n18133 ;
  assign n18136 = n17954 | n18135 ;
  assign n18137 = n71353 & n18136 ;
  assign n18138 = n17960 | n18137 ;
  assign n18140 = n71356 & n18138 ;
  assign n18141 = n17965 | n18140 ;
  assign n18142 = n71359 & n18141 ;
  assign n18143 = n17971 | n18142 ;
  assign n18145 = n71362 & n18143 ;
  assign n18146 = n17976 | n18145 ;
  assign n18147 = n71365 & n18146 ;
  assign n18148 = n17982 | n18147 ;
  assign n18150 = n71368 & n18148 ;
  assign n18151 = n17987 | n18150 ;
  assign n18152 = n71371 & n18151 ;
  assign n18153 = n17993 | n18152 ;
  assign n18155 = n71374 & n18153 ;
  assign n18156 = n17998 | n18155 ;
  assign n18157 = n71377 & n18156 ;
  assign n18158 = n18004 | n18157 ;
  assign n18160 = n71380 & n18158 ;
  assign n18161 = n18009 | n18160 ;
  assign n18162 = n71383 & n18161 ;
  assign n18163 = n18015 | n18162 ;
  assign n18165 = n71386 & n18163 ;
  assign n18166 = n18020 | n18165 ;
  assign n18167 = n71389 & n18166 ;
  assign n18168 = n18026 | n18167 ;
  assign n18170 = n17434 | n18031 ;
  assign n71402 = ~n18170 ;
  assign n18171 = n18168 & n71402 ;
  assign n18172 = n18032 | n18171 ;
  assign n146 = ~n18052 ;
  assign n18173 = n146 & n18172 ;
  assign n18174 = n71392 & n18168 ;
  assign n18175 = n18031 | n18174 ;
  assign n18176 = n71395 & n18175 ;
  assign n18177 = n18049 | n18176 ;
  assign n18178 = n17425 & n71399 ;
  assign n18179 = n18177 & n18178 ;
  assign n18180 = n18173 | n18179 ;
  assign n18181 = n71253 & n18180 ;
  assign n71404 = ~n18179 ;
  assign n18768 = x110 & n71404 ;
  assign n71405 = ~n18173 ;
  assign n18769 = n71405 & n18768 ;
  assign n18770 = n18181 | n18769 ;
  assign n71406 = ~n18167 ;
  assign n18169 = n18026 & n71406 ;
  assign n18182 = n17442 | n18026 ;
  assign n71407 = ~n18182 ;
  assign n18183 = n18022 & n71407 ;
  assign n18184 = n18169 | n18183 ;
  assign n18185 = n146 & n18184 ;
  assign n18186 = n17433 & n71399 ;
  assign n18187 = n18177 & n18186 ;
  assign n18188 = n18185 | n18187 ;
  assign n18189 = n70935 & n18188 ;
  assign n71408 = ~n18017 ;
  assign n18021 = n71408 & n18020 ;
  assign n18190 = n17450 | n18020 ;
  assign n71409 = ~n18190 ;
  assign n18191 = n18163 & n71409 ;
  assign n18192 = n18021 | n18191 ;
  assign n18193 = n146 & n18192 ;
  assign n18194 = n17441 & n71399 ;
  assign n18195 = n18177 & n18194 ;
  assign n18196 = n18193 | n18195 ;
  assign n18197 = n70927 & n18196 ;
  assign n71410 = ~n18195 ;
  assign n18757 = x108 & n71410 ;
  assign n71411 = ~n18193 ;
  assign n18758 = n71411 & n18757 ;
  assign n18759 = n18197 | n18758 ;
  assign n71412 = ~n18162 ;
  assign n18164 = n18015 & n71412 ;
  assign n18198 = n17458 | n18015 ;
  assign n71413 = ~n18198 ;
  assign n18199 = n18011 & n71413 ;
  assign n18200 = n18164 | n18199 ;
  assign n18201 = n146 & n18200 ;
  assign n18202 = n17449 & n71399 ;
  assign n18203 = n18177 & n18202 ;
  assign n18204 = n18201 | n18203 ;
  assign n18205 = n70609 & n18204 ;
  assign n71414 = ~n18006 ;
  assign n18010 = n71414 & n18009 ;
  assign n18206 = n17466 | n18009 ;
  assign n71415 = ~n18206 ;
  assign n18207 = n18158 & n71415 ;
  assign n18208 = n18010 | n18207 ;
  assign n18209 = n146 & n18208 ;
  assign n18210 = n17457 & n71399 ;
  assign n18211 = n18177 & n18210 ;
  assign n18212 = n18209 | n18211 ;
  assign n18213 = n70276 & n18212 ;
  assign n71416 = ~n18211 ;
  assign n18747 = x106 & n71416 ;
  assign n71417 = ~n18209 ;
  assign n18748 = n71417 & n18747 ;
  assign n18749 = n18213 | n18748 ;
  assign n71418 = ~n18157 ;
  assign n18159 = n18004 & n71418 ;
  assign n18214 = n17474 | n18004 ;
  assign n71419 = ~n18214 ;
  assign n18215 = n18000 & n71419 ;
  assign n18216 = n18159 | n18215 ;
  assign n18217 = n146 & n18216 ;
  assign n18218 = n17465 & n71399 ;
  assign n18219 = n18177 & n18218 ;
  assign n18220 = n18217 | n18219 ;
  assign n18221 = n70176 & n18220 ;
  assign n71420 = ~n17995 ;
  assign n17999 = n71420 & n17998 ;
  assign n18222 = n17482 | n17998 ;
  assign n71421 = ~n18222 ;
  assign n18223 = n18153 & n71421 ;
  assign n18224 = n17999 | n18223 ;
  assign n18225 = n146 & n18224 ;
  assign n18226 = n17473 & n71399 ;
  assign n18227 = n18177 & n18226 ;
  assign n18228 = n18225 | n18227 ;
  assign n18229 = n69857 & n18228 ;
  assign n71422 = ~n18227 ;
  assign n18737 = x104 & n71422 ;
  assign n71423 = ~n18225 ;
  assign n18738 = n71423 & n18737 ;
  assign n18739 = n18229 | n18738 ;
  assign n71424 = ~n18152 ;
  assign n18154 = n17993 & n71424 ;
  assign n18230 = n17490 | n17993 ;
  assign n71425 = ~n18230 ;
  assign n18231 = n17989 & n71425 ;
  assign n18232 = n18154 | n18231 ;
  assign n18233 = n146 & n18232 ;
  assign n18234 = n17481 & n71399 ;
  assign n18235 = n18177 & n18234 ;
  assign n18236 = n18233 | n18235 ;
  assign n18237 = n69656 & n18236 ;
  assign n71426 = ~n17984 ;
  assign n17988 = n71426 & n17987 ;
  assign n18238 = n17498 | n17987 ;
  assign n71427 = ~n18238 ;
  assign n18239 = n18148 & n71427 ;
  assign n18240 = n17988 | n18239 ;
  assign n18241 = n146 & n18240 ;
  assign n18242 = n17489 & n71399 ;
  assign n18243 = n18177 & n18242 ;
  assign n18244 = n18241 | n18243 ;
  assign n18245 = n69528 & n18244 ;
  assign n71428 = ~n18243 ;
  assign n18727 = x102 & n71428 ;
  assign n71429 = ~n18241 ;
  assign n18728 = n71429 & n18727 ;
  assign n18729 = n18245 | n18728 ;
  assign n71430 = ~n18147 ;
  assign n18149 = n17982 & n71430 ;
  assign n18246 = n17506 | n17982 ;
  assign n71431 = ~n18246 ;
  assign n18247 = n17978 & n71431 ;
  assign n18248 = n18149 | n18247 ;
  assign n18249 = n146 & n18248 ;
  assign n18250 = n17497 & n71399 ;
  assign n18251 = n18177 & n18250 ;
  assign n18252 = n18249 | n18251 ;
  assign n18253 = n69261 & n18252 ;
  assign n71432 = ~n17973 ;
  assign n17977 = n71432 & n17976 ;
  assign n18254 = n17514 | n17976 ;
  assign n71433 = ~n18254 ;
  assign n18255 = n18143 & n71433 ;
  assign n18256 = n17977 | n18255 ;
  assign n18257 = n146 & n18256 ;
  assign n18258 = n17505 & n71399 ;
  assign n18259 = n18177 & n18258 ;
  assign n18260 = n18257 | n18259 ;
  assign n18261 = n69075 & n18260 ;
  assign n71434 = ~n18259 ;
  assign n18717 = x100 & n71434 ;
  assign n71435 = ~n18257 ;
  assign n18718 = n71435 & n18717 ;
  assign n18719 = n18261 | n18718 ;
  assign n71436 = ~n18142 ;
  assign n18144 = n17971 & n71436 ;
  assign n18262 = n17522 | n17971 ;
  assign n71437 = ~n18262 ;
  assign n18263 = n17967 & n71437 ;
  assign n18264 = n18144 | n18263 ;
  assign n18265 = n146 & n18264 ;
  assign n18266 = n17513 & n71399 ;
  assign n18267 = n18177 & n18266 ;
  assign n18268 = n18265 | n18267 ;
  assign n18269 = n68993 & n18268 ;
  assign n71438 = ~n17962 ;
  assign n17966 = n71438 & n17965 ;
  assign n18270 = n17530 | n17965 ;
  assign n71439 = ~n18270 ;
  assign n18271 = n18138 & n71439 ;
  assign n18272 = n17966 | n18271 ;
  assign n18273 = n146 & n18272 ;
  assign n18274 = n17521 & n71399 ;
  assign n18275 = n18177 & n18274 ;
  assign n18276 = n18273 | n18275 ;
  assign n18277 = n68716 & n18276 ;
  assign n71440 = ~n18275 ;
  assign n18707 = x98 & n71440 ;
  assign n71441 = ~n18273 ;
  assign n18708 = n71441 & n18707 ;
  assign n18709 = n18277 | n18708 ;
  assign n71442 = ~n18137 ;
  assign n18139 = n17960 & n71442 ;
  assign n18278 = n17538 | n17960 ;
  assign n71443 = ~n18278 ;
  assign n18279 = n17956 & n71443 ;
  assign n18280 = n18139 | n18279 ;
  assign n18281 = n146 & n18280 ;
  assign n18282 = n17529 & n71399 ;
  assign n18283 = n18177 & n18282 ;
  assign n18284 = n18281 | n18283 ;
  assign n18285 = n68545 & n18284 ;
  assign n71444 = ~n17951 ;
  assign n17955 = n71444 & n17954 ;
  assign n18286 = n17546 | n17954 ;
  assign n71445 = ~n18286 ;
  assign n18287 = n18133 & n71445 ;
  assign n18288 = n17955 | n18287 ;
  assign n18289 = n146 & n18288 ;
  assign n18290 = n17537 & n71399 ;
  assign n18291 = n18177 & n18290 ;
  assign n18292 = n18289 | n18291 ;
  assign n18293 = n68438 & n18292 ;
  assign n71446 = ~n18291 ;
  assign n18697 = x96 & n71446 ;
  assign n71447 = ~n18289 ;
  assign n18698 = n71447 & n18697 ;
  assign n18699 = n18293 | n18698 ;
  assign n71448 = ~n18132 ;
  assign n18134 = n17949 & n71448 ;
  assign n18294 = n17554 | n17949 ;
  assign n71449 = ~n18294 ;
  assign n18295 = n17945 & n71449 ;
  assign n18296 = n18134 | n18295 ;
  assign n18297 = n146 & n18296 ;
  assign n18298 = n17545 & n71399 ;
  assign n18299 = n18177 & n18298 ;
  assign n18300 = n18297 | n18299 ;
  assign n18301 = n68214 & n18300 ;
  assign n71450 = ~n17940 ;
  assign n17944 = n71450 & n17943 ;
  assign n18302 = n17562 | n17943 ;
  assign n71451 = ~n18302 ;
  assign n18303 = n18128 & n71451 ;
  assign n18304 = n17944 | n18303 ;
  assign n18305 = n146 & n18304 ;
  assign n18306 = n17553 & n71399 ;
  assign n18307 = n18177 & n18306 ;
  assign n18308 = n18305 | n18307 ;
  assign n18309 = n68058 & n18308 ;
  assign n71452 = ~n18307 ;
  assign n18687 = x94 & n71452 ;
  assign n71453 = ~n18305 ;
  assign n18688 = n71453 & n18687 ;
  assign n18689 = n18309 | n18688 ;
  assign n71454 = ~n18127 ;
  assign n18129 = n17938 & n71454 ;
  assign n18310 = n17570 | n17938 ;
  assign n71455 = ~n18310 ;
  assign n18311 = n17934 & n71455 ;
  assign n18312 = n18129 | n18311 ;
  assign n18313 = n146 & n18312 ;
  assign n18314 = n17561 & n71399 ;
  assign n18315 = n18177 & n18314 ;
  assign n18316 = n18313 | n18315 ;
  assign n18317 = n67986 & n18316 ;
  assign n71456 = ~n17929 ;
  assign n17933 = n71456 & n17932 ;
  assign n18318 = n17578 | n17932 ;
  assign n71457 = ~n18318 ;
  assign n18319 = n18123 & n71457 ;
  assign n18320 = n17933 | n18319 ;
  assign n18321 = n146 & n18320 ;
  assign n18322 = n17569 & n71399 ;
  assign n18323 = n18177 & n18322 ;
  assign n18324 = n18321 | n18323 ;
  assign n18325 = n67763 & n18324 ;
  assign n71458 = ~n18323 ;
  assign n18677 = x92 & n71458 ;
  assign n71459 = ~n18321 ;
  assign n18678 = n71459 & n18677 ;
  assign n18679 = n18325 | n18678 ;
  assign n71460 = ~n18122 ;
  assign n18124 = n17927 & n71460 ;
  assign n18326 = n17586 | n17927 ;
  assign n71461 = ~n18326 ;
  assign n18327 = n17923 & n71461 ;
  assign n18328 = n18124 | n18327 ;
  assign n18329 = n146 & n18328 ;
  assign n18330 = n17577 & n71399 ;
  assign n18331 = n18177 & n18330 ;
  assign n18332 = n18329 | n18331 ;
  assign n18333 = n67622 & n18332 ;
  assign n71462 = ~n17918 ;
  assign n17922 = n71462 & n17921 ;
  assign n18334 = n17594 | n17921 ;
  assign n71463 = ~n18334 ;
  assign n18335 = n18118 & n71463 ;
  assign n18336 = n17922 | n18335 ;
  assign n18337 = n146 & n18336 ;
  assign n18338 = n17585 & n71399 ;
  assign n18339 = n18177 & n18338 ;
  assign n18340 = n18337 | n18339 ;
  assign n18341 = n67531 & n18340 ;
  assign n71464 = ~n18339 ;
  assign n18667 = x90 & n71464 ;
  assign n71465 = ~n18337 ;
  assign n18668 = n71465 & n18667 ;
  assign n18669 = n18341 | n18668 ;
  assign n71466 = ~n18117 ;
  assign n18119 = n17916 & n71466 ;
  assign n18342 = n17602 | n17916 ;
  assign n71467 = ~n18342 ;
  assign n18343 = n17912 & n71467 ;
  assign n18344 = n18119 | n18343 ;
  assign n18345 = n146 & n18344 ;
  assign n18346 = n17593 & n71399 ;
  assign n18347 = n18177 & n18346 ;
  assign n18348 = n18345 | n18347 ;
  assign n18349 = n67348 & n18348 ;
  assign n71468 = ~n17907 ;
  assign n17911 = n71468 & n17910 ;
  assign n18350 = n17610 | n17910 ;
  assign n71469 = ~n18350 ;
  assign n18351 = n18113 & n71469 ;
  assign n18352 = n17911 | n18351 ;
  assign n18353 = n146 & n18352 ;
  assign n18354 = n17601 & n71399 ;
  assign n18355 = n18177 & n18354 ;
  assign n18356 = n18353 | n18355 ;
  assign n18357 = n67222 & n18356 ;
  assign n71470 = ~n18355 ;
  assign n18657 = x88 & n71470 ;
  assign n71471 = ~n18353 ;
  assign n18658 = n71471 & n18657 ;
  assign n18659 = n18357 | n18658 ;
  assign n71472 = ~n18112 ;
  assign n18114 = n17905 & n71472 ;
  assign n18358 = n17618 | n17905 ;
  assign n71473 = ~n18358 ;
  assign n18359 = n17901 & n71473 ;
  assign n18360 = n18114 | n18359 ;
  assign n18361 = n146 & n18360 ;
  assign n18362 = n17609 & n71399 ;
  assign n18363 = n18177 & n18362 ;
  assign n18364 = n18361 | n18363 ;
  assign n18365 = n67164 & n18364 ;
  assign n71474 = ~n17896 ;
  assign n17900 = n71474 & n17899 ;
  assign n18366 = n17626 | n17899 ;
  assign n71475 = ~n18366 ;
  assign n18367 = n18108 & n71475 ;
  assign n18368 = n17900 | n18367 ;
  assign n18369 = n146 & n18368 ;
  assign n18370 = n17617 & n71399 ;
  assign n18371 = n18177 & n18370 ;
  assign n18372 = n18369 | n18371 ;
  assign n18373 = n66979 & n18372 ;
  assign n71476 = ~n18371 ;
  assign n18647 = x86 & n71476 ;
  assign n71477 = ~n18369 ;
  assign n18648 = n71477 & n18647 ;
  assign n18649 = n18373 | n18648 ;
  assign n71478 = ~n18107 ;
  assign n18109 = n17894 & n71478 ;
  assign n18374 = n17634 | n17894 ;
  assign n71479 = ~n18374 ;
  assign n18375 = n17890 & n71479 ;
  assign n18376 = n18109 | n18375 ;
  assign n18377 = n146 & n18376 ;
  assign n18378 = n17625 & n71399 ;
  assign n18379 = n18177 & n18378 ;
  assign n18380 = n18377 | n18379 ;
  assign n18381 = n66868 & n18380 ;
  assign n71480 = ~n17885 ;
  assign n17889 = n71480 & n17888 ;
  assign n18382 = n17642 | n17888 ;
  assign n71481 = ~n18382 ;
  assign n18383 = n18103 & n71481 ;
  assign n18384 = n17889 | n18383 ;
  assign n18385 = n146 & n18384 ;
  assign n18386 = n17633 & n71399 ;
  assign n18387 = n18177 & n18386 ;
  assign n18388 = n18385 | n18387 ;
  assign n18389 = n66797 & n18388 ;
  assign n71482 = ~n18387 ;
  assign n18636 = x84 & n71482 ;
  assign n71483 = ~n18385 ;
  assign n18637 = n71483 & n18636 ;
  assign n18638 = n18389 | n18637 ;
  assign n71484 = ~n18102 ;
  assign n18104 = n17883 & n71484 ;
  assign n18390 = n17650 | n17883 ;
  assign n71485 = ~n18390 ;
  assign n18391 = n17879 & n71485 ;
  assign n18392 = n18104 | n18391 ;
  assign n18393 = n146 & n18392 ;
  assign n18394 = n17641 & n71399 ;
  assign n18395 = n18177 & n18394 ;
  assign n18396 = n18393 | n18395 ;
  assign n18397 = n66654 & n18396 ;
  assign n71486 = ~n17874 ;
  assign n17878 = n71486 & n17877 ;
  assign n18398 = n17658 | n17877 ;
  assign n71487 = ~n18398 ;
  assign n18399 = n18098 & n71487 ;
  assign n18400 = n17878 | n18399 ;
  assign n18401 = n146 & n18400 ;
  assign n18402 = n17649 & n71399 ;
  assign n18403 = n18177 & n18402 ;
  assign n18404 = n18401 | n18403 ;
  assign n18405 = n66560 & n18404 ;
  assign n71488 = ~n18403 ;
  assign n18626 = x82 & n71488 ;
  assign n71489 = ~n18401 ;
  assign n18627 = n71489 & n18626 ;
  assign n18628 = n18405 | n18627 ;
  assign n71490 = ~n18097 ;
  assign n18099 = n17872 & n71490 ;
  assign n18406 = n17666 | n17872 ;
  assign n71491 = ~n18406 ;
  assign n18407 = n17868 & n71491 ;
  assign n18408 = n18099 | n18407 ;
  assign n18409 = n146 & n18408 ;
  assign n18410 = n17657 & n71399 ;
  assign n18411 = n18177 & n18410 ;
  assign n18412 = n18409 | n18411 ;
  assign n18413 = n66505 & n18412 ;
  assign n71492 = ~n17863 ;
  assign n17867 = n71492 & n17866 ;
  assign n18414 = n17674 | n17866 ;
  assign n71493 = ~n18414 ;
  assign n18415 = n18093 & n71493 ;
  assign n18416 = n17867 | n18415 ;
  assign n18417 = n146 & n18416 ;
  assign n18418 = n17665 & n71399 ;
  assign n18419 = n18177 & n18418 ;
  assign n18420 = n18417 | n18419 ;
  assign n18421 = n66379 & n18420 ;
  assign n71494 = ~n18419 ;
  assign n18616 = x80 & n71494 ;
  assign n71495 = ~n18417 ;
  assign n18617 = n71495 & n18616 ;
  assign n18618 = n18421 | n18617 ;
  assign n71496 = ~n18092 ;
  assign n18094 = n17861 & n71496 ;
  assign n18422 = n17682 | n17861 ;
  assign n71497 = ~n18422 ;
  assign n18423 = n17857 & n71497 ;
  assign n18424 = n18094 | n18423 ;
  assign n18425 = n146 & n18424 ;
  assign n18426 = n17673 & n71399 ;
  assign n18427 = n18177 & n18426 ;
  assign n18428 = n18425 | n18427 ;
  assign n18429 = n66299 & n18428 ;
  assign n71498 = ~n17852 ;
  assign n17856 = n71498 & n17855 ;
  assign n18430 = n17690 | n17855 ;
  assign n71499 = ~n18430 ;
  assign n18431 = n18088 & n71499 ;
  assign n18432 = n17856 | n18431 ;
  assign n18433 = n146 & n18432 ;
  assign n18434 = n17681 & n71399 ;
  assign n18435 = n18177 & n18434 ;
  assign n18436 = n18433 | n18435 ;
  assign n18437 = n66244 & n18436 ;
  assign n71500 = ~n18435 ;
  assign n18606 = x78 & n71500 ;
  assign n71501 = ~n18433 ;
  assign n18607 = n71501 & n18606 ;
  assign n18608 = n18437 | n18607 ;
  assign n71502 = ~n18087 ;
  assign n18089 = n17850 & n71502 ;
  assign n18438 = n17698 | n17850 ;
  assign n71503 = ~n18438 ;
  assign n18439 = n17846 & n71503 ;
  assign n18440 = n18089 | n18439 ;
  assign n18441 = n146 & n18440 ;
  assign n18442 = n17689 & n71399 ;
  assign n18443 = n18177 & n18442 ;
  assign n18444 = n18441 | n18443 ;
  assign n18445 = n66145 & n18444 ;
  assign n71504 = ~n17841 ;
  assign n17845 = n71504 & n17844 ;
  assign n18446 = n17706 | n17844 ;
  assign n71505 = ~n18446 ;
  assign n18447 = n18083 & n71505 ;
  assign n18448 = n17845 | n18447 ;
  assign n18449 = n146 & n18448 ;
  assign n18450 = n17697 & n71399 ;
  assign n18451 = n18177 & n18450 ;
  assign n18452 = n18449 | n18451 ;
  assign n18453 = n66081 & n18452 ;
  assign n71506 = ~n18451 ;
  assign n18596 = x76 & n71506 ;
  assign n71507 = ~n18449 ;
  assign n18597 = n71507 & n18596 ;
  assign n18598 = n18453 | n18597 ;
  assign n71508 = ~n18082 ;
  assign n18084 = n17839 & n71508 ;
  assign n18454 = n17714 | n17839 ;
  assign n71509 = ~n18454 ;
  assign n18455 = n17835 & n71509 ;
  assign n18456 = n18084 | n18455 ;
  assign n18457 = n146 & n18456 ;
  assign n18458 = n17705 & n71399 ;
  assign n18459 = n18177 & n18458 ;
  assign n18460 = n18457 | n18459 ;
  assign n18461 = n66043 & n18460 ;
  assign n71510 = ~n17830 ;
  assign n17834 = n71510 & n17833 ;
  assign n18462 = n17722 | n17833 ;
  assign n71511 = ~n18462 ;
  assign n18463 = n18078 & n71511 ;
  assign n18464 = n17834 | n18463 ;
  assign n18465 = n146 & n18464 ;
  assign n18466 = n17713 & n71399 ;
  assign n18467 = n18177 & n18466 ;
  assign n18468 = n18465 | n18467 ;
  assign n18469 = n65960 & n18468 ;
  assign n71512 = ~n18467 ;
  assign n18586 = x74 & n71512 ;
  assign n71513 = ~n18465 ;
  assign n18587 = n71513 & n18586 ;
  assign n18588 = n18469 | n18587 ;
  assign n71514 = ~n18077 ;
  assign n18079 = n17828 & n71514 ;
  assign n18470 = n17730 | n17828 ;
  assign n71515 = ~n18470 ;
  assign n18471 = n17824 & n71515 ;
  assign n18472 = n18079 | n18471 ;
  assign n18473 = n146 & n18472 ;
  assign n18474 = n17721 & n71399 ;
  assign n18475 = n18177 & n18474 ;
  assign n18476 = n18473 | n18475 ;
  assign n18477 = n65909 & n18476 ;
  assign n71516 = ~n17819 ;
  assign n17823 = n71516 & n17822 ;
  assign n18478 = n17738 | n17822 ;
  assign n71517 = ~n18478 ;
  assign n18479 = n18073 & n71517 ;
  assign n18480 = n17823 | n18479 ;
  assign n18481 = n146 & n18480 ;
  assign n18482 = n17729 & n71399 ;
  assign n18483 = n18177 & n18482 ;
  assign n18484 = n18481 | n18483 ;
  assign n18485 = n65877 & n18484 ;
  assign n71518 = ~n18483 ;
  assign n18576 = x72 & n71518 ;
  assign n71519 = ~n18481 ;
  assign n18577 = n71519 & n18576 ;
  assign n18578 = n18485 | n18577 ;
  assign n71520 = ~n18072 ;
  assign n18074 = n17817 & n71520 ;
  assign n18486 = n17747 | n17817 ;
  assign n71521 = ~n18486 ;
  assign n18487 = n17813 & n71521 ;
  assign n18488 = n18074 | n18487 ;
  assign n18489 = n146 & n18488 ;
  assign n18490 = n17737 & n71399 ;
  assign n18491 = n18177 & n18490 ;
  assign n18492 = n18489 | n18491 ;
  assign n18493 = n65820 & n18492 ;
  assign n71522 = ~n17809 ;
  assign n18070 = n71522 & n17812 ;
  assign n18494 = n17756 | n17812 ;
  assign n71523 = ~n18494 ;
  assign n18495 = n18068 & n71523 ;
  assign n18496 = n18070 | n18495 ;
  assign n18497 = n146 & n18496 ;
  assign n18498 = n17746 & n71399 ;
  assign n18499 = n18177 & n18498 ;
  assign n18500 = n18497 | n18499 ;
  assign n18501 = n65791 & n18500 ;
  assign n71524 = ~n18499 ;
  assign n18566 = x70 & n71524 ;
  assign n71525 = ~n18497 ;
  assign n18567 = n71525 & n18566 ;
  assign n18568 = n18501 | n18567 ;
  assign n71526 = ~n18066 ;
  assign n18067 = n17807 & n71526 ;
  assign n18502 = n17800 | n18063 ;
  assign n18503 = n17764 | n17807 ;
  assign n71527 = ~n18503 ;
  assign n18504 = n18502 & n71527 ;
  assign n18505 = n18067 | n18504 ;
  assign n18506 = n146 & n18505 ;
  assign n18507 = n17755 & n71399 ;
  assign n18508 = n18177 & n18507 ;
  assign n18509 = n18506 | n18508 ;
  assign n18510 = n65772 & n18509 ;
  assign n71528 = ~n17800 ;
  assign n18064 = n71528 & n18063 ;
  assign n18511 = n17770 | n18063 ;
  assign n71529 = ~n18511 ;
  assign n18512 = n17799 & n71529 ;
  assign n18513 = n18064 | n18512 ;
  assign n18514 = n146 & n18513 ;
  assign n18515 = n17763 & n71399 ;
  assign n18516 = n18177 & n18515 ;
  assign n18517 = n18514 | n18516 ;
  assign n18518 = n65746 & n18517 ;
  assign n71530 = ~n18516 ;
  assign n18556 = x68 & n71530 ;
  assign n71531 = ~n18514 ;
  assign n18557 = n71531 & n18556 ;
  assign n18558 = n18518 | n18557 ;
  assign n71532 = ~n18059 ;
  assign n18060 = n17798 & n71532 ;
  assign n18519 = n17794 | n17798 ;
  assign n71533 = ~n18519 ;
  assign n18520 = n17793 & n71533 ;
  assign n18521 = n18060 | n18520 ;
  assign n18522 = n146 & n18521 ;
  assign n18523 = n17769 & n71399 ;
  assign n18524 = n18177 & n18523 ;
  assign n18525 = n18522 | n18524 ;
  assign n18526 = n65721 & n18525 ;
  assign n18527 = n17790 & n17792 ;
  assign n18528 = n71261 & n18527 ;
  assign n71534 = ~n18528 ;
  assign n18529 = n18058 & n71534 ;
  assign n18530 = n146 & n18529 ;
  assign n18531 = n71399 & n18055 ;
  assign n18532 = n18177 & n18531 ;
  assign n18533 = n18530 | n18532 ;
  assign n18534 = n65686 & n18533 ;
  assign n71535 = ~n18532 ;
  assign n18546 = x66 & n71535 ;
  assign n71536 = ~n18530 ;
  assign n18547 = n71536 & n18546 ;
  assign n18548 = n18534 | n18547 ;
  assign n18054 = n17792 & n146 ;
  assign n18053 = x64 & n146 ;
  assign n71537 = ~n18053 ;
  assign n18535 = x17 & n71537 ;
  assign n18536 = n18054 | n18535 ;
  assign n18537 = x65 & n18536 ;
  assign n18538 = n71399 & n18177 ;
  assign n71538 = ~n18538 ;
  assign n18539 = n17792 & n71538 ;
  assign n18540 = x65 | n18539 ;
  assign n18541 = n18535 | n18540 ;
  assign n71539 = ~n18537 ;
  assign n18542 = n71539 & n18541 ;
  assign n71540 = ~x16 ;
  assign n18543 = n71540 & x64 ;
  assign n18544 = n18542 | n18543 ;
  assign n18545 = n65670 & n18536 ;
  assign n71541 = ~n18545 ;
  assign n18549 = n18544 & n71541 ;
  assign n18550 = n18548 | n18549 ;
  assign n71542 = ~n18534 ;
  assign n18551 = n71542 & n18550 ;
  assign n71543 = ~n18524 ;
  assign n18552 = x67 & n71543 ;
  assign n71544 = ~n18522 ;
  assign n18553 = n71544 & n18552 ;
  assign n18554 = n18526 | n18553 ;
  assign n18555 = n18551 | n18554 ;
  assign n71545 = ~n18526 ;
  assign n18559 = n71545 & n18555 ;
  assign n18560 = n18558 | n18559 ;
  assign n71546 = ~n18518 ;
  assign n18561 = n71546 & n18560 ;
  assign n71547 = ~n18508 ;
  assign n18562 = x69 & n71547 ;
  assign n71548 = ~n18506 ;
  assign n18563 = n71548 & n18562 ;
  assign n18564 = n18510 | n18563 ;
  assign n18565 = n18561 | n18564 ;
  assign n71549 = ~n18510 ;
  assign n18569 = n71549 & n18565 ;
  assign n18570 = n18568 | n18569 ;
  assign n71550 = ~n18501 ;
  assign n18571 = n71550 & n18570 ;
  assign n71551 = ~n18491 ;
  assign n18572 = x71 & n71551 ;
  assign n71552 = ~n18489 ;
  assign n18573 = n71552 & n18572 ;
  assign n18574 = n18493 | n18573 ;
  assign n18575 = n18571 | n18574 ;
  assign n71553 = ~n18493 ;
  assign n18579 = n71553 & n18575 ;
  assign n18580 = n18578 | n18579 ;
  assign n71554 = ~n18485 ;
  assign n18581 = n71554 & n18580 ;
  assign n71555 = ~n18475 ;
  assign n18582 = x73 & n71555 ;
  assign n71556 = ~n18473 ;
  assign n18583 = n71556 & n18582 ;
  assign n18584 = n18477 | n18583 ;
  assign n18585 = n18581 | n18584 ;
  assign n71557 = ~n18477 ;
  assign n18589 = n71557 & n18585 ;
  assign n18590 = n18588 | n18589 ;
  assign n71558 = ~n18469 ;
  assign n18591 = n71558 & n18590 ;
  assign n71559 = ~n18459 ;
  assign n18592 = x75 & n71559 ;
  assign n71560 = ~n18457 ;
  assign n18593 = n71560 & n18592 ;
  assign n18594 = n18461 | n18593 ;
  assign n18595 = n18591 | n18594 ;
  assign n71561 = ~n18461 ;
  assign n18599 = n71561 & n18595 ;
  assign n18600 = n18598 | n18599 ;
  assign n71562 = ~n18453 ;
  assign n18601 = n71562 & n18600 ;
  assign n71563 = ~n18443 ;
  assign n18602 = x77 & n71563 ;
  assign n71564 = ~n18441 ;
  assign n18603 = n71564 & n18602 ;
  assign n18604 = n18445 | n18603 ;
  assign n18605 = n18601 | n18604 ;
  assign n71565 = ~n18445 ;
  assign n18609 = n71565 & n18605 ;
  assign n18610 = n18608 | n18609 ;
  assign n71566 = ~n18437 ;
  assign n18611 = n71566 & n18610 ;
  assign n71567 = ~n18427 ;
  assign n18612 = x79 & n71567 ;
  assign n71568 = ~n18425 ;
  assign n18613 = n71568 & n18612 ;
  assign n18614 = n18429 | n18613 ;
  assign n18615 = n18611 | n18614 ;
  assign n71569 = ~n18429 ;
  assign n18619 = n71569 & n18615 ;
  assign n18620 = n18618 | n18619 ;
  assign n71570 = ~n18421 ;
  assign n18621 = n71570 & n18620 ;
  assign n71571 = ~n18411 ;
  assign n18622 = x81 & n71571 ;
  assign n71572 = ~n18409 ;
  assign n18623 = n71572 & n18622 ;
  assign n18624 = n18413 | n18623 ;
  assign n18625 = n18621 | n18624 ;
  assign n71573 = ~n18413 ;
  assign n18629 = n71573 & n18625 ;
  assign n18630 = n18628 | n18629 ;
  assign n71574 = ~n18405 ;
  assign n18631 = n71574 & n18630 ;
  assign n71575 = ~n18395 ;
  assign n18632 = x83 & n71575 ;
  assign n71576 = ~n18393 ;
  assign n18633 = n71576 & n18632 ;
  assign n18634 = n18397 | n18633 ;
  assign n18635 = n18631 | n18634 ;
  assign n71577 = ~n18397 ;
  assign n18639 = n71577 & n18635 ;
  assign n18640 = n18638 | n18639 ;
  assign n71578 = ~n18389 ;
  assign n18641 = n71578 & n18640 ;
  assign n71579 = ~n18379 ;
  assign n18642 = x85 & n71579 ;
  assign n71580 = ~n18377 ;
  assign n18643 = n71580 & n18642 ;
  assign n18644 = n18381 | n18643 ;
  assign n18646 = n18641 | n18644 ;
  assign n71581 = ~n18381 ;
  assign n18650 = n71581 & n18646 ;
  assign n18651 = n18649 | n18650 ;
  assign n71582 = ~n18373 ;
  assign n18652 = n71582 & n18651 ;
  assign n71583 = ~n18363 ;
  assign n18653 = x87 & n71583 ;
  assign n71584 = ~n18361 ;
  assign n18654 = n71584 & n18653 ;
  assign n18655 = n18365 | n18654 ;
  assign n18656 = n18652 | n18655 ;
  assign n71585 = ~n18365 ;
  assign n18660 = n71585 & n18656 ;
  assign n18661 = n18659 | n18660 ;
  assign n71586 = ~n18357 ;
  assign n18662 = n71586 & n18661 ;
  assign n71587 = ~n18347 ;
  assign n18663 = x89 & n71587 ;
  assign n71588 = ~n18345 ;
  assign n18664 = n71588 & n18663 ;
  assign n18665 = n18349 | n18664 ;
  assign n18666 = n18662 | n18665 ;
  assign n71589 = ~n18349 ;
  assign n18670 = n71589 & n18666 ;
  assign n18671 = n18669 | n18670 ;
  assign n71590 = ~n18341 ;
  assign n18672 = n71590 & n18671 ;
  assign n71591 = ~n18331 ;
  assign n18673 = x91 & n71591 ;
  assign n71592 = ~n18329 ;
  assign n18674 = n71592 & n18673 ;
  assign n18675 = n18333 | n18674 ;
  assign n18676 = n18672 | n18675 ;
  assign n71593 = ~n18333 ;
  assign n18680 = n71593 & n18676 ;
  assign n18681 = n18679 | n18680 ;
  assign n71594 = ~n18325 ;
  assign n18682 = n71594 & n18681 ;
  assign n71595 = ~n18315 ;
  assign n18683 = x93 & n71595 ;
  assign n71596 = ~n18313 ;
  assign n18684 = n71596 & n18683 ;
  assign n18685 = n18317 | n18684 ;
  assign n18686 = n18682 | n18685 ;
  assign n71597 = ~n18317 ;
  assign n18690 = n71597 & n18686 ;
  assign n18691 = n18689 | n18690 ;
  assign n71598 = ~n18309 ;
  assign n18692 = n71598 & n18691 ;
  assign n71599 = ~n18299 ;
  assign n18693 = x95 & n71599 ;
  assign n71600 = ~n18297 ;
  assign n18694 = n71600 & n18693 ;
  assign n18695 = n18301 | n18694 ;
  assign n18696 = n18692 | n18695 ;
  assign n71601 = ~n18301 ;
  assign n18700 = n71601 & n18696 ;
  assign n18701 = n18699 | n18700 ;
  assign n71602 = ~n18293 ;
  assign n18702 = n71602 & n18701 ;
  assign n71603 = ~n18283 ;
  assign n18703 = x97 & n71603 ;
  assign n71604 = ~n18281 ;
  assign n18704 = n71604 & n18703 ;
  assign n18705 = n18285 | n18704 ;
  assign n18706 = n18702 | n18705 ;
  assign n71605 = ~n18285 ;
  assign n18710 = n71605 & n18706 ;
  assign n18711 = n18709 | n18710 ;
  assign n71606 = ~n18277 ;
  assign n18712 = n71606 & n18711 ;
  assign n71607 = ~n18267 ;
  assign n18713 = x99 & n71607 ;
  assign n71608 = ~n18265 ;
  assign n18714 = n71608 & n18713 ;
  assign n18715 = n18269 | n18714 ;
  assign n18716 = n18712 | n18715 ;
  assign n71609 = ~n18269 ;
  assign n18720 = n71609 & n18716 ;
  assign n18721 = n18719 | n18720 ;
  assign n71610 = ~n18261 ;
  assign n18722 = n71610 & n18721 ;
  assign n71611 = ~n18251 ;
  assign n18723 = x101 & n71611 ;
  assign n71612 = ~n18249 ;
  assign n18724 = n71612 & n18723 ;
  assign n18725 = n18253 | n18724 ;
  assign n18726 = n18722 | n18725 ;
  assign n71613 = ~n18253 ;
  assign n18730 = n71613 & n18726 ;
  assign n18731 = n18729 | n18730 ;
  assign n71614 = ~n18245 ;
  assign n18732 = n71614 & n18731 ;
  assign n71615 = ~n18235 ;
  assign n18733 = x103 & n71615 ;
  assign n71616 = ~n18233 ;
  assign n18734 = n71616 & n18733 ;
  assign n18735 = n18237 | n18734 ;
  assign n18736 = n18732 | n18735 ;
  assign n71617 = ~n18237 ;
  assign n18740 = n71617 & n18736 ;
  assign n18741 = n18739 | n18740 ;
  assign n71618 = ~n18229 ;
  assign n18742 = n71618 & n18741 ;
  assign n71619 = ~n18219 ;
  assign n18743 = x105 & n71619 ;
  assign n71620 = ~n18217 ;
  assign n18744 = n71620 & n18743 ;
  assign n18745 = n18221 | n18744 ;
  assign n18746 = n18742 | n18745 ;
  assign n71621 = ~n18221 ;
  assign n18750 = n71621 & n18746 ;
  assign n18751 = n18749 | n18750 ;
  assign n71622 = ~n18213 ;
  assign n18752 = n71622 & n18751 ;
  assign n71623 = ~n18203 ;
  assign n18753 = x107 & n71623 ;
  assign n71624 = ~n18201 ;
  assign n18754 = n71624 & n18753 ;
  assign n18755 = n18205 | n18754 ;
  assign n18756 = n18752 | n18755 ;
  assign n71625 = ~n18205 ;
  assign n18760 = n71625 & n18756 ;
  assign n18761 = n18759 | n18760 ;
  assign n71626 = ~n18197 ;
  assign n18762 = n71626 & n18761 ;
  assign n71627 = ~n18187 ;
  assign n18763 = x109 & n71627 ;
  assign n71628 = ~n18185 ;
  assign n18764 = n71628 & n18763 ;
  assign n18765 = n18189 | n18764 ;
  assign n18767 = n18762 | n18765 ;
  assign n71629 = ~n18189 ;
  assign n18771 = n71629 & n18767 ;
  assign n18772 = n18770 | n18771 ;
  assign n71630 = ~n18181 ;
  assign n18773 = n71630 & n18772 ;
  assign n18774 = n17426 | n18045 ;
  assign n18775 = n18041 | n18774 ;
  assign n71631 = ~n18775 ;
  assign n18776 = n18033 & n71631 ;
  assign n18777 = n18041 | n18045 ;
  assign n71632 = ~n18176 ;
  assign n18778 = n71632 & n18777 ;
  assign n18779 = n18776 | n18778 ;
  assign n18780 = n146 & n18779 ;
  assign n18781 = n17324 & n18040 ;
  assign n18782 = n18177 & n18781 ;
  assign n18783 = n18780 | n18782 ;
  assign n71633 = ~x111 ;
  assign n18784 = n71633 & n18783 ;
  assign n71634 = ~n18782 ;
  assign n18785 = x111 & n71634 ;
  assign n71635 = ~n18780 ;
  assign n18786 = n71635 & n18785 ;
  assign n18787 = n66858 | n18786 ;
  assign n18788 = n18784 | n18787 ;
  assign n18789 = n18773 | n18788 ;
  assign n71636 = ~n18047 ;
  assign n18790 = n71636 & n18783 ;
  assign n71637 = ~n18790 ;
  assign n18791 = n18789 & n71637 ;
  assign n71638 = ~n18771 ;
  assign n18902 = n18770 & n71638 ;
  assign n18795 = x64 & n71538 ;
  assign n71639 = ~n18795 ;
  assign n18796 = x17 & n71639 ;
  assign n18797 = n18054 | n18796 ;
  assign n18798 = x65 & n18797 ;
  assign n71640 = ~n18798 ;
  assign n18799 = n18541 & n71640 ;
  assign n18800 = n18543 | n18799 ;
  assign n18801 = n71541 & n18800 ;
  assign n18803 = n18548 | n18801 ;
  assign n18804 = n71542 & n18803 ;
  assign n18805 = n18554 | n18804 ;
  assign n18806 = n71545 & n18805 ;
  assign n18807 = n18558 | n18806 ;
  assign n18808 = n71546 & n18807 ;
  assign n18809 = n18564 | n18808 ;
  assign n18810 = n71549 & n18809 ;
  assign n18811 = n18568 | n18810 ;
  assign n18812 = n71550 & n18811 ;
  assign n18813 = n18574 | n18812 ;
  assign n18814 = n71553 & n18813 ;
  assign n18815 = n18578 | n18814 ;
  assign n18816 = n71554 & n18815 ;
  assign n18817 = n18584 | n18816 ;
  assign n18818 = n71557 & n18817 ;
  assign n18819 = n18588 | n18818 ;
  assign n18820 = n71558 & n18819 ;
  assign n18821 = n18594 | n18820 ;
  assign n18822 = n71561 & n18821 ;
  assign n18823 = n18598 | n18822 ;
  assign n18824 = n71562 & n18823 ;
  assign n18825 = n18604 | n18824 ;
  assign n18826 = n71565 & n18825 ;
  assign n18827 = n18608 | n18826 ;
  assign n18828 = n71566 & n18827 ;
  assign n18829 = n18614 | n18828 ;
  assign n18830 = n71569 & n18829 ;
  assign n18831 = n18618 | n18830 ;
  assign n18832 = n71570 & n18831 ;
  assign n18833 = n18624 | n18832 ;
  assign n18834 = n71573 & n18833 ;
  assign n18835 = n18628 | n18834 ;
  assign n18836 = n71574 & n18835 ;
  assign n18837 = n18634 | n18836 ;
  assign n18838 = n71577 & n18837 ;
  assign n18839 = n18638 | n18838 ;
  assign n18840 = n71578 & n18839 ;
  assign n18841 = n18644 | n18840 ;
  assign n18842 = n71581 & n18841 ;
  assign n18843 = n18649 | n18842 ;
  assign n18844 = n71582 & n18843 ;
  assign n18845 = n18655 | n18844 ;
  assign n18846 = n71585 & n18845 ;
  assign n18847 = n18659 | n18846 ;
  assign n18848 = n71586 & n18847 ;
  assign n18849 = n18665 | n18848 ;
  assign n18850 = n71589 & n18849 ;
  assign n18851 = n18669 | n18850 ;
  assign n18852 = n71590 & n18851 ;
  assign n18853 = n18675 | n18852 ;
  assign n18854 = n71593 & n18853 ;
  assign n18855 = n18679 | n18854 ;
  assign n18856 = n71594 & n18855 ;
  assign n18857 = n18685 | n18856 ;
  assign n18858 = n71597 & n18857 ;
  assign n18859 = n18689 | n18858 ;
  assign n18860 = n71598 & n18859 ;
  assign n18861 = n18695 | n18860 ;
  assign n18862 = n71601 & n18861 ;
  assign n18863 = n18699 | n18862 ;
  assign n18864 = n71602 & n18863 ;
  assign n18865 = n18705 | n18864 ;
  assign n18866 = n71605 & n18865 ;
  assign n18867 = n18709 | n18866 ;
  assign n18868 = n71606 & n18867 ;
  assign n18869 = n18715 | n18868 ;
  assign n18870 = n71609 & n18869 ;
  assign n18871 = n18719 | n18870 ;
  assign n18872 = n71610 & n18871 ;
  assign n18873 = n18725 | n18872 ;
  assign n18874 = n71613 & n18873 ;
  assign n18875 = n18729 | n18874 ;
  assign n18876 = n71614 & n18875 ;
  assign n18877 = n18735 | n18876 ;
  assign n18878 = n71617 & n18877 ;
  assign n18879 = n18739 | n18878 ;
  assign n18880 = n71618 & n18879 ;
  assign n18881 = n18745 | n18880 ;
  assign n18882 = n71621 & n18881 ;
  assign n18883 = n18749 | n18882 ;
  assign n18884 = n71622 & n18883 ;
  assign n18885 = n18755 | n18884 ;
  assign n18886 = n71625 & n18885 ;
  assign n18887 = n18759 | n18886 ;
  assign n18888 = n71626 & n18887 ;
  assign n18889 = n18765 | n18888 ;
  assign n18903 = n18189 | n18770 ;
  assign n71641 = ~n18903 ;
  assign n18904 = n18889 & n71641 ;
  assign n18905 = n18902 | n18904 ;
  assign n145 = ~n18791 ;
  assign n18906 = n145 & n18905 ;
  assign n18907 = n18180 & n71637 ;
  assign n18908 = n18789 & n18907 ;
  assign n18909 = n18906 | n18908 ;
  assign n18792 = n18181 | n18786 ;
  assign n18793 = n18784 | n18792 ;
  assign n71643 = ~n18793 ;
  assign n18794 = n18772 & n71643 ;
  assign n18890 = n71629 & n18889 ;
  assign n18891 = n18770 | n18890 ;
  assign n18892 = n71630 & n18891 ;
  assign n18893 = n18784 | n18786 ;
  assign n71644 = ~n18892 ;
  assign n18894 = n71644 & n18893 ;
  assign n18895 = n18794 | n18894 ;
  assign n18896 = n145 & n18895 ;
  assign n18897 = n18047 & n18783 ;
  assign n18898 = n18789 & n18897 ;
  assign n18899 = n18896 | n18898 ;
  assign n71645 = ~x112 ;
  assign n18900 = n71645 & n18899 ;
  assign n18910 = n71633 & n18909 ;
  assign n71646 = ~n18888 ;
  assign n18911 = n18765 & n71646 ;
  assign n18766 = n18197 | n18765 ;
  assign n71647 = ~n18766 ;
  assign n18912 = n71647 & n18887 ;
  assign n18913 = n18911 | n18912 ;
  assign n18914 = n145 & n18913 ;
  assign n18915 = n18188 & n71637 ;
  assign n18916 = n18789 & n18915 ;
  assign n18917 = n18914 | n18916 ;
  assign n18918 = n71253 & n18917 ;
  assign n71648 = ~n18760 ;
  assign n18919 = n18759 & n71648 ;
  assign n18920 = n18205 | n18759 ;
  assign n71649 = ~n18920 ;
  assign n18921 = n18885 & n71649 ;
  assign n18922 = n18919 | n18921 ;
  assign n18923 = n145 & n18922 ;
  assign n18924 = n18196 & n71637 ;
  assign n18925 = n18789 & n18924 ;
  assign n18926 = n18923 | n18925 ;
  assign n18927 = n70935 & n18926 ;
  assign n71650 = ~n18884 ;
  assign n18928 = n18755 & n71650 ;
  assign n18929 = n18213 | n18755 ;
  assign n71651 = ~n18929 ;
  assign n18930 = n18751 & n71651 ;
  assign n18931 = n18928 | n18930 ;
  assign n18932 = n145 & n18931 ;
  assign n18933 = n18204 & n71637 ;
  assign n18934 = n18789 & n18933 ;
  assign n18935 = n18932 | n18934 ;
  assign n18936 = n70927 & n18935 ;
  assign n71652 = ~n18750 ;
  assign n18937 = n18749 & n71652 ;
  assign n18938 = n18221 | n18749 ;
  assign n71653 = ~n18938 ;
  assign n18939 = n18881 & n71653 ;
  assign n18940 = n18937 | n18939 ;
  assign n18941 = n145 & n18940 ;
  assign n18942 = n18212 & n71637 ;
  assign n18943 = n18789 & n18942 ;
  assign n18944 = n18941 | n18943 ;
  assign n18945 = n70609 & n18944 ;
  assign n71654 = ~n18880 ;
  assign n18946 = n18745 & n71654 ;
  assign n18947 = n18229 | n18745 ;
  assign n71655 = ~n18947 ;
  assign n18948 = n18741 & n71655 ;
  assign n18949 = n18946 | n18948 ;
  assign n18950 = n145 & n18949 ;
  assign n18951 = n18220 & n71637 ;
  assign n18952 = n18789 & n18951 ;
  assign n18953 = n18950 | n18952 ;
  assign n18954 = n70276 & n18953 ;
  assign n71656 = ~n18740 ;
  assign n18955 = n18739 & n71656 ;
  assign n18956 = n18237 | n18739 ;
  assign n71657 = ~n18956 ;
  assign n18957 = n18877 & n71657 ;
  assign n18958 = n18955 | n18957 ;
  assign n18959 = n145 & n18958 ;
  assign n18960 = n18228 & n71637 ;
  assign n18961 = n18789 & n18960 ;
  assign n18962 = n18959 | n18961 ;
  assign n18963 = n70176 & n18962 ;
  assign n71658 = ~n18876 ;
  assign n18964 = n18735 & n71658 ;
  assign n18965 = n18245 | n18735 ;
  assign n71659 = ~n18965 ;
  assign n18966 = n18731 & n71659 ;
  assign n18967 = n18964 | n18966 ;
  assign n18968 = n145 & n18967 ;
  assign n18969 = n18236 & n71637 ;
  assign n18970 = n18789 & n18969 ;
  assign n18971 = n18968 | n18970 ;
  assign n18972 = n69857 & n18971 ;
  assign n71660 = ~n18730 ;
  assign n18973 = n18729 & n71660 ;
  assign n18974 = n18253 | n18729 ;
  assign n71661 = ~n18974 ;
  assign n18975 = n18873 & n71661 ;
  assign n18976 = n18973 | n18975 ;
  assign n18977 = n145 & n18976 ;
  assign n18978 = n18244 & n71637 ;
  assign n18979 = n18789 & n18978 ;
  assign n18980 = n18977 | n18979 ;
  assign n18981 = n69656 & n18980 ;
  assign n71662 = ~n18872 ;
  assign n18982 = n18725 & n71662 ;
  assign n18983 = n18261 | n18725 ;
  assign n71663 = ~n18983 ;
  assign n18984 = n18721 & n71663 ;
  assign n18985 = n18982 | n18984 ;
  assign n18986 = n145 & n18985 ;
  assign n18987 = n18252 & n71637 ;
  assign n18988 = n18789 & n18987 ;
  assign n18989 = n18986 | n18988 ;
  assign n18990 = n69528 & n18989 ;
  assign n71664 = ~n18720 ;
  assign n18991 = n18719 & n71664 ;
  assign n18992 = n18269 | n18719 ;
  assign n71665 = ~n18992 ;
  assign n18993 = n18869 & n71665 ;
  assign n18994 = n18991 | n18993 ;
  assign n18995 = n145 & n18994 ;
  assign n18996 = n18260 & n71637 ;
  assign n18997 = n18789 & n18996 ;
  assign n18998 = n18995 | n18997 ;
  assign n18999 = n69261 & n18998 ;
  assign n71666 = ~n18868 ;
  assign n19000 = n18715 & n71666 ;
  assign n19001 = n18277 | n18715 ;
  assign n71667 = ~n19001 ;
  assign n19002 = n18711 & n71667 ;
  assign n19003 = n19000 | n19002 ;
  assign n19004 = n145 & n19003 ;
  assign n19005 = n18268 & n71637 ;
  assign n19006 = n18789 & n19005 ;
  assign n19007 = n19004 | n19006 ;
  assign n19008 = n69075 & n19007 ;
  assign n71668 = ~n18710 ;
  assign n19009 = n18709 & n71668 ;
  assign n19010 = n18285 | n18709 ;
  assign n71669 = ~n19010 ;
  assign n19011 = n18865 & n71669 ;
  assign n19012 = n19009 | n19011 ;
  assign n19013 = n145 & n19012 ;
  assign n19014 = n18276 & n71637 ;
  assign n19015 = n18789 & n19014 ;
  assign n19016 = n19013 | n19015 ;
  assign n19017 = n68993 & n19016 ;
  assign n71670 = ~n18864 ;
  assign n19018 = n18705 & n71670 ;
  assign n19019 = n18293 | n18705 ;
  assign n71671 = ~n19019 ;
  assign n19020 = n18701 & n71671 ;
  assign n19021 = n19018 | n19020 ;
  assign n19022 = n145 & n19021 ;
  assign n19023 = n18284 & n71637 ;
  assign n19024 = n18789 & n19023 ;
  assign n19025 = n19022 | n19024 ;
  assign n19026 = n68716 & n19025 ;
  assign n71672 = ~n18700 ;
  assign n19027 = n18699 & n71672 ;
  assign n19028 = n18301 | n18699 ;
  assign n71673 = ~n19028 ;
  assign n19029 = n18861 & n71673 ;
  assign n19030 = n19027 | n19029 ;
  assign n19031 = n145 & n19030 ;
  assign n19032 = n18292 & n71637 ;
  assign n19033 = n18789 & n19032 ;
  assign n19034 = n19031 | n19033 ;
  assign n19035 = n68545 & n19034 ;
  assign n71674 = ~n18860 ;
  assign n19036 = n18695 & n71674 ;
  assign n19037 = n18309 | n18695 ;
  assign n71675 = ~n19037 ;
  assign n19038 = n18691 & n71675 ;
  assign n19039 = n19036 | n19038 ;
  assign n19040 = n145 & n19039 ;
  assign n19041 = n18300 & n71637 ;
  assign n19042 = n18789 & n19041 ;
  assign n19043 = n19040 | n19042 ;
  assign n19044 = n68438 & n19043 ;
  assign n71676 = ~n18690 ;
  assign n19045 = n18689 & n71676 ;
  assign n19046 = n18317 | n18689 ;
  assign n71677 = ~n19046 ;
  assign n19047 = n18857 & n71677 ;
  assign n19048 = n19045 | n19047 ;
  assign n19049 = n145 & n19048 ;
  assign n19050 = n18308 & n71637 ;
  assign n19051 = n18789 & n19050 ;
  assign n19052 = n19049 | n19051 ;
  assign n19053 = n68214 & n19052 ;
  assign n71678 = ~n18856 ;
  assign n19054 = n18685 & n71678 ;
  assign n19055 = n18325 | n18685 ;
  assign n71679 = ~n19055 ;
  assign n19056 = n18681 & n71679 ;
  assign n19057 = n19054 | n19056 ;
  assign n19058 = n145 & n19057 ;
  assign n19059 = n18316 & n71637 ;
  assign n19060 = n18789 & n19059 ;
  assign n19061 = n19058 | n19060 ;
  assign n19062 = n68058 & n19061 ;
  assign n71680 = ~n18680 ;
  assign n19063 = n18679 & n71680 ;
  assign n19064 = n18333 | n18679 ;
  assign n71681 = ~n19064 ;
  assign n19065 = n18853 & n71681 ;
  assign n19066 = n19063 | n19065 ;
  assign n19067 = n145 & n19066 ;
  assign n19068 = n18324 & n71637 ;
  assign n19069 = n18789 & n19068 ;
  assign n19070 = n19067 | n19069 ;
  assign n19071 = n67986 & n19070 ;
  assign n71682 = ~n18852 ;
  assign n19072 = n18675 & n71682 ;
  assign n19073 = n18341 | n18675 ;
  assign n71683 = ~n19073 ;
  assign n19074 = n18671 & n71683 ;
  assign n19075 = n19072 | n19074 ;
  assign n19076 = n145 & n19075 ;
  assign n19077 = n18332 & n71637 ;
  assign n19078 = n18789 & n19077 ;
  assign n19079 = n19076 | n19078 ;
  assign n19080 = n67763 & n19079 ;
  assign n71684 = ~n18670 ;
  assign n19081 = n18669 & n71684 ;
  assign n19082 = n18349 | n18669 ;
  assign n71685 = ~n19082 ;
  assign n19083 = n18849 & n71685 ;
  assign n19084 = n19081 | n19083 ;
  assign n19085 = n145 & n19084 ;
  assign n19086 = n18340 & n71637 ;
  assign n19087 = n18789 & n19086 ;
  assign n19088 = n19085 | n19087 ;
  assign n19089 = n67622 & n19088 ;
  assign n71686 = ~n18848 ;
  assign n19090 = n18665 & n71686 ;
  assign n19091 = n18357 | n18665 ;
  assign n71687 = ~n19091 ;
  assign n19092 = n18661 & n71687 ;
  assign n19093 = n19090 | n19092 ;
  assign n19094 = n145 & n19093 ;
  assign n19095 = n18348 & n71637 ;
  assign n19096 = n18789 & n19095 ;
  assign n19097 = n19094 | n19096 ;
  assign n19098 = n67531 & n19097 ;
  assign n71688 = ~n18660 ;
  assign n19099 = n18659 & n71688 ;
  assign n19100 = n18365 | n18659 ;
  assign n71689 = ~n19100 ;
  assign n19101 = n18845 & n71689 ;
  assign n19102 = n19099 | n19101 ;
  assign n19103 = n145 & n19102 ;
  assign n19104 = n18356 & n71637 ;
  assign n19105 = n18789 & n19104 ;
  assign n19106 = n19103 | n19105 ;
  assign n19107 = n67348 & n19106 ;
  assign n71690 = ~n18844 ;
  assign n19108 = n18655 & n71690 ;
  assign n19109 = n18373 | n18655 ;
  assign n71691 = ~n19109 ;
  assign n19110 = n18651 & n71691 ;
  assign n19111 = n19108 | n19110 ;
  assign n19112 = n145 & n19111 ;
  assign n19113 = n18364 & n71637 ;
  assign n19114 = n18789 & n19113 ;
  assign n19115 = n19112 | n19114 ;
  assign n19116 = n67222 & n19115 ;
  assign n71692 = ~n18650 ;
  assign n19117 = n18649 & n71692 ;
  assign n19118 = n18381 | n18649 ;
  assign n71693 = ~n19118 ;
  assign n19119 = n18841 & n71693 ;
  assign n19120 = n19117 | n19119 ;
  assign n19121 = n145 & n19120 ;
  assign n19122 = n18372 & n71637 ;
  assign n19123 = n18789 & n19122 ;
  assign n19124 = n19121 | n19123 ;
  assign n19125 = n67164 & n19124 ;
  assign n71694 = ~n18840 ;
  assign n19126 = n18644 & n71694 ;
  assign n18645 = n18389 | n18644 ;
  assign n71695 = ~n18645 ;
  assign n19127 = n71695 & n18839 ;
  assign n19128 = n19126 | n19127 ;
  assign n19129 = n145 & n19128 ;
  assign n19130 = n18380 & n71637 ;
  assign n19131 = n18789 & n19130 ;
  assign n19132 = n19129 | n19131 ;
  assign n19133 = n66979 & n19132 ;
  assign n71696 = ~n18639 ;
  assign n19134 = n18638 & n71696 ;
  assign n19135 = n18397 | n18638 ;
  assign n71697 = ~n19135 ;
  assign n19136 = n18837 & n71697 ;
  assign n19137 = n19134 | n19136 ;
  assign n19138 = n145 & n19137 ;
  assign n19139 = n18388 & n71637 ;
  assign n19140 = n18789 & n19139 ;
  assign n19141 = n19138 | n19140 ;
  assign n19142 = n66868 & n19141 ;
  assign n71698 = ~n18836 ;
  assign n19143 = n18634 & n71698 ;
  assign n19144 = n18405 | n18634 ;
  assign n71699 = ~n19144 ;
  assign n19145 = n18630 & n71699 ;
  assign n19146 = n19143 | n19145 ;
  assign n19147 = n145 & n19146 ;
  assign n19148 = n18396 & n71637 ;
  assign n19149 = n18789 & n19148 ;
  assign n19150 = n19147 | n19149 ;
  assign n19151 = n66797 & n19150 ;
  assign n71700 = ~n18629 ;
  assign n19152 = n18628 & n71700 ;
  assign n19153 = n18413 | n18628 ;
  assign n71701 = ~n19153 ;
  assign n19154 = n18833 & n71701 ;
  assign n19155 = n19152 | n19154 ;
  assign n19156 = n145 & n19155 ;
  assign n19157 = n18404 & n71637 ;
  assign n19158 = n18789 & n19157 ;
  assign n19159 = n19156 | n19158 ;
  assign n19160 = n66654 & n19159 ;
  assign n71702 = ~n18832 ;
  assign n19161 = n18624 & n71702 ;
  assign n19162 = n18421 | n18624 ;
  assign n71703 = ~n19162 ;
  assign n19163 = n18620 & n71703 ;
  assign n19164 = n19161 | n19163 ;
  assign n19165 = n145 & n19164 ;
  assign n19166 = n18412 & n71637 ;
  assign n19167 = n18789 & n19166 ;
  assign n19168 = n19165 | n19167 ;
  assign n19169 = n66560 & n19168 ;
  assign n71704 = ~n18619 ;
  assign n19170 = n18618 & n71704 ;
  assign n19171 = n18429 | n18618 ;
  assign n71705 = ~n19171 ;
  assign n19172 = n18829 & n71705 ;
  assign n19173 = n19170 | n19172 ;
  assign n19174 = n145 & n19173 ;
  assign n19175 = n18420 & n71637 ;
  assign n19176 = n18789 & n19175 ;
  assign n19177 = n19174 | n19176 ;
  assign n19178 = n66505 & n19177 ;
  assign n71706 = ~n18828 ;
  assign n19179 = n18614 & n71706 ;
  assign n19180 = n18437 | n18614 ;
  assign n71707 = ~n19180 ;
  assign n19181 = n18610 & n71707 ;
  assign n19182 = n19179 | n19181 ;
  assign n19183 = n145 & n19182 ;
  assign n19184 = n18428 & n71637 ;
  assign n19185 = n18789 & n19184 ;
  assign n19186 = n19183 | n19185 ;
  assign n19187 = n66379 & n19186 ;
  assign n71708 = ~n18609 ;
  assign n19188 = n18608 & n71708 ;
  assign n19189 = n18445 | n18608 ;
  assign n71709 = ~n19189 ;
  assign n19190 = n18825 & n71709 ;
  assign n19191 = n19188 | n19190 ;
  assign n19192 = n145 & n19191 ;
  assign n19193 = n18436 & n71637 ;
  assign n19194 = n18789 & n19193 ;
  assign n19195 = n19192 | n19194 ;
  assign n19196 = n66299 & n19195 ;
  assign n71710 = ~n18824 ;
  assign n19197 = n18604 & n71710 ;
  assign n19198 = n18453 | n18604 ;
  assign n71711 = ~n19198 ;
  assign n19199 = n18600 & n71711 ;
  assign n19200 = n19197 | n19199 ;
  assign n19201 = n145 & n19200 ;
  assign n19202 = n18444 & n71637 ;
  assign n19203 = n18789 & n19202 ;
  assign n19204 = n19201 | n19203 ;
  assign n19205 = n66244 & n19204 ;
  assign n71712 = ~n18599 ;
  assign n19206 = n18598 & n71712 ;
  assign n19207 = n18461 | n18598 ;
  assign n71713 = ~n19207 ;
  assign n19208 = n18821 & n71713 ;
  assign n19209 = n19206 | n19208 ;
  assign n19210 = n145 & n19209 ;
  assign n19211 = n18452 & n71637 ;
  assign n19212 = n18789 & n19211 ;
  assign n19213 = n19210 | n19212 ;
  assign n19214 = n66145 & n19213 ;
  assign n71714 = ~n18820 ;
  assign n19215 = n18594 & n71714 ;
  assign n19216 = n18469 | n18594 ;
  assign n71715 = ~n19216 ;
  assign n19217 = n18590 & n71715 ;
  assign n19218 = n19215 | n19217 ;
  assign n19219 = n145 & n19218 ;
  assign n19220 = n18460 & n71637 ;
  assign n19221 = n18789 & n19220 ;
  assign n19222 = n19219 | n19221 ;
  assign n19223 = n66081 & n19222 ;
  assign n71716 = ~n18589 ;
  assign n19224 = n18588 & n71716 ;
  assign n19225 = n18477 | n18588 ;
  assign n71717 = ~n19225 ;
  assign n19226 = n18817 & n71717 ;
  assign n19227 = n19224 | n19226 ;
  assign n19228 = n145 & n19227 ;
  assign n19229 = n18468 & n71637 ;
  assign n19230 = n18789 & n19229 ;
  assign n19231 = n19228 | n19230 ;
  assign n19232 = n66043 & n19231 ;
  assign n71718 = ~n18816 ;
  assign n19233 = n18584 & n71718 ;
  assign n19234 = n18485 | n18584 ;
  assign n71719 = ~n19234 ;
  assign n19235 = n18580 & n71719 ;
  assign n19236 = n19233 | n19235 ;
  assign n19237 = n145 & n19236 ;
  assign n19238 = n18476 & n71637 ;
  assign n19239 = n18789 & n19238 ;
  assign n19240 = n19237 | n19239 ;
  assign n19241 = n65960 & n19240 ;
  assign n71720 = ~n18579 ;
  assign n19242 = n18578 & n71720 ;
  assign n19243 = n18493 | n18578 ;
  assign n71721 = ~n19243 ;
  assign n19244 = n18813 & n71721 ;
  assign n19245 = n19242 | n19244 ;
  assign n19246 = n145 & n19245 ;
  assign n19247 = n18484 & n71637 ;
  assign n19248 = n18789 & n19247 ;
  assign n19249 = n19246 | n19248 ;
  assign n19250 = n65909 & n19249 ;
  assign n71722 = ~n18812 ;
  assign n19251 = n18574 & n71722 ;
  assign n19252 = n18501 | n18574 ;
  assign n71723 = ~n19252 ;
  assign n19253 = n18570 & n71723 ;
  assign n19254 = n19251 | n19253 ;
  assign n19255 = n145 & n19254 ;
  assign n19256 = n18492 & n71637 ;
  assign n19257 = n18789 & n19256 ;
  assign n19258 = n19255 | n19257 ;
  assign n19259 = n65877 & n19258 ;
  assign n71724 = ~n18569 ;
  assign n19260 = n18568 & n71724 ;
  assign n19261 = n18510 | n18568 ;
  assign n71725 = ~n19261 ;
  assign n19262 = n18809 & n71725 ;
  assign n19263 = n19260 | n19262 ;
  assign n19264 = n145 & n19263 ;
  assign n19265 = n18500 & n71637 ;
  assign n19266 = n18789 & n19265 ;
  assign n19267 = n19264 | n19266 ;
  assign n19268 = n65820 & n19267 ;
  assign n71726 = ~n18808 ;
  assign n19269 = n18564 & n71726 ;
  assign n19270 = n18518 | n18564 ;
  assign n71727 = ~n19270 ;
  assign n19271 = n18560 & n71727 ;
  assign n19272 = n19269 | n19271 ;
  assign n19273 = n145 & n19272 ;
  assign n19274 = n18509 & n71637 ;
  assign n19275 = n18789 & n19274 ;
  assign n19276 = n19273 | n19275 ;
  assign n19277 = n65791 & n19276 ;
  assign n71728 = ~n18559 ;
  assign n19278 = n18558 & n71728 ;
  assign n19279 = n18526 | n18558 ;
  assign n71729 = ~n19279 ;
  assign n19280 = n18805 & n71729 ;
  assign n19281 = n19278 | n19280 ;
  assign n19282 = n145 & n19281 ;
  assign n19283 = n18517 & n71637 ;
  assign n19284 = n18789 & n19283 ;
  assign n19285 = n19282 | n19284 ;
  assign n19286 = n65772 & n19285 ;
  assign n71730 = ~n18804 ;
  assign n19288 = n18554 & n71730 ;
  assign n19287 = n18534 | n18554 ;
  assign n71731 = ~n19287 ;
  assign n19289 = n18803 & n71731 ;
  assign n19290 = n19288 | n19289 ;
  assign n19291 = n145 & n19290 ;
  assign n19292 = n18525 & n71637 ;
  assign n19293 = n18789 & n19292 ;
  assign n19294 = n19291 | n19293 ;
  assign n19295 = n65746 & n19294 ;
  assign n71732 = ~n18549 ;
  assign n19296 = n18548 & n71732 ;
  assign n18802 = n18545 | n18548 ;
  assign n71733 = ~n18802 ;
  assign n19297 = n18544 & n71733 ;
  assign n19298 = n19296 | n19297 ;
  assign n19299 = n145 & n19298 ;
  assign n19300 = n18533 & n71637 ;
  assign n19301 = n18789 & n19300 ;
  assign n19302 = n19299 | n19301 ;
  assign n19303 = n65721 & n19302 ;
  assign n19304 = n18541 & n18543 ;
  assign n19305 = n71539 & n19304 ;
  assign n71734 = ~n19305 ;
  assign n19306 = n18544 & n71734 ;
  assign n19307 = n145 & n19306 ;
  assign n19308 = n18536 & n71637 ;
  assign n19309 = n18789 & n19308 ;
  assign n19310 = n19307 | n19309 ;
  assign n19311 = n65686 & n19310 ;
  assign n18901 = n18543 & n145 ;
  assign n19312 = x64 & n145 ;
  assign n71735 = ~n19312 ;
  assign n19313 = x16 & n71735 ;
  assign n19314 = n18901 | n19313 ;
  assign n19325 = n65670 & n19314 ;
  assign n19315 = n18788 | n18892 ;
  assign n19316 = n71637 & n19315 ;
  assign n71736 = ~n19316 ;
  assign n19317 = x64 & n71736 ;
  assign n71737 = ~n19317 ;
  assign n19318 = x16 & n71737 ;
  assign n19319 = n18901 | n19318 ;
  assign n19320 = x65 & n19319 ;
  assign n19321 = x65 | n18901 ;
  assign n19322 = n19318 | n19321 ;
  assign n71738 = ~n19320 ;
  assign n19323 = n71738 & n19322 ;
  assign n71739 = ~x15 ;
  assign n19324 = n71739 & x64 ;
  assign n19326 = n19323 | n19324 ;
  assign n71740 = ~n19325 ;
  assign n19327 = n71740 & n19326 ;
  assign n71741 = ~n19309 ;
  assign n19328 = x66 & n71741 ;
  assign n71742 = ~n19307 ;
  assign n19329 = n71742 & n19328 ;
  assign n19330 = n19311 | n19329 ;
  assign n19331 = n19327 | n19330 ;
  assign n71743 = ~n19311 ;
  assign n19332 = n71743 & n19331 ;
  assign n71744 = ~n19301 ;
  assign n19333 = x67 & n71744 ;
  assign n71745 = ~n19299 ;
  assign n19334 = n71745 & n19333 ;
  assign n19335 = n19303 | n19334 ;
  assign n19336 = n19332 | n19335 ;
  assign n71746 = ~n19303 ;
  assign n19337 = n71746 & n19336 ;
  assign n71747 = ~n19293 ;
  assign n19338 = x68 & n71747 ;
  assign n71748 = ~n19291 ;
  assign n19339 = n71748 & n19338 ;
  assign n19340 = n19337 | n19339 ;
  assign n71749 = ~n19295 ;
  assign n19341 = n71749 & n19340 ;
  assign n71750 = ~n19284 ;
  assign n19342 = x69 & n71750 ;
  assign n71751 = ~n19282 ;
  assign n19343 = n71751 & n19342 ;
  assign n19344 = n19286 | n19343 ;
  assign n19345 = n19341 | n19344 ;
  assign n71752 = ~n19286 ;
  assign n19346 = n71752 & n19345 ;
  assign n71753 = ~n19275 ;
  assign n19347 = x70 & n71753 ;
  assign n71754 = ~n19273 ;
  assign n19348 = n71754 & n19347 ;
  assign n19349 = n19277 | n19348 ;
  assign n19351 = n19346 | n19349 ;
  assign n71755 = ~n19277 ;
  assign n19352 = n71755 & n19351 ;
  assign n71756 = ~n19266 ;
  assign n19353 = x71 & n71756 ;
  assign n71757 = ~n19264 ;
  assign n19354 = n71757 & n19353 ;
  assign n19355 = n19268 | n19354 ;
  assign n19356 = n19352 | n19355 ;
  assign n71758 = ~n19268 ;
  assign n19357 = n71758 & n19356 ;
  assign n71759 = ~n19257 ;
  assign n19358 = x72 & n71759 ;
  assign n71760 = ~n19255 ;
  assign n19359 = n71760 & n19358 ;
  assign n19360 = n19259 | n19359 ;
  assign n19362 = n19357 | n19360 ;
  assign n71761 = ~n19259 ;
  assign n19363 = n71761 & n19362 ;
  assign n71762 = ~n19248 ;
  assign n19364 = x73 & n71762 ;
  assign n71763 = ~n19246 ;
  assign n19365 = n71763 & n19364 ;
  assign n19366 = n19250 | n19365 ;
  assign n19367 = n19363 | n19366 ;
  assign n71764 = ~n19250 ;
  assign n19368 = n71764 & n19367 ;
  assign n71765 = ~n19239 ;
  assign n19369 = x74 & n71765 ;
  assign n71766 = ~n19237 ;
  assign n19370 = n71766 & n19369 ;
  assign n19371 = n19241 | n19370 ;
  assign n19373 = n19368 | n19371 ;
  assign n71767 = ~n19241 ;
  assign n19374 = n71767 & n19373 ;
  assign n71768 = ~n19230 ;
  assign n19375 = x75 & n71768 ;
  assign n71769 = ~n19228 ;
  assign n19376 = n71769 & n19375 ;
  assign n19377 = n19232 | n19376 ;
  assign n19378 = n19374 | n19377 ;
  assign n71770 = ~n19232 ;
  assign n19379 = n71770 & n19378 ;
  assign n71771 = ~n19221 ;
  assign n19380 = x76 & n71771 ;
  assign n71772 = ~n19219 ;
  assign n19381 = n71772 & n19380 ;
  assign n19382 = n19223 | n19381 ;
  assign n19384 = n19379 | n19382 ;
  assign n71773 = ~n19223 ;
  assign n19385 = n71773 & n19384 ;
  assign n71774 = ~n19212 ;
  assign n19386 = x77 & n71774 ;
  assign n71775 = ~n19210 ;
  assign n19387 = n71775 & n19386 ;
  assign n19388 = n19214 | n19387 ;
  assign n19389 = n19385 | n19388 ;
  assign n71776 = ~n19214 ;
  assign n19390 = n71776 & n19389 ;
  assign n71777 = ~n19203 ;
  assign n19391 = x78 & n71777 ;
  assign n71778 = ~n19201 ;
  assign n19392 = n71778 & n19391 ;
  assign n19393 = n19205 | n19392 ;
  assign n19395 = n19390 | n19393 ;
  assign n71779 = ~n19205 ;
  assign n19396 = n71779 & n19395 ;
  assign n71780 = ~n19194 ;
  assign n19397 = x79 & n71780 ;
  assign n71781 = ~n19192 ;
  assign n19398 = n71781 & n19397 ;
  assign n19399 = n19196 | n19398 ;
  assign n19400 = n19396 | n19399 ;
  assign n71782 = ~n19196 ;
  assign n19401 = n71782 & n19400 ;
  assign n71783 = ~n19185 ;
  assign n19402 = x80 & n71783 ;
  assign n71784 = ~n19183 ;
  assign n19403 = n71784 & n19402 ;
  assign n19404 = n19187 | n19403 ;
  assign n19406 = n19401 | n19404 ;
  assign n71785 = ~n19187 ;
  assign n19407 = n71785 & n19406 ;
  assign n71786 = ~n19176 ;
  assign n19408 = x81 & n71786 ;
  assign n71787 = ~n19174 ;
  assign n19409 = n71787 & n19408 ;
  assign n19410 = n19178 | n19409 ;
  assign n19411 = n19407 | n19410 ;
  assign n71788 = ~n19178 ;
  assign n19412 = n71788 & n19411 ;
  assign n71789 = ~n19167 ;
  assign n19413 = x82 & n71789 ;
  assign n71790 = ~n19165 ;
  assign n19414 = n71790 & n19413 ;
  assign n19415 = n19169 | n19414 ;
  assign n19417 = n19412 | n19415 ;
  assign n71791 = ~n19169 ;
  assign n19418 = n71791 & n19417 ;
  assign n71792 = ~n19158 ;
  assign n19419 = x83 & n71792 ;
  assign n71793 = ~n19156 ;
  assign n19420 = n71793 & n19419 ;
  assign n19421 = n19160 | n19420 ;
  assign n19422 = n19418 | n19421 ;
  assign n71794 = ~n19160 ;
  assign n19423 = n71794 & n19422 ;
  assign n71795 = ~n19149 ;
  assign n19424 = x84 & n71795 ;
  assign n71796 = ~n19147 ;
  assign n19425 = n71796 & n19424 ;
  assign n19426 = n19151 | n19425 ;
  assign n19428 = n19423 | n19426 ;
  assign n71797 = ~n19151 ;
  assign n19429 = n71797 & n19428 ;
  assign n71798 = ~n19140 ;
  assign n19430 = x85 & n71798 ;
  assign n71799 = ~n19138 ;
  assign n19431 = n71799 & n19430 ;
  assign n19432 = n19142 | n19431 ;
  assign n19433 = n19429 | n19432 ;
  assign n71800 = ~n19142 ;
  assign n19434 = n71800 & n19433 ;
  assign n71801 = ~n19131 ;
  assign n19435 = x86 & n71801 ;
  assign n71802 = ~n19129 ;
  assign n19436 = n71802 & n19435 ;
  assign n19437 = n19133 | n19436 ;
  assign n19439 = n19434 | n19437 ;
  assign n71803 = ~n19133 ;
  assign n19440 = n71803 & n19439 ;
  assign n71804 = ~n19123 ;
  assign n19441 = x87 & n71804 ;
  assign n71805 = ~n19121 ;
  assign n19442 = n71805 & n19441 ;
  assign n19443 = n19125 | n19442 ;
  assign n19444 = n19440 | n19443 ;
  assign n71806 = ~n19125 ;
  assign n19445 = n71806 & n19444 ;
  assign n71807 = ~n19114 ;
  assign n19446 = x88 & n71807 ;
  assign n71808 = ~n19112 ;
  assign n19447 = n71808 & n19446 ;
  assign n19448 = n19116 | n19447 ;
  assign n19450 = n19445 | n19448 ;
  assign n71809 = ~n19116 ;
  assign n19451 = n71809 & n19450 ;
  assign n71810 = ~n19105 ;
  assign n19452 = x89 & n71810 ;
  assign n71811 = ~n19103 ;
  assign n19453 = n71811 & n19452 ;
  assign n19454 = n19107 | n19453 ;
  assign n19455 = n19451 | n19454 ;
  assign n71812 = ~n19107 ;
  assign n19456 = n71812 & n19455 ;
  assign n71813 = ~n19096 ;
  assign n19457 = x90 & n71813 ;
  assign n71814 = ~n19094 ;
  assign n19458 = n71814 & n19457 ;
  assign n19459 = n19098 | n19458 ;
  assign n19461 = n19456 | n19459 ;
  assign n71815 = ~n19098 ;
  assign n19462 = n71815 & n19461 ;
  assign n71816 = ~n19087 ;
  assign n19463 = x91 & n71816 ;
  assign n71817 = ~n19085 ;
  assign n19464 = n71817 & n19463 ;
  assign n19465 = n19089 | n19464 ;
  assign n19466 = n19462 | n19465 ;
  assign n71818 = ~n19089 ;
  assign n19467 = n71818 & n19466 ;
  assign n71819 = ~n19078 ;
  assign n19468 = x92 & n71819 ;
  assign n71820 = ~n19076 ;
  assign n19469 = n71820 & n19468 ;
  assign n19470 = n19080 | n19469 ;
  assign n19472 = n19467 | n19470 ;
  assign n71821 = ~n19080 ;
  assign n19473 = n71821 & n19472 ;
  assign n71822 = ~n19069 ;
  assign n19474 = x93 & n71822 ;
  assign n71823 = ~n19067 ;
  assign n19475 = n71823 & n19474 ;
  assign n19476 = n19071 | n19475 ;
  assign n19477 = n19473 | n19476 ;
  assign n71824 = ~n19071 ;
  assign n19478 = n71824 & n19477 ;
  assign n71825 = ~n19060 ;
  assign n19479 = x94 & n71825 ;
  assign n71826 = ~n19058 ;
  assign n19480 = n71826 & n19479 ;
  assign n19481 = n19062 | n19480 ;
  assign n19483 = n19478 | n19481 ;
  assign n71827 = ~n19062 ;
  assign n19484 = n71827 & n19483 ;
  assign n71828 = ~n19051 ;
  assign n19485 = x95 & n71828 ;
  assign n71829 = ~n19049 ;
  assign n19486 = n71829 & n19485 ;
  assign n19487 = n19053 | n19486 ;
  assign n19488 = n19484 | n19487 ;
  assign n71830 = ~n19053 ;
  assign n19489 = n71830 & n19488 ;
  assign n71831 = ~n19042 ;
  assign n19490 = x96 & n71831 ;
  assign n71832 = ~n19040 ;
  assign n19491 = n71832 & n19490 ;
  assign n19492 = n19044 | n19491 ;
  assign n19494 = n19489 | n19492 ;
  assign n71833 = ~n19044 ;
  assign n19495 = n71833 & n19494 ;
  assign n71834 = ~n19033 ;
  assign n19496 = x97 & n71834 ;
  assign n71835 = ~n19031 ;
  assign n19497 = n71835 & n19496 ;
  assign n19498 = n19035 | n19497 ;
  assign n19499 = n19495 | n19498 ;
  assign n71836 = ~n19035 ;
  assign n19500 = n71836 & n19499 ;
  assign n71837 = ~n19024 ;
  assign n19501 = x98 & n71837 ;
  assign n71838 = ~n19022 ;
  assign n19502 = n71838 & n19501 ;
  assign n19503 = n19026 | n19502 ;
  assign n19505 = n19500 | n19503 ;
  assign n71839 = ~n19026 ;
  assign n19506 = n71839 & n19505 ;
  assign n71840 = ~n19015 ;
  assign n19507 = x99 & n71840 ;
  assign n71841 = ~n19013 ;
  assign n19508 = n71841 & n19507 ;
  assign n19509 = n19017 | n19508 ;
  assign n19510 = n19506 | n19509 ;
  assign n71842 = ~n19017 ;
  assign n19511 = n71842 & n19510 ;
  assign n71843 = ~n19006 ;
  assign n19512 = x100 & n71843 ;
  assign n71844 = ~n19004 ;
  assign n19513 = n71844 & n19512 ;
  assign n19514 = n19008 | n19513 ;
  assign n19516 = n19511 | n19514 ;
  assign n71845 = ~n19008 ;
  assign n19517 = n71845 & n19516 ;
  assign n71846 = ~n18997 ;
  assign n19518 = x101 & n71846 ;
  assign n71847 = ~n18995 ;
  assign n19519 = n71847 & n19518 ;
  assign n19520 = n18999 | n19519 ;
  assign n19521 = n19517 | n19520 ;
  assign n71848 = ~n18999 ;
  assign n19522 = n71848 & n19521 ;
  assign n71849 = ~n18988 ;
  assign n19523 = x102 & n71849 ;
  assign n71850 = ~n18986 ;
  assign n19524 = n71850 & n19523 ;
  assign n19525 = n18990 | n19524 ;
  assign n19527 = n19522 | n19525 ;
  assign n71851 = ~n18990 ;
  assign n19528 = n71851 & n19527 ;
  assign n71852 = ~n18979 ;
  assign n19529 = x103 & n71852 ;
  assign n71853 = ~n18977 ;
  assign n19530 = n71853 & n19529 ;
  assign n19531 = n18981 | n19530 ;
  assign n19532 = n19528 | n19531 ;
  assign n71854 = ~n18981 ;
  assign n19533 = n71854 & n19532 ;
  assign n71855 = ~n18970 ;
  assign n19534 = x104 & n71855 ;
  assign n71856 = ~n18968 ;
  assign n19535 = n71856 & n19534 ;
  assign n19536 = n18972 | n19535 ;
  assign n19538 = n19533 | n19536 ;
  assign n71857 = ~n18972 ;
  assign n19539 = n71857 & n19538 ;
  assign n71858 = ~n18961 ;
  assign n19540 = x105 & n71858 ;
  assign n71859 = ~n18959 ;
  assign n19541 = n71859 & n19540 ;
  assign n19542 = n18963 | n19541 ;
  assign n19543 = n19539 | n19542 ;
  assign n71860 = ~n18963 ;
  assign n19544 = n71860 & n19543 ;
  assign n71861 = ~n18952 ;
  assign n19545 = x106 & n71861 ;
  assign n71862 = ~n18950 ;
  assign n19546 = n71862 & n19545 ;
  assign n19547 = n18954 | n19546 ;
  assign n19549 = n19544 | n19547 ;
  assign n71863 = ~n18954 ;
  assign n19550 = n71863 & n19549 ;
  assign n71864 = ~n18943 ;
  assign n19551 = x107 & n71864 ;
  assign n71865 = ~n18941 ;
  assign n19552 = n71865 & n19551 ;
  assign n19553 = n18945 | n19552 ;
  assign n19554 = n19550 | n19553 ;
  assign n71866 = ~n18945 ;
  assign n19555 = n71866 & n19554 ;
  assign n71867 = ~n18934 ;
  assign n19556 = x108 & n71867 ;
  assign n71868 = ~n18932 ;
  assign n19557 = n71868 & n19556 ;
  assign n19558 = n18936 | n19557 ;
  assign n19560 = n19555 | n19558 ;
  assign n71869 = ~n18936 ;
  assign n19561 = n71869 & n19560 ;
  assign n71870 = ~n18925 ;
  assign n19562 = x109 & n71870 ;
  assign n71871 = ~n18923 ;
  assign n19563 = n71871 & n19562 ;
  assign n19564 = n18927 | n19563 ;
  assign n19565 = n19561 | n19564 ;
  assign n71872 = ~n18927 ;
  assign n19566 = n71872 & n19565 ;
  assign n71873 = ~n18916 ;
  assign n19567 = x110 & n71873 ;
  assign n71874 = ~n18914 ;
  assign n19568 = n71874 & n19567 ;
  assign n19569 = n18918 | n19568 ;
  assign n19571 = n19566 | n19569 ;
  assign n71875 = ~n18918 ;
  assign n19572 = n71875 & n19571 ;
  assign n71876 = ~n18908 ;
  assign n19573 = x111 & n71876 ;
  assign n71877 = ~n18906 ;
  assign n19574 = n71877 & n19573 ;
  assign n19575 = n18910 | n19574 ;
  assign n19576 = n19572 | n19575 ;
  assign n71878 = ~n18910 ;
  assign n19577 = n71878 & n19576 ;
  assign n71879 = ~n18898 ;
  assign n19578 = x112 & n71879 ;
  assign n71880 = ~n18896 ;
  assign n19579 = n71880 & n19578 ;
  assign n19580 = n18900 | n19579 ;
  assign n19582 = n19577 | n19580 ;
  assign n71881 = ~n18900 ;
  assign n19583 = n71881 & n19582 ;
  assign n19584 = n279 | n19583 ;
  assign n19585 = n18909 & n19584 ;
  assign n19586 = x65 & n19314 ;
  assign n71882 = ~n19586 ;
  assign n19587 = n19322 & n71882 ;
  assign n19588 = n19324 | n19587 ;
  assign n19589 = n71740 & n19588 ;
  assign n19590 = n19330 | n19589 ;
  assign n19591 = n71743 & n19590 ;
  assign n19592 = n19334 | n19591 ;
  assign n19594 = n71746 & n19592 ;
  assign n19595 = n19295 | n19339 ;
  assign n19597 = n19594 | n19595 ;
  assign n19598 = n71749 & n19597 ;
  assign n19599 = n19343 | n19598 ;
  assign n19601 = n71752 & n19599 ;
  assign n19602 = n19349 | n19601 ;
  assign n19603 = n71755 & n19602 ;
  assign n19604 = n19355 | n19603 ;
  assign n19606 = n71758 & n19604 ;
  assign n19607 = n19360 | n19606 ;
  assign n19608 = n71761 & n19607 ;
  assign n19609 = n19366 | n19608 ;
  assign n19611 = n71764 & n19609 ;
  assign n19612 = n19371 | n19611 ;
  assign n19613 = n71767 & n19612 ;
  assign n19614 = n19377 | n19613 ;
  assign n19616 = n71770 & n19614 ;
  assign n19617 = n19382 | n19616 ;
  assign n19618 = n71773 & n19617 ;
  assign n19619 = n19388 | n19618 ;
  assign n19621 = n71776 & n19619 ;
  assign n19622 = n19393 | n19621 ;
  assign n19623 = n71779 & n19622 ;
  assign n19624 = n19399 | n19623 ;
  assign n19626 = n71782 & n19624 ;
  assign n19627 = n19404 | n19626 ;
  assign n19628 = n71785 & n19627 ;
  assign n19629 = n19410 | n19628 ;
  assign n19631 = n71788 & n19629 ;
  assign n19632 = n19415 | n19631 ;
  assign n19633 = n71791 & n19632 ;
  assign n19634 = n19421 | n19633 ;
  assign n19636 = n71794 & n19634 ;
  assign n19637 = n19426 | n19636 ;
  assign n19638 = n71797 & n19637 ;
  assign n19639 = n19432 | n19638 ;
  assign n19641 = n71800 & n19639 ;
  assign n19642 = n19437 | n19641 ;
  assign n19643 = n71803 & n19642 ;
  assign n19644 = n19443 | n19643 ;
  assign n19646 = n71806 & n19644 ;
  assign n19647 = n19448 | n19646 ;
  assign n19648 = n71809 & n19647 ;
  assign n19649 = n19454 | n19648 ;
  assign n19651 = n71812 & n19649 ;
  assign n19652 = n19459 | n19651 ;
  assign n19653 = n71815 & n19652 ;
  assign n19654 = n19465 | n19653 ;
  assign n19656 = n71818 & n19654 ;
  assign n19657 = n19470 | n19656 ;
  assign n19658 = n71821 & n19657 ;
  assign n19659 = n19476 | n19658 ;
  assign n19661 = n71824 & n19659 ;
  assign n19662 = n19481 | n19661 ;
  assign n19663 = n71827 & n19662 ;
  assign n19664 = n19487 | n19663 ;
  assign n19666 = n71830 & n19664 ;
  assign n19667 = n19492 | n19666 ;
  assign n19668 = n71833 & n19667 ;
  assign n19669 = n19498 | n19668 ;
  assign n19671 = n71836 & n19669 ;
  assign n19672 = n19503 | n19671 ;
  assign n19673 = n71839 & n19672 ;
  assign n19674 = n19509 | n19673 ;
  assign n19676 = n71842 & n19674 ;
  assign n19677 = n19514 | n19676 ;
  assign n19678 = n71845 & n19677 ;
  assign n19679 = n19520 | n19678 ;
  assign n19681 = n71848 & n19679 ;
  assign n19682 = n19525 | n19681 ;
  assign n19683 = n71851 & n19682 ;
  assign n19684 = n19531 | n19683 ;
  assign n19686 = n71854 & n19684 ;
  assign n19687 = n19536 | n19686 ;
  assign n19688 = n71857 & n19687 ;
  assign n19689 = n19542 | n19688 ;
  assign n19691 = n71860 & n19689 ;
  assign n19692 = n19547 | n19691 ;
  assign n19693 = n71863 & n19692 ;
  assign n19694 = n19553 | n19693 ;
  assign n19696 = n71866 & n19694 ;
  assign n19697 = n19558 | n19696 ;
  assign n19698 = n71869 & n19697 ;
  assign n19699 = n19564 | n19698 ;
  assign n19701 = n71872 & n19699 ;
  assign n19702 = n19569 | n19701 ;
  assign n19703 = n71875 & n19702 ;
  assign n71883 = ~n19703 ;
  assign n19704 = n19575 & n71883 ;
  assign n19706 = n18918 | n19575 ;
  assign n71884 = ~n19706 ;
  assign n19707 = n19571 & n71884 ;
  assign n19708 = n19704 | n19707 ;
  assign n19709 = n66715 & n19708 ;
  assign n71885 = ~n19583 ;
  assign n19710 = n71885 & n19709 ;
  assign n19711 = n19585 | n19710 ;
  assign n19712 = n71645 & n19711 ;
  assign n71886 = ~n19710 ;
  assign n20340 = x112 & n71886 ;
  assign n71887 = ~n19585 ;
  assign n20341 = n71887 & n20340 ;
  assign n20342 = n19712 | n20341 ;
  assign n19713 = n18917 & n19584 ;
  assign n71888 = ~n19566 ;
  assign n19570 = n71888 & n19569 ;
  assign n19714 = n18927 | n19569 ;
  assign n71889 = ~n19714 ;
  assign n19715 = n19699 & n71889 ;
  assign n19716 = n19570 | n19715 ;
  assign n19717 = n66715 & n19716 ;
  assign n19718 = n71885 & n19717 ;
  assign n19719 = n19713 | n19718 ;
  assign n19720 = n71633 & n19719 ;
  assign n19721 = n18926 & n19584 ;
  assign n71890 = ~n19698 ;
  assign n19700 = n19564 & n71890 ;
  assign n19722 = n18936 | n19564 ;
  assign n71891 = ~n19722 ;
  assign n19723 = n19560 & n71891 ;
  assign n19724 = n19700 | n19723 ;
  assign n19725 = n66715 & n19724 ;
  assign n19726 = n71885 & n19725 ;
  assign n19727 = n19721 | n19726 ;
  assign n19728 = n71253 & n19727 ;
  assign n71892 = ~n19726 ;
  assign n20329 = x110 & n71892 ;
  assign n71893 = ~n19721 ;
  assign n20330 = n71893 & n20329 ;
  assign n20331 = n19728 | n20330 ;
  assign n19729 = n18935 & n19584 ;
  assign n71894 = ~n19555 ;
  assign n19559 = n71894 & n19558 ;
  assign n19730 = n18945 | n19558 ;
  assign n71895 = ~n19730 ;
  assign n19731 = n19694 & n71895 ;
  assign n19732 = n19559 | n19731 ;
  assign n19733 = n66715 & n19732 ;
  assign n19734 = n71885 & n19733 ;
  assign n19735 = n19729 | n19734 ;
  assign n19736 = n70935 & n19735 ;
  assign n19737 = n18944 & n19584 ;
  assign n71896 = ~n19693 ;
  assign n19695 = n19553 & n71896 ;
  assign n19738 = n18954 | n19553 ;
  assign n71897 = ~n19738 ;
  assign n19739 = n19549 & n71897 ;
  assign n19740 = n19695 | n19739 ;
  assign n19741 = n66715 & n19740 ;
  assign n19742 = n71885 & n19741 ;
  assign n19743 = n19737 | n19742 ;
  assign n19744 = n70927 & n19743 ;
  assign n71898 = ~n19742 ;
  assign n20319 = x108 & n71898 ;
  assign n71899 = ~n19737 ;
  assign n20320 = n71899 & n20319 ;
  assign n20321 = n19744 | n20320 ;
  assign n19745 = n18953 & n19584 ;
  assign n71900 = ~n19544 ;
  assign n19548 = n71900 & n19547 ;
  assign n19746 = n18963 | n19547 ;
  assign n71901 = ~n19746 ;
  assign n19747 = n19689 & n71901 ;
  assign n19748 = n19548 | n19747 ;
  assign n19749 = n66715 & n19748 ;
  assign n19750 = n71885 & n19749 ;
  assign n19751 = n19745 | n19750 ;
  assign n19752 = n70609 & n19751 ;
  assign n19753 = n18962 & n19584 ;
  assign n71902 = ~n19688 ;
  assign n19690 = n19542 & n71902 ;
  assign n19754 = n18972 | n19542 ;
  assign n71903 = ~n19754 ;
  assign n19755 = n19538 & n71903 ;
  assign n19756 = n19690 | n19755 ;
  assign n19757 = n66715 & n19756 ;
  assign n19758 = n71885 & n19757 ;
  assign n19759 = n19753 | n19758 ;
  assign n19760 = n70276 & n19759 ;
  assign n71904 = ~n19758 ;
  assign n20309 = x106 & n71904 ;
  assign n71905 = ~n19753 ;
  assign n20310 = n71905 & n20309 ;
  assign n20311 = n19760 | n20310 ;
  assign n19761 = n18971 & n19584 ;
  assign n71906 = ~n19533 ;
  assign n19537 = n71906 & n19536 ;
  assign n19762 = n18981 | n19536 ;
  assign n71907 = ~n19762 ;
  assign n19763 = n19684 & n71907 ;
  assign n19764 = n19537 | n19763 ;
  assign n19765 = n66715 & n19764 ;
  assign n19766 = n71885 & n19765 ;
  assign n19767 = n19761 | n19766 ;
  assign n19768 = n70176 & n19767 ;
  assign n19769 = n18980 & n19584 ;
  assign n71908 = ~n19683 ;
  assign n19685 = n19531 & n71908 ;
  assign n19770 = n18990 | n19531 ;
  assign n71909 = ~n19770 ;
  assign n19771 = n19527 & n71909 ;
  assign n19772 = n19685 | n19771 ;
  assign n19773 = n66715 & n19772 ;
  assign n19774 = n71885 & n19773 ;
  assign n19775 = n19769 | n19774 ;
  assign n19776 = n69857 & n19775 ;
  assign n71910 = ~n19774 ;
  assign n20299 = x104 & n71910 ;
  assign n71911 = ~n19769 ;
  assign n20300 = n71911 & n20299 ;
  assign n20301 = n19776 | n20300 ;
  assign n19777 = n18989 & n19584 ;
  assign n71912 = ~n19522 ;
  assign n19526 = n71912 & n19525 ;
  assign n19778 = n18999 | n19525 ;
  assign n71913 = ~n19778 ;
  assign n19779 = n19679 & n71913 ;
  assign n19780 = n19526 | n19779 ;
  assign n19781 = n66715 & n19780 ;
  assign n19782 = n71885 & n19781 ;
  assign n19783 = n19777 | n19782 ;
  assign n19784 = n69656 & n19783 ;
  assign n19785 = n18998 & n19584 ;
  assign n71914 = ~n19678 ;
  assign n19680 = n19520 & n71914 ;
  assign n19786 = n19008 | n19520 ;
  assign n71915 = ~n19786 ;
  assign n19787 = n19516 & n71915 ;
  assign n19788 = n19680 | n19787 ;
  assign n19789 = n66715 & n19788 ;
  assign n19790 = n71885 & n19789 ;
  assign n19791 = n19785 | n19790 ;
  assign n19792 = n69528 & n19791 ;
  assign n71916 = ~n19790 ;
  assign n20289 = x102 & n71916 ;
  assign n71917 = ~n19785 ;
  assign n20290 = n71917 & n20289 ;
  assign n20291 = n19792 | n20290 ;
  assign n19793 = n19007 & n19584 ;
  assign n71918 = ~n19511 ;
  assign n19515 = n71918 & n19514 ;
  assign n19794 = n19017 | n19514 ;
  assign n71919 = ~n19794 ;
  assign n19795 = n19674 & n71919 ;
  assign n19796 = n19515 | n19795 ;
  assign n19797 = n66715 & n19796 ;
  assign n19798 = n71885 & n19797 ;
  assign n19799 = n19793 | n19798 ;
  assign n19800 = n69261 & n19799 ;
  assign n19801 = n19016 & n19584 ;
  assign n71920 = ~n19673 ;
  assign n19675 = n19509 & n71920 ;
  assign n19802 = n19026 | n19509 ;
  assign n71921 = ~n19802 ;
  assign n19803 = n19505 & n71921 ;
  assign n19804 = n19675 | n19803 ;
  assign n19805 = n66715 & n19804 ;
  assign n19806 = n71885 & n19805 ;
  assign n19807 = n19801 | n19806 ;
  assign n19808 = n69075 & n19807 ;
  assign n71922 = ~n19806 ;
  assign n20279 = x100 & n71922 ;
  assign n71923 = ~n19801 ;
  assign n20280 = n71923 & n20279 ;
  assign n20281 = n19808 | n20280 ;
  assign n19809 = n19025 & n19584 ;
  assign n71924 = ~n19500 ;
  assign n19504 = n71924 & n19503 ;
  assign n19810 = n19035 | n19503 ;
  assign n71925 = ~n19810 ;
  assign n19811 = n19669 & n71925 ;
  assign n19812 = n19504 | n19811 ;
  assign n19813 = n66715 & n19812 ;
  assign n19814 = n71885 & n19813 ;
  assign n19815 = n19809 | n19814 ;
  assign n19816 = n68993 & n19815 ;
  assign n19817 = n19034 & n19584 ;
  assign n71926 = ~n19668 ;
  assign n19670 = n19498 & n71926 ;
  assign n19818 = n19044 | n19498 ;
  assign n71927 = ~n19818 ;
  assign n19819 = n19494 & n71927 ;
  assign n19820 = n19670 | n19819 ;
  assign n19821 = n66715 & n19820 ;
  assign n19822 = n71885 & n19821 ;
  assign n19823 = n19817 | n19822 ;
  assign n19824 = n68716 & n19823 ;
  assign n71928 = ~n19822 ;
  assign n20269 = x98 & n71928 ;
  assign n71929 = ~n19817 ;
  assign n20270 = n71929 & n20269 ;
  assign n20271 = n19824 | n20270 ;
  assign n19825 = n19043 & n19584 ;
  assign n71930 = ~n19489 ;
  assign n19493 = n71930 & n19492 ;
  assign n19826 = n19053 | n19492 ;
  assign n71931 = ~n19826 ;
  assign n19827 = n19664 & n71931 ;
  assign n19828 = n19493 | n19827 ;
  assign n19829 = n66715 & n19828 ;
  assign n19830 = n71885 & n19829 ;
  assign n19831 = n19825 | n19830 ;
  assign n19832 = n68545 & n19831 ;
  assign n19833 = n19052 & n19584 ;
  assign n71932 = ~n19663 ;
  assign n19665 = n19487 & n71932 ;
  assign n19834 = n19062 | n19487 ;
  assign n71933 = ~n19834 ;
  assign n19835 = n19483 & n71933 ;
  assign n19836 = n19665 | n19835 ;
  assign n19837 = n66715 & n19836 ;
  assign n19838 = n71885 & n19837 ;
  assign n19839 = n19833 | n19838 ;
  assign n19840 = n68438 & n19839 ;
  assign n71934 = ~n19838 ;
  assign n20259 = x96 & n71934 ;
  assign n71935 = ~n19833 ;
  assign n20260 = n71935 & n20259 ;
  assign n20261 = n19840 | n20260 ;
  assign n19841 = n19061 & n19584 ;
  assign n71936 = ~n19478 ;
  assign n19482 = n71936 & n19481 ;
  assign n19842 = n19071 | n19481 ;
  assign n71937 = ~n19842 ;
  assign n19843 = n19659 & n71937 ;
  assign n19844 = n19482 | n19843 ;
  assign n19845 = n66715 & n19844 ;
  assign n19846 = n71885 & n19845 ;
  assign n19847 = n19841 | n19846 ;
  assign n19848 = n68214 & n19847 ;
  assign n19849 = n19070 & n19584 ;
  assign n71938 = ~n19658 ;
  assign n19660 = n19476 & n71938 ;
  assign n19850 = n19080 | n19476 ;
  assign n71939 = ~n19850 ;
  assign n19851 = n19472 & n71939 ;
  assign n19852 = n19660 | n19851 ;
  assign n19853 = n66715 & n19852 ;
  assign n19854 = n71885 & n19853 ;
  assign n19855 = n19849 | n19854 ;
  assign n19856 = n68058 & n19855 ;
  assign n71940 = ~n19854 ;
  assign n20249 = x94 & n71940 ;
  assign n71941 = ~n19849 ;
  assign n20250 = n71941 & n20249 ;
  assign n20251 = n19856 | n20250 ;
  assign n19857 = n19079 & n19584 ;
  assign n71942 = ~n19467 ;
  assign n19471 = n71942 & n19470 ;
  assign n19858 = n19089 | n19470 ;
  assign n71943 = ~n19858 ;
  assign n19859 = n19654 & n71943 ;
  assign n19860 = n19471 | n19859 ;
  assign n19861 = n66715 & n19860 ;
  assign n19862 = n71885 & n19861 ;
  assign n19863 = n19857 | n19862 ;
  assign n19864 = n67986 & n19863 ;
  assign n19865 = n19088 & n19584 ;
  assign n71944 = ~n19653 ;
  assign n19655 = n19465 & n71944 ;
  assign n19866 = n19098 | n19465 ;
  assign n71945 = ~n19866 ;
  assign n19867 = n19461 & n71945 ;
  assign n19868 = n19655 | n19867 ;
  assign n19869 = n66715 & n19868 ;
  assign n19870 = n71885 & n19869 ;
  assign n19871 = n19865 | n19870 ;
  assign n19872 = n67763 & n19871 ;
  assign n71946 = ~n19870 ;
  assign n20239 = x92 & n71946 ;
  assign n71947 = ~n19865 ;
  assign n20240 = n71947 & n20239 ;
  assign n20241 = n19872 | n20240 ;
  assign n19873 = n19097 & n19584 ;
  assign n71948 = ~n19456 ;
  assign n19460 = n71948 & n19459 ;
  assign n19874 = n19107 | n19459 ;
  assign n71949 = ~n19874 ;
  assign n19875 = n19649 & n71949 ;
  assign n19876 = n19460 | n19875 ;
  assign n19877 = n66715 & n19876 ;
  assign n19878 = n71885 & n19877 ;
  assign n19879 = n19873 | n19878 ;
  assign n19880 = n67622 & n19879 ;
  assign n19881 = n19106 & n19584 ;
  assign n71950 = ~n19648 ;
  assign n19650 = n19454 & n71950 ;
  assign n19882 = n19116 | n19454 ;
  assign n71951 = ~n19882 ;
  assign n19883 = n19450 & n71951 ;
  assign n19884 = n19650 | n19883 ;
  assign n19885 = n66715 & n19884 ;
  assign n19886 = n71885 & n19885 ;
  assign n19887 = n19881 | n19886 ;
  assign n19888 = n67531 & n19887 ;
  assign n71952 = ~n19886 ;
  assign n20229 = x90 & n71952 ;
  assign n71953 = ~n19881 ;
  assign n20230 = n71953 & n20229 ;
  assign n20231 = n19888 | n20230 ;
  assign n19889 = n19115 & n19584 ;
  assign n71954 = ~n19445 ;
  assign n19449 = n71954 & n19448 ;
  assign n19890 = n19125 | n19448 ;
  assign n71955 = ~n19890 ;
  assign n19891 = n19644 & n71955 ;
  assign n19892 = n19449 | n19891 ;
  assign n19893 = n66715 & n19892 ;
  assign n19894 = n71885 & n19893 ;
  assign n19895 = n19889 | n19894 ;
  assign n19896 = n67348 & n19895 ;
  assign n19897 = n19124 & n19584 ;
  assign n71956 = ~n19643 ;
  assign n19645 = n19443 & n71956 ;
  assign n19898 = n19133 | n19443 ;
  assign n71957 = ~n19898 ;
  assign n19899 = n19439 & n71957 ;
  assign n19900 = n19645 | n19899 ;
  assign n19901 = n66715 & n19900 ;
  assign n19902 = n71885 & n19901 ;
  assign n19903 = n19897 | n19902 ;
  assign n19904 = n67222 & n19903 ;
  assign n71958 = ~n19902 ;
  assign n20219 = x88 & n71958 ;
  assign n71959 = ~n19897 ;
  assign n20220 = n71959 & n20219 ;
  assign n20221 = n19904 | n20220 ;
  assign n19905 = n19132 & n19584 ;
  assign n71960 = ~n19434 ;
  assign n19438 = n71960 & n19437 ;
  assign n19906 = n19142 | n19437 ;
  assign n71961 = ~n19906 ;
  assign n19907 = n19639 & n71961 ;
  assign n19908 = n19438 | n19907 ;
  assign n19909 = n66715 & n19908 ;
  assign n19910 = n71885 & n19909 ;
  assign n19911 = n19905 | n19910 ;
  assign n19912 = n67164 & n19911 ;
  assign n19913 = n19141 & n19584 ;
  assign n71962 = ~n19638 ;
  assign n19640 = n19432 & n71962 ;
  assign n19914 = n19151 | n19432 ;
  assign n71963 = ~n19914 ;
  assign n19915 = n19428 & n71963 ;
  assign n19916 = n19640 | n19915 ;
  assign n19917 = n66715 & n19916 ;
  assign n19918 = n71885 & n19917 ;
  assign n19919 = n19913 | n19918 ;
  assign n19920 = n66979 & n19919 ;
  assign n71964 = ~n19918 ;
  assign n20208 = x86 & n71964 ;
  assign n71965 = ~n19913 ;
  assign n20209 = n71965 & n20208 ;
  assign n20210 = n19920 | n20209 ;
  assign n19921 = n19150 & n19584 ;
  assign n71966 = ~n19423 ;
  assign n19427 = n71966 & n19426 ;
  assign n19922 = n19160 | n19426 ;
  assign n71967 = ~n19922 ;
  assign n19923 = n19634 & n71967 ;
  assign n19924 = n19427 | n19923 ;
  assign n19925 = n66715 & n19924 ;
  assign n19926 = n71885 & n19925 ;
  assign n19927 = n19921 | n19926 ;
  assign n19928 = n66868 & n19927 ;
  assign n19929 = n19159 & n19584 ;
  assign n71968 = ~n19633 ;
  assign n19635 = n19421 & n71968 ;
  assign n19930 = n19169 | n19421 ;
  assign n71969 = ~n19930 ;
  assign n19931 = n19417 & n71969 ;
  assign n19932 = n19635 | n19931 ;
  assign n19933 = n66715 & n19932 ;
  assign n19934 = n71885 & n19933 ;
  assign n19935 = n19929 | n19934 ;
  assign n19936 = n66797 & n19935 ;
  assign n71970 = ~n19934 ;
  assign n20198 = x84 & n71970 ;
  assign n71971 = ~n19929 ;
  assign n20199 = n71971 & n20198 ;
  assign n20200 = n19936 | n20199 ;
  assign n19937 = n19168 & n19584 ;
  assign n71972 = ~n19412 ;
  assign n19416 = n71972 & n19415 ;
  assign n19938 = n19178 | n19415 ;
  assign n71973 = ~n19938 ;
  assign n19939 = n19629 & n71973 ;
  assign n19940 = n19416 | n19939 ;
  assign n19941 = n66715 & n19940 ;
  assign n19942 = n71885 & n19941 ;
  assign n19943 = n19937 | n19942 ;
  assign n19944 = n66654 & n19943 ;
  assign n19945 = n19177 & n19584 ;
  assign n71974 = ~n19628 ;
  assign n19630 = n19410 & n71974 ;
  assign n19946 = n19187 | n19410 ;
  assign n71975 = ~n19946 ;
  assign n19947 = n19406 & n71975 ;
  assign n19948 = n19630 | n19947 ;
  assign n19949 = n66715 & n19948 ;
  assign n19950 = n71885 & n19949 ;
  assign n19951 = n19945 | n19950 ;
  assign n19952 = n66560 & n19951 ;
  assign n71976 = ~n19950 ;
  assign n20187 = x82 & n71976 ;
  assign n71977 = ~n19945 ;
  assign n20188 = n71977 & n20187 ;
  assign n20189 = n19952 | n20188 ;
  assign n19953 = n19186 & n19584 ;
  assign n71978 = ~n19401 ;
  assign n19405 = n71978 & n19404 ;
  assign n19954 = n19196 | n19404 ;
  assign n71979 = ~n19954 ;
  assign n19955 = n19624 & n71979 ;
  assign n19956 = n19405 | n19955 ;
  assign n19957 = n66715 & n19956 ;
  assign n19958 = n71885 & n19957 ;
  assign n19959 = n19953 | n19958 ;
  assign n19960 = n66505 & n19959 ;
  assign n19961 = n19195 & n19584 ;
  assign n71980 = ~n19623 ;
  assign n19625 = n19399 & n71980 ;
  assign n19962 = n19205 | n19399 ;
  assign n71981 = ~n19962 ;
  assign n19963 = n19395 & n71981 ;
  assign n19964 = n19625 | n19963 ;
  assign n19965 = n66715 & n19964 ;
  assign n19966 = n71885 & n19965 ;
  assign n19967 = n19961 | n19966 ;
  assign n19968 = n66379 & n19967 ;
  assign n71982 = ~n19966 ;
  assign n20176 = x80 & n71982 ;
  assign n71983 = ~n19961 ;
  assign n20177 = n71983 & n20176 ;
  assign n20178 = n19968 | n20177 ;
  assign n19969 = n19204 & n19584 ;
  assign n71984 = ~n19390 ;
  assign n19394 = n71984 & n19393 ;
  assign n19970 = n19214 | n19393 ;
  assign n71985 = ~n19970 ;
  assign n19971 = n19619 & n71985 ;
  assign n19972 = n19394 | n19971 ;
  assign n19973 = n66715 & n19972 ;
  assign n19974 = n71885 & n19973 ;
  assign n19975 = n19969 | n19974 ;
  assign n19976 = n66299 & n19975 ;
  assign n19977 = n19213 & n19584 ;
  assign n71986 = ~n19618 ;
  assign n19620 = n19388 & n71986 ;
  assign n19978 = n19223 | n19388 ;
  assign n71987 = ~n19978 ;
  assign n19979 = n19384 & n71987 ;
  assign n19980 = n19620 | n19979 ;
  assign n19981 = n66715 & n19980 ;
  assign n19982 = n71885 & n19981 ;
  assign n19983 = n19977 | n19982 ;
  assign n19984 = n66244 & n19983 ;
  assign n71988 = ~n19982 ;
  assign n20166 = x78 & n71988 ;
  assign n71989 = ~n19977 ;
  assign n20167 = n71989 & n20166 ;
  assign n20168 = n19984 | n20167 ;
  assign n19985 = n19222 & n19584 ;
  assign n71990 = ~n19379 ;
  assign n19383 = n71990 & n19382 ;
  assign n19986 = n19232 | n19382 ;
  assign n71991 = ~n19986 ;
  assign n19987 = n19614 & n71991 ;
  assign n19988 = n19383 | n19987 ;
  assign n19989 = n66715 & n19988 ;
  assign n19990 = n71885 & n19989 ;
  assign n19991 = n19985 | n19990 ;
  assign n19992 = n66145 & n19991 ;
  assign n19993 = n19231 & n19584 ;
  assign n71992 = ~n19613 ;
  assign n19615 = n19377 & n71992 ;
  assign n19994 = n19241 | n19377 ;
  assign n71993 = ~n19994 ;
  assign n19995 = n19373 & n71993 ;
  assign n19996 = n19615 | n19995 ;
  assign n19997 = n66715 & n19996 ;
  assign n19998 = n71885 & n19997 ;
  assign n19999 = n19993 | n19998 ;
  assign n20000 = n66081 & n19999 ;
  assign n71994 = ~n19998 ;
  assign n20156 = x76 & n71994 ;
  assign n71995 = ~n19993 ;
  assign n20157 = n71995 & n20156 ;
  assign n20158 = n20000 | n20157 ;
  assign n20001 = n19240 & n19584 ;
  assign n71996 = ~n19368 ;
  assign n19372 = n71996 & n19371 ;
  assign n20002 = n19250 | n19371 ;
  assign n71997 = ~n20002 ;
  assign n20003 = n19609 & n71997 ;
  assign n20004 = n19372 | n20003 ;
  assign n20005 = n66715 & n20004 ;
  assign n20006 = n71885 & n20005 ;
  assign n20007 = n20001 | n20006 ;
  assign n20008 = n66043 & n20007 ;
  assign n20009 = n19249 & n19584 ;
  assign n71998 = ~n19608 ;
  assign n19610 = n19366 & n71998 ;
  assign n20010 = n19259 | n19366 ;
  assign n71999 = ~n20010 ;
  assign n20011 = n19362 & n71999 ;
  assign n20012 = n19610 | n20011 ;
  assign n20013 = n66715 & n20012 ;
  assign n20014 = n71885 & n20013 ;
  assign n20015 = n20009 | n20014 ;
  assign n20016 = n65960 & n20015 ;
  assign n72000 = ~n20014 ;
  assign n20146 = x74 & n72000 ;
  assign n72001 = ~n20009 ;
  assign n20147 = n72001 & n20146 ;
  assign n20148 = n20016 | n20147 ;
  assign n20017 = n19258 & n19584 ;
  assign n72002 = ~n19357 ;
  assign n19361 = n72002 & n19360 ;
  assign n20018 = n19268 | n19360 ;
  assign n72003 = ~n20018 ;
  assign n20019 = n19604 & n72003 ;
  assign n20020 = n19361 | n20019 ;
  assign n20021 = n66715 & n20020 ;
  assign n20022 = n71885 & n20021 ;
  assign n20023 = n20017 | n20022 ;
  assign n20024 = n65909 & n20023 ;
  assign n20025 = n19267 & n19584 ;
  assign n72004 = ~n19603 ;
  assign n19605 = n19355 & n72004 ;
  assign n20026 = n19277 | n19355 ;
  assign n72005 = ~n20026 ;
  assign n20027 = n19351 & n72005 ;
  assign n20028 = n19605 | n20027 ;
  assign n20029 = n66715 & n20028 ;
  assign n20030 = n71885 & n20029 ;
  assign n20031 = n20025 | n20030 ;
  assign n20032 = n65877 & n20031 ;
  assign n72006 = ~n20030 ;
  assign n20136 = x72 & n72006 ;
  assign n72007 = ~n20025 ;
  assign n20137 = n72007 & n20136 ;
  assign n20138 = n20032 | n20137 ;
  assign n20033 = n19276 & n19584 ;
  assign n72008 = ~n19346 ;
  assign n19350 = n72008 & n19349 ;
  assign n20034 = n19344 | n19598 ;
  assign n20035 = n19286 | n19349 ;
  assign n72009 = ~n20035 ;
  assign n20036 = n20034 & n72009 ;
  assign n20037 = n19350 | n20036 ;
  assign n20038 = n66715 & n20037 ;
  assign n20039 = n71885 & n20038 ;
  assign n20040 = n20033 | n20039 ;
  assign n20041 = n65820 & n20040 ;
  assign n20042 = n19285 & n19584 ;
  assign n72010 = ~n19598 ;
  assign n19600 = n19344 & n72010 ;
  assign n20043 = n19337 | n19595 ;
  assign n20044 = n19295 | n19344 ;
  assign n72011 = ~n20044 ;
  assign n20045 = n20043 & n72011 ;
  assign n20046 = n19600 | n20045 ;
  assign n20047 = n66715 & n20046 ;
  assign n20048 = n71885 & n20047 ;
  assign n20049 = n20042 | n20048 ;
  assign n20050 = n65791 & n20049 ;
  assign n72012 = ~n20048 ;
  assign n20125 = x70 & n72012 ;
  assign n72013 = ~n20042 ;
  assign n20126 = n72013 & n20125 ;
  assign n20127 = n20050 | n20126 ;
  assign n20051 = n19294 & n19584 ;
  assign n72014 = ~n19337 ;
  assign n19596 = n72014 & n19595 ;
  assign n20052 = n19335 | n19591 ;
  assign n20053 = n19303 | n19595 ;
  assign n72015 = ~n20053 ;
  assign n20054 = n20052 & n72015 ;
  assign n20055 = n19596 | n20054 ;
  assign n20056 = n66715 & n20055 ;
  assign n20057 = n71885 & n20056 ;
  assign n20058 = n20051 | n20057 ;
  assign n20059 = n65772 & n20058 ;
  assign n20060 = n19302 & n19584 ;
  assign n72016 = ~n19591 ;
  assign n19593 = n19335 & n72016 ;
  assign n20061 = n19311 | n19335 ;
  assign n72017 = ~n20061 ;
  assign n20062 = n19590 & n72017 ;
  assign n20063 = n19593 | n20062 ;
  assign n20064 = n66715 & n20063 ;
  assign n20065 = n71885 & n20064 ;
  assign n20066 = n20060 | n20065 ;
  assign n20067 = n65746 & n20066 ;
  assign n72018 = ~n20065 ;
  assign n20115 = x68 & n72018 ;
  assign n72019 = ~n20060 ;
  assign n20116 = n72019 & n20115 ;
  assign n20117 = n20067 | n20116 ;
  assign n20068 = n19310 & n19584 ;
  assign n20069 = n19325 | n19330 ;
  assign n72020 = ~n20069 ;
  assign n20070 = n19588 & n72020 ;
  assign n72021 = ~n19327 ;
  assign n20071 = n72021 & n19330 ;
  assign n20072 = n20070 | n20071 ;
  assign n20073 = n66715 & n20072 ;
  assign n20074 = n71885 & n20073 ;
  assign n20075 = n20068 | n20074 ;
  assign n20076 = n65721 & n20075 ;
  assign n20077 = n19319 & n19584 ;
  assign n20078 = n19322 & n19324 ;
  assign n20079 = n71882 & n20078 ;
  assign n20080 = n279 | n20079 ;
  assign n72022 = ~n20080 ;
  assign n20081 = n19588 & n72022 ;
  assign n20082 = n71885 & n20081 ;
  assign n20083 = n20077 | n20082 ;
  assign n20084 = n65686 & n20083 ;
  assign n72023 = ~n20082 ;
  assign n20105 = x66 & n72023 ;
  assign n72024 = ~n20077 ;
  assign n20106 = n72024 & n20105 ;
  assign n20107 = n20084 | n20106 ;
  assign n19705 = n19575 | n19703 ;
  assign n20085 = n71878 & n19705 ;
  assign n20086 = n19580 | n20085 ;
  assign n20087 = n71881 & n20086 ;
  assign n72025 = ~x113 ;
  assign n20088 = x64 & n72025 ;
  assign n72026 = ~n65497 ;
  assign n20089 = n72026 & n20088 ;
  assign n72027 = ~n65414 ;
  assign n20090 = n72027 & n20089 ;
  assign n20091 = n65681 & n20090 ;
  assign n72028 = ~n20087 ;
  assign n20092 = n72028 & n20091 ;
  assign n72029 = ~n20092 ;
  assign n20093 = x15 & n72029 ;
  assign n20094 = n71255 & n19324 ;
  assign n20095 = n67026 & n20094 ;
  assign n20096 = n71885 & n20095 ;
  assign n20097 = n20093 | n20096 ;
  assign n20098 = x65 & n20097 ;
  assign n20099 = x65 | n20096 ;
  assign n20100 = n20093 | n20099 ;
  assign n72030 = ~n20098 ;
  assign n20101 = n72030 & n20100 ;
  assign n72031 = ~x14 ;
  assign n20102 = n72031 & x64 ;
  assign n20103 = n20101 | n20102 ;
  assign n20104 = n65670 & n20097 ;
  assign n72032 = ~n20104 ;
  assign n20108 = n20103 & n72032 ;
  assign n20109 = n20107 | n20108 ;
  assign n72033 = ~n20084 ;
  assign n20110 = n72033 & n20109 ;
  assign n72034 = ~n20074 ;
  assign n20111 = x67 & n72034 ;
  assign n72035 = ~n20068 ;
  assign n20112 = n72035 & n20111 ;
  assign n20113 = n20076 | n20112 ;
  assign n20114 = n20110 | n20113 ;
  assign n72036 = ~n20076 ;
  assign n20118 = n72036 & n20114 ;
  assign n20119 = n20117 | n20118 ;
  assign n72037 = ~n20067 ;
  assign n20120 = n72037 & n20119 ;
  assign n72038 = ~n20057 ;
  assign n20121 = x69 & n72038 ;
  assign n72039 = ~n20051 ;
  assign n20122 = n72039 & n20121 ;
  assign n20123 = n20059 | n20122 ;
  assign n20124 = n20120 | n20123 ;
  assign n72040 = ~n20059 ;
  assign n20128 = n72040 & n20124 ;
  assign n20129 = n20127 | n20128 ;
  assign n72041 = ~n20050 ;
  assign n20130 = n72041 & n20129 ;
  assign n72042 = ~n20039 ;
  assign n20131 = x71 & n72042 ;
  assign n72043 = ~n20033 ;
  assign n20132 = n72043 & n20131 ;
  assign n20133 = n20041 | n20132 ;
  assign n20135 = n20130 | n20133 ;
  assign n72044 = ~n20041 ;
  assign n20139 = n72044 & n20135 ;
  assign n20140 = n20138 | n20139 ;
  assign n72045 = ~n20032 ;
  assign n20141 = n72045 & n20140 ;
  assign n72046 = ~n20022 ;
  assign n20142 = x73 & n72046 ;
  assign n72047 = ~n20017 ;
  assign n20143 = n72047 & n20142 ;
  assign n20144 = n20024 | n20143 ;
  assign n20145 = n20141 | n20144 ;
  assign n72048 = ~n20024 ;
  assign n20149 = n72048 & n20145 ;
  assign n20150 = n20148 | n20149 ;
  assign n72049 = ~n20016 ;
  assign n20151 = n72049 & n20150 ;
  assign n72050 = ~n20006 ;
  assign n20152 = x75 & n72050 ;
  assign n72051 = ~n20001 ;
  assign n20153 = n72051 & n20152 ;
  assign n20154 = n20008 | n20153 ;
  assign n20155 = n20151 | n20154 ;
  assign n72052 = ~n20008 ;
  assign n20159 = n72052 & n20155 ;
  assign n20160 = n20158 | n20159 ;
  assign n72053 = ~n20000 ;
  assign n20161 = n72053 & n20160 ;
  assign n72054 = ~n19990 ;
  assign n20162 = x77 & n72054 ;
  assign n72055 = ~n19985 ;
  assign n20163 = n72055 & n20162 ;
  assign n20164 = n19992 | n20163 ;
  assign n20165 = n20161 | n20164 ;
  assign n72056 = ~n19992 ;
  assign n20169 = n72056 & n20165 ;
  assign n20170 = n20168 | n20169 ;
  assign n72057 = ~n19984 ;
  assign n20171 = n72057 & n20170 ;
  assign n72058 = ~n19974 ;
  assign n20172 = x79 & n72058 ;
  assign n72059 = ~n19969 ;
  assign n20173 = n72059 & n20172 ;
  assign n20174 = n19976 | n20173 ;
  assign n20175 = n20171 | n20174 ;
  assign n72060 = ~n19976 ;
  assign n20180 = n72060 & n20175 ;
  assign n20181 = n20178 | n20180 ;
  assign n72061 = ~n19968 ;
  assign n20182 = n72061 & n20181 ;
  assign n72062 = ~n19958 ;
  assign n20183 = x81 & n72062 ;
  assign n72063 = ~n19953 ;
  assign n20184 = n72063 & n20183 ;
  assign n20185 = n19960 | n20184 ;
  assign n20186 = n20182 | n20185 ;
  assign n72064 = ~n19960 ;
  assign n20191 = n72064 & n20186 ;
  assign n20192 = n20189 | n20191 ;
  assign n72065 = ~n19952 ;
  assign n20193 = n72065 & n20192 ;
  assign n72066 = ~n19942 ;
  assign n20194 = x83 & n72066 ;
  assign n72067 = ~n19937 ;
  assign n20195 = n72067 & n20194 ;
  assign n20196 = n19944 | n20195 ;
  assign n20197 = n20193 | n20196 ;
  assign n72068 = ~n19944 ;
  assign n20201 = n72068 & n20197 ;
  assign n20202 = n20200 | n20201 ;
  assign n72069 = ~n19936 ;
  assign n20203 = n72069 & n20202 ;
  assign n72070 = ~n19926 ;
  assign n20204 = x85 & n72070 ;
  assign n72071 = ~n19921 ;
  assign n20205 = n72071 & n20204 ;
  assign n20206 = n19928 | n20205 ;
  assign n20207 = n20203 | n20206 ;
  assign n72072 = ~n19928 ;
  assign n20212 = n72072 & n20207 ;
  assign n20213 = n20210 | n20212 ;
  assign n72073 = ~n19920 ;
  assign n20214 = n72073 & n20213 ;
  assign n72074 = ~n19910 ;
  assign n20215 = x87 & n72074 ;
  assign n72075 = ~n19905 ;
  assign n20216 = n72075 & n20215 ;
  assign n20217 = n19912 | n20216 ;
  assign n20218 = n20214 | n20217 ;
  assign n72076 = ~n19912 ;
  assign n20222 = n72076 & n20218 ;
  assign n20223 = n20221 | n20222 ;
  assign n72077 = ~n19904 ;
  assign n20224 = n72077 & n20223 ;
  assign n72078 = ~n19894 ;
  assign n20225 = x89 & n72078 ;
  assign n72079 = ~n19889 ;
  assign n20226 = n72079 & n20225 ;
  assign n20227 = n19896 | n20226 ;
  assign n20228 = n20224 | n20227 ;
  assign n72080 = ~n19896 ;
  assign n20232 = n72080 & n20228 ;
  assign n20233 = n20231 | n20232 ;
  assign n72081 = ~n19888 ;
  assign n20234 = n72081 & n20233 ;
  assign n72082 = ~n19878 ;
  assign n20235 = x91 & n72082 ;
  assign n72083 = ~n19873 ;
  assign n20236 = n72083 & n20235 ;
  assign n20237 = n19880 | n20236 ;
  assign n20238 = n20234 | n20237 ;
  assign n72084 = ~n19880 ;
  assign n20242 = n72084 & n20238 ;
  assign n20243 = n20241 | n20242 ;
  assign n72085 = ~n19872 ;
  assign n20244 = n72085 & n20243 ;
  assign n72086 = ~n19862 ;
  assign n20245 = x93 & n72086 ;
  assign n72087 = ~n19857 ;
  assign n20246 = n72087 & n20245 ;
  assign n20247 = n19864 | n20246 ;
  assign n20248 = n20244 | n20247 ;
  assign n72088 = ~n19864 ;
  assign n20252 = n72088 & n20248 ;
  assign n20253 = n20251 | n20252 ;
  assign n72089 = ~n19856 ;
  assign n20254 = n72089 & n20253 ;
  assign n72090 = ~n19846 ;
  assign n20255 = x95 & n72090 ;
  assign n72091 = ~n19841 ;
  assign n20256 = n72091 & n20255 ;
  assign n20257 = n19848 | n20256 ;
  assign n20258 = n20254 | n20257 ;
  assign n72092 = ~n19848 ;
  assign n20262 = n72092 & n20258 ;
  assign n20263 = n20261 | n20262 ;
  assign n72093 = ~n19840 ;
  assign n20264 = n72093 & n20263 ;
  assign n72094 = ~n19830 ;
  assign n20265 = x97 & n72094 ;
  assign n72095 = ~n19825 ;
  assign n20266 = n72095 & n20265 ;
  assign n20267 = n19832 | n20266 ;
  assign n20268 = n20264 | n20267 ;
  assign n72096 = ~n19832 ;
  assign n20272 = n72096 & n20268 ;
  assign n20273 = n20271 | n20272 ;
  assign n72097 = ~n19824 ;
  assign n20274 = n72097 & n20273 ;
  assign n72098 = ~n19814 ;
  assign n20275 = x99 & n72098 ;
  assign n72099 = ~n19809 ;
  assign n20276 = n72099 & n20275 ;
  assign n20277 = n19816 | n20276 ;
  assign n20278 = n20274 | n20277 ;
  assign n72100 = ~n19816 ;
  assign n20282 = n72100 & n20278 ;
  assign n20283 = n20281 | n20282 ;
  assign n72101 = ~n19808 ;
  assign n20284 = n72101 & n20283 ;
  assign n72102 = ~n19798 ;
  assign n20285 = x101 & n72102 ;
  assign n72103 = ~n19793 ;
  assign n20286 = n72103 & n20285 ;
  assign n20287 = n19800 | n20286 ;
  assign n20288 = n20284 | n20287 ;
  assign n72104 = ~n19800 ;
  assign n20292 = n72104 & n20288 ;
  assign n20293 = n20291 | n20292 ;
  assign n72105 = ~n19792 ;
  assign n20294 = n72105 & n20293 ;
  assign n72106 = ~n19782 ;
  assign n20295 = x103 & n72106 ;
  assign n72107 = ~n19777 ;
  assign n20296 = n72107 & n20295 ;
  assign n20297 = n19784 | n20296 ;
  assign n20298 = n20294 | n20297 ;
  assign n72108 = ~n19784 ;
  assign n20302 = n72108 & n20298 ;
  assign n20303 = n20301 | n20302 ;
  assign n72109 = ~n19776 ;
  assign n20304 = n72109 & n20303 ;
  assign n72110 = ~n19766 ;
  assign n20305 = x105 & n72110 ;
  assign n72111 = ~n19761 ;
  assign n20306 = n72111 & n20305 ;
  assign n20307 = n19768 | n20306 ;
  assign n20308 = n20304 | n20307 ;
  assign n72112 = ~n19768 ;
  assign n20312 = n72112 & n20308 ;
  assign n20313 = n20311 | n20312 ;
  assign n72113 = ~n19760 ;
  assign n20314 = n72113 & n20313 ;
  assign n72114 = ~n19750 ;
  assign n20315 = x107 & n72114 ;
  assign n72115 = ~n19745 ;
  assign n20316 = n72115 & n20315 ;
  assign n20317 = n19752 | n20316 ;
  assign n20318 = n20314 | n20317 ;
  assign n72116 = ~n19752 ;
  assign n20322 = n72116 & n20318 ;
  assign n20323 = n20321 | n20322 ;
  assign n72117 = ~n19744 ;
  assign n20324 = n72117 & n20323 ;
  assign n72118 = ~n19734 ;
  assign n20325 = x109 & n72118 ;
  assign n72119 = ~n19729 ;
  assign n20326 = n72119 & n20325 ;
  assign n20327 = n19736 | n20326 ;
  assign n20328 = n20324 | n20327 ;
  assign n72120 = ~n19736 ;
  assign n20332 = n72120 & n20328 ;
  assign n20333 = n20331 | n20332 ;
  assign n72121 = ~n19728 ;
  assign n20334 = n72121 & n20333 ;
  assign n72122 = ~n19718 ;
  assign n20335 = x111 & n72122 ;
  assign n72123 = ~n19713 ;
  assign n20336 = n72123 & n20335 ;
  assign n20337 = n19720 | n20336 ;
  assign n20339 = n20334 | n20337 ;
  assign n72124 = ~n19720 ;
  assign n20343 = n72124 & n20339 ;
  assign n20344 = n20342 | n20343 ;
  assign n72125 = ~n19712 ;
  assign n20345 = n72125 & n20344 ;
  assign n72126 = ~n19577 ;
  assign n19581 = n72126 & n19580 ;
  assign n20346 = n18910 | n19580 ;
  assign n72127 = ~n20346 ;
  assign n20347 = n19705 & n72127 ;
  assign n20348 = n19581 | n20347 ;
  assign n20349 = n19584 | n20348 ;
  assign n72128 = ~n18899 ;
  assign n20350 = n72128 & n19584 ;
  assign n72129 = ~n20350 ;
  assign n20351 = n20349 & n72129 ;
  assign n20352 = n72025 & n20351 ;
  assign n144 = ~n19584 ;
  assign n20353 = n144 & n20348 ;
  assign n20354 = n18899 & n19584 ;
  assign n72131 = ~n20354 ;
  assign n20355 = x113 & n72131 ;
  assign n72132 = ~n20353 ;
  assign n20356 = n72132 & n20355 ;
  assign n20359 = n20356 | n20358 ;
  assign n20360 = n20352 | n20359 ;
  assign n20361 = n20345 | n20360 ;
  assign n20362 = n66715 & n20351 ;
  assign n72133 = ~n20362 ;
  assign n20363 = n20361 & n72133 ;
  assign n21170 = n19712 | n20356 ;
  assign n21171 = n20352 | n21170 ;
  assign n72134 = ~n21171 ;
  assign n21172 = n20344 & n72134 ;
  assign n20365 = n71885 & n20091 ;
  assign n72135 = ~n20365 ;
  assign n20366 = x15 & n72135 ;
  assign n20367 = n20096 | n20366 ;
  assign n20368 = x65 & n20367 ;
  assign n72136 = ~n20368 ;
  assign n20369 = n20100 & n72136 ;
  assign n20370 = n20102 | n20369 ;
  assign n20371 = n72032 & n20370 ;
  assign n20372 = n20107 | n20371 ;
  assign n20373 = n72033 & n20372 ;
  assign n20374 = n20113 | n20373 ;
  assign n20375 = n72036 & n20374 ;
  assign n20376 = n20117 | n20375 ;
  assign n20377 = n72037 & n20376 ;
  assign n20378 = n20123 | n20377 ;
  assign n20379 = n72040 & n20378 ;
  assign n20380 = n20127 | n20379 ;
  assign n20381 = n72041 & n20380 ;
  assign n20382 = n20133 | n20381 ;
  assign n20383 = n72044 & n20382 ;
  assign n20384 = n20138 | n20383 ;
  assign n20385 = n72045 & n20384 ;
  assign n20386 = n20144 | n20385 ;
  assign n20387 = n72048 & n20386 ;
  assign n20388 = n20148 | n20387 ;
  assign n20389 = n72049 & n20388 ;
  assign n20390 = n20154 | n20389 ;
  assign n20391 = n72052 & n20390 ;
  assign n20392 = n20158 | n20391 ;
  assign n20393 = n72053 & n20392 ;
  assign n20394 = n20164 | n20393 ;
  assign n20395 = n72056 & n20394 ;
  assign n20396 = n20168 | n20395 ;
  assign n20397 = n72057 & n20396 ;
  assign n20398 = n20174 | n20397 ;
  assign n20399 = n72060 & n20398 ;
  assign n20400 = n20178 | n20399 ;
  assign n20401 = n72061 & n20400 ;
  assign n20402 = n20185 | n20401 ;
  assign n20403 = n72064 & n20402 ;
  assign n20404 = n20189 | n20403 ;
  assign n20405 = n72065 & n20404 ;
  assign n20406 = n20196 | n20405 ;
  assign n20407 = n72068 & n20406 ;
  assign n20408 = n20200 | n20407 ;
  assign n20409 = n72069 & n20408 ;
  assign n20410 = n20206 | n20409 ;
  assign n20411 = n72072 & n20410 ;
  assign n20412 = n20210 | n20411 ;
  assign n20413 = n72073 & n20412 ;
  assign n20414 = n20217 | n20413 ;
  assign n20415 = n72076 & n20414 ;
  assign n20416 = n20221 | n20415 ;
  assign n20417 = n72077 & n20416 ;
  assign n20418 = n20227 | n20417 ;
  assign n20419 = n72080 & n20418 ;
  assign n20420 = n20231 | n20419 ;
  assign n20421 = n72081 & n20420 ;
  assign n20422 = n20237 | n20421 ;
  assign n20423 = n72084 & n20422 ;
  assign n20424 = n20241 | n20423 ;
  assign n20425 = n72085 & n20424 ;
  assign n20426 = n20247 | n20425 ;
  assign n20427 = n72088 & n20426 ;
  assign n20428 = n20251 | n20427 ;
  assign n20429 = n72089 & n20428 ;
  assign n20430 = n20257 | n20429 ;
  assign n20431 = n72092 & n20430 ;
  assign n20432 = n20261 | n20431 ;
  assign n20433 = n72093 & n20432 ;
  assign n20434 = n20267 | n20433 ;
  assign n20435 = n72096 & n20434 ;
  assign n20436 = n20271 | n20435 ;
  assign n20437 = n72097 & n20436 ;
  assign n20438 = n20277 | n20437 ;
  assign n20439 = n72100 & n20438 ;
  assign n20440 = n20281 | n20439 ;
  assign n20441 = n72101 & n20440 ;
  assign n20442 = n20287 | n20441 ;
  assign n20443 = n72104 & n20442 ;
  assign n20444 = n20291 | n20443 ;
  assign n20445 = n72105 & n20444 ;
  assign n20446 = n20297 | n20445 ;
  assign n20447 = n72108 & n20446 ;
  assign n20448 = n20301 | n20447 ;
  assign n20449 = n72109 & n20448 ;
  assign n20450 = n20307 | n20449 ;
  assign n20451 = n72112 & n20450 ;
  assign n20452 = n20311 | n20451 ;
  assign n20453 = n72113 & n20452 ;
  assign n20454 = n20317 | n20453 ;
  assign n20455 = n72116 & n20454 ;
  assign n20456 = n20321 | n20455 ;
  assign n20457 = n72117 & n20456 ;
  assign n20458 = n20327 | n20457 ;
  assign n20459 = n72120 & n20458 ;
  assign n20460 = n20331 | n20459 ;
  assign n20461 = n72121 & n20460 ;
  assign n20462 = n20337 | n20461 ;
  assign n20463 = n72124 & n20462 ;
  assign n20890 = n20342 | n20463 ;
  assign n20891 = n72125 & n20890 ;
  assign n21173 = n20352 | n20356 ;
  assign n72137 = ~n20891 ;
  assign n21174 = n72137 & n21173 ;
  assign n21175 = n21172 | n21174 ;
  assign n143 = ~n20363 ;
  assign n21176 = n143 & n21175 ;
  assign n21177 = n279 & n18899 ;
  assign n21178 = n20361 & n21177 ;
  assign n21179 = n21176 | n21178 ;
  assign n72139 = ~n20358 ;
  assign n21187 = n72139 & n21179 ;
  assign n72140 = ~n20343 ;
  assign n20464 = n20342 & n72140 ;
  assign n20465 = n19720 | n20342 ;
  assign n72141 = ~n20465 ;
  assign n20466 = n20462 & n72141 ;
  assign n20467 = n20464 | n20466 ;
  assign n20468 = n143 & n20467 ;
  assign n20469 = n19711 & n72133 ;
  assign n20470 = n20361 & n20469 ;
  assign n20471 = n20468 | n20470 ;
  assign n20472 = n72025 & n20471 ;
  assign n72142 = ~n20461 ;
  assign n20473 = n20337 & n72142 ;
  assign n20338 = n19728 | n20337 ;
  assign n72143 = ~n20338 ;
  assign n20474 = n72143 & n20460 ;
  assign n20475 = n20473 | n20474 ;
  assign n20476 = n143 & n20475 ;
  assign n20477 = n19719 & n72133 ;
  assign n20478 = n20361 & n20477 ;
  assign n20479 = n20476 | n20478 ;
  assign n20480 = n71645 & n20479 ;
  assign n72144 = ~n20332 ;
  assign n20481 = n20331 & n72144 ;
  assign n20482 = n19736 | n20331 ;
  assign n72145 = ~n20482 ;
  assign n20483 = n20458 & n72145 ;
  assign n20484 = n20481 | n20483 ;
  assign n20485 = n143 & n20484 ;
  assign n20486 = n19727 & n72133 ;
  assign n20487 = n20361 & n20486 ;
  assign n20488 = n20485 | n20487 ;
  assign n20489 = n71633 & n20488 ;
  assign n72146 = ~n20457 ;
  assign n20490 = n20327 & n72146 ;
  assign n20491 = n19744 | n20327 ;
  assign n72147 = ~n20491 ;
  assign n20492 = n20323 & n72147 ;
  assign n20493 = n20490 | n20492 ;
  assign n20494 = n143 & n20493 ;
  assign n20495 = n19735 & n72133 ;
  assign n20496 = n20361 & n20495 ;
  assign n20497 = n20494 | n20496 ;
  assign n20498 = n71253 & n20497 ;
  assign n72148 = ~n20322 ;
  assign n20499 = n20321 & n72148 ;
  assign n20500 = n19752 | n20321 ;
  assign n72149 = ~n20500 ;
  assign n20501 = n20454 & n72149 ;
  assign n20502 = n20499 | n20501 ;
  assign n20503 = n143 & n20502 ;
  assign n20504 = n19743 & n72133 ;
  assign n20505 = n20361 & n20504 ;
  assign n20506 = n20503 | n20505 ;
  assign n20507 = n70935 & n20506 ;
  assign n72150 = ~n20453 ;
  assign n20508 = n20317 & n72150 ;
  assign n20509 = n19760 | n20317 ;
  assign n72151 = ~n20509 ;
  assign n20510 = n20313 & n72151 ;
  assign n20511 = n20508 | n20510 ;
  assign n20512 = n143 & n20511 ;
  assign n20513 = n19751 & n72133 ;
  assign n20514 = n20361 & n20513 ;
  assign n20515 = n20512 | n20514 ;
  assign n20516 = n70927 & n20515 ;
  assign n72152 = ~n20312 ;
  assign n20517 = n20311 & n72152 ;
  assign n20518 = n19768 | n20311 ;
  assign n72153 = ~n20518 ;
  assign n20519 = n20450 & n72153 ;
  assign n20520 = n20517 | n20519 ;
  assign n20521 = n143 & n20520 ;
  assign n20522 = n19759 & n72133 ;
  assign n20523 = n20361 & n20522 ;
  assign n20524 = n20521 | n20523 ;
  assign n20525 = n70609 & n20524 ;
  assign n72154 = ~n20449 ;
  assign n20526 = n20307 & n72154 ;
  assign n20527 = n19776 | n20307 ;
  assign n72155 = ~n20527 ;
  assign n20528 = n20303 & n72155 ;
  assign n20529 = n20526 | n20528 ;
  assign n20530 = n143 & n20529 ;
  assign n20531 = n19767 & n72133 ;
  assign n20532 = n20361 & n20531 ;
  assign n20533 = n20530 | n20532 ;
  assign n20534 = n70276 & n20533 ;
  assign n72156 = ~n20302 ;
  assign n20535 = n20301 & n72156 ;
  assign n20536 = n19784 | n20301 ;
  assign n72157 = ~n20536 ;
  assign n20537 = n20446 & n72157 ;
  assign n20538 = n20535 | n20537 ;
  assign n20539 = n143 & n20538 ;
  assign n20540 = n19775 & n72133 ;
  assign n20541 = n20361 & n20540 ;
  assign n20542 = n20539 | n20541 ;
  assign n20543 = n70176 & n20542 ;
  assign n72158 = ~n20445 ;
  assign n20544 = n20297 & n72158 ;
  assign n20545 = n19792 | n20297 ;
  assign n72159 = ~n20545 ;
  assign n20546 = n20293 & n72159 ;
  assign n20547 = n20544 | n20546 ;
  assign n20548 = n143 & n20547 ;
  assign n20549 = n19783 & n72133 ;
  assign n20550 = n20361 & n20549 ;
  assign n20551 = n20548 | n20550 ;
  assign n20552 = n69857 & n20551 ;
  assign n72160 = ~n20292 ;
  assign n20553 = n20291 & n72160 ;
  assign n20554 = n19800 | n20291 ;
  assign n72161 = ~n20554 ;
  assign n20555 = n20442 & n72161 ;
  assign n20556 = n20553 | n20555 ;
  assign n20557 = n143 & n20556 ;
  assign n20558 = n19791 & n72133 ;
  assign n20559 = n20361 & n20558 ;
  assign n20560 = n20557 | n20559 ;
  assign n20561 = n69656 & n20560 ;
  assign n72162 = ~n20441 ;
  assign n20562 = n20287 & n72162 ;
  assign n20563 = n19808 | n20287 ;
  assign n72163 = ~n20563 ;
  assign n20564 = n20283 & n72163 ;
  assign n20565 = n20562 | n20564 ;
  assign n20566 = n143 & n20565 ;
  assign n20567 = n19799 & n72133 ;
  assign n20568 = n20361 & n20567 ;
  assign n20569 = n20566 | n20568 ;
  assign n20570 = n69528 & n20569 ;
  assign n72164 = ~n20282 ;
  assign n20571 = n20281 & n72164 ;
  assign n20572 = n19816 | n20281 ;
  assign n72165 = ~n20572 ;
  assign n20573 = n20438 & n72165 ;
  assign n20574 = n20571 | n20573 ;
  assign n20575 = n143 & n20574 ;
  assign n20576 = n19807 & n72133 ;
  assign n20577 = n20361 & n20576 ;
  assign n20578 = n20575 | n20577 ;
  assign n20579 = n69261 & n20578 ;
  assign n72166 = ~n20437 ;
  assign n20580 = n20277 & n72166 ;
  assign n20581 = n19824 | n20277 ;
  assign n72167 = ~n20581 ;
  assign n20582 = n20273 & n72167 ;
  assign n20583 = n20580 | n20582 ;
  assign n20584 = n143 & n20583 ;
  assign n20585 = n19815 & n72133 ;
  assign n20586 = n20361 & n20585 ;
  assign n20587 = n20584 | n20586 ;
  assign n20588 = n69075 & n20587 ;
  assign n72168 = ~n20272 ;
  assign n20589 = n20271 & n72168 ;
  assign n20590 = n19832 | n20271 ;
  assign n72169 = ~n20590 ;
  assign n20591 = n20434 & n72169 ;
  assign n20592 = n20589 | n20591 ;
  assign n20593 = n143 & n20592 ;
  assign n20594 = n19823 & n72133 ;
  assign n20595 = n20361 & n20594 ;
  assign n20596 = n20593 | n20595 ;
  assign n20597 = n68993 & n20596 ;
  assign n72170 = ~n20433 ;
  assign n20598 = n20267 & n72170 ;
  assign n20599 = n19840 | n20267 ;
  assign n72171 = ~n20599 ;
  assign n20600 = n20263 & n72171 ;
  assign n20601 = n20598 | n20600 ;
  assign n20602 = n143 & n20601 ;
  assign n20603 = n19831 & n72133 ;
  assign n20604 = n20361 & n20603 ;
  assign n20605 = n20602 | n20604 ;
  assign n20606 = n68716 & n20605 ;
  assign n72172 = ~n20262 ;
  assign n20607 = n20261 & n72172 ;
  assign n20608 = n19848 | n20261 ;
  assign n72173 = ~n20608 ;
  assign n20609 = n20430 & n72173 ;
  assign n20610 = n20607 | n20609 ;
  assign n20611 = n143 & n20610 ;
  assign n20612 = n19839 & n72133 ;
  assign n20613 = n20361 & n20612 ;
  assign n20614 = n20611 | n20613 ;
  assign n20615 = n68545 & n20614 ;
  assign n72174 = ~n20429 ;
  assign n20616 = n20257 & n72174 ;
  assign n20617 = n19856 | n20257 ;
  assign n72175 = ~n20617 ;
  assign n20618 = n20253 & n72175 ;
  assign n20619 = n20616 | n20618 ;
  assign n20620 = n143 & n20619 ;
  assign n20621 = n19847 & n72133 ;
  assign n20622 = n20361 & n20621 ;
  assign n20623 = n20620 | n20622 ;
  assign n20624 = n68438 & n20623 ;
  assign n72176 = ~n20252 ;
  assign n20625 = n20251 & n72176 ;
  assign n20626 = n19864 | n20251 ;
  assign n72177 = ~n20626 ;
  assign n20627 = n20426 & n72177 ;
  assign n20628 = n20625 | n20627 ;
  assign n20629 = n143 & n20628 ;
  assign n20630 = n19855 & n72133 ;
  assign n20631 = n20361 & n20630 ;
  assign n20632 = n20629 | n20631 ;
  assign n20633 = n68214 & n20632 ;
  assign n72178 = ~n20425 ;
  assign n20634 = n20247 & n72178 ;
  assign n20635 = n19872 | n20247 ;
  assign n72179 = ~n20635 ;
  assign n20636 = n20243 & n72179 ;
  assign n20637 = n20634 | n20636 ;
  assign n20638 = n143 & n20637 ;
  assign n20639 = n19863 & n72133 ;
  assign n20640 = n20361 & n20639 ;
  assign n20641 = n20638 | n20640 ;
  assign n20642 = n68058 & n20641 ;
  assign n72180 = ~n20242 ;
  assign n20643 = n20241 & n72180 ;
  assign n20644 = n19880 | n20241 ;
  assign n72181 = ~n20644 ;
  assign n20645 = n20422 & n72181 ;
  assign n20646 = n20643 | n20645 ;
  assign n20647 = n143 & n20646 ;
  assign n20648 = n19871 & n72133 ;
  assign n20649 = n20361 & n20648 ;
  assign n20650 = n20647 | n20649 ;
  assign n20651 = n67986 & n20650 ;
  assign n72182 = ~n20421 ;
  assign n20652 = n20237 & n72182 ;
  assign n20653 = n19888 | n20237 ;
  assign n72183 = ~n20653 ;
  assign n20654 = n20233 & n72183 ;
  assign n20655 = n20652 | n20654 ;
  assign n20656 = n143 & n20655 ;
  assign n20657 = n19879 & n72133 ;
  assign n20658 = n20361 & n20657 ;
  assign n20659 = n20656 | n20658 ;
  assign n20660 = n67763 & n20659 ;
  assign n72184 = ~n20232 ;
  assign n20661 = n20231 & n72184 ;
  assign n20662 = n19896 | n20231 ;
  assign n72185 = ~n20662 ;
  assign n20663 = n20418 & n72185 ;
  assign n20664 = n20661 | n20663 ;
  assign n20665 = n143 & n20664 ;
  assign n20666 = n19887 & n72133 ;
  assign n20667 = n20361 & n20666 ;
  assign n20668 = n20665 | n20667 ;
  assign n20669 = n67622 & n20668 ;
  assign n72186 = ~n20417 ;
  assign n20670 = n20227 & n72186 ;
  assign n20671 = n19904 | n20227 ;
  assign n72187 = ~n20671 ;
  assign n20672 = n20223 & n72187 ;
  assign n20673 = n20670 | n20672 ;
  assign n20674 = n143 & n20673 ;
  assign n20675 = n19895 & n72133 ;
  assign n20676 = n20361 & n20675 ;
  assign n20677 = n20674 | n20676 ;
  assign n20678 = n67531 & n20677 ;
  assign n72188 = ~n20222 ;
  assign n20679 = n20221 & n72188 ;
  assign n20680 = n19912 | n20221 ;
  assign n72189 = ~n20680 ;
  assign n20681 = n20414 & n72189 ;
  assign n20682 = n20679 | n20681 ;
  assign n20683 = n143 & n20682 ;
  assign n20684 = n19903 & n72133 ;
  assign n20685 = n20361 & n20684 ;
  assign n20686 = n20683 | n20685 ;
  assign n20687 = n67348 & n20686 ;
  assign n72190 = ~n20413 ;
  assign n20688 = n20217 & n72190 ;
  assign n20689 = n19920 | n20217 ;
  assign n72191 = ~n20689 ;
  assign n20690 = n20213 & n72191 ;
  assign n20691 = n20688 | n20690 ;
  assign n20692 = n143 & n20691 ;
  assign n20693 = n19911 & n72133 ;
  assign n20694 = n20361 & n20693 ;
  assign n20695 = n20692 | n20694 ;
  assign n20696 = n67222 & n20695 ;
  assign n72192 = ~n20212 ;
  assign n20697 = n20210 & n72192 ;
  assign n20211 = n19928 | n20210 ;
  assign n72193 = ~n20211 ;
  assign n20698 = n20207 & n72193 ;
  assign n20699 = n20697 | n20698 ;
  assign n20700 = n143 & n20699 ;
  assign n20701 = n19919 & n72133 ;
  assign n20702 = n20361 & n20701 ;
  assign n20703 = n20700 | n20702 ;
  assign n20704 = n67164 & n20703 ;
  assign n72194 = ~n20409 ;
  assign n20705 = n20206 & n72194 ;
  assign n20706 = n19936 | n20206 ;
  assign n72195 = ~n20706 ;
  assign n20707 = n20202 & n72195 ;
  assign n20708 = n20705 | n20707 ;
  assign n20709 = n143 & n20708 ;
  assign n20710 = n19927 & n72133 ;
  assign n20711 = n20361 & n20710 ;
  assign n20712 = n20709 | n20711 ;
  assign n20713 = n66979 & n20712 ;
  assign n72196 = ~n20201 ;
  assign n20714 = n20200 & n72196 ;
  assign n20715 = n19944 | n20200 ;
  assign n72197 = ~n20715 ;
  assign n20716 = n20406 & n72197 ;
  assign n20717 = n20714 | n20716 ;
  assign n20718 = n143 & n20717 ;
  assign n20719 = n19935 & n72133 ;
  assign n20720 = n20361 & n20719 ;
  assign n20721 = n20718 | n20720 ;
  assign n20722 = n66868 & n20721 ;
  assign n72198 = ~n20405 ;
  assign n20723 = n20196 & n72198 ;
  assign n20724 = n19952 | n20196 ;
  assign n72199 = ~n20724 ;
  assign n20725 = n20192 & n72199 ;
  assign n20726 = n20723 | n20725 ;
  assign n20727 = n143 & n20726 ;
  assign n20728 = n19943 & n72133 ;
  assign n20729 = n20361 & n20728 ;
  assign n20730 = n20727 | n20729 ;
  assign n20731 = n66797 & n20730 ;
  assign n72200 = ~n20191 ;
  assign n20732 = n20189 & n72200 ;
  assign n20190 = n19960 | n20189 ;
  assign n72201 = ~n20190 ;
  assign n20733 = n20186 & n72201 ;
  assign n20734 = n20732 | n20733 ;
  assign n20735 = n143 & n20734 ;
  assign n20736 = n19951 & n72133 ;
  assign n20737 = n20361 & n20736 ;
  assign n20738 = n20735 | n20737 ;
  assign n20739 = n66654 & n20738 ;
  assign n72202 = ~n20401 ;
  assign n20740 = n20185 & n72202 ;
  assign n20741 = n19968 | n20185 ;
  assign n72203 = ~n20741 ;
  assign n20742 = n20181 & n72203 ;
  assign n20743 = n20740 | n20742 ;
  assign n20744 = n143 & n20743 ;
  assign n20745 = n19959 & n72133 ;
  assign n20746 = n20361 & n20745 ;
  assign n20747 = n20744 | n20746 ;
  assign n20748 = n66560 & n20747 ;
  assign n72204 = ~n20180 ;
  assign n20749 = n20178 & n72204 ;
  assign n20179 = n19976 | n20178 ;
  assign n72205 = ~n20179 ;
  assign n20750 = n20175 & n72205 ;
  assign n20751 = n20749 | n20750 ;
  assign n20752 = n143 & n20751 ;
  assign n20753 = n19967 & n72133 ;
  assign n20754 = n20361 & n20753 ;
  assign n20755 = n20752 | n20754 ;
  assign n20756 = n66505 & n20755 ;
  assign n72206 = ~n20397 ;
  assign n20757 = n20174 & n72206 ;
  assign n20758 = n19984 | n20174 ;
  assign n72207 = ~n20758 ;
  assign n20759 = n20170 & n72207 ;
  assign n20760 = n20757 | n20759 ;
  assign n20761 = n143 & n20760 ;
  assign n20762 = n19975 & n72133 ;
  assign n20763 = n20361 & n20762 ;
  assign n20764 = n20761 | n20763 ;
  assign n20765 = n66379 & n20764 ;
  assign n72208 = ~n20169 ;
  assign n20766 = n20168 & n72208 ;
  assign n20767 = n19992 | n20168 ;
  assign n72209 = ~n20767 ;
  assign n20768 = n20394 & n72209 ;
  assign n20769 = n20766 | n20768 ;
  assign n20770 = n143 & n20769 ;
  assign n20771 = n19983 & n72133 ;
  assign n20772 = n20361 & n20771 ;
  assign n20773 = n20770 | n20772 ;
  assign n20774 = n66299 & n20773 ;
  assign n72210 = ~n20393 ;
  assign n20775 = n20164 & n72210 ;
  assign n20776 = n20000 | n20164 ;
  assign n72211 = ~n20776 ;
  assign n20777 = n20160 & n72211 ;
  assign n20778 = n20775 | n20777 ;
  assign n20779 = n143 & n20778 ;
  assign n20780 = n19991 & n72133 ;
  assign n20781 = n20361 & n20780 ;
  assign n20782 = n20779 | n20781 ;
  assign n20783 = n66244 & n20782 ;
  assign n72212 = ~n20159 ;
  assign n20784 = n20158 & n72212 ;
  assign n20785 = n20008 | n20158 ;
  assign n72213 = ~n20785 ;
  assign n20786 = n20390 & n72213 ;
  assign n20787 = n20784 | n20786 ;
  assign n20788 = n143 & n20787 ;
  assign n20789 = n19999 & n72133 ;
  assign n20790 = n20361 & n20789 ;
  assign n20791 = n20788 | n20790 ;
  assign n20792 = n66145 & n20791 ;
  assign n72214 = ~n20389 ;
  assign n20793 = n20154 & n72214 ;
  assign n20794 = n20016 | n20154 ;
  assign n72215 = ~n20794 ;
  assign n20795 = n20150 & n72215 ;
  assign n20796 = n20793 | n20795 ;
  assign n20797 = n143 & n20796 ;
  assign n20798 = n20007 & n72133 ;
  assign n20799 = n20361 & n20798 ;
  assign n20800 = n20797 | n20799 ;
  assign n20801 = n66081 & n20800 ;
  assign n72216 = ~n20149 ;
  assign n20802 = n20148 & n72216 ;
  assign n20803 = n20024 | n20148 ;
  assign n72217 = ~n20803 ;
  assign n20804 = n20386 & n72217 ;
  assign n20805 = n20802 | n20804 ;
  assign n20806 = n143 & n20805 ;
  assign n20807 = n20015 & n72133 ;
  assign n20808 = n20361 & n20807 ;
  assign n20809 = n20806 | n20808 ;
  assign n20810 = n66043 & n20809 ;
  assign n72218 = ~n20385 ;
  assign n20811 = n20144 & n72218 ;
  assign n20812 = n20032 | n20144 ;
  assign n72219 = ~n20812 ;
  assign n20813 = n20140 & n72219 ;
  assign n20814 = n20811 | n20813 ;
  assign n20815 = n143 & n20814 ;
  assign n20816 = n20023 & n72133 ;
  assign n20817 = n20361 & n20816 ;
  assign n20818 = n20815 | n20817 ;
  assign n20819 = n65960 & n20818 ;
  assign n72220 = ~n20139 ;
  assign n20820 = n20138 & n72220 ;
  assign n20821 = n20041 | n20138 ;
  assign n72221 = ~n20821 ;
  assign n20822 = n20382 & n72221 ;
  assign n20823 = n20820 | n20822 ;
  assign n20824 = n143 & n20823 ;
  assign n20825 = n20031 & n72133 ;
  assign n20826 = n20361 & n20825 ;
  assign n20827 = n20824 | n20826 ;
  assign n20828 = n65909 & n20827 ;
  assign n72222 = ~n20381 ;
  assign n20829 = n20133 & n72222 ;
  assign n20134 = n20050 | n20133 ;
  assign n72223 = ~n20134 ;
  assign n20830 = n72223 & n20380 ;
  assign n20831 = n20829 | n20830 ;
  assign n20832 = n143 & n20831 ;
  assign n20833 = n20040 & n72133 ;
  assign n20834 = n20361 & n20833 ;
  assign n20835 = n20832 | n20834 ;
  assign n20836 = n65877 & n20835 ;
  assign n72224 = ~n20128 ;
  assign n20837 = n20127 & n72224 ;
  assign n20838 = n20059 | n20127 ;
  assign n72225 = ~n20838 ;
  assign n20839 = n20378 & n72225 ;
  assign n20840 = n20837 | n20839 ;
  assign n20841 = n143 & n20840 ;
  assign n20842 = n20049 & n72133 ;
  assign n20843 = n20361 & n20842 ;
  assign n20844 = n20841 | n20843 ;
  assign n20845 = n65820 & n20844 ;
  assign n72226 = ~n20377 ;
  assign n20846 = n20123 & n72226 ;
  assign n20847 = n20067 | n20123 ;
  assign n72227 = ~n20847 ;
  assign n20848 = n20119 & n72227 ;
  assign n20849 = n20846 | n20848 ;
  assign n20850 = n143 & n20849 ;
  assign n20851 = n20058 & n72133 ;
  assign n20852 = n20361 & n20851 ;
  assign n20853 = n20850 | n20852 ;
  assign n20854 = n65791 & n20853 ;
  assign n72228 = ~n20118 ;
  assign n20856 = n20117 & n72228 ;
  assign n20855 = n20076 | n20117 ;
  assign n72229 = ~n20855 ;
  assign n20857 = n20114 & n72229 ;
  assign n20858 = n20856 | n20857 ;
  assign n20859 = n143 & n20858 ;
  assign n20860 = n20066 & n72133 ;
  assign n20861 = n20361 & n20860 ;
  assign n20862 = n20859 | n20861 ;
  assign n20863 = n65772 & n20862 ;
  assign n72230 = ~n20373 ;
  assign n20865 = n20113 & n72230 ;
  assign n20864 = n20084 | n20113 ;
  assign n72231 = ~n20864 ;
  assign n20866 = n20372 & n72231 ;
  assign n20867 = n20865 | n20866 ;
  assign n20868 = n143 & n20867 ;
  assign n20869 = n20075 & n72133 ;
  assign n20870 = n20361 & n20869 ;
  assign n20871 = n20868 | n20870 ;
  assign n20872 = n65746 & n20871 ;
  assign n72232 = ~n20108 ;
  assign n20874 = n20107 & n72232 ;
  assign n20873 = n20104 | n20107 ;
  assign n72233 = ~n20873 ;
  assign n20875 = n20103 & n72233 ;
  assign n20876 = n20874 | n20875 ;
  assign n20877 = n143 & n20876 ;
  assign n20878 = n20083 & n72133 ;
  assign n20879 = n20361 & n20878 ;
  assign n20880 = n20877 | n20879 ;
  assign n20881 = n65721 & n20880 ;
  assign n20882 = n20100 & n20102 ;
  assign n20883 = n72030 & n20882 ;
  assign n72234 = ~n20883 ;
  assign n20884 = n20103 & n72234 ;
  assign n20885 = n143 & n20884 ;
  assign n20886 = n20097 & n72133 ;
  assign n20887 = n20361 & n20886 ;
  assign n20888 = n20885 | n20887 ;
  assign n20889 = n65686 & n20888 ;
  assign n20364 = n20102 & n143 ;
  assign n20896 = x64 & n143 ;
  assign n72235 = ~n20896 ;
  assign n20897 = x14 & n72235 ;
  assign n20898 = n20364 | n20897 ;
  assign n20900 = x65 & n20898 ;
  assign n20892 = n20360 | n20891 ;
  assign n20893 = n72133 & n20892 ;
  assign n72236 = ~n20893 ;
  assign n20894 = x64 & n72236 ;
  assign n72237 = ~n20894 ;
  assign n20895 = x14 & n72237 ;
  assign n20899 = x65 | n20364 ;
  assign n20901 = n20895 | n20899 ;
  assign n72238 = ~n20900 ;
  assign n20902 = n72238 & n20901 ;
  assign n72239 = ~x13 ;
  assign n20903 = n72239 & x64 ;
  assign n20904 = n20902 | n20903 ;
  assign n20905 = n65670 & n20898 ;
  assign n72240 = ~n20905 ;
  assign n20906 = n20904 & n72240 ;
  assign n72241 = ~n20887 ;
  assign n20907 = x66 & n72241 ;
  assign n72242 = ~n20885 ;
  assign n20908 = n72242 & n20907 ;
  assign n20909 = n20889 | n20908 ;
  assign n20910 = n20906 | n20909 ;
  assign n72243 = ~n20889 ;
  assign n20911 = n72243 & n20910 ;
  assign n72244 = ~n20879 ;
  assign n20912 = x67 & n72244 ;
  assign n72245 = ~n20877 ;
  assign n20913 = n72245 & n20912 ;
  assign n20914 = n20881 | n20913 ;
  assign n20915 = n20911 | n20914 ;
  assign n72246 = ~n20881 ;
  assign n20916 = n72246 & n20915 ;
  assign n72247 = ~n20870 ;
  assign n20917 = x68 & n72247 ;
  assign n72248 = ~n20868 ;
  assign n20918 = n72248 & n20917 ;
  assign n20919 = n20872 | n20918 ;
  assign n20920 = n20916 | n20919 ;
  assign n72249 = ~n20872 ;
  assign n20921 = n72249 & n20920 ;
  assign n72250 = ~n20861 ;
  assign n20922 = x69 & n72250 ;
  assign n72251 = ~n20859 ;
  assign n20923 = n72251 & n20922 ;
  assign n20924 = n20863 | n20923 ;
  assign n20926 = n20921 | n20924 ;
  assign n72252 = ~n20863 ;
  assign n20927 = n72252 & n20926 ;
  assign n72253 = ~n20852 ;
  assign n20928 = x70 & n72253 ;
  assign n72254 = ~n20850 ;
  assign n20929 = n72254 & n20928 ;
  assign n20930 = n20854 | n20929 ;
  assign n20931 = n20927 | n20930 ;
  assign n72255 = ~n20854 ;
  assign n20932 = n72255 & n20931 ;
  assign n72256 = ~n20843 ;
  assign n20933 = x71 & n72256 ;
  assign n72257 = ~n20841 ;
  assign n20934 = n72257 & n20933 ;
  assign n20935 = n20845 | n20934 ;
  assign n20937 = n20932 | n20935 ;
  assign n72258 = ~n20845 ;
  assign n20938 = n72258 & n20937 ;
  assign n72259 = ~n20834 ;
  assign n20939 = x72 & n72259 ;
  assign n72260 = ~n20832 ;
  assign n20940 = n72260 & n20939 ;
  assign n20941 = n20836 | n20940 ;
  assign n20942 = n20938 | n20941 ;
  assign n72261 = ~n20836 ;
  assign n20943 = n72261 & n20942 ;
  assign n72262 = ~n20826 ;
  assign n20944 = x73 & n72262 ;
  assign n72263 = ~n20824 ;
  assign n20945 = n72263 & n20944 ;
  assign n20946 = n20828 | n20945 ;
  assign n20948 = n20943 | n20946 ;
  assign n72264 = ~n20828 ;
  assign n20949 = n72264 & n20948 ;
  assign n72265 = ~n20817 ;
  assign n20950 = x74 & n72265 ;
  assign n72266 = ~n20815 ;
  assign n20951 = n72266 & n20950 ;
  assign n20952 = n20819 | n20951 ;
  assign n20953 = n20949 | n20952 ;
  assign n72267 = ~n20819 ;
  assign n20954 = n72267 & n20953 ;
  assign n72268 = ~n20808 ;
  assign n20955 = x75 & n72268 ;
  assign n72269 = ~n20806 ;
  assign n20956 = n72269 & n20955 ;
  assign n20957 = n20810 | n20956 ;
  assign n20959 = n20954 | n20957 ;
  assign n72270 = ~n20810 ;
  assign n20960 = n72270 & n20959 ;
  assign n72271 = ~n20799 ;
  assign n20961 = x76 & n72271 ;
  assign n72272 = ~n20797 ;
  assign n20962 = n72272 & n20961 ;
  assign n20963 = n20801 | n20962 ;
  assign n20964 = n20960 | n20963 ;
  assign n72273 = ~n20801 ;
  assign n20965 = n72273 & n20964 ;
  assign n72274 = ~n20790 ;
  assign n20966 = x77 & n72274 ;
  assign n72275 = ~n20788 ;
  assign n20967 = n72275 & n20966 ;
  assign n20968 = n20792 | n20967 ;
  assign n20970 = n20965 | n20968 ;
  assign n72276 = ~n20792 ;
  assign n20971 = n72276 & n20970 ;
  assign n72277 = ~n20781 ;
  assign n20972 = x78 & n72277 ;
  assign n72278 = ~n20779 ;
  assign n20973 = n72278 & n20972 ;
  assign n20974 = n20783 | n20973 ;
  assign n20975 = n20971 | n20974 ;
  assign n72279 = ~n20783 ;
  assign n20976 = n72279 & n20975 ;
  assign n72280 = ~n20772 ;
  assign n20977 = x79 & n72280 ;
  assign n72281 = ~n20770 ;
  assign n20978 = n72281 & n20977 ;
  assign n20979 = n20774 | n20978 ;
  assign n20981 = n20976 | n20979 ;
  assign n72282 = ~n20774 ;
  assign n20982 = n72282 & n20981 ;
  assign n72283 = ~n20763 ;
  assign n20983 = x80 & n72283 ;
  assign n72284 = ~n20761 ;
  assign n20984 = n72284 & n20983 ;
  assign n20985 = n20765 | n20984 ;
  assign n20986 = n20982 | n20985 ;
  assign n72285 = ~n20765 ;
  assign n20987 = n72285 & n20986 ;
  assign n72286 = ~n20754 ;
  assign n20988 = x81 & n72286 ;
  assign n72287 = ~n20752 ;
  assign n20989 = n72287 & n20988 ;
  assign n20990 = n20756 | n20989 ;
  assign n20992 = n20987 | n20990 ;
  assign n72288 = ~n20756 ;
  assign n20993 = n72288 & n20992 ;
  assign n72289 = ~n20746 ;
  assign n20994 = x82 & n72289 ;
  assign n72290 = ~n20744 ;
  assign n20995 = n72290 & n20994 ;
  assign n20996 = n20748 | n20995 ;
  assign n20997 = n20993 | n20996 ;
  assign n72291 = ~n20748 ;
  assign n20998 = n72291 & n20997 ;
  assign n72292 = ~n20737 ;
  assign n20999 = x83 & n72292 ;
  assign n72293 = ~n20735 ;
  assign n21000 = n72293 & n20999 ;
  assign n21001 = n20739 | n21000 ;
  assign n21003 = n20998 | n21001 ;
  assign n72294 = ~n20739 ;
  assign n21004 = n72294 & n21003 ;
  assign n72295 = ~n20729 ;
  assign n21005 = x84 & n72295 ;
  assign n72296 = ~n20727 ;
  assign n21006 = n72296 & n21005 ;
  assign n21007 = n20731 | n21006 ;
  assign n21008 = n21004 | n21007 ;
  assign n72297 = ~n20731 ;
  assign n21009 = n72297 & n21008 ;
  assign n72298 = ~n20720 ;
  assign n21010 = x85 & n72298 ;
  assign n72299 = ~n20718 ;
  assign n21011 = n72299 & n21010 ;
  assign n21012 = n20722 | n21011 ;
  assign n21014 = n21009 | n21012 ;
  assign n72300 = ~n20722 ;
  assign n21015 = n72300 & n21014 ;
  assign n72301 = ~n20711 ;
  assign n21016 = x86 & n72301 ;
  assign n72302 = ~n20709 ;
  assign n21017 = n72302 & n21016 ;
  assign n21018 = n20713 | n21017 ;
  assign n21019 = n21015 | n21018 ;
  assign n72303 = ~n20713 ;
  assign n21020 = n72303 & n21019 ;
  assign n72304 = ~n20702 ;
  assign n21021 = x87 & n72304 ;
  assign n72305 = ~n20700 ;
  assign n21022 = n72305 & n21021 ;
  assign n21023 = n20704 | n21022 ;
  assign n21025 = n21020 | n21023 ;
  assign n72306 = ~n20704 ;
  assign n21026 = n72306 & n21025 ;
  assign n72307 = ~n20694 ;
  assign n21027 = x88 & n72307 ;
  assign n72308 = ~n20692 ;
  assign n21028 = n72308 & n21027 ;
  assign n21029 = n20696 | n21028 ;
  assign n21030 = n21026 | n21029 ;
  assign n72309 = ~n20696 ;
  assign n21031 = n72309 & n21030 ;
  assign n72310 = ~n20685 ;
  assign n21032 = x89 & n72310 ;
  assign n72311 = ~n20683 ;
  assign n21033 = n72311 & n21032 ;
  assign n21034 = n20687 | n21033 ;
  assign n21036 = n21031 | n21034 ;
  assign n72312 = ~n20687 ;
  assign n21037 = n72312 & n21036 ;
  assign n72313 = ~n20676 ;
  assign n21038 = x90 & n72313 ;
  assign n72314 = ~n20674 ;
  assign n21039 = n72314 & n21038 ;
  assign n21040 = n20678 | n21039 ;
  assign n21041 = n21037 | n21040 ;
  assign n72315 = ~n20678 ;
  assign n21042 = n72315 & n21041 ;
  assign n72316 = ~n20667 ;
  assign n21043 = x91 & n72316 ;
  assign n72317 = ~n20665 ;
  assign n21044 = n72317 & n21043 ;
  assign n21045 = n20669 | n21044 ;
  assign n21047 = n21042 | n21045 ;
  assign n72318 = ~n20669 ;
  assign n21048 = n72318 & n21047 ;
  assign n72319 = ~n20658 ;
  assign n21049 = x92 & n72319 ;
  assign n72320 = ~n20656 ;
  assign n21050 = n72320 & n21049 ;
  assign n21051 = n20660 | n21050 ;
  assign n21052 = n21048 | n21051 ;
  assign n72321 = ~n20660 ;
  assign n21053 = n72321 & n21052 ;
  assign n72322 = ~n20649 ;
  assign n21054 = x93 & n72322 ;
  assign n72323 = ~n20647 ;
  assign n21055 = n72323 & n21054 ;
  assign n21056 = n20651 | n21055 ;
  assign n21058 = n21053 | n21056 ;
  assign n72324 = ~n20651 ;
  assign n21059 = n72324 & n21058 ;
  assign n72325 = ~n20640 ;
  assign n21060 = x94 & n72325 ;
  assign n72326 = ~n20638 ;
  assign n21061 = n72326 & n21060 ;
  assign n21062 = n20642 | n21061 ;
  assign n21063 = n21059 | n21062 ;
  assign n72327 = ~n20642 ;
  assign n21064 = n72327 & n21063 ;
  assign n72328 = ~n20631 ;
  assign n21065 = x95 & n72328 ;
  assign n72329 = ~n20629 ;
  assign n21066 = n72329 & n21065 ;
  assign n21067 = n20633 | n21066 ;
  assign n21069 = n21064 | n21067 ;
  assign n72330 = ~n20633 ;
  assign n21070 = n72330 & n21069 ;
  assign n72331 = ~n20622 ;
  assign n21071 = x96 & n72331 ;
  assign n72332 = ~n20620 ;
  assign n21072 = n72332 & n21071 ;
  assign n21073 = n20624 | n21072 ;
  assign n21074 = n21070 | n21073 ;
  assign n72333 = ~n20624 ;
  assign n21075 = n72333 & n21074 ;
  assign n72334 = ~n20613 ;
  assign n21076 = x97 & n72334 ;
  assign n72335 = ~n20611 ;
  assign n21077 = n72335 & n21076 ;
  assign n21078 = n20615 | n21077 ;
  assign n21080 = n21075 | n21078 ;
  assign n72336 = ~n20615 ;
  assign n21081 = n72336 & n21080 ;
  assign n72337 = ~n20604 ;
  assign n21082 = x98 & n72337 ;
  assign n72338 = ~n20602 ;
  assign n21083 = n72338 & n21082 ;
  assign n21084 = n20606 | n21083 ;
  assign n21085 = n21081 | n21084 ;
  assign n72339 = ~n20606 ;
  assign n21086 = n72339 & n21085 ;
  assign n72340 = ~n20595 ;
  assign n21087 = x99 & n72340 ;
  assign n72341 = ~n20593 ;
  assign n21088 = n72341 & n21087 ;
  assign n21089 = n20597 | n21088 ;
  assign n21091 = n21086 | n21089 ;
  assign n72342 = ~n20597 ;
  assign n21092 = n72342 & n21091 ;
  assign n72343 = ~n20586 ;
  assign n21093 = x100 & n72343 ;
  assign n72344 = ~n20584 ;
  assign n21094 = n72344 & n21093 ;
  assign n21095 = n20588 | n21094 ;
  assign n21096 = n21092 | n21095 ;
  assign n72345 = ~n20588 ;
  assign n21097 = n72345 & n21096 ;
  assign n72346 = ~n20577 ;
  assign n21098 = x101 & n72346 ;
  assign n72347 = ~n20575 ;
  assign n21099 = n72347 & n21098 ;
  assign n21100 = n20579 | n21099 ;
  assign n21102 = n21097 | n21100 ;
  assign n72348 = ~n20579 ;
  assign n21103 = n72348 & n21102 ;
  assign n72349 = ~n20568 ;
  assign n21104 = x102 & n72349 ;
  assign n72350 = ~n20566 ;
  assign n21105 = n72350 & n21104 ;
  assign n21106 = n20570 | n21105 ;
  assign n21107 = n21103 | n21106 ;
  assign n72351 = ~n20570 ;
  assign n21108 = n72351 & n21107 ;
  assign n72352 = ~n20559 ;
  assign n21109 = x103 & n72352 ;
  assign n72353 = ~n20557 ;
  assign n21110 = n72353 & n21109 ;
  assign n21111 = n20561 | n21110 ;
  assign n21113 = n21108 | n21111 ;
  assign n72354 = ~n20561 ;
  assign n21114 = n72354 & n21113 ;
  assign n72355 = ~n20550 ;
  assign n21115 = x104 & n72355 ;
  assign n72356 = ~n20548 ;
  assign n21116 = n72356 & n21115 ;
  assign n21117 = n20552 | n21116 ;
  assign n21118 = n21114 | n21117 ;
  assign n72357 = ~n20552 ;
  assign n21119 = n72357 & n21118 ;
  assign n72358 = ~n20541 ;
  assign n21120 = x105 & n72358 ;
  assign n72359 = ~n20539 ;
  assign n21121 = n72359 & n21120 ;
  assign n21122 = n20543 | n21121 ;
  assign n21124 = n21119 | n21122 ;
  assign n72360 = ~n20543 ;
  assign n21125 = n72360 & n21124 ;
  assign n72361 = ~n20532 ;
  assign n21126 = x106 & n72361 ;
  assign n72362 = ~n20530 ;
  assign n21127 = n72362 & n21126 ;
  assign n21128 = n20534 | n21127 ;
  assign n21129 = n21125 | n21128 ;
  assign n72363 = ~n20534 ;
  assign n21130 = n72363 & n21129 ;
  assign n72364 = ~n20523 ;
  assign n21131 = x107 & n72364 ;
  assign n72365 = ~n20521 ;
  assign n21132 = n72365 & n21131 ;
  assign n21133 = n20525 | n21132 ;
  assign n21135 = n21130 | n21133 ;
  assign n72366 = ~n20525 ;
  assign n21136 = n72366 & n21135 ;
  assign n72367 = ~n20514 ;
  assign n21137 = x108 & n72367 ;
  assign n72368 = ~n20512 ;
  assign n21138 = n72368 & n21137 ;
  assign n21139 = n20516 | n21138 ;
  assign n21140 = n21136 | n21139 ;
  assign n72369 = ~n20516 ;
  assign n21141 = n72369 & n21140 ;
  assign n72370 = ~n20505 ;
  assign n21142 = x109 & n72370 ;
  assign n72371 = ~n20503 ;
  assign n21143 = n72371 & n21142 ;
  assign n21144 = n20507 | n21143 ;
  assign n21146 = n21141 | n21144 ;
  assign n72372 = ~n20507 ;
  assign n21147 = n72372 & n21146 ;
  assign n72373 = ~n20496 ;
  assign n21148 = x110 & n72373 ;
  assign n72374 = ~n20494 ;
  assign n21149 = n72374 & n21148 ;
  assign n21150 = n20498 | n21149 ;
  assign n21151 = n21147 | n21150 ;
  assign n72375 = ~n20498 ;
  assign n21152 = n72375 & n21151 ;
  assign n72376 = ~n20487 ;
  assign n21153 = x111 & n72376 ;
  assign n72377 = ~n20485 ;
  assign n21154 = n72377 & n21153 ;
  assign n21155 = n20489 | n21154 ;
  assign n21157 = n21152 | n21155 ;
  assign n72378 = ~n20489 ;
  assign n21158 = n72378 & n21157 ;
  assign n72379 = ~n20478 ;
  assign n21159 = x112 & n72379 ;
  assign n72380 = ~n20476 ;
  assign n21160 = n72380 & n21159 ;
  assign n21161 = n20480 | n21160 ;
  assign n21162 = n21158 | n21161 ;
  assign n72381 = ~n20480 ;
  assign n21163 = n72381 & n21162 ;
  assign n72382 = ~n20470 ;
  assign n21164 = x113 & n72382 ;
  assign n72383 = ~n20468 ;
  assign n21165 = n72383 & n21164 ;
  assign n21166 = n20472 | n21165 ;
  assign n21168 = n21163 | n21166 ;
  assign n72384 = ~n20472 ;
  assign n21169 = n72384 & n21168 ;
  assign n72385 = ~x114 ;
  assign n21180 = n72385 & n21179 ;
  assign n72386 = ~n21178 ;
  assign n21181 = x114 & n72386 ;
  assign n72387 = ~n21176 ;
  assign n21182 = n72387 & n21181 ;
  assign n21183 = n268 | n270 ;
  assign n21184 = n278 | n21183 ;
  assign n21185 = n21182 | n21184 ;
  assign n21186 = n21180 | n21185 ;
  assign n21188 = n21169 | n21186 ;
  assign n72388 = ~n21187 ;
  assign n21189 = n72388 & n21188 ;
  assign n21318 = n20472 | n21182 ;
  assign n21319 = n21180 | n21318 ;
  assign n72389 = ~n21319 ;
  assign n21320 = n21168 & n72389 ;
  assign n21192 = n20364 | n20895 ;
  assign n21193 = x65 & n21192 ;
  assign n72390 = ~n21193 ;
  assign n21194 = n20901 & n72390 ;
  assign n21195 = n20903 | n21194 ;
  assign n21196 = n72240 & n21195 ;
  assign n21197 = n20909 | n21196 ;
  assign n21198 = n72243 & n21197 ;
  assign n21200 = n20914 | n21198 ;
  assign n21201 = n72246 & n21200 ;
  assign n21203 = n20919 | n21201 ;
  assign n21204 = n72249 & n21203 ;
  assign n21205 = n20924 | n21204 ;
  assign n21206 = n72252 & n21205 ;
  assign n21207 = n20930 | n21206 ;
  assign n21209 = n72255 & n21207 ;
  assign n21210 = n20935 | n21209 ;
  assign n21211 = n72258 & n21210 ;
  assign n21212 = n20941 | n21211 ;
  assign n21214 = n72261 & n21212 ;
  assign n21215 = n20946 | n21214 ;
  assign n21216 = n72264 & n21215 ;
  assign n21217 = n20952 | n21216 ;
  assign n21219 = n72267 & n21217 ;
  assign n21220 = n20957 | n21219 ;
  assign n21221 = n72270 & n21220 ;
  assign n21222 = n20963 | n21221 ;
  assign n21224 = n72273 & n21222 ;
  assign n21225 = n20968 | n21224 ;
  assign n21226 = n72276 & n21225 ;
  assign n21227 = n20974 | n21226 ;
  assign n21229 = n72279 & n21227 ;
  assign n21230 = n20979 | n21229 ;
  assign n21231 = n72282 & n21230 ;
  assign n21232 = n20985 | n21231 ;
  assign n21234 = n72285 & n21232 ;
  assign n21235 = n20990 | n21234 ;
  assign n21236 = n72288 & n21235 ;
  assign n21237 = n20996 | n21236 ;
  assign n21239 = n72291 & n21237 ;
  assign n21240 = n21001 | n21239 ;
  assign n21241 = n72294 & n21240 ;
  assign n21242 = n21007 | n21241 ;
  assign n21244 = n72297 & n21242 ;
  assign n21245 = n21012 | n21244 ;
  assign n21246 = n72300 & n21245 ;
  assign n21247 = n21018 | n21246 ;
  assign n21249 = n72303 & n21247 ;
  assign n21250 = n21023 | n21249 ;
  assign n21251 = n72306 & n21250 ;
  assign n21252 = n21029 | n21251 ;
  assign n21254 = n72309 & n21252 ;
  assign n21255 = n21034 | n21254 ;
  assign n21256 = n72312 & n21255 ;
  assign n21257 = n21040 | n21256 ;
  assign n21259 = n72315 & n21257 ;
  assign n21260 = n21045 | n21259 ;
  assign n21261 = n72318 & n21260 ;
  assign n21262 = n21051 | n21261 ;
  assign n21264 = n72321 & n21262 ;
  assign n21265 = n21056 | n21264 ;
  assign n21266 = n72324 & n21265 ;
  assign n21267 = n21062 | n21266 ;
  assign n21269 = n72327 & n21267 ;
  assign n21270 = n21067 | n21269 ;
  assign n21271 = n72330 & n21270 ;
  assign n21272 = n21073 | n21271 ;
  assign n21274 = n72333 & n21272 ;
  assign n21275 = n21078 | n21274 ;
  assign n21276 = n72336 & n21275 ;
  assign n21277 = n21084 | n21276 ;
  assign n21279 = n72339 & n21277 ;
  assign n21280 = n21089 | n21279 ;
  assign n21281 = n72342 & n21280 ;
  assign n21282 = n21095 | n21281 ;
  assign n21284 = n72345 & n21282 ;
  assign n21285 = n21100 | n21284 ;
  assign n21286 = n72348 & n21285 ;
  assign n21287 = n21106 | n21286 ;
  assign n21289 = n72351 & n21287 ;
  assign n21290 = n21111 | n21289 ;
  assign n21291 = n72354 & n21290 ;
  assign n21292 = n21117 | n21291 ;
  assign n21294 = n72357 & n21292 ;
  assign n21295 = n21122 | n21294 ;
  assign n21296 = n72360 & n21295 ;
  assign n21297 = n21128 | n21296 ;
  assign n21299 = n72363 & n21297 ;
  assign n21300 = n21133 | n21299 ;
  assign n21301 = n72366 & n21300 ;
  assign n21302 = n21139 | n21301 ;
  assign n21304 = n72369 & n21302 ;
  assign n21305 = n21144 | n21304 ;
  assign n21306 = n72372 & n21305 ;
  assign n21307 = n21150 | n21306 ;
  assign n21309 = n72375 & n21307 ;
  assign n21310 = n21155 | n21309 ;
  assign n21311 = n72378 & n21310 ;
  assign n21312 = n21161 | n21311 ;
  assign n21314 = n72381 & n21312 ;
  assign n21315 = n21166 | n21314 ;
  assign n21316 = n72384 & n21315 ;
  assign n21321 = n21180 | n21182 ;
  assign n72391 = ~n21316 ;
  assign n21322 = n72391 & n21321 ;
  assign n21323 = n21320 | n21322 ;
  assign n142 = ~n21189 ;
  assign n21324 = n142 & n21323 ;
  assign n21317 = n21186 | n21316 ;
  assign n21325 = n20358 & n21179 ;
  assign n21326 = n21317 & n21325 ;
  assign n21327 = n21324 | n21326 ;
  assign n72393 = ~x115 ;
  assign n21328 = n72393 & n21327 ;
  assign n72394 = ~n21326 ;
  assign n22026 = x115 & n72394 ;
  assign n72395 = ~n21324 ;
  assign n22027 = n72395 & n22026 ;
  assign n22028 = n21328 | n22027 ;
  assign n72396 = ~n21163 ;
  assign n21167 = n72396 & n21166 ;
  assign n21329 = n20480 | n21166 ;
  assign n72397 = ~n21329 ;
  assign n21330 = n21312 & n72397 ;
  assign n21331 = n21167 | n21330 ;
  assign n21332 = n142 & n21331 ;
  assign n21333 = n20471 & n72388 ;
  assign n21334 = n21317 & n21333 ;
  assign n21335 = n21332 | n21334 ;
  assign n21336 = n72385 & n21335 ;
  assign n72398 = ~n21311 ;
  assign n21313 = n21161 & n72398 ;
  assign n21337 = n20489 | n21161 ;
  assign n72399 = ~n21337 ;
  assign n21338 = n21157 & n72399 ;
  assign n21339 = n21313 | n21338 ;
  assign n21340 = n142 & n21339 ;
  assign n21341 = n20479 & n72388 ;
  assign n21342 = n21317 & n21341 ;
  assign n21343 = n21340 | n21342 ;
  assign n21344 = n72025 & n21343 ;
  assign n72400 = ~n21342 ;
  assign n22014 = x113 & n72400 ;
  assign n72401 = ~n21340 ;
  assign n22015 = n72401 & n22014 ;
  assign n22016 = n21344 | n22015 ;
  assign n72402 = ~n21152 ;
  assign n21156 = n72402 & n21155 ;
  assign n21345 = n20498 | n21155 ;
  assign n72403 = ~n21345 ;
  assign n21346 = n21307 & n72403 ;
  assign n21347 = n21156 | n21346 ;
  assign n21348 = n142 & n21347 ;
  assign n21349 = n20488 & n72388 ;
  assign n21350 = n21317 & n21349 ;
  assign n21351 = n21348 | n21350 ;
  assign n21352 = n71645 & n21351 ;
  assign n72404 = ~n21306 ;
  assign n21308 = n21150 & n72404 ;
  assign n21353 = n20507 | n21150 ;
  assign n72405 = ~n21353 ;
  assign n21354 = n21146 & n72405 ;
  assign n21355 = n21308 | n21354 ;
  assign n21356 = n142 & n21355 ;
  assign n21357 = n20497 & n72388 ;
  assign n21358 = n21317 & n21357 ;
  assign n21359 = n21356 | n21358 ;
  assign n21360 = n71633 & n21359 ;
  assign n72406 = ~n21358 ;
  assign n22002 = x111 & n72406 ;
  assign n72407 = ~n21356 ;
  assign n22003 = n72407 & n22002 ;
  assign n22004 = n21360 | n22003 ;
  assign n72408 = ~n21141 ;
  assign n21145 = n72408 & n21144 ;
  assign n21361 = n20516 | n21144 ;
  assign n72409 = ~n21361 ;
  assign n21362 = n21302 & n72409 ;
  assign n21363 = n21145 | n21362 ;
  assign n21364 = n142 & n21363 ;
  assign n21365 = n20506 & n72388 ;
  assign n21366 = n21317 & n21365 ;
  assign n21367 = n21364 | n21366 ;
  assign n21368 = n71253 & n21367 ;
  assign n72410 = ~n21301 ;
  assign n21303 = n21139 & n72410 ;
  assign n21369 = n20525 | n21139 ;
  assign n72411 = ~n21369 ;
  assign n21370 = n21135 & n72411 ;
  assign n21371 = n21303 | n21370 ;
  assign n21372 = n142 & n21371 ;
  assign n21373 = n20515 & n72388 ;
  assign n21374 = n21317 & n21373 ;
  assign n21375 = n21372 | n21374 ;
  assign n21376 = n70935 & n21375 ;
  assign n72412 = ~n21374 ;
  assign n21990 = x109 & n72412 ;
  assign n72413 = ~n21372 ;
  assign n21991 = n72413 & n21990 ;
  assign n21992 = n21376 | n21991 ;
  assign n72414 = ~n21130 ;
  assign n21134 = n72414 & n21133 ;
  assign n21377 = n20534 | n21133 ;
  assign n72415 = ~n21377 ;
  assign n21378 = n21297 & n72415 ;
  assign n21379 = n21134 | n21378 ;
  assign n21380 = n142 & n21379 ;
  assign n21381 = n20524 & n72388 ;
  assign n21382 = n21317 & n21381 ;
  assign n21383 = n21380 | n21382 ;
  assign n21384 = n70927 & n21383 ;
  assign n72416 = ~n21296 ;
  assign n21298 = n21128 & n72416 ;
  assign n21385 = n20543 | n21128 ;
  assign n72417 = ~n21385 ;
  assign n21386 = n21124 & n72417 ;
  assign n21387 = n21298 | n21386 ;
  assign n21388 = n142 & n21387 ;
  assign n21389 = n20533 & n72388 ;
  assign n21390 = n21317 & n21389 ;
  assign n21391 = n21388 | n21390 ;
  assign n21392 = n70609 & n21391 ;
  assign n72418 = ~n21390 ;
  assign n21978 = x107 & n72418 ;
  assign n72419 = ~n21388 ;
  assign n21979 = n72419 & n21978 ;
  assign n21980 = n21392 | n21979 ;
  assign n72420 = ~n21119 ;
  assign n21123 = n72420 & n21122 ;
  assign n21393 = n20552 | n21122 ;
  assign n72421 = ~n21393 ;
  assign n21394 = n21292 & n72421 ;
  assign n21395 = n21123 | n21394 ;
  assign n21396 = n142 & n21395 ;
  assign n21397 = n20542 & n72388 ;
  assign n21398 = n21317 & n21397 ;
  assign n21399 = n21396 | n21398 ;
  assign n21400 = n70276 & n21399 ;
  assign n72422 = ~n21291 ;
  assign n21293 = n21117 & n72422 ;
  assign n21401 = n20561 | n21117 ;
  assign n72423 = ~n21401 ;
  assign n21402 = n21113 & n72423 ;
  assign n21403 = n21293 | n21402 ;
  assign n21404 = n142 & n21403 ;
  assign n21405 = n20551 & n72388 ;
  assign n21406 = n21317 & n21405 ;
  assign n21407 = n21404 | n21406 ;
  assign n21408 = n70176 & n21407 ;
  assign n72424 = ~n21406 ;
  assign n21966 = x105 & n72424 ;
  assign n72425 = ~n21404 ;
  assign n21967 = n72425 & n21966 ;
  assign n21968 = n21408 | n21967 ;
  assign n72426 = ~n21108 ;
  assign n21112 = n72426 & n21111 ;
  assign n21409 = n20570 | n21111 ;
  assign n72427 = ~n21409 ;
  assign n21410 = n21287 & n72427 ;
  assign n21411 = n21112 | n21410 ;
  assign n21412 = n142 & n21411 ;
  assign n21413 = n20560 & n72388 ;
  assign n21414 = n21317 & n21413 ;
  assign n21415 = n21412 | n21414 ;
  assign n21416 = n69857 & n21415 ;
  assign n72428 = ~n21286 ;
  assign n21288 = n21106 & n72428 ;
  assign n21417 = n20579 | n21106 ;
  assign n72429 = ~n21417 ;
  assign n21418 = n21102 & n72429 ;
  assign n21419 = n21288 | n21418 ;
  assign n21420 = n142 & n21419 ;
  assign n21421 = n20569 & n72388 ;
  assign n21422 = n21317 & n21421 ;
  assign n21423 = n21420 | n21422 ;
  assign n21424 = n69656 & n21423 ;
  assign n72430 = ~n21422 ;
  assign n21954 = x103 & n72430 ;
  assign n72431 = ~n21420 ;
  assign n21955 = n72431 & n21954 ;
  assign n21956 = n21424 | n21955 ;
  assign n72432 = ~n21097 ;
  assign n21101 = n72432 & n21100 ;
  assign n21425 = n20588 | n21100 ;
  assign n72433 = ~n21425 ;
  assign n21426 = n21282 & n72433 ;
  assign n21427 = n21101 | n21426 ;
  assign n21428 = n142 & n21427 ;
  assign n21429 = n20578 & n72388 ;
  assign n21430 = n21317 & n21429 ;
  assign n21431 = n21428 | n21430 ;
  assign n21432 = n69528 & n21431 ;
  assign n72434 = ~n21281 ;
  assign n21283 = n21095 & n72434 ;
  assign n21433 = n20597 | n21095 ;
  assign n72435 = ~n21433 ;
  assign n21434 = n21091 & n72435 ;
  assign n21435 = n21283 | n21434 ;
  assign n21436 = n142 & n21435 ;
  assign n21437 = n20587 & n72388 ;
  assign n21438 = n21317 & n21437 ;
  assign n21439 = n21436 | n21438 ;
  assign n21440 = n69261 & n21439 ;
  assign n72436 = ~n21438 ;
  assign n21942 = x101 & n72436 ;
  assign n72437 = ~n21436 ;
  assign n21943 = n72437 & n21942 ;
  assign n21944 = n21440 | n21943 ;
  assign n72438 = ~n21086 ;
  assign n21090 = n72438 & n21089 ;
  assign n21441 = n20606 | n21089 ;
  assign n72439 = ~n21441 ;
  assign n21442 = n21277 & n72439 ;
  assign n21443 = n21090 | n21442 ;
  assign n21444 = n142 & n21443 ;
  assign n21445 = n20596 & n72388 ;
  assign n21446 = n21317 & n21445 ;
  assign n21447 = n21444 | n21446 ;
  assign n21448 = n69075 & n21447 ;
  assign n72440 = ~n21276 ;
  assign n21278 = n21084 & n72440 ;
  assign n21449 = n20615 | n21084 ;
  assign n72441 = ~n21449 ;
  assign n21450 = n21080 & n72441 ;
  assign n21451 = n21278 | n21450 ;
  assign n21452 = n142 & n21451 ;
  assign n21453 = n20605 & n72388 ;
  assign n21454 = n21317 & n21453 ;
  assign n21455 = n21452 | n21454 ;
  assign n21456 = n68993 & n21455 ;
  assign n72442 = ~n21454 ;
  assign n21930 = x99 & n72442 ;
  assign n72443 = ~n21452 ;
  assign n21931 = n72443 & n21930 ;
  assign n21932 = n21456 | n21931 ;
  assign n72444 = ~n21075 ;
  assign n21079 = n72444 & n21078 ;
  assign n21457 = n20624 | n21078 ;
  assign n72445 = ~n21457 ;
  assign n21458 = n21272 & n72445 ;
  assign n21459 = n21079 | n21458 ;
  assign n21460 = n142 & n21459 ;
  assign n21461 = n20614 & n72388 ;
  assign n21462 = n21317 & n21461 ;
  assign n21463 = n21460 | n21462 ;
  assign n21464 = n68716 & n21463 ;
  assign n72446 = ~n21271 ;
  assign n21273 = n21073 & n72446 ;
  assign n21465 = n20633 | n21073 ;
  assign n72447 = ~n21465 ;
  assign n21466 = n21069 & n72447 ;
  assign n21467 = n21273 | n21466 ;
  assign n21468 = n142 & n21467 ;
  assign n21469 = n20623 & n72388 ;
  assign n21470 = n21317 & n21469 ;
  assign n21471 = n21468 | n21470 ;
  assign n21472 = n68545 & n21471 ;
  assign n72448 = ~n21470 ;
  assign n21918 = x97 & n72448 ;
  assign n72449 = ~n21468 ;
  assign n21919 = n72449 & n21918 ;
  assign n21920 = n21472 | n21919 ;
  assign n72450 = ~n21064 ;
  assign n21068 = n72450 & n21067 ;
  assign n21473 = n20642 | n21067 ;
  assign n72451 = ~n21473 ;
  assign n21474 = n21267 & n72451 ;
  assign n21475 = n21068 | n21474 ;
  assign n21476 = n142 & n21475 ;
  assign n21477 = n20632 & n72388 ;
  assign n21478 = n21317 & n21477 ;
  assign n21479 = n21476 | n21478 ;
  assign n21480 = n68438 & n21479 ;
  assign n72452 = ~n21266 ;
  assign n21268 = n21062 & n72452 ;
  assign n21481 = n20651 | n21062 ;
  assign n72453 = ~n21481 ;
  assign n21482 = n21058 & n72453 ;
  assign n21483 = n21268 | n21482 ;
  assign n21484 = n142 & n21483 ;
  assign n21485 = n20641 & n72388 ;
  assign n21486 = n21317 & n21485 ;
  assign n21487 = n21484 | n21486 ;
  assign n21488 = n68214 & n21487 ;
  assign n72454 = ~n21486 ;
  assign n21906 = x95 & n72454 ;
  assign n72455 = ~n21484 ;
  assign n21907 = n72455 & n21906 ;
  assign n21908 = n21488 | n21907 ;
  assign n72456 = ~n21053 ;
  assign n21057 = n72456 & n21056 ;
  assign n21489 = n20660 | n21056 ;
  assign n72457 = ~n21489 ;
  assign n21490 = n21262 & n72457 ;
  assign n21491 = n21057 | n21490 ;
  assign n21492 = n142 & n21491 ;
  assign n21493 = n20650 & n72388 ;
  assign n21494 = n21317 & n21493 ;
  assign n21495 = n21492 | n21494 ;
  assign n21496 = n68058 & n21495 ;
  assign n72458 = ~n21261 ;
  assign n21263 = n21051 & n72458 ;
  assign n21497 = n20669 | n21051 ;
  assign n72459 = ~n21497 ;
  assign n21498 = n21047 & n72459 ;
  assign n21499 = n21263 | n21498 ;
  assign n21500 = n142 & n21499 ;
  assign n21501 = n20659 & n72388 ;
  assign n21502 = n21317 & n21501 ;
  assign n21503 = n21500 | n21502 ;
  assign n21504 = n67986 & n21503 ;
  assign n72460 = ~n21502 ;
  assign n21894 = x93 & n72460 ;
  assign n72461 = ~n21500 ;
  assign n21895 = n72461 & n21894 ;
  assign n21896 = n21504 | n21895 ;
  assign n72462 = ~n21042 ;
  assign n21046 = n72462 & n21045 ;
  assign n21505 = n20678 | n21045 ;
  assign n72463 = ~n21505 ;
  assign n21506 = n21257 & n72463 ;
  assign n21507 = n21046 | n21506 ;
  assign n21508 = n142 & n21507 ;
  assign n21509 = n20668 & n72388 ;
  assign n21510 = n21317 & n21509 ;
  assign n21511 = n21508 | n21510 ;
  assign n21512 = n67763 & n21511 ;
  assign n72464 = ~n21256 ;
  assign n21258 = n21040 & n72464 ;
  assign n21513 = n20687 | n21040 ;
  assign n72465 = ~n21513 ;
  assign n21514 = n21036 & n72465 ;
  assign n21515 = n21258 | n21514 ;
  assign n21516 = n142 & n21515 ;
  assign n21517 = n20677 & n72388 ;
  assign n21518 = n21317 & n21517 ;
  assign n21519 = n21516 | n21518 ;
  assign n21520 = n67622 & n21519 ;
  assign n72466 = ~n21518 ;
  assign n21882 = x91 & n72466 ;
  assign n72467 = ~n21516 ;
  assign n21883 = n72467 & n21882 ;
  assign n21884 = n21520 | n21883 ;
  assign n72468 = ~n21031 ;
  assign n21035 = n72468 & n21034 ;
  assign n21521 = n20696 | n21034 ;
  assign n72469 = ~n21521 ;
  assign n21522 = n21252 & n72469 ;
  assign n21523 = n21035 | n21522 ;
  assign n21524 = n142 & n21523 ;
  assign n21525 = n20686 & n72388 ;
  assign n21526 = n21317 & n21525 ;
  assign n21527 = n21524 | n21526 ;
  assign n21528 = n67531 & n21527 ;
  assign n72470 = ~n21251 ;
  assign n21253 = n21029 & n72470 ;
  assign n21529 = n20704 | n21029 ;
  assign n72471 = ~n21529 ;
  assign n21530 = n21025 & n72471 ;
  assign n21531 = n21253 | n21530 ;
  assign n21532 = n142 & n21531 ;
  assign n21533 = n20695 & n72388 ;
  assign n21534 = n21317 & n21533 ;
  assign n21535 = n21532 | n21534 ;
  assign n21536 = n67348 & n21535 ;
  assign n72472 = ~n21534 ;
  assign n21870 = x89 & n72472 ;
  assign n72473 = ~n21532 ;
  assign n21871 = n72473 & n21870 ;
  assign n21872 = n21536 | n21871 ;
  assign n72474 = ~n21020 ;
  assign n21024 = n72474 & n21023 ;
  assign n21537 = n20713 | n21023 ;
  assign n72475 = ~n21537 ;
  assign n21538 = n21247 & n72475 ;
  assign n21539 = n21024 | n21538 ;
  assign n21540 = n142 & n21539 ;
  assign n21541 = n20703 & n72388 ;
  assign n21542 = n21317 & n21541 ;
  assign n21543 = n21540 | n21542 ;
  assign n21544 = n67222 & n21543 ;
  assign n72476 = ~n21246 ;
  assign n21248 = n21018 & n72476 ;
  assign n21545 = n20722 | n21018 ;
  assign n72477 = ~n21545 ;
  assign n21546 = n21014 & n72477 ;
  assign n21547 = n21248 | n21546 ;
  assign n21548 = n142 & n21547 ;
  assign n21549 = n20712 & n72388 ;
  assign n21550 = n21317 & n21549 ;
  assign n21551 = n21548 | n21550 ;
  assign n21552 = n67164 & n21551 ;
  assign n72478 = ~n21550 ;
  assign n21858 = x87 & n72478 ;
  assign n72479 = ~n21548 ;
  assign n21859 = n72479 & n21858 ;
  assign n21860 = n21552 | n21859 ;
  assign n72480 = ~n21009 ;
  assign n21013 = n72480 & n21012 ;
  assign n21553 = n20731 | n21012 ;
  assign n72481 = ~n21553 ;
  assign n21554 = n21242 & n72481 ;
  assign n21555 = n21013 | n21554 ;
  assign n21556 = n142 & n21555 ;
  assign n21557 = n20721 & n72388 ;
  assign n21558 = n21317 & n21557 ;
  assign n21559 = n21556 | n21558 ;
  assign n21560 = n66979 & n21559 ;
  assign n72482 = ~n21241 ;
  assign n21243 = n21007 & n72482 ;
  assign n21561 = n20739 | n21007 ;
  assign n72483 = ~n21561 ;
  assign n21562 = n21003 & n72483 ;
  assign n21563 = n21243 | n21562 ;
  assign n21564 = n142 & n21563 ;
  assign n21565 = n20730 & n72388 ;
  assign n21566 = n21317 & n21565 ;
  assign n21567 = n21564 | n21566 ;
  assign n21568 = n66868 & n21567 ;
  assign n72484 = ~n21566 ;
  assign n21846 = x85 & n72484 ;
  assign n72485 = ~n21564 ;
  assign n21847 = n72485 & n21846 ;
  assign n21848 = n21568 | n21847 ;
  assign n72486 = ~n20998 ;
  assign n21002 = n72486 & n21001 ;
  assign n21569 = n20748 | n21001 ;
  assign n72487 = ~n21569 ;
  assign n21570 = n21237 & n72487 ;
  assign n21571 = n21002 | n21570 ;
  assign n21572 = n142 & n21571 ;
  assign n21573 = n20738 & n72388 ;
  assign n21574 = n21317 & n21573 ;
  assign n21575 = n21572 | n21574 ;
  assign n21576 = n66797 & n21575 ;
  assign n72488 = ~n21236 ;
  assign n21238 = n20996 & n72488 ;
  assign n21577 = n20756 | n20996 ;
  assign n72489 = ~n21577 ;
  assign n21578 = n20992 & n72489 ;
  assign n21579 = n21238 | n21578 ;
  assign n21580 = n142 & n21579 ;
  assign n21581 = n20747 & n72388 ;
  assign n21582 = n21317 & n21581 ;
  assign n21583 = n21580 | n21582 ;
  assign n21584 = n66654 & n21583 ;
  assign n72490 = ~n21582 ;
  assign n21834 = x83 & n72490 ;
  assign n72491 = ~n21580 ;
  assign n21835 = n72491 & n21834 ;
  assign n21836 = n21584 | n21835 ;
  assign n72492 = ~n20987 ;
  assign n20991 = n72492 & n20990 ;
  assign n21585 = n20765 | n20990 ;
  assign n72493 = ~n21585 ;
  assign n21586 = n21232 & n72493 ;
  assign n21587 = n20991 | n21586 ;
  assign n21588 = n142 & n21587 ;
  assign n21589 = n20755 & n72388 ;
  assign n21590 = n21317 & n21589 ;
  assign n21591 = n21588 | n21590 ;
  assign n21592 = n66560 & n21591 ;
  assign n72494 = ~n21231 ;
  assign n21233 = n20985 & n72494 ;
  assign n21593 = n20774 | n20985 ;
  assign n72495 = ~n21593 ;
  assign n21594 = n20981 & n72495 ;
  assign n21595 = n21233 | n21594 ;
  assign n21596 = n142 & n21595 ;
  assign n21597 = n20764 & n72388 ;
  assign n21598 = n21317 & n21597 ;
  assign n21599 = n21596 | n21598 ;
  assign n21600 = n66505 & n21599 ;
  assign n72496 = ~n21598 ;
  assign n21822 = x81 & n72496 ;
  assign n72497 = ~n21596 ;
  assign n21823 = n72497 & n21822 ;
  assign n21824 = n21600 | n21823 ;
  assign n72498 = ~n20976 ;
  assign n20980 = n72498 & n20979 ;
  assign n21601 = n20783 | n20979 ;
  assign n72499 = ~n21601 ;
  assign n21602 = n21227 & n72499 ;
  assign n21603 = n20980 | n21602 ;
  assign n21604 = n142 & n21603 ;
  assign n21605 = n20773 & n72388 ;
  assign n21606 = n21317 & n21605 ;
  assign n21607 = n21604 | n21606 ;
  assign n21608 = n66379 & n21607 ;
  assign n72500 = ~n21226 ;
  assign n21228 = n20974 & n72500 ;
  assign n21609 = n20792 | n20974 ;
  assign n72501 = ~n21609 ;
  assign n21610 = n20970 & n72501 ;
  assign n21611 = n21228 | n21610 ;
  assign n21612 = n142 & n21611 ;
  assign n21613 = n20782 & n72388 ;
  assign n21614 = n21317 & n21613 ;
  assign n21615 = n21612 | n21614 ;
  assign n21616 = n66299 & n21615 ;
  assign n72502 = ~n21614 ;
  assign n21810 = x79 & n72502 ;
  assign n72503 = ~n21612 ;
  assign n21811 = n72503 & n21810 ;
  assign n21812 = n21616 | n21811 ;
  assign n72504 = ~n20965 ;
  assign n20969 = n72504 & n20968 ;
  assign n21617 = n20801 | n20968 ;
  assign n72505 = ~n21617 ;
  assign n21618 = n21222 & n72505 ;
  assign n21619 = n20969 | n21618 ;
  assign n21620 = n142 & n21619 ;
  assign n21621 = n20791 & n72388 ;
  assign n21622 = n21317 & n21621 ;
  assign n21623 = n21620 | n21622 ;
  assign n21624 = n66244 & n21623 ;
  assign n72506 = ~n21221 ;
  assign n21223 = n20963 & n72506 ;
  assign n21625 = n20810 | n20963 ;
  assign n72507 = ~n21625 ;
  assign n21626 = n20959 & n72507 ;
  assign n21627 = n21223 | n21626 ;
  assign n21628 = n142 & n21627 ;
  assign n21629 = n20800 & n72388 ;
  assign n21630 = n21317 & n21629 ;
  assign n21631 = n21628 | n21630 ;
  assign n21632 = n66145 & n21631 ;
  assign n72508 = ~n21630 ;
  assign n21798 = x77 & n72508 ;
  assign n72509 = ~n21628 ;
  assign n21799 = n72509 & n21798 ;
  assign n21800 = n21632 | n21799 ;
  assign n72510 = ~n20954 ;
  assign n20958 = n72510 & n20957 ;
  assign n21633 = n20819 | n20957 ;
  assign n72511 = ~n21633 ;
  assign n21634 = n21217 & n72511 ;
  assign n21635 = n20958 | n21634 ;
  assign n21636 = n142 & n21635 ;
  assign n21637 = n20809 & n72388 ;
  assign n21638 = n21317 & n21637 ;
  assign n21639 = n21636 | n21638 ;
  assign n21640 = n66081 & n21639 ;
  assign n72512 = ~n21216 ;
  assign n21218 = n20952 & n72512 ;
  assign n21641 = n20828 | n20952 ;
  assign n72513 = ~n21641 ;
  assign n21642 = n20948 & n72513 ;
  assign n21643 = n21218 | n21642 ;
  assign n21644 = n142 & n21643 ;
  assign n21645 = n20818 & n72388 ;
  assign n21646 = n21317 & n21645 ;
  assign n21647 = n21644 | n21646 ;
  assign n21648 = n66043 & n21647 ;
  assign n72514 = ~n21646 ;
  assign n21786 = x75 & n72514 ;
  assign n72515 = ~n21644 ;
  assign n21787 = n72515 & n21786 ;
  assign n21788 = n21648 | n21787 ;
  assign n72516 = ~n20943 ;
  assign n20947 = n72516 & n20946 ;
  assign n21649 = n20836 | n20946 ;
  assign n72517 = ~n21649 ;
  assign n21650 = n21212 & n72517 ;
  assign n21651 = n20947 | n21650 ;
  assign n21652 = n142 & n21651 ;
  assign n21653 = n20827 & n72388 ;
  assign n21654 = n21317 & n21653 ;
  assign n21655 = n21652 | n21654 ;
  assign n21656 = n65960 & n21655 ;
  assign n72518 = ~n21211 ;
  assign n21213 = n20941 & n72518 ;
  assign n21657 = n20845 | n20941 ;
  assign n72519 = ~n21657 ;
  assign n21658 = n20937 & n72519 ;
  assign n21659 = n21213 | n21658 ;
  assign n21660 = n142 & n21659 ;
  assign n21661 = n20835 & n72388 ;
  assign n21662 = n21317 & n21661 ;
  assign n21663 = n21660 | n21662 ;
  assign n21664 = n65909 & n21663 ;
  assign n72520 = ~n21662 ;
  assign n21774 = x73 & n72520 ;
  assign n72521 = ~n21660 ;
  assign n21775 = n72521 & n21774 ;
  assign n21776 = n21664 | n21775 ;
  assign n72522 = ~n20932 ;
  assign n20936 = n72522 & n20935 ;
  assign n21665 = n20854 | n20935 ;
  assign n72523 = ~n21665 ;
  assign n21666 = n21207 & n72523 ;
  assign n21667 = n20936 | n21666 ;
  assign n21668 = n142 & n21667 ;
  assign n21669 = n20844 & n72388 ;
  assign n21670 = n21317 & n21669 ;
  assign n21671 = n21668 | n21670 ;
  assign n21672 = n65877 & n21671 ;
  assign n72524 = ~n21206 ;
  assign n21208 = n20930 & n72524 ;
  assign n21673 = n20863 | n20930 ;
  assign n72525 = ~n21673 ;
  assign n21674 = n20926 & n72525 ;
  assign n21675 = n21208 | n21674 ;
  assign n21676 = n142 & n21675 ;
  assign n21677 = n20853 & n72388 ;
  assign n21678 = n21317 & n21677 ;
  assign n21679 = n21676 | n21678 ;
  assign n21680 = n65820 & n21679 ;
  assign n72526 = ~n21678 ;
  assign n21762 = x71 & n72526 ;
  assign n72527 = ~n21676 ;
  assign n21763 = n72527 & n21762 ;
  assign n21764 = n21680 | n21763 ;
  assign n72528 = ~n20921 ;
  assign n20925 = n72528 & n20924 ;
  assign n21681 = n20872 | n20924 ;
  assign n72529 = ~n21681 ;
  assign n21682 = n21203 & n72529 ;
  assign n21683 = n20925 | n21682 ;
  assign n21684 = n142 & n21683 ;
  assign n21685 = n20862 & n72388 ;
  assign n21686 = n21317 & n21685 ;
  assign n21687 = n21684 | n21686 ;
  assign n21688 = n65791 & n21687 ;
  assign n72530 = ~n21201 ;
  assign n21202 = n20919 & n72530 ;
  assign n21689 = n20881 | n20919 ;
  assign n72531 = ~n21689 ;
  assign n21690 = n20915 & n72531 ;
  assign n21691 = n21202 | n21690 ;
  assign n21692 = n142 & n21691 ;
  assign n21693 = n20871 & n72388 ;
  assign n21694 = n21317 & n21693 ;
  assign n21695 = n21692 | n21694 ;
  assign n21696 = n65772 & n21695 ;
  assign n72532 = ~n21694 ;
  assign n21751 = x69 & n72532 ;
  assign n72533 = ~n21692 ;
  assign n21752 = n72533 & n21751 ;
  assign n21753 = n21696 | n21752 ;
  assign n72534 = ~n20911 ;
  assign n21199 = n72534 & n20914 ;
  assign n21697 = n20889 | n20914 ;
  assign n72535 = ~n21697 ;
  assign n21698 = n20910 & n72535 ;
  assign n21699 = n21199 | n21698 ;
  assign n21700 = n142 & n21699 ;
  assign n21701 = n20880 & n72388 ;
  assign n21702 = n21317 & n21701 ;
  assign n21703 = n21700 | n21702 ;
  assign n21704 = n65746 & n21703 ;
  assign n72536 = ~n20906 ;
  assign n21706 = n72536 & n20909 ;
  assign n21705 = n20905 | n20909 ;
  assign n72537 = ~n21705 ;
  assign n21707 = n20904 & n72537 ;
  assign n21708 = n21706 | n21707 ;
  assign n21709 = n142 & n21708 ;
  assign n21710 = n20888 & n72388 ;
  assign n21711 = n21317 & n21710 ;
  assign n21712 = n21709 | n21711 ;
  assign n21713 = n65721 & n21712 ;
  assign n72538 = ~n21711 ;
  assign n21741 = x67 & n72538 ;
  assign n72539 = ~n21709 ;
  assign n21742 = n72539 & n21741 ;
  assign n21743 = n21713 | n21742 ;
  assign n21714 = n20901 & n20903 ;
  assign n21715 = n72238 & n21714 ;
  assign n72540 = ~n21715 ;
  assign n21716 = n21195 & n72540 ;
  assign n21717 = n142 & n21716 ;
  assign n21718 = n20898 & n72388 ;
  assign n21719 = n21317 & n21718 ;
  assign n21720 = n21717 | n21719 ;
  assign n21721 = n65686 & n21720 ;
  assign n72541 = ~x12 ;
  assign n21731 = n72541 & x64 ;
  assign n21190 = n20903 & n142 ;
  assign n21722 = n72388 & n21317 ;
  assign n72542 = ~n21722 ;
  assign n21723 = x64 & n72542 ;
  assign n72543 = ~n21723 ;
  assign n21724 = x13 & n72543 ;
  assign n21725 = n21190 | n21724 ;
  assign n21726 = x65 & n21725 ;
  assign n21191 = x64 & n142 ;
  assign n72544 = ~n21191 ;
  assign n21727 = x13 & n72544 ;
  assign n21728 = n20903 & n72542 ;
  assign n21729 = x65 | n21728 ;
  assign n21730 = n21727 | n21729 ;
  assign n72545 = ~n21726 ;
  assign n21732 = n72545 & n21730 ;
  assign n21733 = n21731 | n21732 ;
  assign n21734 = n21190 | n21727 ;
  assign n21735 = n65670 & n21734 ;
  assign n72546 = ~n21735 ;
  assign n21736 = n21733 & n72546 ;
  assign n72547 = ~n21719 ;
  assign n21737 = x66 & n72547 ;
  assign n72548 = ~n21717 ;
  assign n21738 = n72548 & n21737 ;
  assign n21739 = n21721 | n21738 ;
  assign n21740 = n21736 | n21739 ;
  assign n72549 = ~n21721 ;
  assign n21744 = n72549 & n21740 ;
  assign n21745 = n21743 | n21744 ;
  assign n72550 = ~n21713 ;
  assign n21746 = n72550 & n21745 ;
  assign n72551 = ~n21702 ;
  assign n21747 = x68 & n72551 ;
  assign n72552 = ~n21700 ;
  assign n21748 = n72552 & n21747 ;
  assign n21749 = n21704 | n21748 ;
  assign n21750 = n21746 | n21749 ;
  assign n72553 = ~n21704 ;
  assign n21754 = n72553 & n21750 ;
  assign n21755 = n21753 | n21754 ;
  assign n72554 = ~n21696 ;
  assign n21756 = n72554 & n21755 ;
  assign n72555 = ~n21686 ;
  assign n21757 = x70 & n72555 ;
  assign n72556 = ~n21684 ;
  assign n21758 = n72556 & n21757 ;
  assign n21759 = n21688 | n21758 ;
  assign n21761 = n21756 | n21759 ;
  assign n72557 = ~n21688 ;
  assign n21766 = n72557 & n21761 ;
  assign n21767 = n21764 | n21766 ;
  assign n72558 = ~n21680 ;
  assign n21768 = n72558 & n21767 ;
  assign n72559 = ~n21670 ;
  assign n21769 = x72 & n72559 ;
  assign n72560 = ~n21668 ;
  assign n21770 = n72560 & n21769 ;
  assign n21771 = n21672 | n21770 ;
  assign n21773 = n21768 | n21771 ;
  assign n72561 = ~n21672 ;
  assign n21778 = n72561 & n21773 ;
  assign n21779 = n21776 | n21778 ;
  assign n72562 = ~n21664 ;
  assign n21780 = n72562 & n21779 ;
  assign n72563 = ~n21654 ;
  assign n21781 = x74 & n72563 ;
  assign n72564 = ~n21652 ;
  assign n21782 = n72564 & n21781 ;
  assign n21783 = n21656 | n21782 ;
  assign n21785 = n21780 | n21783 ;
  assign n72565 = ~n21656 ;
  assign n21790 = n72565 & n21785 ;
  assign n21791 = n21788 | n21790 ;
  assign n72566 = ~n21648 ;
  assign n21792 = n72566 & n21791 ;
  assign n72567 = ~n21638 ;
  assign n21793 = x76 & n72567 ;
  assign n72568 = ~n21636 ;
  assign n21794 = n72568 & n21793 ;
  assign n21795 = n21640 | n21794 ;
  assign n21797 = n21792 | n21795 ;
  assign n72569 = ~n21640 ;
  assign n21802 = n72569 & n21797 ;
  assign n21803 = n21800 | n21802 ;
  assign n72570 = ~n21632 ;
  assign n21804 = n72570 & n21803 ;
  assign n72571 = ~n21622 ;
  assign n21805 = x78 & n72571 ;
  assign n72572 = ~n21620 ;
  assign n21806 = n72572 & n21805 ;
  assign n21807 = n21624 | n21806 ;
  assign n21809 = n21804 | n21807 ;
  assign n72573 = ~n21624 ;
  assign n21814 = n72573 & n21809 ;
  assign n21815 = n21812 | n21814 ;
  assign n72574 = ~n21616 ;
  assign n21816 = n72574 & n21815 ;
  assign n72575 = ~n21606 ;
  assign n21817 = x80 & n72575 ;
  assign n72576 = ~n21604 ;
  assign n21818 = n72576 & n21817 ;
  assign n21819 = n21608 | n21818 ;
  assign n21821 = n21816 | n21819 ;
  assign n72577 = ~n21608 ;
  assign n21826 = n72577 & n21821 ;
  assign n21827 = n21824 | n21826 ;
  assign n72578 = ~n21600 ;
  assign n21828 = n72578 & n21827 ;
  assign n72579 = ~n21590 ;
  assign n21829 = x82 & n72579 ;
  assign n72580 = ~n21588 ;
  assign n21830 = n72580 & n21829 ;
  assign n21831 = n21592 | n21830 ;
  assign n21833 = n21828 | n21831 ;
  assign n72581 = ~n21592 ;
  assign n21838 = n72581 & n21833 ;
  assign n21839 = n21836 | n21838 ;
  assign n72582 = ~n21584 ;
  assign n21840 = n72582 & n21839 ;
  assign n72583 = ~n21574 ;
  assign n21841 = x84 & n72583 ;
  assign n72584 = ~n21572 ;
  assign n21842 = n72584 & n21841 ;
  assign n21843 = n21576 | n21842 ;
  assign n21845 = n21840 | n21843 ;
  assign n72585 = ~n21576 ;
  assign n21850 = n72585 & n21845 ;
  assign n21851 = n21848 | n21850 ;
  assign n72586 = ~n21568 ;
  assign n21852 = n72586 & n21851 ;
  assign n72587 = ~n21558 ;
  assign n21853 = x86 & n72587 ;
  assign n72588 = ~n21556 ;
  assign n21854 = n72588 & n21853 ;
  assign n21855 = n21560 | n21854 ;
  assign n21857 = n21852 | n21855 ;
  assign n72589 = ~n21560 ;
  assign n21862 = n72589 & n21857 ;
  assign n21863 = n21860 | n21862 ;
  assign n72590 = ~n21552 ;
  assign n21864 = n72590 & n21863 ;
  assign n72591 = ~n21542 ;
  assign n21865 = x88 & n72591 ;
  assign n72592 = ~n21540 ;
  assign n21866 = n72592 & n21865 ;
  assign n21867 = n21544 | n21866 ;
  assign n21869 = n21864 | n21867 ;
  assign n72593 = ~n21544 ;
  assign n21874 = n72593 & n21869 ;
  assign n21875 = n21872 | n21874 ;
  assign n72594 = ~n21536 ;
  assign n21876 = n72594 & n21875 ;
  assign n72595 = ~n21526 ;
  assign n21877 = x90 & n72595 ;
  assign n72596 = ~n21524 ;
  assign n21878 = n72596 & n21877 ;
  assign n21879 = n21528 | n21878 ;
  assign n21881 = n21876 | n21879 ;
  assign n72597 = ~n21528 ;
  assign n21886 = n72597 & n21881 ;
  assign n21887 = n21884 | n21886 ;
  assign n72598 = ~n21520 ;
  assign n21888 = n72598 & n21887 ;
  assign n72599 = ~n21510 ;
  assign n21889 = x92 & n72599 ;
  assign n72600 = ~n21508 ;
  assign n21890 = n72600 & n21889 ;
  assign n21891 = n21512 | n21890 ;
  assign n21893 = n21888 | n21891 ;
  assign n72601 = ~n21512 ;
  assign n21898 = n72601 & n21893 ;
  assign n21899 = n21896 | n21898 ;
  assign n72602 = ~n21504 ;
  assign n21900 = n72602 & n21899 ;
  assign n72603 = ~n21494 ;
  assign n21901 = x94 & n72603 ;
  assign n72604 = ~n21492 ;
  assign n21902 = n72604 & n21901 ;
  assign n21903 = n21496 | n21902 ;
  assign n21905 = n21900 | n21903 ;
  assign n72605 = ~n21496 ;
  assign n21910 = n72605 & n21905 ;
  assign n21911 = n21908 | n21910 ;
  assign n72606 = ~n21488 ;
  assign n21912 = n72606 & n21911 ;
  assign n72607 = ~n21478 ;
  assign n21913 = x96 & n72607 ;
  assign n72608 = ~n21476 ;
  assign n21914 = n72608 & n21913 ;
  assign n21915 = n21480 | n21914 ;
  assign n21917 = n21912 | n21915 ;
  assign n72609 = ~n21480 ;
  assign n21922 = n72609 & n21917 ;
  assign n21923 = n21920 | n21922 ;
  assign n72610 = ~n21472 ;
  assign n21924 = n72610 & n21923 ;
  assign n72611 = ~n21462 ;
  assign n21925 = x98 & n72611 ;
  assign n72612 = ~n21460 ;
  assign n21926 = n72612 & n21925 ;
  assign n21927 = n21464 | n21926 ;
  assign n21929 = n21924 | n21927 ;
  assign n72613 = ~n21464 ;
  assign n21934 = n72613 & n21929 ;
  assign n21935 = n21932 | n21934 ;
  assign n72614 = ~n21456 ;
  assign n21936 = n72614 & n21935 ;
  assign n72615 = ~n21446 ;
  assign n21937 = x100 & n72615 ;
  assign n72616 = ~n21444 ;
  assign n21938 = n72616 & n21937 ;
  assign n21939 = n21448 | n21938 ;
  assign n21941 = n21936 | n21939 ;
  assign n72617 = ~n21448 ;
  assign n21946 = n72617 & n21941 ;
  assign n21947 = n21944 | n21946 ;
  assign n72618 = ~n21440 ;
  assign n21948 = n72618 & n21947 ;
  assign n72619 = ~n21430 ;
  assign n21949 = x102 & n72619 ;
  assign n72620 = ~n21428 ;
  assign n21950 = n72620 & n21949 ;
  assign n21951 = n21432 | n21950 ;
  assign n21953 = n21948 | n21951 ;
  assign n72621 = ~n21432 ;
  assign n21958 = n72621 & n21953 ;
  assign n21959 = n21956 | n21958 ;
  assign n72622 = ~n21424 ;
  assign n21960 = n72622 & n21959 ;
  assign n72623 = ~n21414 ;
  assign n21961 = x104 & n72623 ;
  assign n72624 = ~n21412 ;
  assign n21962 = n72624 & n21961 ;
  assign n21963 = n21416 | n21962 ;
  assign n21965 = n21960 | n21963 ;
  assign n72625 = ~n21416 ;
  assign n21970 = n72625 & n21965 ;
  assign n21971 = n21968 | n21970 ;
  assign n72626 = ~n21408 ;
  assign n21972 = n72626 & n21971 ;
  assign n72627 = ~n21398 ;
  assign n21973 = x106 & n72627 ;
  assign n72628 = ~n21396 ;
  assign n21974 = n72628 & n21973 ;
  assign n21975 = n21400 | n21974 ;
  assign n21977 = n21972 | n21975 ;
  assign n72629 = ~n21400 ;
  assign n21982 = n72629 & n21977 ;
  assign n21983 = n21980 | n21982 ;
  assign n72630 = ~n21392 ;
  assign n21984 = n72630 & n21983 ;
  assign n72631 = ~n21382 ;
  assign n21985 = x108 & n72631 ;
  assign n72632 = ~n21380 ;
  assign n21986 = n72632 & n21985 ;
  assign n21987 = n21384 | n21986 ;
  assign n21989 = n21984 | n21987 ;
  assign n72633 = ~n21384 ;
  assign n21994 = n72633 & n21989 ;
  assign n21995 = n21992 | n21994 ;
  assign n72634 = ~n21376 ;
  assign n21996 = n72634 & n21995 ;
  assign n72635 = ~n21366 ;
  assign n21997 = x110 & n72635 ;
  assign n72636 = ~n21364 ;
  assign n21998 = n72636 & n21997 ;
  assign n21999 = n21368 | n21998 ;
  assign n22001 = n21996 | n21999 ;
  assign n72637 = ~n21368 ;
  assign n22006 = n72637 & n22001 ;
  assign n22007 = n22004 | n22006 ;
  assign n72638 = ~n21360 ;
  assign n22008 = n72638 & n22007 ;
  assign n72639 = ~n21350 ;
  assign n22009 = x112 & n72639 ;
  assign n72640 = ~n21348 ;
  assign n22010 = n72640 & n22009 ;
  assign n22011 = n21352 | n22010 ;
  assign n22013 = n22008 | n22011 ;
  assign n72641 = ~n21352 ;
  assign n22018 = n72641 & n22013 ;
  assign n22019 = n22016 | n22018 ;
  assign n72642 = ~n21344 ;
  assign n22020 = n72642 & n22019 ;
  assign n72643 = ~n21334 ;
  assign n22021 = x114 & n72643 ;
  assign n72644 = ~n21332 ;
  assign n22022 = n72644 & n22021 ;
  assign n22023 = n21336 | n22022 ;
  assign n22025 = n22020 | n22023 ;
  assign n72645 = ~n21336 ;
  assign n22029 = n72645 & n22025 ;
  assign n22030 = n22028 | n22029 ;
  assign n72646 = ~n21328 ;
  assign n22031 = n72646 & n22030 ;
  assign n22032 = n65429 | n22031 ;
  assign n72647 = ~n21327 ;
  assign n22033 = n72647 & n22032 ;
  assign n72648 = ~n22029 ;
  assign n22833 = n22028 & n72648 ;
  assign n22037 = x65 & n21734 ;
  assign n72649 = ~n22037 ;
  assign n22038 = n21730 & n72649 ;
  assign n22040 = n21731 | n22038 ;
  assign n22042 = n72546 & n22040 ;
  assign n22043 = n21739 | n22042 ;
  assign n22044 = n72549 & n22043 ;
  assign n22045 = n21743 | n22044 ;
  assign n22046 = n72550 & n22045 ;
  assign n22047 = n21749 | n22046 ;
  assign n22048 = n72553 & n22047 ;
  assign n22049 = n21753 | n22048 ;
  assign n22050 = n72554 & n22049 ;
  assign n22051 = n21759 | n22050 ;
  assign n22052 = n72557 & n22051 ;
  assign n22053 = n21764 | n22052 ;
  assign n22054 = n72558 & n22053 ;
  assign n22055 = n21771 | n22054 ;
  assign n22056 = n72561 & n22055 ;
  assign n22057 = n21776 | n22056 ;
  assign n22058 = n72562 & n22057 ;
  assign n22059 = n21783 | n22058 ;
  assign n22060 = n72565 & n22059 ;
  assign n22061 = n21788 | n22060 ;
  assign n22062 = n72566 & n22061 ;
  assign n22063 = n21795 | n22062 ;
  assign n22064 = n72569 & n22063 ;
  assign n22065 = n21800 | n22064 ;
  assign n22066 = n72570 & n22065 ;
  assign n22067 = n21807 | n22066 ;
  assign n22068 = n72573 & n22067 ;
  assign n22069 = n21812 | n22068 ;
  assign n22070 = n72574 & n22069 ;
  assign n22071 = n21819 | n22070 ;
  assign n22072 = n72577 & n22071 ;
  assign n22073 = n21824 | n22072 ;
  assign n22074 = n72578 & n22073 ;
  assign n22075 = n21831 | n22074 ;
  assign n22076 = n72581 & n22075 ;
  assign n22077 = n21836 | n22076 ;
  assign n22078 = n72582 & n22077 ;
  assign n22079 = n21843 | n22078 ;
  assign n22080 = n72585 & n22079 ;
  assign n22081 = n21848 | n22080 ;
  assign n22082 = n72586 & n22081 ;
  assign n22083 = n21855 | n22082 ;
  assign n22084 = n72589 & n22083 ;
  assign n22085 = n21860 | n22084 ;
  assign n22086 = n72590 & n22085 ;
  assign n22087 = n21867 | n22086 ;
  assign n22088 = n72593 & n22087 ;
  assign n22089 = n21872 | n22088 ;
  assign n22090 = n72594 & n22089 ;
  assign n22091 = n21879 | n22090 ;
  assign n22092 = n72597 & n22091 ;
  assign n22093 = n21884 | n22092 ;
  assign n22094 = n72598 & n22093 ;
  assign n22095 = n21891 | n22094 ;
  assign n22096 = n72601 & n22095 ;
  assign n22097 = n21896 | n22096 ;
  assign n22098 = n72602 & n22097 ;
  assign n22099 = n21903 | n22098 ;
  assign n22100 = n72605 & n22099 ;
  assign n22101 = n21908 | n22100 ;
  assign n22102 = n72606 & n22101 ;
  assign n22103 = n21915 | n22102 ;
  assign n22104 = n72609 & n22103 ;
  assign n22105 = n21920 | n22104 ;
  assign n22106 = n72610 & n22105 ;
  assign n22107 = n21927 | n22106 ;
  assign n22108 = n72613 & n22107 ;
  assign n22109 = n21932 | n22108 ;
  assign n22110 = n72614 & n22109 ;
  assign n22111 = n21939 | n22110 ;
  assign n22112 = n72617 & n22111 ;
  assign n22113 = n21944 | n22112 ;
  assign n22114 = n72618 & n22113 ;
  assign n22115 = n21951 | n22114 ;
  assign n22116 = n72621 & n22115 ;
  assign n22117 = n21956 | n22116 ;
  assign n22118 = n72622 & n22117 ;
  assign n22119 = n21963 | n22118 ;
  assign n22120 = n72625 & n22119 ;
  assign n22121 = n21968 | n22120 ;
  assign n22122 = n72626 & n22121 ;
  assign n22123 = n21975 | n22122 ;
  assign n22124 = n72629 & n22123 ;
  assign n22125 = n21980 | n22124 ;
  assign n22126 = n72630 & n22125 ;
  assign n22127 = n21987 | n22126 ;
  assign n22128 = n72633 & n22127 ;
  assign n22129 = n21992 | n22128 ;
  assign n22130 = n72634 & n22129 ;
  assign n22131 = n21999 | n22130 ;
  assign n22132 = n72637 & n22131 ;
  assign n22133 = n22004 | n22132 ;
  assign n22134 = n72638 & n22133 ;
  assign n22135 = n22011 | n22134 ;
  assign n22136 = n72641 & n22135 ;
  assign n22137 = n22016 | n22136 ;
  assign n22139 = n72642 & n22137 ;
  assign n22543 = n22023 | n22139 ;
  assign n22834 = n21336 | n22028 ;
  assign n72650 = ~n22834 ;
  assign n22835 = n22543 & n72650 ;
  assign n22836 = n22833 | n22835 ;
  assign n22837 = n22032 | n22836 ;
  assign n72651 = ~n22033 ;
  assign n22838 = n72651 & n22837 ;
  assign n22846 = n67021 & n22838 ;
  assign n22035 = n21335 & n22032 ;
  assign n22024 = n21344 | n22023 ;
  assign n72652 = ~n22024 ;
  assign n22138 = n72652 & n22137 ;
  assign n72653 = ~n22139 ;
  assign n22140 = n22023 & n72653 ;
  assign n22141 = n22138 | n22140 ;
  assign n22142 = n67021 & n22141 ;
  assign n72654 = ~n22031 ;
  assign n22143 = n72654 & n22142 ;
  assign n22144 = n22035 | n22143 ;
  assign n22145 = n72393 & n22144 ;
  assign n22146 = n21343 & n22032 ;
  assign n22017 = n21352 | n22016 ;
  assign n72655 = ~n22017 ;
  assign n22147 = n22013 & n72655 ;
  assign n72656 = ~n22018 ;
  assign n22148 = n22016 & n72656 ;
  assign n22149 = n22147 | n22148 ;
  assign n22150 = n67021 & n22149 ;
  assign n22151 = n72654 & n22150 ;
  assign n22152 = n22146 | n22151 ;
  assign n22153 = n72385 & n22152 ;
  assign n22154 = n21351 & n22032 ;
  assign n22012 = n21360 | n22011 ;
  assign n72657 = ~n22012 ;
  assign n22155 = n72657 & n22133 ;
  assign n72658 = ~n22134 ;
  assign n22156 = n22011 & n72658 ;
  assign n22157 = n22155 | n22156 ;
  assign n22158 = n67021 & n22157 ;
  assign n22159 = n72654 & n22158 ;
  assign n22160 = n22154 | n22159 ;
  assign n22161 = n72025 & n22160 ;
  assign n22162 = n21359 & n22032 ;
  assign n22005 = n21368 | n22004 ;
  assign n72659 = ~n22005 ;
  assign n22163 = n22001 & n72659 ;
  assign n72660 = ~n22006 ;
  assign n22164 = n22004 & n72660 ;
  assign n22165 = n22163 | n22164 ;
  assign n22166 = n67021 & n22165 ;
  assign n22167 = n72654 & n22166 ;
  assign n22168 = n22162 | n22167 ;
  assign n22169 = n71645 & n22168 ;
  assign n22170 = n21367 & n22032 ;
  assign n22000 = n21376 | n21999 ;
  assign n72661 = ~n22000 ;
  assign n22171 = n72661 & n22129 ;
  assign n72662 = ~n22130 ;
  assign n22172 = n21999 & n72662 ;
  assign n22173 = n22171 | n22172 ;
  assign n22174 = n67021 & n22173 ;
  assign n22175 = n72654 & n22174 ;
  assign n22176 = n22170 | n22175 ;
  assign n22177 = n71633 & n22176 ;
  assign n22178 = n21375 & n22032 ;
  assign n21993 = n21384 | n21992 ;
  assign n72663 = ~n21993 ;
  assign n22179 = n21989 & n72663 ;
  assign n72664 = ~n21994 ;
  assign n22180 = n21992 & n72664 ;
  assign n22181 = n22179 | n22180 ;
  assign n22182 = n67021 & n22181 ;
  assign n22183 = n72654 & n22182 ;
  assign n22184 = n22178 | n22183 ;
  assign n22185 = n71253 & n22184 ;
  assign n22186 = n21383 & n22032 ;
  assign n21988 = n21392 | n21987 ;
  assign n72665 = ~n21988 ;
  assign n22187 = n72665 & n22125 ;
  assign n72666 = ~n22126 ;
  assign n22188 = n21987 & n72666 ;
  assign n22189 = n22187 | n22188 ;
  assign n22190 = n67021 & n22189 ;
  assign n22191 = n72654 & n22190 ;
  assign n22192 = n22186 | n22191 ;
  assign n22193 = n70935 & n22192 ;
  assign n22194 = n21391 & n22032 ;
  assign n21981 = n21400 | n21980 ;
  assign n72667 = ~n21981 ;
  assign n22195 = n21977 & n72667 ;
  assign n72668 = ~n21982 ;
  assign n22196 = n21980 & n72668 ;
  assign n22197 = n22195 | n22196 ;
  assign n22198 = n67021 & n22197 ;
  assign n22199 = n72654 & n22198 ;
  assign n22200 = n22194 | n22199 ;
  assign n22201 = n70927 & n22200 ;
  assign n22202 = n21399 & n22032 ;
  assign n21976 = n21408 | n21975 ;
  assign n72669 = ~n21976 ;
  assign n22203 = n72669 & n22121 ;
  assign n72670 = ~n22122 ;
  assign n22204 = n21975 & n72670 ;
  assign n22205 = n22203 | n22204 ;
  assign n22206 = n67021 & n22205 ;
  assign n22207 = n72654 & n22206 ;
  assign n22208 = n22202 | n22207 ;
  assign n22209 = n70609 & n22208 ;
  assign n22210 = n21407 & n22032 ;
  assign n21969 = n21416 | n21968 ;
  assign n72671 = ~n21969 ;
  assign n22211 = n21965 & n72671 ;
  assign n72672 = ~n21970 ;
  assign n22212 = n21968 & n72672 ;
  assign n22213 = n22211 | n22212 ;
  assign n22214 = n67021 & n22213 ;
  assign n22215 = n72654 & n22214 ;
  assign n22216 = n22210 | n22215 ;
  assign n22217 = n70276 & n22216 ;
  assign n22218 = n21415 & n22032 ;
  assign n21964 = n21424 | n21963 ;
  assign n72673 = ~n21964 ;
  assign n22219 = n72673 & n22117 ;
  assign n72674 = ~n22118 ;
  assign n22220 = n21963 & n72674 ;
  assign n22221 = n22219 | n22220 ;
  assign n22222 = n67021 & n22221 ;
  assign n22223 = n72654 & n22222 ;
  assign n22224 = n22218 | n22223 ;
  assign n22225 = n70176 & n22224 ;
  assign n22226 = n21423 & n22032 ;
  assign n21957 = n21432 | n21956 ;
  assign n72675 = ~n21957 ;
  assign n22227 = n21953 & n72675 ;
  assign n72676 = ~n21958 ;
  assign n22228 = n21956 & n72676 ;
  assign n22229 = n22227 | n22228 ;
  assign n22230 = n67021 & n22229 ;
  assign n22231 = n72654 & n22230 ;
  assign n22232 = n22226 | n22231 ;
  assign n22233 = n69857 & n22232 ;
  assign n22234 = n21431 & n22032 ;
  assign n21952 = n21440 | n21951 ;
  assign n72677 = ~n21952 ;
  assign n22235 = n72677 & n22113 ;
  assign n72678 = ~n22114 ;
  assign n22236 = n21951 & n72678 ;
  assign n22237 = n22235 | n22236 ;
  assign n22238 = n67021 & n22237 ;
  assign n22239 = n72654 & n22238 ;
  assign n22240 = n22234 | n22239 ;
  assign n22241 = n69656 & n22240 ;
  assign n22242 = n21439 & n22032 ;
  assign n21945 = n21448 | n21944 ;
  assign n72679 = ~n21945 ;
  assign n22243 = n21941 & n72679 ;
  assign n72680 = ~n21946 ;
  assign n22244 = n21944 & n72680 ;
  assign n22245 = n22243 | n22244 ;
  assign n22246 = n67021 & n22245 ;
  assign n22247 = n72654 & n22246 ;
  assign n22248 = n22242 | n22247 ;
  assign n22249 = n69528 & n22248 ;
  assign n22250 = n21447 & n22032 ;
  assign n21940 = n21456 | n21939 ;
  assign n72681 = ~n21940 ;
  assign n22251 = n72681 & n22109 ;
  assign n72682 = ~n22110 ;
  assign n22252 = n21939 & n72682 ;
  assign n22253 = n22251 | n22252 ;
  assign n22254 = n67021 & n22253 ;
  assign n22255 = n72654 & n22254 ;
  assign n22256 = n22250 | n22255 ;
  assign n22257 = n69261 & n22256 ;
  assign n22258 = n21455 & n22032 ;
  assign n21933 = n21464 | n21932 ;
  assign n72683 = ~n21933 ;
  assign n22259 = n21929 & n72683 ;
  assign n72684 = ~n21934 ;
  assign n22260 = n21932 & n72684 ;
  assign n22261 = n22259 | n22260 ;
  assign n22262 = n67021 & n22261 ;
  assign n22263 = n72654 & n22262 ;
  assign n22264 = n22258 | n22263 ;
  assign n22265 = n69075 & n22264 ;
  assign n22266 = n21463 & n22032 ;
  assign n21928 = n21472 | n21927 ;
  assign n72685 = ~n21928 ;
  assign n22267 = n72685 & n22105 ;
  assign n72686 = ~n22106 ;
  assign n22268 = n21927 & n72686 ;
  assign n22269 = n22267 | n22268 ;
  assign n22270 = n67021 & n22269 ;
  assign n22271 = n72654 & n22270 ;
  assign n22272 = n22266 | n22271 ;
  assign n22273 = n68993 & n22272 ;
  assign n22274 = n21471 & n22032 ;
  assign n21921 = n21480 | n21920 ;
  assign n72687 = ~n21921 ;
  assign n22275 = n21917 & n72687 ;
  assign n72688 = ~n21922 ;
  assign n22276 = n21920 & n72688 ;
  assign n22277 = n22275 | n22276 ;
  assign n22278 = n67021 & n22277 ;
  assign n22279 = n72654 & n22278 ;
  assign n22280 = n22274 | n22279 ;
  assign n22281 = n68716 & n22280 ;
  assign n22282 = n21479 & n22032 ;
  assign n21916 = n21488 | n21915 ;
  assign n72689 = ~n21916 ;
  assign n22283 = n72689 & n22101 ;
  assign n72690 = ~n22102 ;
  assign n22284 = n21915 & n72690 ;
  assign n22285 = n22283 | n22284 ;
  assign n22286 = n67021 & n22285 ;
  assign n22287 = n72654 & n22286 ;
  assign n22288 = n22282 | n22287 ;
  assign n22289 = n68545 & n22288 ;
  assign n22290 = n21487 & n22032 ;
  assign n21909 = n21496 | n21908 ;
  assign n72691 = ~n21909 ;
  assign n22291 = n21905 & n72691 ;
  assign n72692 = ~n21910 ;
  assign n22292 = n21908 & n72692 ;
  assign n22293 = n22291 | n22292 ;
  assign n22294 = n67021 & n22293 ;
  assign n22295 = n72654 & n22294 ;
  assign n22296 = n22290 | n22295 ;
  assign n22297 = n68438 & n22296 ;
  assign n22298 = n21495 & n22032 ;
  assign n21904 = n21504 | n21903 ;
  assign n72693 = ~n21904 ;
  assign n22299 = n72693 & n22097 ;
  assign n72694 = ~n22098 ;
  assign n22300 = n21903 & n72694 ;
  assign n22301 = n22299 | n22300 ;
  assign n22302 = n67021 & n22301 ;
  assign n22303 = n72654 & n22302 ;
  assign n22304 = n22298 | n22303 ;
  assign n22305 = n68214 & n22304 ;
  assign n22306 = n21503 & n22032 ;
  assign n21897 = n21512 | n21896 ;
  assign n72695 = ~n21897 ;
  assign n22307 = n21893 & n72695 ;
  assign n72696 = ~n21898 ;
  assign n22308 = n21896 & n72696 ;
  assign n22309 = n22307 | n22308 ;
  assign n22310 = n67021 & n22309 ;
  assign n22311 = n72654 & n22310 ;
  assign n22312 = n22306 | n22311 ;
  assign n22313 = n68058 & n22312 ;
  assign n22314 = n21511 & n22032 ;
  assign n21892 = n21520 | n21891 ;
  assign n72697 = ~n21892 ;
  assign n22315 = n72697 & n22093 ;
  assign n72698 = ~n22094 ;
  assign n22316 = n21891 & n72698 ;
  assign n22317 = n22315 | n22316 ;
  assign n22318 = n67021 & n22317 ;
  assign n22319 = n72654 & n22318 ;
  assign n22320 = n22314 | n22319 ;
  assign n22321 = n67986 & n22320 ;
  assign n22322 = n21519 & n22032 ;
  assign n21885 = n21528 | n21884 ;
  assign n72699 = ~n21885 ;
  assign n22323 = n21881 & n72699 ;
  assign n72700 = ~n21886 ;
  assign n22324 = n21884 & n72700 ;
  assign n22325 = n22323 | n22324 ;
  assign n22326 = n67021 & n22325 ;
  assign n22327 = n72654 & n22326 ;
  assign n22328 = n22322 | n22327 ;
  assign n22329 = n67763 & n22328 ;
  assign n22330 = n21527 & n22032 ;
  assign n21880 = n21536 | n21879 ;
  assign n72701 = ~n21880 ;
  assign n22331 = n72701 & n22089 ;
  assign n72702 = ~n22090 ;
  assign n22332 = n21879 & n72702 ;
  assign n22333 = n22331 | n22332 ;
  assign n22334 = n67021 & n22333 ;
  assign n22335 = n72654 & n22334 ;
  assign n22336 = n22330 | n22335 ;
  assign n22337 = n67622 & n22336 ;
  assign n22338 = n21535 & n22032 ;
  assign n21873 = n21544 | n21872 ;
  assign n72703 = ~n21873 ;
  assign n22339 = n21869 & n72703 ;
  assign n72704 = ~n21874 ;
  assign n22340 = n21872 & n72704 ;
  assign n22341 = n22339 | n22340 ;
  assign n22342 = n67021 & n22341 ;
  assign n22343 = n72654 & n22342 ;
  assign n22344 = n22338 | n22343 ;
  assign n22345 = n67531 & n22344 ;
  assign n22346 = n21543 & n22032 ;
  assign n21868 = n21552 | n21867 ;
  assign n72705 = ~n21868 ;
  assign n22347 = n72705 & n22085 ;
  assign n72706 = ~n22086 ;
  assign n22348 = n21867 & n72706 ;
  assign n22349 = n22347 | n22348 ;
  assign n22350 = n67021 & n22349 ;
  assign n22351 = n72654 & n22350 ;
  assign n22352 = n22346 | n22351 ;
  assign n22353 = n67348 & n22352 ;
  assign n22354 = n21551 & n22032 ;
  assign n21861 = n21560 | n21860 ;
  assign n72707 = ~n21861 ;
  assign n22355 = n21857 & n72707 ;
  assign n72708 = ~n21862 ;
  assign n22356 = n21860 & n72708 ;
  assign n22357 = n22355 | n22356 ;
  assign n22358 = n67021 & n22357 ;
  assign n22359 = n72654 & n22358 ;
  assign n22360 = n22354 | n22359 ;
  assign n22361 = n67222 & n22360 ;
  assign n22362 = n21559 & n22032 ;
  assign n21856 = n21568 | n21855 ;
  assign n72709 = ~n21856 ;
  assign n22363 = n72709 & n22081 ;
  assign n72710 = ~n22082 ;
  assign n22364 = n21855 & n72710 ;
  assign n22365 = n22363 | n22364 ;
  assign n22366 = n67021 & n22365 ;
  assign n22367 = n72654 & n22366 ;
  assign n22368 = n22362 | n22367 ;
  assign n22369 = n67164 & n22368 ;
  assign n22370 = n21567 & n22032 ;
  assign n21849 = n21576 | n21848 ;
  assign n72711 = ~n21849 ;
  assign n22371 = n21845 & n72711 ;
  assign n72712 = ~n21850 ;
  assign n22372 = n21848 & n72712 ;
  assign n22373 = n22371 | n22372 ;
  assign n22374 = n67021 & n22373 ;
  assign n22375 = n72654 & n22374 ;
  assign n22376 = n22370 | n22375 ;
  assign n22377 = n66979 & n22376 ;
  assign n22378 = n21575 & n22032 ;
  assign n21844 = n21584 | n21843 ;
  assign n72713 = ~n21844 ;
  assign n22379 = n72713 & n22077 ;
  assign n72714 = ~n22078 ;
  assign n22380 = n21843 & n72714 ;
  assign n22381 = n22379 | n22380 ;
  assign n22382 = n67021 & n22381 ;
  assign n22383 = n72654 & n22382 ;
  assign n22384 = n22378 | n22383 ;
  assign n22385 = n66868 & n22384 ;
  assign n22386 = n21583 & n22032 ;
  assign n21837 = n21592 | n21836 ;
  assign n72715 = ~n21837 ;
  assign n22387 = n21833 & n72715 ;
  assign n72716 = ~n21838 ;
  assign n22388 = n21836 & n72716 ;
  assign n22389 = n22387 | n22388 ;
  assign n22390 = n67021 & n22389 ;
  assign n22391 = n72654 & n22390 ;
  assign n22392 = n22386 | n22391 ;
  assign n22393 = n66797 & n22392 ;
  assign n22394 = n21591 & n22032 ;
  assign n21832 = n21600 | n21831 ;
  assign n72717 = ~n21832 ;
  assign n22395 = n72717 & n22073 ;
  assign n72718 = ~n22074 ;
  assign n22396 = n21831 & n72718 ;
  assign n22397 = n22395 | n22396 ;
  assign n22398 = n67021 & n22397 ;
  assign n22399 = n72654 & n22398 ;
  assign n22400 = n22394 | n22399 ;
  assign n22401 = n66654 & n22400 ;
  assign n22402 = n21599 & n22032 ;
  assign n21825 = n21608 | n21824 ;
  assign n72719 = ~n21825 ;
  assign n22403 = n21821 & n72719 ;
  assign n72720 = ~n21826 ;
  assign n22404 = n21824 & n72720 ;
  assign n22405 = n22403 | n22404 ;
  assign n22406 = n67021 & n22405 ;
  assign n22407 = n72654 & n22406 ;
  assign n22408 = n22402 | n22407 ;
  assign n22409 = n66560 & n22408 ;
  assign n22410 = n21607 & n22032 ;
  assign n21820 = n21616 | n21819 ;
  assign n72721 = ~n21820 ;
  assign n22411 = n72721 & n22069 ;
  assign n72722 = ~n22070 ;
  assign n22412 = n21819 & n72722 ;
  assign n22413 = n22411 | n22412 ;
  assign n22414 = n67021 & n22413 ;
  assign n22415 = n72654 & n22414 ;
  assign n22416 = n22410 | n22415 ;
  assign n22417 = n66505 & n22416 ;
  assign n22418 = n21615 & n22032 ;
  assign n21813 = n21624 | n21812 ;
  assign n72723 = ~n21813 ;
  assign n22419 = n21809 & n72723 ;
  assign n72724 = ~n21814 ;
  assign n22420 = n21812 & n72724 ;
  assign n22421 = n22419 | n22420 ;
  assign n22422 = n67021 & n22421 ;
  assign n22423 = n72654 & n22422 ;
  assign n22424 = n22418 | n22423 ;
  assign n22425 = n66379 & n22424 ;
  assign n22426 = n21623 & n22032 ;
  assign n21808 = n21632 | n21807 ;
  assign n72725 = ~n21808 ;
  assign n22427 = n72725 & n22065 ;
  assign n72726 = ~n22066 ;
  assign n22428 = n21807 & n72726 ;
  assign n22429 = n22427 | n22428 ;
  assign n22430 = n67021 & n22429 ;
  assign n22431 = n72654 & n22430 ;
  assign n22432 = n22426 | n22431 ;
  assign n22433 = n66299 & n22432 ;
  assign n22434 = n21631 & n22032 ;
  assign n21801 = n21640 | n21800 ;
  assign n72727 = ~n21801 ;
  assign n22435 = n21797 & n72727 ;
  assign n72728 = ~n21802 ;
  assign n22436 = n21800 & n72728 ;
  assign n22437 = n22435 | n22436 ;
  assign n22438 = n67021 & n22437 ;
  assign n22439 = n72654 & n22438 ;
  assign n22440 = n22434 | n22439 ;
  assign n22441 = n66244 & n22440 ;
  assign n22442 = n21639 & n22032 ;
  assign n21796 = n21648 | n21795 ;
  assign n72729 = ~n21796 ;
  assign n22443 = n72729 & n22061 ;
  assign n72730 = ~n22062 ;
  assign n22444 = n21795 & n72730 ;
  assign n22445 = n22443 | n22444 ;
  assign n22446 = n67021 & n22445 ;
  assign n22447 = n72654 & n22446 ;
  assign n22448 = n22442 | n22447 ;
  assign n22449 = n66145 & n22448 ;
  assign n22450 = n21647 & n22032 ;
  assign n21789 = n21656 | n21788 ;
  assign n72731 = ~n21789 ;
  assign n22451 = n21785 & n72731 ;
  assign n72732 = ~n21790 ;
  assign n22452 = n21788 & n72732 ;
  assign n22453 = n22451 | n22452 ;
  assign n22454 = n67021 & n22453 ;
  assign n22455 = n72654 & n22454 ;
  assign n22456 = n22450 | n22455 ;
  assign n22457 = n66081 & n22456 ;
  assign n22458 = n21655 & n22032 ;
  assign n21784 = n21664 | n21783 ;
  assign n72733 = ~n21784 ;
  assign n22459 = n72733 & n22057 ;
  assign n72734 = ~n22058 ;
  assign n22460 = n21783 & n72734 ;
  assign n22461 = n22459 | n22460 ;
  assign n22462 = n67021 & n22461 ;
  assign n22463 = n72654 & n22462 ;
  assign n22464 = n22458 | n22463 ;
  assign n22465 = n66043 & n22464 ;
  assign n22466 = n21663 & n22032 ;
  assign n21777 = n21672 | n21776 ;
  assign n72735 = ~n21777 ;
  assign n22467 = n21773 & n72735 ;
  assign n72736 = ~n21778 ;
  assign n22468 = n21776 & n72736 ;
  assign n22469 = n22467 | n22468 ;
  assign n22470 = n67021 & n22469 ;
  assign n22471 = n72654 & n22470 ;
  assign n22472 = n22466 | n22471 ;
  assign n22473 = n65960 & n22472 ;
  assign n22474 = n21671 & n22032 ;
  assign n21772 = n21680 | n21771 ;
  assign n72737 = ~n21772 ;
  assign n22475 = n72737 & n22053 ;
  assign n72738 = ~n22054 ;
  assign n22476 = n21771 & n72738 ;
  assign n22477 = n22475 | n22476 ;
  assign n22478 = n67021 & n22477 ;
  assign n22479 = n72654 & n22478 ;
  assign n22480 = n22474 | n22479 ;
  assign n22481 = n65909 & n22480 ;
  assign n22482 = n21679 & n22032 ;
  assign n21765 = n21688 | n21764 ;
  assign n72739 = ~n21765 ;
  assign n22483 = n21761 & n72739 ;
  assign n72740 = ~n21766 ;
  assign n22484 = n21764 & n72740 ;
  assign n22485 = n22483 | n22484 ;
  assign n22486 = n67021 & n22485 ;
  assign n22487 = n72654 & n22486 ;
  assign n22488 = n22482 | n22487 ;
  assign n22489 = n65877 & n22488 ;
  assign n22490 = n21687 & n22032 ;
  assign n21760 = n21696 | n21759 ;
  assign n72741 = ~n21760 ;
  assign n22491 = n72741 & n22049 ;
  assign n72742 = ~n22050 ;
  assign n22492 = n21759 & n72742 ;
  assign n22493 = n22491 | n22492 ;
  assign n22494 = n67021 & n22493 ;
  assign n22495 = n72654 & n22494 ;
  assign n22496 = n22490 | n22495 ;
  assign n22497 = n65820 & n22496 ;
  assign n22498 = n21695 & n22032 ;
  assign n22036 = n21704 | n21753 ;
  assign n72743 = ~n22036 ;
  assign n22499 = n21750 & n72743 ;
  assign n72744 = ~n21754 ;
  assign n22500 = n21753 & n72744 ;
  assign n22501 = n22499 | n22500 ;
  assign n22502 = n67021 & n22501 ;
  assign n22503 = n72654 & n22502 ;
  assign n22504 = n22498 | n22503 ;
  assign n22505 = n65791 & n22504 ;
  assign n22506 = n21703 & n22032 ;
  assign n22507 = n21713 | n21749 ;
  assign n72745 = ~n22507 ;
  assign n22508 = n22045 & n72745 ;
  assign n72746 = ~n22046 ;
  assign n22509 = n21749 & n72746 ;
  assign n22510 = n22508 | n22509 ;
  assign n22511 = n67021 & n22510 ;
  assign n22512 = n72654 & n22511 ;
  assign n22513 = n22506 | n22512 ;
  assign n22514 = n65772 & n22513 ;
  assign n22515 = n21712 & n22032 ;
  assign n22516 = n21721 | n21743 ;
  assign n72747 = ~n22516 ;
  assign n22517 = n22043 & n72747 ;
  assign n72748 = ~n21744 ;
  assign n22518 = n21743 & n72748 ;
  assign n22519 = n22517 | n22518 ;
  assign n22520 = n67021 & n22519 ;
  assign n22521 = n72654 & n22520 ;
  assign n22522 = n22515 | n22521 ;
  assign n22523 = n65746 & n22522 ;
  assign n22524 = n21720 & n22032 ;
  assign n22041 = n21735 | n21739 ;
  assign n72749 = ~n22041 ;
  assign n22525 = n21733 & n72749 ;
  assign n72750 = ~n22042 ;
  assign n22526 = n21739 & n72750 ;
  assign n22527 = n22525 | n22526 ;
  assign n22528 = n67021 & n22527 ;
  assign n22529 = n72654 & n22528 ;
  assign n22530 = n22524 | n22529 ;
  assign n22531 = n65721 & n22530 ;
  assign n22034 = n21734 & n22032 ;
  assign n22039 = n21730 & n21731 ;
  assign n22532 = n72545 & n22039 ;
  assign n22533 = n65429 | n22532 ;
  assign n72751 = ~n22533 ;
  assign n22534 = n21733 & n72751 ;
  assign n22535 = n72654 & n22534 ;
  assign n22536 = n22034 | n22535 ;
  assign n22537 = n65686 & n22536 ;
  assign n72752 = ~x116 ;
  assign n22538 = x64 & n72752 ;
  assign n72753 = ~n268 ;
  assign n22539 = n72753 & n22538 ;
  assign n22540 = n65709 & n22539 ;
  assign n22544 = n72645 & n22543 ;
  assign n22545 = n22028 | n22544 ;
  assign n22546 = n72646 & n22545 ;
  assign n72754 = ~n22546 ;
  assign n22547 = n22540 & n72754 ;
  assign n72755 = ~n22547 ;
  assign n22548 = x12 & n72755 ;
  assign n22549 = n72027 & n21731 ;
  assign n22550 = n65681 & n22549 ;
  assign n22551 = n72654 & n22550 ;
  assign n22552 = n22548 | n22551 ;
  assign n22554 = x65 & n22552 ;
  assign n22541 = n72654 & n22540 ;
  assign n72756 = ~n22541 ;
  assign n22542 = x12 & n72756 ;
  assign n22553 = x65 | n22551 ;
  assign n22555 = n22542 | n22553 ;
  assign n72757 = ~n22554 ;
  assign n22556 = n72757 & n22555 ;
  assign n72758 = ~x11 ;
  assign n22557 = n72758 & x64 ;
  assign n22558 = n22556 | n22557 ;
  assign n22559 = n65670 & n22552 ;
  assign n72759 = ~n22559 ;
  assign n22560 = n22558 & n72759 ;
  assign n72760 = ~n22535 ;
  assign n22561 = x66 & n72760 ;
  assign n72761 = ~n22034 ;
  assign n22562 = n72761 & n22561 ;
  assign n22563 = n22537 | n22562 ;
  assign n22564 = n22560 | n22563 ;
  assign n72762 = ~n22537 ;
  assign n22565 = n72762 & n22564 ;
  assign n72763 = ~n22529 ;
  assign n22566 = x67 & n72763 ;
  assign n72764 = ~n22524 ;
  assign n22567 = n72764 & n22566 ;
  assign n22568 = n22565 | n22567 ;
  assign n72765 = ~n22531 ;
  assign n22569 = n72765 & n22568 ;
  assign n72766 = ~n22521 ;
  assign n22570 = x68 & n72766 ;
  assign n72767 = ~n22515 ;
  assign n22571 = n72767 & n22570 ;
  assign n22572 = n22523 | n22571 ;
  assign n22573 = n22569 | n22572 ;
  assign n72768 = ~n22523 ;
  assign n22574 = n72768 & n22573 ;
  assign n72769 = ~n22512 ;
  assign n22575 = x69 & n72769 ;
  assign n72770 = ~n22506 ;
  assign n22576 = n72770 & n22575 ;
  assign n22577 = n22514 | n22576 ;
  assign n22578 = n22574 | n22577 ;
  assign n72771 = ~n22514 ;
  assign n22579 = n72771 & n22578 ;
  assign n72772 = ~n22503 ;
  assign n22580 = x70 & n72772 ;
  assign n72773 = ~n22498 ;
  assign n22581 = n72773 & n22580 ;
  assign n22582 = n22505 | n22581 ;
  assign n22583 = n22579 | n22582 ;
  assign n72774 = ~n22505 ;
  assign n22584 = n72774 & n22583 ;
  assign n72775 = ~n22495 ;
  assign n22585 = x71 & n72775 ;
  assign n72776 = ~n22490 ;
  assign n22586 = n72776 & n22585 ;
  assign n22587 = n22497 | n22586 ;
  assign n22589 = n22584 | n22587 ;
  assign n72777 = ~n22497 ;
  assign n22590 = n72777 & n22589 ;
  assign n72778 = ~n22487 ;
  assign n22591 = x72 & n72778 ;
  assign n72779 = ~n22482 ;
  assign n22592 = n72779 & n22591 ;
  assign n22593 = n22489 | n22592 ;
  assign n22594 = n22590 | n22593 ;
  assign n72780 = ~n22489 ;
  assign n22595 = n72780 & n22594 ;
  assign n72781 = ~n22479 ;
  assign n22596 = x73 & n72781 ;
  assign n72782 = ~n22474 ;
  assign n22597 = n72782 & n22596 ;
  assign n22598 = n22481 | n22597 ;
  assign n22600 = n22595 | n22598 ;
  assign n72783 = ~n22481 ;
  assign n22601 = n72783 & n22600 ;
  assign n72784 = ~n22471 ;
  assign n22602 = x74 & n72784 ;
  assign n72785 = ~n22466 ;
  assign n22603 = n72785 & n22602 ;
  assign n22604 = n22473 | n22603 ;
  assign n22605 = n22601 | n22604 ;
  assign n72786 = ~n22473 ;
  assign n22606 = n72786 & n22605 ;
  assign n72787 = ~n22463 ;
  assign n22607 = x75 & n72787 ;
  assign n72788 = ~n22458 ;
  assign n22608 = n72788 & n22607 ;
  assign n22609 = n22465 | n22608 ;
  assign n22611 = n22606 | n22609 ;
  assign n72789 = ~n22465 ;
  assign n22612 = n72789 & n22611 ;
  assign n72790 = ~n22455 ;
  assign n22613 = x76 & n72790 ;
  assign n72791 = ~n22450 ;
  assign n22614 = n72791 & n22613 ;
  assign n22615 = n22457 | n22614 ;
  assign n22616 = n22612 | n22615 ;
  assign n72792 = ~n22457 ;
  assign n22617 = n72792 & n22616 ;
  assign n72793 = ~n22447 ;
  assign n22618 = x77 & n72793 ;
  assign n72794 = ~n22442 ;
  assign n22619 = n72794 & n22618 ;
  assign n22620 = n22449 | n22619 ;
  assign n22622 = n22617 | n22620 ;
  assign n72795 = ~n22449 ;
  assign n22623 = n72795 & n22622 ;
  assign n72796 = ~n22439 ;
  assign n22624 = x78 & n72796 ;
  assign n72797 = ~n22434 ;
  assign n22625 = n72797 & n22624 ;
  assign n22626 = n22441 | n22625 ;
  assign n22627 = n22623 | n22626 ;
  assign n72798 = ~n22441 ;
  assign n22628 = n72798 & n22627 ;
  assign n72799 = ~n22431 ;
  assign n22629 = x79 & n72799 ;
  assign n72800 = ~n22426 ;
  assign n22630 = n72800 & n22629 ;
  assign n22631 = n22433 | n22630 ;
  assign n22633 = n22628 | n22631 ;
  assign n72801 = ~n22433 ;
  assign n22634 = n72801 & n22633 ;
  assign n72802 = ~n22423 ;
  assign n22635 = x80 & n72802 ;
  assign n72803 = ~n22418 ;
  assign n22636 = n72803 & n22635 ;
  assign n22637 = n22425 | n22636 ;
  assign n22638 = n22634 | n22637 ;
  assign n72804 = ~n22425 ;
  assign n22639 = n72804 & n22638 ;
  assign n72805 = ~n22415 ;
  assign n22640 = x81 & n72805 ;
  assign n72806 = ~n22410 ;
  assign n22641 = n72806 & n22640 ;
  assign n22642 = n22417 | n22641 ;
  assign n22644 = n22639 | n22642 ;
  assign n72807 = ~n22417 ;
  assign n22645 = n72807 & n22644 ;
  assign n72808 = ~n22407 ;
  assign n22646 = x82 & n72808 ;
  assign n72809 = ~n22402 ;
  assign n22647 = n72809 & n22646 ;
  assign n22648 = n22409 | n22647 ;
  assign n22649 = n22645 | n22648 ;
  assign n72810 = ~n22409 ;
  assign n22650 = n72810 & n22649 ;
  assign n72811 = ~n22399 ;
  assign n22651 = x83 & n72811 ;
  assign n72812 = ~n22394 ;
  assign n22652 = n72812 & n22651 ;
  assign n22653 = n22401 | n22652 ;
  assign n22655 = n22650 | n22653 ;
  assign n72813 = ~n22401 ;
  assign n22656 = n72813 & n22655 ;
  assign n72814 = ~n22391 ;
  assign n22657 = x84 & n72814 ;
  assign n72815 = ~n22386 ;
  assign n22658 = n72815 & n22657 ;
  assign n22659 = n22393 | n22658 ;
  assign n22660 = n22656 | n22659 ;
  assign n72816 = ~n22393 ;
  assign n22661 = n72816 & n22660 ;
  assign n72817 = ~n22383 ;
  assign n22662 = x85 & n72817 ;
  assign n72818 = ~n22378 ;
  assign n22663 = n72818 & n22662 ;
  assign n22664 = n22385 | n22663 ;
  assign n22666 = n22661 | n22664 ;
  assign n72819 = ~n22385 ;
  assign n22667 = n72819 & n22666 ;
  assign n72820 = ~n22375 ;
  assign n22668 = x86 & n72820 ;
  assign n72821 = ~n22370 ;
  assign n22669 = n72821 & n22668 ;
  assign n22670 = n22377 | n22669 ;
  assign n22671 = n22667 | n22670 ;
  assign n72822 = ~n22377 ;
  assign n22672 = n72822 & n22671 ;
  assign n72823 = ~n22367 ;
  assign n22673 = x87 & n72823 ;
  assign n72824 = ~n22362 ;
  assign n22674 = n72824 & n22673 ;
  assign n22675 = n22369 | n22674 ;
  assign n22677 = n22672 | n22675 ;
  assign n72825 = ~n22369 ;
  assign n22678 = n72825 & n22677 ;
  assign n72826 = ~n22359 ;
  assign n22679 = x88 & n72826 ;
  assign n72827 = ~n22354 ;
  assign n22680 = n72827 & n22679 ;
  assign n22681 = n22361 | n22680 ;
  assign n22682 = n22678 | n22681 ;
  assign n72828 = ~n22361 ;
  assign n22683 = n72828 & n22682 ;
  assign n72829 = ~n22351 ;
  assign n22684 = x89 & n72829 ;
  assign n72830 = ~n22346 ;
  assign n22685 = n72830 & n22684 ;
  assign n22686 = n22353 | n22685 ;
  assign n22688 = n22683 | n22686 ;
  assign n72831 = ~n22353 ;
  assign n22689 = n72831 & n22688 ;
  assign n72832 = ~n22343 ;
  assign n22690 = x90 & n72832 ;
  assign n72833 = ~n22338 ;
  assign n22691 = n72833 & n22690 ;
  assign n22692 = n22345 | n22691 ;
  assign n22693 = n22689 | n22692 ;
  assign n72834 = ~n22345 ;
  assign n22694 = n72834 & n22693 ;
  assign n72835 = ~n22335 ;
  assign n22695 = x91 & n72835 ;
  assign n72836 = ~n22330 ;
  assign n22696 = n72836 & n22695 ;
  assign n22697 = n22337 | n22696 ;
  assign n22699 = n22694 | n22697 ;
  assign n72837 = ~n22337 ;
  assign n22700 = n72837 & n22699 ;
  assign n72838 = ~n22327 ;
  assign n22701 = x92 & n72838 ;
  assign n72839 = ~n22322 ;
  assign n22702 = n72839 & n22701 ;
  assign n22703 = n22329 | n22702 ;
  assign n22704 = n22700 | n22703 ;
  assign n72840 = ~n22329 ;
  assign n22705 = n72840 & n22704 ;
  assign n72841 = ~n22319 ;
  assign n22706 = x93 & n72841 ;
  assign n72842 = ~n22314 ;
  assign n22707 = n72842 & n22706 ;
  assign n22708 = n22321 | n22707 ;
  assign n22710 = n22705 | n22708 ;
  assign n72843 = ~n22321 ;
  assign n22711 = n72843 & n22710 ;
  assign n72844 = ~n22311 ;
  assign n22712 = x94 & n72844 ;
  assign n72845 = ~n22306 ;
  assign n22713 = n72845 & n22712 ;
  assign n22714 = n22313 | n22713 ;
  assign n22715 = n22711 | n22714 ;
  assign n72846 = ~n22313 ;
  assign n22716 = n72846 & n22715 ;
  assign n72847 = ~n22303 ;
  assign n22717 = x95 & n72847 ;
  assign n72848 = ~n22298 ;
  assign n22718 = n72848 & n22717 ;
  assign n22719 = n22305 | n22718 ;
  assign n22721 = n22716 | n22719 ;
  assign n72849 = ~n22305 ;
  assign n22722 = n72849 & n22721 ;
  assign n72850 = ~n22295 ;
  assign n22723 = x96 & n72850 ;
  assign n72851 = ~n22290 ;
  assign n22724 = n72851 & n22723 ;
  assign n22725 = n22297 | n22724 ;
  assign n22726 = n22722 | n22725 ;
  assign n72852 = ~n22297 ;
  assign n22727 = n72852 & n22726 ;
  assign n72853 = ~n22287 ;
  assign n22728 = x97 & n72853 ;
  assign n72854 = ~n22282 ;
  assign n22729 = n72854 & n22728 ;
  assign n22730 = n22289 | n22729 ;
  assign n22732 = n22727 | n22730 ;
  assign n72855 = ~n22289 ;
  assign n22733 = n72855 & n22732 ;
  assign n72856 = ~n22279 ;
  assign n22734 = x98 & n72856 ;
  assign n72857 = ~n22274 ;
  assign n22735 = n72857 & n22734 ;
  assign n22736 = n22281 | n22735 ;
  assign n22737 = n22733 | n22736 ;
  assign n72858 = ~n22281 ;
  assign n22738 = n72858 & n22737 ;
  assign n72859 = ~n22271 ;
  assign n22739 = x99 & n72859 ;
  assign n72860 = ~n22266 ;
  assign n22740 = n72860 & n22739 ;
  assign n22741 = n22273 | n22740 ;
  assign n22743 = n22738 | n22741 ;
  assign n72861 = ~n22273 ;
  assign n22744 = n72861 & n22743 ;
  assign n72862 = ~n22263 ;
  assign n22745 = x100 & n72862 ;
  assign n72863 = ~n22258 ;
  assign n22746 = n72863 & n22745 ;
  assign n22747 = n22265 | n22746 ;
  assign n22748 = n22744 | n22747 ;
  assign n72864 = ~n22265 ;
  assign n22749 = n72864 & n22748 ;
  assign n72865 = ~n22255 ;
  assign n22750 = x101 & n72865 ;
  assign n72866 = ~n22250 ;
  assign n22751 = n72866 & n22750 ;
  assign n22752 = n22257 | n22751 ;
  assign n22754 = n22749 | n22752 ;
  assign n72867 = ~n22257 ;
  assign n22755 = n72867 & n22754 ;
  assign n72868 = ~n22247 ;
  assign n22756 = x102 & n72868 ;
  assign n72869 = ~n22242 ;
  assign n22757 = n72869 & n22756 ;
  assign n22758 = n22249 | n22757 ;
  assign n22759 = n22755 | n22758 ;
  assign n72870 = ~n22249 ;
  assign n22760 = n72870 & n22759 ;
  assign n72871 = ~n22239 ;
  assign n22761 = x103 & n72871 ;
  assign n72872 = ~n22234 ;
  assign n22762 = n72872 & n22761 ;
  assign n22763 = n22241 | n22762 ;
  assign n22765 = n22760 | n22763 ;
  assign n72873 = ~n22241 ;
  assign n22766 = n72873 & n22765 ;
  assign n72874 = ~n22231 ;
  assign n22767 = x104 & n72874 ;
  assign n72875 = ~n22226 ;
  assign n22768 = n72875 & n22767 ;
  assign n22769 = n22233 | n22768 ;
  assign n22770 = n22766 | n22769 ;
  assign n72876 = ~n22233 ;
  assign n22771 = n72876 & n22770 ;
  assign n72877 = ~n22223 ;
  assign n22772 = x105 & n72877 ;
  assign n72878 = ~n22218 ;
  assign n22773 = n72878 & n22772 ;
  assign n22774 = n22225 | n22773 ;
  assign n22776 = n22771 | n22774 ;
  assign n72879 = ~n22225 ;
  assign n22777 = n72879 & n22776 ;
  assign n72880 = ~n22215 ;
  assign n22778 = x106 & n72880 ;
  assign n72881 = ~n22210 ;
  assign n22779 = n72881 & n22778 ;
  assign n22780 = n22217 | n22779 ;
  assign n22781 = n22777 | n22780 ;
  assign n72882 = ~n22217 ;
  assign n22782 = n72882 & n22781 ;
  assign n72883 = ~n22207 ;
  assign n22783 = x107 & n72883 ;
  assign n72884 = ~n22202 ;
  assign n22784 = n72884 & n22783 ;
  assign n22785 = n22209 | n22784 ;
  assign n22787 = n22782 | n22785 ;
  assign n72885 = ~n22209 ;
  assign n22788 = n72885 & n22787 ;
  assign n72886 = ~n22199 ;
  assign n22789 = x108 & n72886 ;
  assign n72887 = ~n22194 ;
  assign n22790 = n72887 & n22789 ;
  assign n22791 = n22201 | n22790 ;
  assign n22792 = n22788 | n22791 ;
  assign n72888 = ~n22201 ;
  assign n22793 = n72888 & n22792 ;
  assign n72889 = ~n22191 ;
  assign n22794 = x109 & n72889 ;
  assign n72890 = ~n22186 ;
  assign n22795 = n72890 & n22794 ;
  assign n22796 = n22193 | n22795 ;
  assign n22798 = n22793 | n22796 ;
  assign n72891 = ~n22193 ;
  assign n22799 = n72891 & n22798 ;
  assign n72892 = ~n22183 ;
  assign n22800 = x110 & n72892 ;
  assign n72893 = ~n22178 ;
  assign n22801 = n72893 & n22800 ;
  assign n22802 = n22185 | n22801 ;
  assign n22803 = n22799 | n22802 ;
  assign n72894 = ~n22185 ;
  assign n22804 = n72894 & n22803 ;
  assign n72895 = ~n22175 ;
  assign n22805 = x111 & n72895 ;
  assign n72896 = ~n22170 ;
  assign n22806 = n72896 & n22805 ;
  assign n22807 = n22177 | n22806 ;
  assign n22809 = n22804 | n22807 ;
  assign n72897 = ~n22177 ;
  assign n22810 = n72897 & n22809 ;
  assign n72898 = ~n22167 ;
  assign n22811 = x112 & n72898 ;
  assign n72899 = ~n22162 ;
  assign n22812 = n72899 & n22811 ;
  assign n22813 = n22169 | n22812 ;
  assign n22814 = n22810 | n22813 ;
  assign n72900 = ~n22169 ;
  assign n22815 = n72900 & n22814 ;
  assign n72901 = ~n22159 ;
  assign n22816 = x113 & n72901 ;
  assign n72902 = ~n22154 ;
  assign n22817 = n72902 & n22816 ;
  assign n22818 = n22161 | n22817 ;
  assign n22820 = n22815 | n22818 ;
  assign n72903 = ~n22161 ;
  assign n22821 = n72903 & n22820 ;
  assign n72904 = ~n22151 ;
  assign n22822 = x114 & n72904 ;
  assign n72905 = ~n22146 ;
  assign n22823 = n72905 & n22822 ;
  assign n22824 = n22153 | n22823 ;
  assign n22825 = n22821 | n22824 ;
  assign n72906 = ~n22153 ;
  assign n22826 = n72906 & n22825 ;
  assign n72907 = ~n22143 ;
  assign n22827 = x115 & n72907 ;
  assign n72908 = ~n22035 ;
  assign n22828 = n72908 & n22827 ;
  assign n22829 = n22145 | n22828 ;
  assign n22831 = n22826 | n22829 ;
  assign n72909 = ~n22145 ;
  assign n22832 = n72909 & n22831 ;
  assign n22839 = n72752 & n22838 ;
  assign n141 = ~n22032 ;
  assign n22840 = n141 & n22836 ;
  assign n22841 = n21327 & n22032 ;
  assign n72911 = ~n22841 ;
  assign n22842 = x116 & n72911 ;
  assign n72912 = ~n22840 ;
  assign n22843 = n72912 & n22842 ;
  assign n22844 = n465 | n22843 ;
  assign n22845 = n22839 | n22844 ;
  assign n22847 = n22832 | n22845 ;
  assign n72913 = ~n22846 ;
  assign n22848 = n72913 & n22847 ;
  assign n72914 = ~n22826 ;
  assign n22830 = n72914 & n22829 ;
  assign n22851 = n22542 | n22551 ;
  assign n22852 = x65 & n22851 ;
  assign n72915 = ~n22852 ;
  assign n22853 = n22555 & n72915 ;
  assign n22854 = n22557 | n22853 ;
  assign n22855 = n72759 & n22854 ;
  assign n22857 = n22562 | n22855 ;
  assign n22858 = n72762 & n22857 ;
  assign n22859 = n22531 | n22567 ;
  assign n22861 = n22858 | n22859 ;
  assign n22862 = n72765 & n22861 ;
  assign n22864 = n22572 | n22862 ;
  assign n22865 = n72768 & n22864 ;
  assign n22867 = n22577 | n22865 ;
  assign n22868 = n72771 & n22867 ;
  assign n22869 = n22582 | n22868 ;
  assign n22871 = n72774 & n22869 ;
  assign n22872 = n22587 | n22871 ;
  assign n22873 = n72777 & n22872 ;
  assign n22874 = n22593 | n22873 ;
  assign n22876 = n72780 & n22874 ;
  assign n22877 = n22598 | n22876 ;
  assign n22878 = n72783 & n22877 ;
  assign n22879 = n22604 | n22878 ;
  assign n22881 = n72786 & n22879 ;
  assign n22882 = n22609 | n22881 ;
  assign n22883 = n72789 & n22882 ;
  assign n22884 = n22615 | n22883 ;
  assign n22886 = n72792 & n22884 ;
  assign n22887 = n22620 | n22886 ;
  assign n22888 = n72795 & n22887 ;
  assign n22889 = n22626 | n22888 ;
  assign n22891 = n72798 & n22889 ;
  assign n22892 = n22631 | n22891 ;
  assign n22893 = n72801 & n22892 ;
  assign n22894 = n22637 | n22893 ;
  assign n22896 = n72804 & n22894 ;
  assign n22897 = n22642 | n22896 ;
  assign n22898 = n72807 & n22897 ;
  assign n22899 = n22648 | n22898 ;
  assign n22901 = n72810 & n22899 ;
  assign n22902 = n22653 | n22901 ;
  assign n22903 = n72813 & n22902 ;
  assign n22904 = n22659 | n22903 ;
  assign n22906 = n72816 & n22904 ;
  assign n22907 = n22664 | n22906 ;
  assign n22908 = n72819 & n22907 ;
  assign n22909 = n22670 | n22908 ;
  assign n22911 = n72822 & n22909 ;
  assign n22912 = n22675 | n22911 ;
  assign n22913 = n72825 & n22912 ;
  assign n22914 = n22681 | n22913 ;
  assign n22916 = n72828 & n22914 ;
  assign n22917 = n22686 | n22916 ;
  assign n22918 = n72831 & n22917 ;
  assign n22919 = n22692 | n22918 ;
  assign n22921 = n72834 & n22919 ;
  assign n22922 = n22697 | n22921 ;
  assign n22923 = n72837 & n22922 ;
  assign n22924 = n22703 | n22923 ;
  assign n22926 = n72840 & n22924 ;
  assign n22927 = n22708 | n22926 ;
  assign n22928 = n72843 & n22927 ;
  assign n22929 = n22714 | n22928 ;
  assign n22931 = n72846 & n22929 ;
  assign n22932 = n22719 | n22931 ;
  assign n22933 = n72849 & n22932 ;
  assign n22934 = n22725 | n22933 ;
  assign n22936 = n72852 & n22934 ;
  assign n22937 = n22730 | n22936 ;
  assign n22938 = n72855 & n22937 ;
  assign n22939 = n22736 | n22938 ;
  assign n22941 = n72858 & n22939 ;
  assign n22942 = n22741 | n22941 ;
  assign n22943 = n72861 & n22942 ;
  assign n22944 = n22747 | n22943 ;
  assign n22946 = n72864 & n22944 ;
  assign n22947 = n22752 | n22946 ;
  assign n22948 = n72867 & n22947 ;
  assign n22949 = n22758 | n22948 ;
  assign n22951 = n72870 & n22949 ;
  assign n22952 = n22763 | n22951 ;
  assign n22953 = n72873 & n22952 ;
  assign n22954 = n22769 | n22953 ;
  assign n22956 = n72876 & n22954 ;
  assign n22957 = n22774 | n22956 ;
  assign n22958 = n72879 & n22957 ;
  assign n22959 = n22780 | n22958 ;
  assign n22961 = n72882 & n22959 ;
  assign n22962 = n22785 | n22961 ;
  assign n22963 = n72885 & n22962 ;
  assign n22964 = n22791 | n22963 ;
  assign n22966 = n72888 & n22964 ;
  assign n22967 = n22796 | n22966 ;
  assign n22968 = n72891 & n22967 ;
  assign n22969 = n22802 | n22968 ;
  assign n22971 = n72894 & n22969 ;
  assign n22972 = n22807 | n22971 ;
  assign n22973 = n72897 & n22972 ;
  assign n22974 = n22813 | n22973 ;
  assign n22976 = n72900 & n22974 ;
  assign n22977 = n22818 | n22976 ;
  assign n22978 = n72903 & n22977 ;
  assign n22980 = n22824 | n22978 ;
  assign n22981 = n22153 | n22829 ;
  assign n72916 = ~n22981 ;
  assign n22982 = n22980 & n72916 ;
  assign n22983 = n22830 | n22982 ;
  assign n140 = ~n22848 ;
  assign n22984 = n140 & n22983 ;
  assign n22985 = n72906 & n22980 ;
  assign n22986 = n22829 | n22985 ;
  assign n22987 = n72909 & n22986 ;
  assign n22988 = n22845 | n22987 ;
  assign n22989 = n22144 & n72913 ;
  assign n22990 = n22988 & n22989 ;
  assign n22991 = n22984 | n22990 ;
  assign n22992 = n72752 & n22991 ;
  assign n72918 = ~n22990 ;
  assign n23664 = x116 & n72918 ;
  assign n72919 = ~n22984 ;
  assign n23665 = n72919 & n23664 ;
  assign n23666 = n22992 | n23665 ;
  assign n72920 = ~n22978 ;
  assign n22979 = n22824 & n72920 ;
  assign n22993 = n22161 | n22824 ;
  assign n72921 = ~n22993 ;
  assign n22994 = n22820 & n72921 ;
  assign n22995 = n22979 | n22994 ;
  assign n22996 = n140 & n22995 ;
  assign n22997 = n22152 & n72913 ;
  assign n22998 = n22988 & n22997 ;
  assign n22999 = n22996 | n22998 ;
  assign n23000 = n72393 & n22999 ;
  assign n72922 = ~n22815 ;
  assign n22819 = n72922 & n22818 ;
  assign n23001 = n22169 | n22818 ;
  assign n72923 = ~n23001 ;
  assign n23002 = n22974 & n72923 ;
  assign n23003 = n22819 | n23002 ;
  assign n23004 = n140 & n23003 ;
  assign n23005 = n22160 & n72913 ;
  assign n23006 = n22988 & n23005 ;
  assign n23007 = n23004 | n23006 ;
  assign n23008 = n72385 & n23007 ;
  assign n72924 = ~n23006 ;
  assign n23654 = x114 & n72924 ;
  assign n72925 = ~n23004 ;
  assign n23655 = n72925 & n23654 ;
  assign n23656 = n23008 | n23655 ;
  assign n72926 = ~n22973 ;
  assign n22975 = n22813 & n72926 ;
  assign n23009 = n22177 | n22813 ;
  assign n72927 = ~n23009 ;
  assign n23010 = n22809 & n72927 ;
  assign n23011 = n22975 | n23010 ;
  assign n23012 = n140 & n23011 ;
  assign n23013 = n22168 & n72913 ;
  assign n23014 = n22988 & n23013 ;
  assign n23015 = n23012 | n23014 ;
  assign n23016 = n72025 & n23015 ;
  assign n72928 = ~n22804 ;
  assign n22808 = n72928 & n22807 ;
  assign n23017 = n22185 | n22807 ;
  assign n72929 = ~n23017 ;
  assign n23018 = n22969 & n72929 ;
  assign n23019 = n22808 | n23018 ;
  assign n23020 = n140 & n23019 ;
  assign n23021 = n22176 & n72913 ;
  assign n23022 = n22988 & n23021 ;
  assign n23023 = n23020 | n23022 ;
  assign n23024 = n71645 & n23023 ;
  assign n72930 = ~n23022 ;
  assign n23643 = x112 & n72930 ;
  assign n72931 = ~n23020 ;
  assign n23644 = n72931 & n23643 ;
  assign n23645 = n23024 | n23644 ;
  assign n72932 = ~n22968 ;
  assign n22970 = n22802 & n72932 ;
  assign n23025 = n22193 | n22802 ;
  assign n72933 = ~n23025 ;
  assign n23026 = n22798 & n72933 ;
  assign n23027 = n22970 | n23026 ;
  assign n23028 = n140 & n23027 ;
  assign n23029 = n22184 & n72913 ;
  assign n23030 = n22988 & n23029 ;
  assign n23031 = n23028 | n23030 ;
  assign n23032 = n71633 & n23031 ;
  assign n72934 = ~n22793 ;
  assign n22797 = n72934 & n22796 ;
  assign n23033 = n22201 | n22796 ;
  assign n72935 = ~n23033 ;
  assign n23034 = n22964 & n72935 ;
  assign n23035 = n22797 | n23034 ;
  assign n23036 = n140 & n23035 ;
  assign n23037 = n22192 & n72913 ;
  assign n23038 = n22988 & n23037 ;
  assign n23039 = n23036 | n23038 ;
  assign n23040 = n71253 & n23039 ;
  assign n72936 = ~n23038 ;
  assign n23633 = x110 & n72936 ;
  assign n72937 = ~n23036 ;
  assign n23634 = n72937 & n23633 ;
  assign n23635 = n23040 | n23634 ;
  assign n72938 = ~n22963 ;
  assign n22965 = n22791 & n72938 ;
  assign n23041 = n22209 | n22791 ;
  assign n72939 = ~n23041 ;
  assign n23042 = n22787 & n72939 ;
  assign n23043 = n22965 | n23042 ;
  assign n23044 = n140 & n23043 ;
  assign n23045 = n22200 & n72913 ;
  assign n23046 = n22988 & n23045 ;
  assign n23047 = n23044 | n23046 ;
  assign n23048 = n70935 & n23047 ;
  assign n72940 = ~n22782 ;
  assign n22786 = n72940 & n22785 ;
  assign n23049 = n22217 | n22785 ;
  assign n72941 = ~n23049 ;
  assign n23050 = n22959 & n72941 ;
  assign n23051 = n22786 | n23050 ;
  assign n23052 = n140 & n23051 ;
  assign n23053 = n22208 & n72913 ;
  assign n23054 = n22988 & n23053 ;
  assign n23055 = n23052 | n23054 ;
  assign n23056 = n70927 & n23055 ;
  assign n72942 = ~n23054 ;
  assign n23622 = x108 & n72942 ;
  assign n72943 = ~n23052 ;
  assign n23623 = n72943 & n23622 ;
  assign n23624 = n23056 | n23623 ;
  assign n72944 = ~n22958 ;
  assign n22960 = n22780 & n72944 ;
  assign n23057 = n22225 | n22780 ;
  assign n72945 = ~n23057 ;
  assign n23058 = n22776 & n72945 ;
  assign n23059 = n22960 | n23058 ;
  assign n23060 = n140 & n23059 ;
  assign n23061 = n22216 & n72913 ;
  assign n23062 = n22988 & n23061 ;
  assign n23063 = n23060 | n23062 ;
  assign n23064 = n70609 & n23063 ;
  assign n72946 = ~n22771 ;
  assign n22775 = n72946 & n22774 ;
  assign n23065 = n22233 | n22774 ;
  assign n72947 = ~n23065 ;
  assign n23066 = n22954 & n72947 ;
  assign n23067 = n22775 | n23066 ;
  assign n23068 = n140 & n23067 ;
  assign n23069 = n22224 & n72913 ;
  assign n23070 = n22988 & n23069 ;
  assign n23071 = n23068 | n23070 ;
  assign n23072 = n70276 & n23071 ;
  assign n72948 = ~n23070 ;
  assign n23612 = x106 & n72948 ;
  assign n72949 = ~n23068 ;
  assign n23613 = n72949 & n23612 ;
  assign n23614 = n23072 | n23613 ;
  assign n72950 = ~n22953 ;
  assign n22955 = n22769 & n72950 ;
  assign n23073 = n22241 | n22769 ;
  assign n72951 = ~n23073 ;
  assign n23074 = n22765 & n72951 ;
  assign n23075 = n22955 | n23074 ;
  assign n23076 = n140 & n23075 ;
  assign n23077 = n22232 & n72913 ;
  assign n23078 = n22988 & n23077 ;
  assign n23079 = n23076 | n23078 ;
  assign n23080 = n70176 & n23079 ;
  assign n72952 = ~n22760 ;
  assign n22764 = n72952 & n22763 ;
  assign n23081 = n22249 | n22763 ;
  assign n72953 = ~n23081 ;
  assign n23082 = n22949 & n72953 ;
  assign n23083 = n22764 | n23082 ;
  assign n23084 = n140 & n23083 ;
  assign n23085 = n22240 & n72913 ;
  assign n23086 = n22988 & n23085 ;
  assign n23087 = n23084 | n23086 ;
  assign n23088 = n69857 & n23087 ;
  assign n72954 = ~n23086 ;
  assign n23601 = x104 & n72954 ;
  assign n72955 = ~n23084 ;
  assign n23602 = n72955 & n23601 ;
  assign n23603 = n23088 | n23602 ;
  assign n72956 = ~n22948 ;
  assign n22950 = n22758 & n72956 ;
  assign n23089 = n22257 | n22758 ;
  assign n72957 = ~n23089 ;
  assign n23090 = n22754 & n72957 ;
  assign n23091 = n22950 | n23090 ;
  assign n23092 = n140 & n23091 ;
  assign n23093 = n22248 & n72913 ;
  assign n23094 = n22988 & n23093 ;
  assign n23095 = n23092 | n23094 ;
  assign n23096 = n69656 & n23095 ;
  assign n72958 = ~n22749 ;
  assign n22753 = n72958 & n22752 ;
  assign n23097 = n22265 | n22752 ;
  assign n72959 = ~n23097 ;
  assign n23098 = n22944 & n72959 ;
  assign n23099 = n22753 | n23098 ;
  assign n23100 = n140 & n23099 ;
  assign n23101 = n22256 & n72913 ;
  assign n23102 = n22988 & n23101 ;
  assign n23103 = n23100 | n23102 ;
  assign n23104 = n69528 & n23103 ;
  assign n72960 = ~n23102 ;
  assign n23591 = x102 & n72960 ;
  assign n72961 = ~n23100 ;
  assign n23592 = n72961 & n23591 ;
  assign n23593 = n23104 | n23592 ;
  assign n72962 = ~n22943 ;
  assign n22945 = n22747 & n72962 ;
  assign n23105 = n22273 | n22747 ;
  assign n72963 = ~n23105 ;
  assign n23106 = n22743 & n72963 ;
  assign n23107 = n22945 | n23106 ;
  assign n23108 = n140 & n23107 ;
  assign n23109 = n22264 & n72913 ;
  assign n23110 = n22988 & n23109 ;
  assign n23111 = n23108 | n23110 ;
  assign n23112 = n69261 & n23111 ;
  assign n72964 = ~n22738 ;
  assign n22742 = n72964 & n22741 ;
  assign n23113 = n22281 | n22741 ;
  assign n72965 = ~n23113 ;
  assign n23114 = n22939 & n72965 ;
  assign n23115 = n22742 | n23114 ;
  assign n23116 = n140 & n23115 ;
  assign n23117 = n22272 & n72913 ;
  assign n23118 = n22988 & n23117 ;
  assign n23119 = n23116 | n23118 ;
  assign n23120 = n69075 & n23119 ;
  assign n72966 = ~n23118 ;
  assign n23581 = x100 & n72966 ;
  assign n72967 = ~n23116 ;
  assign n23582 = n72967 & n23581 ;
  assign n23583 = n23120 | n23582 ;
  assign n72968 = ~n22938 ;
  assign n22940 = n22736 & n72968 ;
  assign n23121 = n22289 | n22736 ;
  assign n72969 = ~n23121 ;
  assign n23122 = n22732 & n72969 ;
  assign n23123 = n22940 | n23122 ;
  assign n23124 = n140 & n23123 ;
  assign n23125 = n22280 & n72913 ;
  assign n23126 = n22988 & n23125 ;
  assign n23127 = n23124 | n23126 ;
  assign n23128 = n68993 & n23127 ;
  assign n72970 = ~n22727 ;
  assign n22731 = n72970 & n22730 ;
  assign n23129 = n22297 | n22730 ;
  assign n72971 = ~n23129 ;
  assign n23130 = n22934 & n72971 ;
  assign n23131 = n22731 | n23130 ;
  assign n23132 = n140 & n23131 ;
  assign n23133 = n22288 & n72913 ;
  assign n23134 = n22988 & n23133 ;
  assign n23135 = n23132 | n23134 ;
  assign n23136 = n68716 & n23135 ;
  assign n72972 = ~n23134 ;
  assign n23571 = x98 & n72972 ;
  assign n72973 = ~n23132 ;
  assign n23572 = n72973 & n23571 ;
  assign n23573 = n23136 | n23572 ;
  assign n72974 = ~n22933 ;
  assign n22935 = n22725 & n72974 ;
  assign n23137 = n22305 | n22725 ;
  assign n72975 = ~n23137 ;
  assign n23138 = n22721 & n72975 ;
  assign n23139 = n22935 | n23138 ;
  assign n23140 = n140 & n23139 ;
  assign n23141 = n22296 & n72913 ;
  assign n23142 = n22988 & n23141 ;
  assign n23143 = n23140 | n23142 ;
  assign n23144 = n68545 & n23143 ;
  assign n72976 = ~n22716 ;
  assign n22720 = n72976 & n22719 ;
  assign n23145 = n22313 | n22719 ;
  assign n72977 = ~n23145 ;
  assign n23146 = n22929 & n72977 ;
  assign n23147 = n22720 | n23146 ;
  assign n23148 = n140 & n23147 ;
  assign n23149 = n22304 & n72913 ;
  assign n23150 = n22988 & n23149 ;
  assign n23151 = n23148 | n23150 ;
  assign n23152 = n68438 & n23151 ;
  assign n72978 = ~n23150 ;
  assign n23561 = x96 & n72978 ;
  assign n72979 = ~n23148 ;
  assign n23562 = n72979 & n23561 ;
  assign n23563 = n23152 | n23562 ;
  assign n72980 = ~n22928 ;
  assign n22930 = n22714 & n72980 ;
  assign n23153 = n22321 | n22714 ;
  assign n72981 = ~n23153 ;
  assign n23154 = n22710 & n72981 ;
  assign n23155 = n22930 | n23154 ;
  assign n23156 = n140 & n23155 ;
  assign n23157 = n22312 & n72913 ;
  assign n23158 = n22988 & n23157 ;
  assign n23159 = n23156 | n23158 ;
  assign n23160 = n68214 & n23159 ;
  assign n72982 = ~n22705 ;
  assign n22709 = n72982 & n22708 ;
  assign n23161 = n22329 | n22708 ;
  assign n72983 = ~n23161 ;
  assign n23162 = n22924 & n72983 ;
  assign n23163 = n22709 | n23162 ;
  assign n23164 = n140 & n23163 ;
  assign n23165 = n22320 & n72913 ;
  assign n23166 = n22988 & n23165 ;
  assign n23167 = n23164 | n23166 ;
  assign n23168 = n68058 & n23167 ;
  assign n72984 = ~n23166 ;
  assign n23551 = x94 & n72984 ;
  assign n72985 = ~n23164 ;
  assign n23552 = n72985 & n23551 ;
  assign n23553 = n23168 | n23552 ;
  assign n72986 = ~n22923 ;
  assign n22925 = n22703 & n72986 ;
  assign n23169 = n22337 | n22703 ;
  assign n72987 = ~n23169 ;
  assign n23170 = n22699 & n72987 ;
  assign n23171 = n22925 | n23170 ;
  assign n23172 = n140 & n23171 ;
  assign n23173 = n22328 & n72913 ;
  assign n23174 = n22988 & n23173 ;
  assign n23175 = n23172 | n23174 ;
  assign n23176 = n67986 & n23175 ;
  assign n72988 = ~n22694 ;
  assign n22698 = n72988 & n22697 ;
  assign n23177 = n22345 | n22697 ;
  assign n72989 = ~n23177 ;
  assign n23178 = n22919 & n72989 ;
  assign n23179 = n22698 | n23178 ;
  assign n23180 = n140 & n23179 ;
  assign n23181 = n22336 & n72913 ;
  assign n23182 = n22988 & n23181 ;
  assign n23183 = n23180 | n23182 ;
  assign n23184 = n67763 & n23183 ;
  assign n72990 = ~n23182 ;
  assign n23541 = x92 & n72990 ;
  assign n72991 = ~n23180 ;
  assign n23542 = n72991 & n23541 ;
  assign n23543 = n23184 | n23542 ;
  assign n72992 = ~n22918 ;
  assign n22920 = n22692 & n72992 ;
  assign n23185 = n22353 | n22692 ;
  assign n72993 = ~n23185 ;
  assign n23186 = n22688 & n72993 ;
  assign n23187 = n22920 | n23186 ;
  assign n23188 = n140 & n23187 ;
  assign n23189 = n22344 & n72913 ;
  assign n23190 = n22988 & n23189 ;
  assign n23191 = n23188 | n23190 ;
  assign n23192 = n67622 & n23191 ;
  assign n72994 = ~n22683 ;
  assign n22687 = n72994 & n22686 ;
  assign n23193 = n22361 | n22686 ;
  assign n72995 = ~n23193 ;
  assign n23194 = n22914 & n72995 ;
  assign n23195 = n22687 | n23194 ;
  assign n23196 = n140 & n23195 ;
  assign n23197 = n22352 & n72913 ;
  assign n23198 = n22988 & n23197 ;
  assign n23199 = n23196 | n23198 ;
  assign n23200 = n67531 & n23199 ;
  assign n72996 = ~n23198 ;
  assign n23531 = x90 & n72996 ;
  assign n72997 = ~n23196 ;
  assign n23532 = n72997 & n23531 ;
  assign n23533 = n23200 | n23532 ;
  assign n72998 = ~n22913 ;
  assign n22915 = n22681 & n72998 ;
  assign n23201 = n22369 | n22681 ;
  assign n72999 = ~n23201 ;
  assign n23202 = n22677 & n72999 ;
  assign n23203 = n22915 | n23202 ;
  assign n23204 = n140 & n23203 ;
  assign n23205 = n22360 & n72913 ;
  assign n23206 = n22988 & n23205 ;
  assign n23207 = n23204 | n23206 ;
  assign n23208 = n67348 & n23207 ;
  assign n73000 = ~n22672 ;
  assign n22676 = n73000 & n22675 ;
  assign n23209 = n22377 | n22675 ;
  assign n73001 = ~n23209 ;
  assign n23210 = n22909 & n73001 ;
  assign n23211 = n22676 | n23210 ;
  assign n23212 = n140 & n23211 ;
  assign n23213 = n22368 & n72913 ;
  assign n23214 = n22988 & n23213 ;
  assign n23215 = n23212 | n23214 ;
  assign n23216 = n67222 & n23215 ;
  assign n73002 = ~n23214 ;
  assign n23520 = x88 & n73002 ;
  assign n73003 = ~n23212 ;
  assign n23521 = n73003 & n23520 ;
  assign n23522 = n23216 | n23521 ;
  assign n73004 = ~n22908 ;
  assign n22910 = n22670 & n73004 ;
  assign n23217 = n22385 | n22670 ;
  assign n73005 = ~n23217 ;
  assign n23218 = n22666 & n73005 ;
  assign n23219 = n22910 | n23218 ;
  assign n23220 = n140 & n23219 ;
  assign n23221 = n22376 & n72913 ;
  assign n23222 = n22988 & n23221 ;
  assign n23223 = n23220 | n23222 ;
  assign n23224 = n67164 & n23223 ;
  assign n73006 = ~n22661 ;
  assign n22665 = n73006 & n22664 ;
  assign n23225 = n22393 | n22664 ;
  assign n73007 = ~n23225 ;
  assign n23226 = n22904 & n73007 ;
  assign n23227 = n22665 | n23226 ;
  assign n23228 = n140 & n23227 ;
  assign n23229 = n22384 & n72913 ;
  assign n23230 = n22988 & n23229 ;
  assign n23231 = n23228 | n23230 ;
  assign n23232 = n66979 & n23231 ;
  assign n73008 = ~n23230 ;
  assign n23510 = x86 & n73008 ;
  assign n73009 = ~n23228 ;
  assign n23511 = n73009 & n23510 ;
  assign n23512 = n23232 | n23511 ;
  assign n73010 = ~n22903 ;
  assign n22905 = n22659 & n73010 ;
  assign n23233 = n22401 | n22659 ;
  assign n73011 = ~n23233 ;
  assign n23234 = n22655 & n73011 ;
  assign n23235 = n22905 | n23234 ;
  assign n23236 = n140 & n23235 ;
  assign n23237 = n22392 & n72913 ;
  assign n23238 = n22988 & n23237 ;
  assign n23239 = n23236 | n23238 ;
  assign n23240 = n66868 & n23239 ;
  assign n73012 = ~n22650 ;
  assign n22654 = n73012 & n22653 ;
  assign n23241 = n22409 | n22653 ;
  assign n73013 = ~n23241 ;
  assign n23242 = n22899 & n73013 ;
  assign n23243 = n22654 | n23242 ;
  assign n23244 = n140 & n23243 ;
  assign n23245 = n22400 & n72913 ;
  assign n23246 = n22988 & n23245 ;
  assign n23247 = n23244 | n23246 ;
  assign n23248 = n66797 & n23247 ;
  assign n73014 = ~n23246 ;
  assign n23498 = x84 & n73014 ;
  assign n73015 = ~n23244 ;
  assign n23499 = n73015 & n23498 ;
  assign n23500 = n23248 | n23499 ;
  assign n73016 = ~n22898 ;
  assign n22900 = n22648 & n73016 ;
  assign n23249 = n22417 | n22648 ;
  assign n73017 = ~n23249 ;
  assign n23250 = n22644 & n73017 ;
  assign n23251 = n22900 | n23250 ;
  assign n23252 = n140 & n23251 ;
  assign n23253 = n22408 & n72913 ;
  assign n23254 = n22988 & n23253 ;
  assign n23255 = n23252 | n23254 ;
  assign n23256 = n66654 & n23255 ;
  assign n73018 = ~n22639 ;
  assign n22643 = n73018 & n22642 ;
  assign n23257 = n22425 | n22642 ;
  assign n73019 = ~n23257 ;
  assign n23258 = n22894 & n73019 ;
  assign n23259 = n22643 | n23258 ;
  assign n23260 = n140 & n23259 ;
  assign n23261 = n22416 & n72913 ;
  assign n23262 = n22988 & n23261 ;
  assign n23263 = n23260 | n23262 ;
  assign n23264 = n66560 & n23263 ;
  assign n73020 = ~n23262 ;
  assign n23488 = x82 & n73020 ;
  assign n73021 = ~n23260 ;
  assign n23489 = n73021 & n23488 ;
  assign n23490 = n23264 | n23489 ;
  assign n73022 = ~n22893 ;
  assign n22895 = n22637 & n73022 ;
  assign n23265 = n22433 | n22637 ;
  assign n73023 = ~n23265 ;
  assign n23266 = n22633 & n73023 ;
  assign n23267 = n22895 | n23266 ;
  assign n23268 = n140 & n23267 ;
  assign n23269 = n22424 & n72913 ;
  assign n23270 = n22988 & n23269 ;
  assign n23271 = n23268 | n23270 ;
  assign n23272 = n66505 & n23271 ;
  assign n73024 = ~n22628 ;
  assign n22632 = n73024 & n22631 ;
  assign n23273 = n22441 | n22631 ;
  assign n73025 = ~n23273 ;
  assign n23274 = n22889 & n73025 ;
  assign n23275 = n22632 | n23274 ;
  assign n23276 = n140 & n23275 ;
  assign n23277 = n22432 & n72913 ;
  assign n23278 = n22988 & n23277 ;
  assign n23279 = n23276 | n23278 ;
  assign n23280 = n66379 & n23279 ;
  assign n73026 = ~n23278 ;
  assign n23477 = x80 & n73026 ;
  assign n73027 = ~n23276 ;
  assign n23478 = n73027 & n23477 ;
  assign n23479 = n23280 | n23478 ;
  assign n73028 = ~n22888 ;
  assign n22890 = n22626 & n73028 ;
  assign n23281 = n22449 | n22626 ;
  assign n73029 = ~n23281 ;
  assign n23282 = n22622 & n73029 ;
  assign n23283 = n22890 | n23282 ;
  assign n23284 = n140 & n23283 ;
  assign n23285 = n22440 & n72913 ;
  assign n23286 = n22988 & n23285 ;
  assign n23287 = n23284 | n23286 ;
  assign n23288 = n66299 & n23287 ;
  assign n73030 = ~n22617 ;
  assign n22621 = n73030 & n22620 ;
  assign n23289 = n22457 | n22620 ;
  assign n73031 = ~n23289 ;
  assign n23290 = n22884 & n73031 ;
  assign n23291 = n22621 | n23290 ;
  assign n23292 = n140 & n23291 ;
  assign n23293 = n22448 & n72913 ;
  assign n23294 = n22988 & n23293 ;
  assign n23295 = n23292 | n23294 ;
  assign n23296 = n66244 & n23295 ;
  assign n73032 = ~n23294 ;
  assign n23466 = x78 & n73032 ;
  assign n73033 = ~n23292 ;
  assign n23467 = n73033 & n23466 ;
  assign n23468 = n23296 | n23467 ;
  assign n73034 = ~n22883 ;
  assign n22885 = n22615 & n73034 ;
  assign n23297 = n22465 | n22615 ;
  assign n73035 = ~n23297 ;
  assign n23298 = n22611 & n73035 ;
  assign n23299 = n22885 | n23298 ;
  assign n23300 = n140 & n23299 ;
  assign n23301 = n22456 & n72913 ;
  assign n23302 = n22988 & n23301 ;
  assign n23303 = n23300 | n23302 ;
  assign n23304 = n66145 & n23303 ;
  assign n73036 = ~n22606 ;
  assign n22610 = n73036 & n22609 ;
  assign n23305 = n22473 | n22609 ;
  assign n73037 = ~n23305 ;
  assign n23306 = n22879 & n73037 ;
  assign n23307 = n22610 | n23306 ;
  assign n23308 = n140 & n23307 ;
  assign n23309 = n22464 & n72913 ;
  assign n23310 = n22988 & n23309 ;
  assign n23311 = n23308 | n23310 ;
  assign n23312 = n66081 & n23311 ;
  assign n73038 = ~n23310 ;
  assign n23456 = x76 & n73038 ;
  assign n73039 = ~n23308 ;
  assign n23457 = n73039 & n23456 ;
  assign n23458 = n23312 | n23457 ;
  assign n73040 = ~n22878 ;
  assign n22880 = n22604 & n73040 ;
  assign n23313 = n22481 | n22604 ;
  assign n73041 = ~n23313 ;
  assign n23314 = n22600 & n73041 ;
  assign n23315 = n22880 | n23314 ;
  assign n23316 = n140 & n23315 ;
  assign n23317 = n22472 & n72913 ;
  assign n23318 = n22988 & n23317 ;
  assign n23319 = n23316 | n23318 ;
  assign n23320 = n66043 & n23319 ;
  assign n73042 = ~n22595 ;
  assign n22599 = n73042 & n22598 ;
  assign n23321 = n22489 | n22598 ;
  assign n73043 = ~n23321 ;
  assign n23322 = n22874 & n73043 ;
  assign n23323 = n22599 | n23322 ;
  assign n23324 = n140 & n23323 ;
  assign n23325 = n22480 & n72913 ;
  assign n23326 = n22988 & n23325 ;
  assign n23327 = n23324 | n23326 ;
  assign n23328 = n65960 & n23327 ;
  assign n73044 = ~n23326 ;
  assign n23446 = x74 & n73044 ;
  assign n73045 = ~n23324 ;
  assign n23447 = n73045 & n23446 ;
  assign n23448 = n23328 | n23447 ;
  assign n73046 = ~n22873 ;
  assign n22875 = n22593 & n73046 ;
  assign n23329 = n22497 | n22593 ;
  assign n73047 = ~n23329 ;
  assign n23330 = n22589 & n73047 ;
  assign n23331 = n22875 | n23330 ;
  assign n23332 = n140 & n23331 ;
  assign n23333 = n22488 & n72913 ;
  assign n23334 = n22988 & n23333 ;
  assign n23335 = n23332 | n23334 ;
  assign n23336 = n65909 & n23335 ;
  assign n73048 = ~n22584 ;
  assign n22588 = n73048 & n22587 ;
  assign n23337 = n22505 | n22587 ;
  assign n73049 = ~n23337 ;
  assign n23338 = n22869 & n73049 ;
  assign n23339 = n22588 | n23338 ;
  assign n23340 = n140 & n23339 ;
  assign n23341 = n22496 & n72913 ;
  assign n23342 = n22988 & n23341 ;
  assign n23343 = n23340 | n23342 ;
  assign n23344 = n65877 & n23343 ;
  assign n73050 = ~n23342 ;
  assign n23435 = x72 & n73050 ;
  assign n73051 = ~n23340 ;
  assign n23436 = n73051 & n23435 ;
  assign n23437 = n23344 | n23436 ;
  assign n73052 = ~n22868 ;
  assign n22870 = n22582 & n73052 ;
  assign n23345 = n22514 | n22582 ;
  assign n73053 = ~n23345 ;
  assign n23346 = n22578 & n73053 ;
  assign n23347 = n22870 | n23346 ;
  assign n23348 = n140 & n23347 ;
  assign n23349 = n22504 & n72913 ;
  assign n23350 = n22988 & n23349 ;
  assign n23351 = n23348 | n23350 ;
  assign n23352 = n65820 & n23351 ;
  assign n73054 = ~n22574 ;
  assign n22866 = n73054 & n22577 ;
  assign n23353 = n22523 | n22577 ;
  assign n73055 = ~n23353 ;
  assign n23354 = n22864 & n73055 ;
  assign n23355 = n22866 | n23354 ;
  assign n23356 = n140 & n23355 ;
  assign n23357 = n22513 & n72913 ;
  assign n23358 = n22988 & n23357 ;
  assign n23359 = n23356 | n23358 ;
  assign n23360 = n65791 & n23359 ;
  assign n73056 = ~n23358 ;
  assign n23425 = x70 & n73056 ;
  assign n73057 = ~n23356 ;
  assign n23426 = n73057 & n23425 ;
  assign n23427 = n23360 | n23426 ;
  assign n73058 = ~n22862 ;
  assign n22863 = n22572 & n73058 ;
  assign n23361 = n22565 | n22859 ;
  assign n23362 = n22531 | n22572 ;
  assign n73059 = ~n23362 ;
  assign n23363 = n23361 & n73059 ;
  assign n23364 = n22863 | n23363 ;
  assign n23365 = n140 & n23364 ;
  assign n23366 = n22522 & n72913 ;
  assign n23367 = n22988 & n23366 ;
  assign n23368 = n23365 | n23367 ;
  assign n23369 = n65772 & n23368 ;
  assign n73060 = ~n22565 ;
  assign n22860 = n73060 & n22859 ;
  assign n23370 = n22537 | n22859 ;
  assign n73061 = ~n23370 ;
  assign n23371 = n22564 & n73061 ;
  assign n23372 = n22860 | n23371 ;
  assign n23373 = n140 & n23372 ;
  assign n23374 = n22530 & n72913 ;
  assign n23375 = n22988 & n23374 ;
  assign n23376 = n23373 | n23375 ;
  assign n23377 = n65746 & n23376 ;
  assign n73062 = ~n23375 ;
  assign n23415 = x68 & n73062 ;
  assign n73063 = ~n23373 ;
  assign n23416 = n73063 & n23415 ;
  assign n23417 = n23377 | n23416 ;
  assign n73064 = ~n22855 ;
  assign n22856 = n22563 & n73064 ;
  assign n23378 = n22559 | n22563 ;
  assign n73065 = ~n23378 ;
  assign n23379 = n22558 & n73065 ;
  assign n23380 = n22856 | n23379 ;
  assign n23381 = n140 & n23380 ;
  assign n23382 = n22536 & n72913 ;
  assign n23383 = n22988 & n23382 ;
  assign n23384 = n23381 | n23383 ;
  assign n23385 = n65721 & n23384 ;
  assign n23386 = n22555 & n22557 ;
  assign n23387 = n72757 & n23386 ;
  assign n73066 = ~n23387 ;
  assign n23388 = n22854 & n73066 ;
  assign n23389 = n140 & n23388 ;
  assign n23390 = n72913 & n22851 ;
  assign n23391 = n22988 & n23390 ;
  assign n23392 = n23389 | n23391 ;
  assign n23393 = n65686 & n23392 ;
  assign n73067 = ~n23391 ;
  assign n23405 = x66 & n73067 ;
  assign n73068 = ~n23389 ;
  assign n23406 = n73068 & n23405 ;
  assign n23407 = n23393 | n23406 ;
  assign n22850 = n22557 & n140 ;
  assign n22849 = x64 & n140 ;
  assign n73069 = ~n22849 ;
  assign n23394 = x11 & n73069 ;
  assign n23395 = n22850 | n23394 ;
  assign n23396 = x65 & n23395 ;
  assign n23397 = n72913 & n22988 ;
  assign n73070 = ~n23397 ;
  assign n23398 = n22557 & n73070 ;
  assign n23399 = x65 | n23398 ;
  assign n23400 = n23394 | n23399 ;
  assign n73071 = ~n23396 ;
  assign n23401 = n73071 & n23400 ;
  assign n73072 = ~x10 ;
  assign n23402 = n73072 & x64 ;
  assign n23403 = n23401 | n23402 ;
  assign n23404 = n65670 & n23395 ;
  assign n73073 = ~n23404 ;
  assign n23408 = n23403 & n73073 ;
  assign n23409 = n23407 | n23408 ;
  assign n73074 = ~n23393 ;
  assign n23410 = n73074 & n23409 ;
  assign n73075 = ~n23383 ;
  assign n23411 = x67 & n73075 ;
  assign n73076 = ~n23381 ;
  assign n23412 = n73076 & n23411 ;
  assign n23413 = n23385 | n23412 ;
  assign n23414 = n23410 | n23413 ;
  assign n73077 = ~n23385 ;
  assign n23418 = n73077 & n23414 ;
  assign n23419 = n23417 | n23418 ;
  assign n73078 = ~n23377 ;
  assign n23420 = n73078 & n23419 ;
  assign n73079 = ~n23367 ;
  assign n23421 = x69 & n73079 ;
  assign n73080 = ~n23365 ;
  assign n23422 = n73080 & n23421 ;
  assign n23423 = n23369 | n23422 ;
  assign n23424 = n23420 | n23423 ;
  assign n73081 = ~n23369 ;
  assign n23428 = n73081 & n23424 ;
  assign n23429 = n23427 | n23428 ;
  assign n73082 = ~n23360 ;
  assign n23430 = n73082 & n23429 ;
  assign n73083 = ~n23350 ;
  assign n23431 = x71 & n73083 ;
  assign n73084 = ~n23348 ;
  assign n23432 = n73084 & n23431 ;
  assign n23433 = n23352 | n23432 ;
  assign n23434 = n23430 | n23433 ;
  assign n73085 = ~n23352 ;
  assign n23438 = n73085 & n23434 ;
  assign n23439 = n23437 | n23438 ;
  assign n73086 = ~n23344 ;
  assign n23440 = n73086 & n23439 ;
  assign n73087 = ~n23334 ;
  assign n23441 = x73 & n73087 ;
  assign n73088 = ~n23332 ;
  assign n23442 = n73088 & n23441 ;
  assign n23443 = n23336 | n23442 ;
  assign n23445 = n23440 | n23443 ;
  assign n73089 = ~n23336 ;
  assign n23449 = n73089 & n23445 ;
  assign n23450 = n23448 | n23449 ;
  assign n73090 = ~n23328 ;
  assign n23451 = n73090 & n23450 ;
  assign n73091 = ~n23318 ;
  assign n23452 = x75 & n73091 ;
  assign n73092 = ~n23316 ;
  assign n23453 = n73092 & n23452 ;
  assign n23454 = n23320 | n23453 ;
  assign n23455 = n23451 | n23454 ;
  assign n73093 = ~n23320 ;
  assign n23459 = n73093 & n23455 ;
  assign n23460 = n23458 | n23459 ;
  assign n73094 = ~n23312 ;
  assign n23461 = n73094 & n23460 ;
  assign n73095 = ~n23302 ;
  assign n23462 = x77 & n73095 ;
  assign n73096 = ~n23300 ;
  assign n23463 = n73096 & n23462 ;
  assign n23464 = n23304 | n23463 ;
  assign n23465 = n23461 | n23464 ;
  assign n73097 = ~n23304 ;
  assign n23469 = n73097 & n23465 ;
  assign n23470 = n23468 | n23469 ;
  assign n73098 = ~n23296 ;
  assign n23471 = n73098 & n23470 ;
  assign n73099 = ~n23286 ;
  assign n23472 = x79 & n73099 ;
  assign n73100 = ~n23284 ;
  assign n23473 = n73100 & n23472 ;
  assign n23474 = n23288 | n23473 ;
  assign n23476 = n23471 | n23474 ;
  assign n73101 = ~n23288 ;
  assign n23481 = n73101 & n23476 ;
  assign n23482 = n23479 | n23481 ;
  assign n73102 = ~n23280 ;
  assign n23483 = n73102 & n23482 ;
  assign n73103 = ~n23270 ;
  assign n23484 = x81 & n73103 ;
  assign n73104 = ~n23268 ;
  assign n23485 = n73104 & n23484 ;
  assign n23486 = n23272 | n23485 ;
  assign n23487 = n23483 | n23486 ;
  assign n73105 = ~n23272 ;
  assign n23491 = n73105 & n23487 ;
  assign n23492 = n23490 | n23491 ;
  assign n73106 = ~n23264 ;
  assign n23493 = n73106 & n23492 ;
  assign n73107 = ~n23254 ;
  assign n23494 = x83 & n73107 ;
  assign n73108 = ~n23252 ;
  assign n23495 = n73108 & n23494 ;
  assign n23496 = n23256 | n23495 ;
  assign n23497 = n23493 | n23496 ;
  assign n73109 = ~n23256 ;
  assign n23502 = n73109 & n23497 ;
  assign n23503 = n23500 | n23502 ;
  assign n73110 = ~n23248 ;
  assign n23504 = n73110 & n23503 ;
  assign n73111 = ~n23238 ;
  assign n23505 = x85 & n73111 ;
  assign n73112 = ~n23236 ;
  assign n23506 = n73112 & n23505 ;
  assign n23507 = n23240 | n23506 ;
  assign n23509 = n23504 | n23507 ;
  assign n73113 = ~n23240 ;
  assign n23513 = n73113 & n23509 ;
  assign n23514 = n23512 | n23513 ;
  assign n73114 = ~n23232 ;
  assign n23515 = n73114 & n23514 ;
  assign n73115 = ~n23222 ;
  assign n23516 = x87 & n73115 ;
  assign n73116 = ~n23220 ;
  assign n23517 = n73116 & n23516 ;
  assign n23518 = n23224 | n23517 ;
  assign n23519 = n23515 | n23518 ;
  assign n73117 = ~n23224 ;
  assign n23524 = n73117 & n23519 ;
  assign n23525 = n23522 | n23524 ;
  assign n73118 = ~n23216 ;
  assign n23526 = n73118 & n23525 ;
  assign n73119 = ~n23206 ;
  assign n23527 = x89 & n73119 ;
  assign n73120 = ~n23204 ;
  assign n23528 = n73120 & n23527 ;
  assign n23529 = n23208 | n23528 ;
  assign n23530 = n23526 | n23529 ;
  assign n73121 = ~n23208 ;
  assign n23534 = n73121 & n23530 ;
  assign n23535 = n23533 | n23534 ;
  assign n73122 = ~n23200 ;
  assign n23536 = n73122 & n23535 ;
  assign n73123 = ~n23190 ;
  assign n23537 = x91 & n73123 ;
  assign n73124 = ~n23188 ;
  assign n23538 = n73124 & n23537 ;
  assign n23539 = n23192 | n23538 ;
  assign n23540 = n23536 | n23539 ;
  assign n73125 = ~n23192 ;
  assign n23544 = n73125 & n23540 ;
  assign n23545 = n23543 | n23544 ;
  assign n73126 = ~n23184 ;
  assign n23546 = n73126 & n23545 ;
  assign n73127 = ~n23174 ;
  assign n23547 = x93 & n73127 ;
  assign n73128 = ~n23172 ;
  assign n23548 = n73128 & n23547 ;
  assign n23549 = n23176 | n23548 ;
  assign n23550 = n23546 | n23549 ;
  assign n73129 = ~n23176 ;
  assign n23554 = n73129 & n23550 ;
  assign n23555 = n23553 | n23554 ;
  assign n73130 = ~n23168 ;
  assign n23556 = n73130 & n23555 ;
  assign n73131 = ~n23158 ;
  assign n23557 = x95 & n73131 ;
  assign n73132 = ~n23156 ;
  assign n23558 = n73132 & n23557 ;
  assign n23559 = n23160 | n23558 ;
  assign n23560 = n23556 | n23559 ;
  assign n73133 = ~n23160 ;
  assign n23564 = n73133 & n23560 ;
  assign n23565 = n23563 | n23564 ;
  assign n73134 = ~n23152 ;
  assign n23566 = n73134 & n23565 ;
  assign n73135 = ~n23142 ;
  assign n23567 = x97 & n73135 ;
  assign n73136 = ~n23140 ;
  assign n23568 = n73136 & n23567 ;
  assign n23569 = n23144 | n23568 ;
  assign n23570 = n23566 | n23569 ;
  assign n73137 = ~n23144 ;
  assign n23574 = n73137 & n23570 ;
  assign n23575 = n23573 | n23574 ;
  assign n73138 = ~n23136 ;
  assign n23576 = n73138 & n23575 ;
  assign n73139 = ~n23126 ;
  assign n23577 = x99 & n73139 ;
  assign n73140 = ~n23124 ;
  assign n23578 = n73140 & n23577 ;
  assign n23579 = n23128 | n23578 ;
  assign n23580 = n23576 | n23579 ;
  assign n73141 = ~n23128 ;
  assign n23584 = n73141 & n23580 ;
  assign n23585 = n23583 | n23584 ;
  assign n73142 = ~n23120 ;
  assign n23586 = n73142 & n23585 ;
  assign n73143 = ~n23110 ;
  assign n23587 = x101 & n73143 ;
  assign n73144 = ~n23108 ;
  assign n23588 = n73144 & n23587 ;
  assign n23589 = n23112 | n23588 ;
  assign n23590 = n23586 | n23589 ;
  assign n73145 = ~n23112 ;
  assign n23594 = n73145 & n23590 ;
  assign n23595 = n23593 | n23594 ;
  assign n73146 = ~n23104 ;
  assign n23596 = n73146 & n23595 ;
  assign n73147 = ~n23094 ;
  assign n23597 = x103 & n73147 ;
  assign n73148 = ~n23092 ;
  assign n23598 = n73148 & n23597 ;
  assign n23599 = n23096 | n23598 ;
  assign n23600 = n23596 | n23599 ;
  assign n73149 = ~n23096 ;
  assign n23605 = n73149 & n23600 ;
  assign n23606 = n23603 | n23605 ;
  assign n73150 = ~n23088 ;
  assign n23607 = n73150 & n23606 ;
  assign n73151 = ~n23078 ;
  assign n23608 = x105 & n73151 ;
  assign n73152 = ~n23076 ;
  assign n23609 = n73152 & n23608 ;
  assign n23610 = n23080 | n23609 ;
  assign n23611 = n23607 | n23610 ;
  assign n73153 = ~n23080 ;
  assign n23615 = n73153 & n23611 ;
  assign n23616 = n23614 | n23615 ;
  assign n73154 = ~n23072 ;
  assign n23617 = n73154 & n23616 ;
  assign n73155 = ~n23062 ;
  assign n23618 = x107 & n73155 ;
  assign n73156 = ~n23060 ;
  assign n23619 = n73156 & n23618 ;
  assign n23620 = n23064 | n23619 ;
  assign n23621 = n23617 | n23620 ;
  assign n73157 = ~n23064 ;
  assign n23626 = n73157 & n23621 ;
  assign n23627 = n23624 | n23626 ;
  assign n73158 = ~n23056 ;
  assign n23628 = n73158 & n23627 ;
  assign n73159 = ~n23046 ;
  assign n23629 = x109 & n73159 ;
  assign n73160 = ~n23044 ;
  assign n23630 = n73160 & n23629 ;
  assign n23631 = n23048 | n23630 ;
  assign n23632 = n23628 | n23631 ;
  assign n73161 = ~n23048 ;
  assign n23636 = n73161 & n23632 ;
  assign n23637 = n23635 | n23636 ;
  assign n73162 = ~n23040 ;
  assign n23638 = n73162 & n23637 ;
  assign n73163 = ~n23030 ;
  assign n23639 = x111 & n73163 ;
  assign n73164 = ~n23028 ;
  assign n23640 = n73164 & n23639 ;
  assign n23641 = n23032 | n23640 ;
  assign n23642 = n23638 | n23641 ;
  assign n73165 = ~n23032 ;
  assign n23646 = n73165 & n23642 ;
  assign n23647 = n23645 | n23646 ;
  assign n73166 = ~n23024 ;
  assign n23648 = n73166 & n23647 ;
  assign n73167 = ~n23014 ;
  assign n23649 = x113 & n73167 ;
  assign n73168 = ~n23012 ;
  assign n23650 = n73168 & n23649 ;
  assign n23651 = n23016 | n23650 ;
  assign n23653 = n23648 | n23651 ;
  assign n73169 = ~n23016 ;
  assign n23657 = n73169 & n23653 ;
  assign n23658 = n23656 | n23657 ;
  assign n73170 = ~n23008 ;
  assign n23659 = n73170 & n23658 ;
  assign n73171 = ~n22998 ;
  assign n23660 = x115 & n73171 ;
  assign n73172 = ~n22996 ;
  assign n23661 = n73172 & n23660 ;
  assign n23662 = n23000 | n23661 ;
  assign n23663 = n23659 | n23662 ;
  assign n73173 = ~n23000 ;
  assign n23667 = n73173 & n23663 ;
  assign n23668 = n23666 | n23667 ;
  assign n73174 = ~n22992 ;
  assign n23669 = n73174 & n23668 ;
  assign n23670 = n22145 | n22843 ;
  assign n23671 = n22839 | n23670 ;
  assign n73175 = ~n23671 ;
  assign n23672 = n22831 & n73175 ;
  assign n23673 = n22839 | n22843 ;
  assign n73176 = ~n22987 ;
  assign n23674 = n73176 & n23673 ;
  assign n23675 = n23672 | n23674 ;
  assign n23676 = n140 & n23675 ;
  assign n23677 = n65429 & n21327 ;
  assign n23678 = n22988 & n23677 ;
  assign n23679 = n23676 | n23678 ;
  assign n73177 = ~x117 ;
  assign n23680 = n73177 & n23679 ;
  assign n73178 = ~n23678 ;
  assign n23681 = x117 & n73178 ;
  assign n73179 = ~n23676 ;
  assign n23682 = n73179 & n23681 ;
  assign n23683 = n65392 | n65407 ;
  assign n23684 = n65369 | n23683 ;
  assign n23685 = n23682 | n23684 ;
  assign n23686 = n23680 | n23685 ;
  assign n23687 = n23669 | n23686 ;
  assign n23688 = n67026 & n23679 ;
  assign n73180 = ~n23688 ;
  assign n23689 = n23687 & n73180 ;
  assign n73181 = ~n23667 ;
  assign n23810 = n23666 & n73181 ;
  assign n23702 = x64 & n73070 ;
  assign n73182 = ~n23702 ;
  assign n23703 = x11 & n73182 ;
  assign n23704 = n22850 | n23703 ;
  assign n23705 = x65 & n23704 ;
  assign n73183 = ~n23705 ;
  assign n23706 = n23400 & n73183 ;
  assign n23707 = n23402 | n23706 ;
  assign n23708 = n73073 & n23707 ;
  assign n23710 = n23407 | n23708 ;
  assign n23711 = n73074 & n23710 ;
  assign n23712 = n23413 | n23711 ;
  assign n23713 = n73077 & n23712 ;
  assign n23714 = n23417 | n23713 ;
  assign n23715 = n73078 & n23714 ;
  assign n23716 = n23423 | n23715 ;
  assign n23717 = n73081 & n23716 ;
  assign n23718 = n23427 | n23717 ;
  assign n23719 = n73082 & n23718 ;
  assign n23720 = n23433 | n23719 ;
  assign n23721 = n73085 & n23720 ;
  assign n23722 = n23437 | n23721 ;
  assign n23723 = n73086 & n23722 ;
  assign n23724 = n23443 | n23723 ;
  assign n23725 = n73089 & n23724 ;
  assign n23726 = n23448 | n23725 ;
  assign n23727 = n73090 & n23726 ;
  assign n23728 = n23454 | n23727 ;
  assign n23729 = n73093 & n23728 ;
  assign n23730 = n23458 | n23729 ;
  assign n23731 = n73094 & n23730 ;
  assign n23732 = n23464 | n23731 ;
  assign n23733 = n73097 & n23732 ;
  assign n23734 = n23468 | n23733 ;
  assign n23735 = n73098 & n23734 ;
  assign n23736 = n23474 | n23735 ;
  assign n23737 = n73101 & n23736 ;
  assign n23738 = n23479 | n23737 ;
  assign n23739 = n73102 & n23738 ;
  assign n23740 = n23486 | n23739 ;
  assign n23741 = n73105 & n23740 ;
  assign n23742 = n23490 | n23741 ;
  assign n23743 = n73106 & n23742 ;
  assign n23744 = n23496 | n23743 ;
  assign n23745 = n73109 & n23744 ;
  assign n23746 = n23500 | n23745 ;
  assign n23747 = n73110 & n23746 ;
  assign n23748 = n23507 | n23747 ;
  assign n23749 = n73113 & n23748 ;
  assign n23750 = n23512 | n23749 ;
  assign n23751 = n73114 & n23750 ;
  assign n23752 = n23518 | n23751 ;
  assign n23753 = n73117 & n23752 ;
  assign n23754 = n23522 | n23753 ;
  assign n23755 = n73118 & n23754 ;
  assign n23756 = n23529 | n23755 ;
  assign n23757 = n73121 & n23756 ;
  assign n23758 = n23533 | n23757 ;
  assign n23759 = n73122 & n23758 ;
  assign n23760 = n23539 | n23759 ;
  assign n23761 = n73125 & n23760 ;
  assign n23762 = n23543 | n23761 ;
  assign n23763 = n73126 & n23762 ;
  assign n23764 = n23549 | n23763 ;
  assign n23765 = n73129 & n23764 ;
  assign n23766 = n23553 | n23765 ;
  assign n23767 = n73130 & n23766 ;
  assign n23768 = n23559 | n23767 ;
  assign n23769 = n73133 & n23768 ;
  assign n23770 = n23563 | n23769 ;
  assign n23771 = n73134 & n23770 ;
  assign n23772 = n23569 | n23771 ;
  assign n23773 = n73137 & n23772 ;
  assign n23774 = n23573 | n23773 ;
  assign n23775 = n73138 & n23774 ;
  assign n23776 = n23579 | n23775 ;
  assign n23777 = n73141 & n23776 ;
  assign n23778 = n23583 | n23777 ;
  assign n23779 = n73142 & n23778 ;
  assign n23780 = n23589 | n23779 ;
  assign n23781 = n73145 & n23780 ;
  assign n23782 = n23593 | n23781 ;
  assign n23783 = n73146 & n23782 ;
  assign n23784 = n23599 | n23783 ;
  assign n23785 = n73149 & n23784 ;
  assign n23786 = n23603 | n23785 ;
  assign n23787 = n73150 & n23786 ;
  assign n23788 = n23610 | n23787 ;
  assign n23789 = n73153 & n23788 ;
  assign n23790 = n23614 | n23789 ;
  assign n23791 = n73154 & n23790 ;
  assign n23792 = n23620 | n23791 ;
  assign n23793 = n73157 & n23792 ;
  assign n23794 = n23624 | n23793 ;
  assign n23795 = n73158 & n23794 ;
  assign n23796 = n23631 | n23795 ;
  assign n23797 = n73161 & n23796 ;
  assign n23798 = n23635 | n23797 ;
  assign n23799 = n73162 & n23798 ;
  assign n23800 = n23641 | n23799 ;
  assign n23801 = n73165 & n23800 ;
  assign n23802 = n23645 | n23801 ;
  assign n23803 = n73166 & n23802 ;
  assign n23804 = n23651 | n23803 ;
  assign n23805 = n73169 & n23804 ;
  assign n23806 = n23656 | n23805 ;
  assign n23807 = n73170 & n23806 ;
  assign n23808 = n23662 | n23807 ;
  assign n23811 = n23000 | n23666 ;
  assign n73184 = ~n23811 ;
  assign n23812 = n23808 & n73184 ;
  assign n23813 = n23810 | n23812 ;
  assign n139 = ~n23689 ;
  assign n23814 = n139 & n23813 ;
  assign n23815 = n22991 & n73180 ;
  assign n23816 = n23687 & n23815 ;
  assign n23817 = n23814 | n23816 ;
  assign n23691 = n22992 | n23682 ;
  assign n23692 = n23680 | n23691 ;
  assign n73186 = ~n23692 ;
  assign n23693 = n23668 & n73186 ;
  assign n23694 = n23680 | n23682 ;
  assign n73187 = ~n23669 ;
  assign n23695 = n73187 & n23694 ;
  assign n23696 = n23693 | n23695 ;
  assign n23697 = n139 & n23696 ;
  assign n23698 = n465 & n23679 ;
  assign n23699 = n23687 & n23698 ;
  assign n23700 = n23697 | n23699 ;
  assign n73188 = ~x118 ;
  assign n23701 = n73188 & n23700 ;
  assign n23818 = n73177 & n23817 ;
  assign n73189 = ~n23807 ;
  assign n23819 = n23662 & n73189 ;
  assign n23820 = n23008 | n23662 ;
  assign n73190 = ~n23820 ;
  assign n23821 = n23658 & n73190 ;
  assign n23822 = n23819 | n23821 ;
  assign n23823 = n139 & n23822 ;
  assign n23824 = n22999 & n73180 ;
  assign n23825 = n23687 & n23824 ;
  assign n23826 = n23823 | n23825 ;
  assign n23827 = n72752 & n23826 ;
  assign n73191 = ~n23657 ;
  assign n23828 = n23656 & n73191 ;
  assign n23829 = n23016 | n23656 ;
  assign n73192 = ~n23829 ;
  assign n23830 = n23804 & n73192 ;
  assign n23831 = n23828 | n23830 ;
  assign n23832 = n139 & n23831 ;
  assign n23833 = n23007 & n73180 ;
  assign n23834 = n23687 & n23833 ;
  assign n23835 = n23832 | n23834 ;
  assign n23836 = n72393 & n23835 ;
  assign n73193 = ~n23803 ;
  assign n23837 = n23651 & n73193 ;
  assign n23652 = n23024 | n23651 ;
  assign n73194 = ~n23652 ;
  assign n23838 = n73194 & n23802 ;
  assign n23839 = n23837 | n23838 ;
  assign n23840 = n139 & n23839 ;
  assign n23841 = n23015 & n73180 ;
  assign n23842 = n23687 & n23841 ;
  assign n23843 = n23840 | n23842 ;
  assign n23844 = n72385 & n23843 ;
  assign n73195 = ~n23646 ;
  assign n23845 = n23645 & n73195 ;
  assign n23846 = n23032 | n23645 ;
  assign n73196 = ~n23846 ;
  assign n23847 = n23800 & n73196 ;
  assign n23848 = n23845 | n23847 ;
  assign n23849 = n139 & n23848 ;
  assign n23850 = n23023 & n73180 ;
  assign n23851 = n23687 & n23850 ;
  assign n23852 = n23849 | n23851 ;
  assign n23853 = n72025 & n23852 ;
  assign n73197 = ~n23799 ;
  assign n23854 = n23641 & n73197 ;
  assign n23855 = n23040 | n23641 ;
  assign n73198 = ~n23855 ;
  assign n23856 = n23637 & n73198 ;
  assign n23857 = n23854 | n23856 ;
  assign n23858 = n139 & n23857 ;
  assign n23859 = n23031 & n73180 ;
  assign n23860 = n23687 & n23859 ;
  assign n23861 = n23858 | n23860 ;
  assign n23862 = n71645 & n23861 ;
  assign n73199 = ~n23636 ;
  assign n23863 = n23635 & n73199 ;
  assign n23864 = n23048 | n23635 ;
  assign n73200 = ~n23864 ;
  assign n23865 = n23796 & n73200 ;
  assign n23866 = n23863 | n23865 ;
  assign n23867 = n139 & n23866 ;
  assign n23868 = n23039 & n73180 ;
  assign n23869 = n23687 & n23868 ;
  assign n23870 = n23867 | n23869 ;
  assign n23871 = n71633 & n23870 ;
  assign n73201 = ~n23795 ;
  assign n23872 = n23631 & n73201 ;
  assign n23873 = n23056 | n23631 ;
  assign n73202 = ~n23873 ;
  assign n23874 = n23627 & n73202 ;
  assign n23875 = n23872 | n23874 ;
  assign n23876 = n139 & n23875 ;
  assign n23877 = n23047 & n73180 ;
  assign n23878 = n23687 & n23877 ;
  assign n23879 = n23876 | n23878 ;
  assign n23880 = n71253 & n23879 ;
  assign n73203 = ~n23626 ;
  assign n23881 = n23624 & n73203 ;
  assign n23625 = n23064 | n23624 ;
  assign n73204 = ~n23625 ;
  assign n23882 = n23621 & n73204 ;
  assign n23883 = n23881 | n23882 ;
  assign n23884 = n139 & n23883 ;
  assign n23885 = n23055 & n73180 ;
  assign n23886 = n23687 & n23885 ;
  assign n23887 = n23884 | n23886 ;
  assign n23888 = n70935 & n23887 ;
  assign n73205 = ~n23791 ;
  assign n23889 = n23620 & n73205 ;
  assign n23890 = n23072 | n23620 ;
  assign n73206 = ~n23890 ;
  assign n23891 = n23616 & n73206 ;
  assign n23892 = n23889 | n23891 ;
  assign n23893 = n139 & n23892 ;
  assign n23894 = n23063 & n73180 ;
  assign n23895 = n23687 & n23894 ;
  assign n23896 = n23893 | n23895 ;
  assign n23897 = n70927 & n23896 ;
  assign n73207 = ~n23615 ;
  assign n23898 = n23614 & n73207 ;
  assign n23899 = n23080 | n23614 ;
  assign n73208 = ~n23899 ;
  assign n23900 = n23788 & n73208 ;
  assign n23901 = n23898 | n23900 ;
  assign n23902 = n139 & n23901 ;
  assign n23903 = n23071 & n73180 ;
  assign n23904 = n23687 & n23903 ;
  assign n23905 = n23902 | n23904 ;
  assign n23906 = n70609 & n23905 ;
  assign n73209 = ~n23787 ;
  assign n23907 = n23610 & n73209 ;
  assign n23908 = n23088 | n23610 ;
  assign n73210 = ~n23908 ;
  assign n23909 = n23606 & n73210 ;
  assign n23910 = n23907 | n23909 ;
  assign n23911 = n139 & n23910 ;
  assign n23912 = n23079 & n73180 ;
  assign n23913 = n23687 & n23912 ;
  assign n23914 = n23911 | n23913 ;
  assign n23915 = n70276 & n23914 ;
  assign n73211 = ~n23605 ;
  assign n23916 = n23603 & n73211 ;
  assign n23604 = n23096 | n23603 ;
  assign n73212 = ~n23604 ;
  assign n23917 = n23600 & n73212 ;
  assign n23918 = n23916 | n23917 ;
  assign n23919 = n139 & n23918 ;
  assign n23920 = n23087 & n73180 ;
  assign n23921 = n23687 & n23920 ;
  assign n23922 = n23919 | n23921 ;
  assign n23923 = n70176 & n23922 ;
  assign n73213 = ~n23783 ;
  assign n23924 = n23599 & n73213 ;
  assign n23925 = n23104 | n23599 ;
  assign n73214 = ~n23925 ;
  assign n23926 = n23595 & n73214 ;
  assign n23927 = n23924 | n23926 ;
  assign n23928 = n139 & n23927 ;
  assign n23929 = n23095 & n73180 ;
  assign n23930 = n23687 & n23929 ;
  assign n23931 = n23928 | n23930 ;
  assign n23932 = n69857 & n23931 ;
  assign n73215 = ~n23594 ;
  assign n23933 = n23593 & n73215 ;
  assign n23934 = n23112 | n23593 ;
  assign n73216 = ~n23934 ;
  assign n23935 = n23780 & n73216 ;
  assign n23936 = n23933 | n23935 ;
  assign n23937 = n139 & n23936 ;
  assign n23938 = n23103 & n73180 ;
  assign n23939 = n23687 & n23938 ;
  assign n23940 = n23937 | n23939 ;
  assign n23941 = n69656 & n23940 ;
  assign n73217 = ~n23779 ;
  assign n23942 = n23589 & n73217 ;
  assign n23943 = n23120 | n23589 ;
  assign n73218 = ~n23943 ;
  assign n23944 = n23585 & n73218 ;
  assign n23945 = n23942 | n23944 ;
  assign n23946 = n139 & n23945 ;
  assign n23947 = n23111 & n73180 ;
  assign n23948 = n23687 & n23947 ;
  assign n23949 = n23946 | n23948 ;
  assign n23950 = n69528 & n23949 ;
  assign n73219 = ~n23584 ;
  assign n23951 = n23583 & n73219 ;
  assign n23952 = n23128 | n23583 ;
  assign n73220 = ~n23952 ;
  assign n23953 = n23776 & n73220 ;
  assign n23954 = n23951 | n23953 ;
  assign n23955 = n139 & n23954 ;
  assign n23956 = n23119 & n73180 ;
  assign n23957 = n23687 & n23956 ;
  assign n23958 = n23955 | n23957 ;
  assign n23959 = n69261 & n23958 ;
  assign n73221 = ~n23775 ;
  assign n23960 = n23579 & n73221 ;
  assign n23961 = n23136 | n23579 ;
  assign n73222 = ~n23961 ;
  assign n23962 = n23575 & n73222 ;
  assign n23963 = n23960 | n23962 ;
  assign n23964 = n139 & n23963 ;
  assign n23965 = n23127 & n73180 ;
  assign n23966 = n23687 & n23965 ;
  assign n23967 = n23964 | n23966 ;
  assign n23968 = n69075 & n23967 ;
  assign n73223 = ~n23574 ;
  assign n23969 = n23573 & n73223 ;
  assign n23970 = n23144 | n23573 ;
  assign n73224 = ~n23970 ;
  assign n23971 = n23772 & n73224 ;
  assign n23972 = n23969 | n23971 ;
  assign n23973 = n139 & n23972 ;
  assign n23974 = n23135 & n73180 ;
  assign n23975 = n23687 & n23974 ;
  assign n23976 = n23973 | n23975 ;
  assign n23977 = n68993 & n23976 ;
  assign n73225 = ~n23771 ;
  assign n23978 = n23569 & n73225 ;
  assign n23979 = n23152 | n23569 ;
  assign n73226 = ~n23979 ;
  assign n23980 = n23565 & n73226 ;
  assign n23981 = n23978 | n23980 ;
  assign n23982 = n139 & n23981 ;
  assign n23983 = n23143 & n73180 ;
  assign n23984 = n23687 & n23983 ;
  assign n23985 = n23982 | n23984 ;
  assign n23986 = n68716 & n23985 ;
  assign n73227 = ~n23564 ;
  assign n23987 = n23563 & n73227 ;
  assign n23988 = n23160 | n23563 ;
  assign n73228 = ~n23988 ;
  assign n23989 = n23768 & n73228 ;
  assign n23990 = n23987 | n23989 ;
  assign n23991 = n139 & n23990 ;
  assign n23992 = n23151 & n73180 ;
  assign n23993 = n23687 & n23992 ;
  assign n23994 = n23991 | n23993 ;
  assign n23995 = n68545 & n23994 ;
  assign n73229 = ~n23767 ;
  assign n23996 = n23559 & n73229 ;
  assign n23997 = n23168 | n23559 ;
  assign n73230 = ~n23997 ;
  assign n23998 = n23555 & n73230 ;
  assign n23999 = n23996 | n23998 ;
  assign n24000 = n139 & n23999 ;
  assign n24001 = n23159 & n73180 ;
  assign n24002 = n23687 & n24001 ;
  assign n24003 = n24000 | n24002 ;
  assign n24004 = n68438 & n24003 ;
  assign n73231 = ~n23554 ;
  assign n24005 = n23553 & n73231 ;
  assign n24006 = n23176 | n23553 ;
  assign n73232 = ~n24006 ;
  assign n24007 = n23764 & n73232 ;
  assign n24008 = n24005 | n24007 ;
  assign n24009 = n139 & n24008 ;
  assign n24010 = n23167 & n73180 ;
  assign n24011 = n23687 & n24010 ;
  assign n24012 = n24009 | n24011 ;
  assign n24013 = n68214 & n24012 ;
  assign n73233 = ~n23763 ;
  assign n24014 = n23549 & n73233 ;
  assign n24015 = n23184 | n23549 ;
  assign n73234 = ~n24015 ;
  assign n24016 = n23545 & n73234 ;
  assign n24017 = n24014 | n24016 ;
  assign n24018 = n139 & n24017 ;
  assign n24019 = n23175 & n73180 ;
  assign n24020 = n23687 & n24019 ;
  assign n24021 = n24018 | n24020 ;
  assign n24022 = n68058 & n24021 ;
  assign n73235 = ~n23544 ;
  assign n24023 = n23543 & n73235 ;
  assign n24024 = n23192 | n23543 ;
  assign n73236 = ~n24024 ;
  assign n24025 = n23760 & n73236 ;
  assign n24026 = n24023 | n24025 ;
  assign n24027 = n139 & n24026 ;
  assign n24028 = n23183 & n73180 ;
  assign n24029 = n23687 & n24028 ;
  assign n24030 = n24027 | n24029 ;
  assign n24031 = n67986 & n24030 ;
  assign n73237 = ~n23759 ;
  assign n24032 = n23539 & n73237 ;
  assign n24033 = n23200 | n23539 ;
  assign n73238 = ~n24033 ;
  assign n24034 = n23535 & n73238 ;
  assign n24035 = n24032 | n24034 ;
  assign n24036 = n139 & n24035 ;
  assign n24037 = n23191 & n73180 ;
  assign n24038 = n23687 & n24037 ;
  assign n24039 = n24036 | n24038 ;
  assign n24040 = n67763 & n24039 ;
  assign n73239 = ~n23534 ;
  assign n24041 = n23533 & n73239 ;
  assign n24042 = n23208 | n23533 ;
  assign n73240 = ~n24042 ;
  assign n24043 = n23756 & n73240 ;
  assign n24044 = n24041 | n24043 ;
  assign n24045 = n139 & n24044 ;
  assign n24046 = n23199 & n73180 ;
  assign n24047 = n23687 & n24046 ;
  assign n24048 = n24045 | n24047 ;
  assign n24049 = n67622 & n24048 ;
  assign n73241 = ~n23755 ;
  assign n24050 = n23529 & n73241 ;
  assign n24051 = n23216 | n23529 ;
  assign n73242 = ~n24051 ;
  assign n24052 = n23525 & n73242 ;
  assign n24053 = n24050 | n24052 ;
  assign n24054 = n139 & n24053 ;
  assign n24055 = n23207 & n73180 ;
  assign n24056 = n23687 & n24055 ;
  assign n24057 = n24054 | n24056 ;
  assign n24058 = n67531 & n24057 ;
  assign n73243 = ~n23524 ;
  assign n24059 = n23522 & n73243 ;
  assign n23523 = n23224 | n23522 ;
  assign n73244 = ~n23523 ;
  assign n24060 = n23519 & n73244 ;
  assign n24061 = n24059 | n24060 ;
  assign n24062 = n139 & n24061 ;
  assign n24063 = n23215 & n73180 ;
  assign n24064 = n23687 & n24063 ;
  assign n24065 = n24062 | n24064 ;
  assign n24066 = n67348 & n24065 ;
  assign n73245 = ~n23751 ;
  assign n24067 = n23518 & n73245 ;
  assign n24068 = n23232 | n23518 ;
  assign n73246 = ~n24068 ;
  assign n24069 = n23514 & n73246 ;
  assign n24070 = n24067 | n24069 ;
  assign n24071 = n139 & n24070 ;
  assign n24072 = n23223 & n73180 ;
  assign n24073 = n23687 & n24072 ;
  assign n24074 = n24071 | n24073 ;
  assign n24075 = n67222 & n24074 ;
  assign n73247 = ~n23513 ;
  assign n24076 = n23512 & n73247 ;
  assign n24077 = n23240 | n23512 ;
  assign n73248 = ~n24077 ;
  assign n24078 = n23748 & n73248 ;
  assign n24079 = n24076 | n24078 ;
  assign n24080 = n139 & n24079 ;
  assign n24081 = n23231 & n73180 ;
  assign n24082 = n23687 & n24081 ;
  assign n24083 = n24080 | n24082 ;
  assign n24084 = n67164 & n24083 ;
  assign n73249 = ~n23747 ;
  assign n24085 = n23507 & n73249 ;
  assign n23508 = n23248 | n23507 ;
  assign n73250 = ~n23508 ;
  assign n24086 = n73250 & n23746 ;
  assign n24087 = n24085 | n24086 ;
  assign n24088 = n139 & n24087 ;
  assign n24089 = n23239 & n73180 ;
  assign n24090 = n23687 & n24089 ;
  assign n24091 = n24088 | n24090 ;
  assign n24092 = n66979 & n24091 ;
  assign n73251 = ~n23502 ;
  assign n24093 = n23500 & n73251 ;
  assign n23501 = n23256 | n23500 ;
  assign n73252 = ~n23501 ;
  assign n24094 = n23497 & n73252 ;
  assign n24095 = n24093 | n24094 ;
  assign n24096 = n139 & n24095 ;
  assign n24097 = n23247 & n73180 ;
  assign n24098 = n23687 & n24097 ;
  assign n24099 = n24096 | n24098 ;
  assign n24100 = n66868 & n24099 ;
  assign n73253 = ~n23743 ;
  assign n24101 = n23496 & n73253 ;
  assign n24102 = n23264 | n23496 ;
  assign n73254 = ~n24102 ;
  assign n24103 = n23492 & n73254 ;
  assign n24104 = n24101 | n24103 ;
  assign n24105 = n139 & n24104 ;
  assign n24106 = n23255 & n73180 ;
  assign n24107 = n23687 & n24106 ;
  assign n24108 = n24105 | n24107 ;
  assign n24109 = n66797 & n24108 ;
  assign n73255 = ~n23491 ;
  assign n24110 = n23490 & n73255 ;
  assign n24111 = n23272 | n23490 ;
  assign n73256 = ~n24111 ;
  assign n24112 = n23740 & n73256 ;
  assign n24113 = n24110 | n24112 ;
  assign n24114 = n139 & n24113 ;
  assign n24115 = n23263 & n73180 ;
  assign n24116 = n23687 & n24115 ;
  assign n24117 = n24114 | n24116 ;
  assign n24118 = n66654 & n24117 ;
  assign n73257 = ~n23739 ;
  assign n24119 = n23486 & n73257 ;
  assign n24120 = n23280 | n23486 ;
  assign n73258 = ~n24120 ;
  assign n24121 = n23482 & n73258 ;
  assign n24122 = n24119 | n24121 ;
  assign n24123 = n139 & n24122 ;
  assign n24124 = n23271 & n73180 ;
  assign n24125 = n23687 & n24124 ;
  assign n24126 = n24123 | n24125 ;
  assign n24127 = n66560 & n24126 ;
  assign n73259 = ~n23481 ;
  assign n24128 = n23479 & n73259 ;
  assign n23480 = n23288 | n23479 ;
  assign n73260 = ~n23480 ;
  assign n24129 = n23476 & n73260 ;
  assign n24130 = n24128 | n24129 ;
  assign n24131 = n139 & n24130 ;
  assign n24132 = n23279 & n73180 ;
  assign n24133 = n23687 & n24132 ;
  assign n24134 = n24131 | n24133 ;
  assign n24135 = n66505 & n24134 ;
  assign n73261 = ~n23735 ;
  assign n24136 = n23474 & n73261 ;
  assign n23475 = n23296 | n23474 ;
  assign n73262 = ~n23475 ;
  assign n24137 = n73262 & n23734 ;
  assign n24138 = n24136 | n24137 ;
  assign n24139 = n139 & n24138 ;
  assign n24140 = n23287 & n73180 ;
  assign n24141 = n23687 & n24140 ;
  assign n24142 = n24139 | n24141 ;
  assign n24143 = n66379 & n24142 ;
  assign n73263 = ~n23469 ;
  assign n24144 = n23468 & n73263 ;
  assign n24145 = n23304 | n23468 ;
  assign n73264 = ~n24145 ;
  assign n24146 = n23732 & n73264 ;
  assign n24147 = n24144 | n24146 ;
  assign n24148 = n139 & n24147 ;
  assign n24149 = n23295 & n73180 ;
  assign n24150 = n23687 & n24149 ;
  assign n24151 = n24148 | n24150 ;
  assign n24152 = n66299 & n24151 ;
  assign n73265 = ~n23731 ;
  assign n24153 = n23464 & n73265 ;
  assign n24154 = n23312 | n23464 ;
  assign n73266 = ~n24154 ;
  assign n24155 = n23460 & n73266 ;
  assign n24156 = n24153 | n24155 ;
  assign n24157 = n139 & n24156 ;
  assign n24158 = n23303 & n73180 ;
  assign n24159 = n23687 & n24158 ;
  assign n24160 = n24157 | n24159 ;
  assign n24161 = n66244 & n24160 ;
  assign n73267 = ~n23459 ;
  assign n24162 = n23458 & n73267 ;
  assign n24163 = n23320 | n23458 ;
  assign n73268 = ~n24163 ;
  assign n24164 = n23728 & n73268 ;
  assign n24165 = n24162 | n24164 ;
  assign n24166 = n139 & n24165 ;
  assign n24167 = n23311 & n73180 ;
  assign n24168 = n23687 & n24167 ;
  assign n24169 = n24166 | n24168 ;
  assign n24170 = n66145 & n24169 ;
  assign n73269 = ~n23727 ;
  assign n24171 = n23454 & n73269 ;
  assign n24172 = n23328 | n23454 ;
  assign n73270 = ~n24172 ;
  assign n24173 = n23450 & n73270 ;
  assign n24174 = n24171 | n24173 ;
  assign n24175 = n139 & n24174 ;
  assign n24176 = n23319 & n73180 ;
  assign n24177 = n23687 & n24176 ;
  assign n24178 = n24175 | n24177 ;
  assign n24179 = n66081 & n24178 ;
  assign n73271 = ~n23449 ;
  assign n24180 = n23448 & n73271 ;
  assign n24181 = n23336 | n23448 ;
  assign n73272 = ~n24181 ;
  assign n24182 = n23724 & n73272 ;
  assign n24183 = n24180 | n24182 ;
  assign n24184 = n139 & n24183 ;
  assign n24185 = n23327 & n73180 ;
  assign n24186 = n23687 & n24185 ;
  assign n24187 = n24184 | n24186 ;
  assign n24188 = n66043 & n24187 ;
  assign n73273 = ~n23723 ;
  assign n24189 = n23443 & n73273 ;
  assign n23444 = n23344 | n23443 ;
  assign n73274 = ~n23444 ;
  assign n24190 = n73274 & n23722 ;
  assign n24191 = n24189 | n24190 ;
  assign n24192 = n139 & n24191 ;
  assign n24193 = n23335 & n73180 ;
  assign n24194 = n23687 & n24193 ;
  assign n24195 = n24192 | n24194 ;
  assign n24196 = n65960 & n24195 ;
  assign n73275 = ~n23438 ;
  assign n24197 = n23437 & n73275 ;
  assign n24198 = n23352 | n23437 ;
  assign n73276 = ~n24198 ;
  assign n24199 = n23720 & n73276 ;
  assign n24200 = n24197 | n24199 ;
  assign n24201 = n139 & n24200 ;
  assign n24202 = n23343 & n73180 ;
  assign n24203 = n23687 & n24202 ;
  assign n24204 = n24201 | n24203 ;
  assign n24205 = n65909 & n24204 ;
  assign n73277 = ~n23719 ;
  assign n24206 = n23433 & n73277 ;
  assign n24207 = n23360 | n23433 ;
  assign n73278 = ~n24207 ;
  assign n24208 = n23429 & n73278 ;
  assign n24209 = n24206 | n24208 ;
  assign n24210 = n139 & n24209 ;
  assign n24211 = n23351 & n73180 ;
  assign n24212 = n23687 & n24211 ;
  assign n24213 = n24210 | n24212 ;
  assign n24214 = n65877 & n24213 ;
  assign n73279 = ~n23428 ;
  assign n24215 = n23427 & n73279 ;
  assign n24216 = n23369 | n23427 ;
  assign n73280 = ~n24216 ;
  assign n24217 = n23716 & n73280 ;
  assign n24218 = n24215 | n24217 ;
  assign n24219 = n139 & n24218 ;
  assign n24220 = n23359 & n73180 ;
  assign n24221 = n23687 & n24220 ;
  assign n24222 = n24219 | n24221 ;
  assign n24223 = n65820 & n24222 ;
  assign n73281 = ~n23715 ;
  assign n24224 = n23423 & n73281 ;
  assign n24225 = n23377 | n23423 ;
  assign n73282 = ~n24225 ;
  assign n24226 = n23419 & n73282 ;
  assign n24227 = n24224 | n24226 ;
  assign n24228 = n139 & n24227 ;
  assign n24229 = n23368 & n73180 ;
  assign n24230 = n23687 & n24229 ;
  assign n24231 = n24228 | n24230 ;
  assign n24232 = n65791 & n24231 ;
  assign n73283 = ~n23418 ;
  assign n24234 = n23417 & n73283 ;
  assign n24233 = n23385 | n23417 ;
  assign n73284 = ~n24233 ;
  assign n24235 = n23414 & n73284 ;
  assign n24236 = n24234 | n24235 ;
  assign n24237 = n139 & n24236 ;
  assign n24238 = n23376 & n73180 ;
  assign n24239 = n23687 & n24238 ;
  assign n24240 = n24237 | n24239 ;
  assign n24241 = n65772 & n24240 ;
  assign n73285 = ~n23711 ;
  assign n24242 = n23413 & n73285 ;
  assign n24243 = n23393 | n23413 ;
  assign n73286 = ~n24243 ;
  assign n24244 = n23409 & n73286 ;
  assign n24245 = n24242 | n24244 ;
  assign n24246 = n139 & n24245 ;
  assign n24247 = n23384 & n73180 ;
  assign n24248 = n23687 & n24247 ;
  assign n24249 = n24246 | n24248 ;
  assign n24250 = n65746 & n24249 ;
  assign n73287 = ~n23408 ;
  assign n24251 = n23407 & n73287 ;
  assign n23709 = n23404 | n23407 ;
  assign n73288 = ~n23709 ;
  assign n24252 = n23403 & n73288 ;
  assign n24253 = n24251 | n24252 ;
  assign n24254 = n139 & n24253 ;
  assign n24255 = n23392 & n73180 ;
  assign n24256 = n23687 & n24255 ;
  assign n24257 = n24254 | n24256 ;
  assign n24258 = n65721 & n24257 ;
  assign n24259 = n23400 & n23402 ;
  assign n24260 = n73071 & n24259 ;
  assign n73289 = ~n24260 ;
  assign n24261 = n23403 & n73289 ;
  assign n24262 = n139 & n24261 ;
  assign n24263 = n23395 & n73180 ;
  assign n24264 = n23687 & n24263 ;
  assign n24265 = n24262 | n24264 ;
  assign n24266 = n65686 & n24265 ;
  assign n23690 = n23402 & n139 ;
  assign n24267 = x64 & n139 ;
  assign n73290 = ~n24267 ;
  assign n24268 = x10 & n73290 ;
  assign n24269 = n23690 | n24268 ;
  assign n24282 = n65670 & n24269 ;
  assign n23809 = n73173 & n23808 ;
  assign n24270 = n23666 | n23809 ;
  assign n24271 = n73174 & n24270 ;
  assign n24272 = n23686 | n24271 ;
  assign n24273 = n73180 & n24272 ;
  assign n73291 = ~n24273 ;
  assign n24274 = x64 & n73291 ;
  assign n73292 = ~n24274 ;
  assign n24275 = x10 & n73292 ;
  assign n24276 = n23690 | n24275 ;
  assign n24277 = x65 & n24276 ;
  assign n24278 = x65 | n23690 ;
  assign n24279 = n24275 | n24278 ;
  assign n73293 = ~n24277 ;
  assign n24280 = n73293 & n24279 ;
  assign n73294 = ~x9 ;
  assign n24281 = n73294 & x64 ;
  assign n24283 = n24280 | n24281 ;
  assign n73295 = ~n24282 ;
  assign n24284 = n73295 & n24283 ;
  assign n73296 = ~n24264 ;
  assign n24285 = x66 & n73296 ;
  assign n73297 = ~n24262 ;
  assign n24286 = n73297 & n24285 ;
  assign n24287 = n24266 | n24286 ;
  assign n24288 = n24284 | n24287 ;
  assign n73298 = ~n24266 ;
  assign n24289 = n73298 & n24288 ;
  assign n73299 = ~n24256 ;
  assign n24290 = x67 & n73299 ;
  assign n73300 = ~n24254 ;
  assign n24291 = n73300 & n24290 ;
  assign n24292 = n24258 | n24291 ;
  assign n24293 = n24289 | n24292 ;
  assign n73301 = ~n24258 ;
  assign n24294 = n73301 & n24293 ;
  assign n73302 = ~n24248 ;
  assign n24295 = x68 & n73302 ;
  assign n73303 = ~n24246 ;
  assign n24296 = n73303 & n24295 ;
  assign n24297 = n24294 | n24296 ;
  assign n73304 = ~n24250 ;
  assign n24298 = n73304 & n24297 ;
  assign n73305 = ~n24239 ;
  assign n24299 = x69 & n73305 ;
  assign n73306 = ~n24237 ;
  assign n24300 = n73306 & n24299 ;
  assign n24301 = n24241 | n24300 ;
  assign n24302 = n24298 | n24301 ;
  assign n73307 = ~n24241 ;
  assign n24303 = n73307 & n24302 ;
  assign n73308 = ~n24230 ;
  assign n24304 = x70 & n73308 ;
  assign n73309 = ~n24228 ;
  assign n24305 = n73309 & n24304 ;
  assign n24306 = n24232 | n24305 ;
  assign n24308 = n24303 | n24306 ;
  assign n73310 = ~n24232 ;
  assign n24310 = n73310 & n24308 ;
  assign n73311 = ~n24221 ;
  assign n24311 = x71 & n73311 ;
  assign n73312 = ~n24219 ;
  assign n24312 = n73312 & n24311 ;
  assign n24313 = n24223 | n24312 ;
  assign n24314 = n24310 | n24313 ;
  assign n73313 = ~n24223 ;
  assign n24315 = n73313 & n24314 ;
  assign n73314 = ~n24212 ;
  assign n24316 = x72 & n73314 ;
  assign n73315 = ~n24210 ;
  assign n24317 = n73315 & n24316 ;
  assign n24318 = n24214 | n24317 ;
  assign n24320 = n24315 | n24318 ;
  assign n73316 = ~n24214 ;
  assign n24321 = n73316 & n24320 ;
  assign n73317 = ~n24203 ;
  assign n24322 = x73 & n73317 ;
  assign n73318 = ~n24201 ;
  assign n24323 = n73318 & n24322 ;
  assign n24324 = n24205 | n24323 ;
  assign n24325 = n24321 | n24324 ;
  assign n73319 = ~n24205 ;
  assign n24326 = n73319 & n24325 ;
  assign n73320 = ~n24194 ;
  assign n24327 = x74 & n73320 ;
  assign n73321 = ~n24192 ;
  assign n24328 = n73321 & n24327 ;
  assign n24329 = n24196 | n24328 ;
  assign n24331 = n24326 | n24329 ;
  assign n73322 = ~n24196 ;
  assign n24332 = n73322 & n24331 ;
  assign n73323 = ~n24186 ;
  assign n24333 = x75 & n73323 ;
  assign n73324 = ~n24184 ;
  assign n24334 = n73324 & n24333 ;
  assign n24335 = n24188 | n24334 ;
  assign n24336 = n24332 | n24335 ;
  assign n73325 = ~n24188 ;
  assign n24337 = n73325 & n24336 ;
  assign n73326 = ~n24177 ;
  assign n24338 = x76 & n73326 ;
  assign n73327 = ~n24175 ;
  assign n24339 = n73327 & n24338 ;
  assign n24340 = n24179 | n24339 ;
  assign n24342 = n24337 | n24340 ;
  assign n73328 = ~n24179 ;
  assign n24343 = n73328 & n24342 ;
  assign n73329 = ~n24168 ;
  assign n24344 = x77 & n73329 ;
  assign n73330 = ~n24166 ;
  assign n24345 = n73330 & n24344 ;
  assign n24346 = n24170 | n24345 ;
  assign n24347 = n24343 | n24346 ;
  assign n73331 = ~n24170 ;
  assign n24348 = n73331 & n24347 ;
  assign n73332 = ~n24159 ;
  assign n24349 = x78 & n73332 ;
  assign n73333 = ~n24157 ;
  assign n24350 = n73333 & n24349 ;
  assign n24351 = n24161 | n24350 ;
  assign n24353 = n24348 | n24351 ;
  assign n73334 = ~n24161 ;
  assign n24354 = n73334 & n24353 ;
  assign n73335 = ~n24150 ;
  assign n24355 = x79 & n73335 ;
  assign n73336 = ~n24148 ;
  assign n24356 = n73336 & n24355 ;
  assign n24357 = n24152 | n24356 ;
  assign n24358 = n24354 | n24357 ;
  assign n73337 = ~n24152 ;
  assign n24359 = n73337 & n24358 ;
  assign n73338 = ~n24141 ;
  assign n24360 = x80 & n73338 ;
  assign n73339 = ~n24139 ;
  assign n24361 = n73339 & n24360 ;
  assign n24362 = n24143 | n24361 ;
  assign n24364 = n24359 | n24362 ;
  assign n73340 = ~n24143 ;
  assign n24365 = n73340 & n24364 ;
  assign n73341 = ~n24133 ;
  assign n24366 = x81 & n73341 ;
  assign n73342 = ~n24131 ;
  assign n24367 = n73342 & n24366 ;
  assign n24368 = n24135 | n24367 ;
  assign n24369 = n24365 | n24368 ;
  assign n73343 = ~n24135 ;
  assign n24370 = n73343 & n24369 ;
  assign n73344 = ~n24125 ;
  assign n24371 = x82 & n73344 ;
  assign n73345 = ~n24123 ;
  assign n24372 = n73345 & n24371 ;
  assign n24373 = n24127 | n24372 ;
  assign n24375 = n24370 | n24373 ;
  assign n73346 = ~n24127 ;
  assign n24376 = n73346 & n24375 ;
  assign n73347 = ~n24116 ;
  assign n24377 = x83 & n73347 ;
  assign n73348 = ~n24114 ;
  assign n24378 = n73348 & n24377 ;
  assign n24379 = n24118 | n24378 ;
  assign n24380 = n24376 | n24379 ;
  assign n73349 = ~n24118 ;
  assign n24381 = n73349 & n24380 ;
  assign n73350 = ~n24107 ;
  assign n24382 = x84 & n73350 ;
  assign n73351 = ~n24105 ;
  assign n24383 = n73351 & n24382 ;
  assign n24384 = n24109 | n24383 ;
  assign n24386 = n24381 | n24384 ;
  assign n73352 = ~n24109 ;
  assign n24387 = n73352 & n24386 ;
  assign n73353 = ~n24098 ;
  assign n24388 = x85 & n73353 ;
  assign n73354 = ~n24096 ;
  assign n24389 = n73354 & n24388 ;
  assign n24390 = n24100 | n24389 ;
  assign n24391 = n24387 | n24390 ;
  assign n73355 = ~n24100 ;
  assign n24392 = n73355 & n24391 ;
  assign n73356 = ~n24090 ;
  assign n24393 = x86 & n73356 ;
  assign n73357 = ~n24088 ;
  assign n24394 = n73357 & n24393 ;
  assign n24395 = n24092 | n24394 ;
  assign n24397 = n24392 | n24395 ;
  assign n73358 = ~n24092 ;
  assign n24398 = n73358 & n24397 ;
  assign n73359 = ~n24082 ;
  assign n24399 = x87 & n73359 ;
  assign n73360 = ~n24080 ;
  assign n24400 = n73360 & n24399 ;
  assign n24401 = n24084 | n24400 ;
  assign n24402 = n24398 | n24401 ;
  assign n73361 = ~n24084 ;
  assign n24403 = n73361 & n24402 ;
  assign n73362 = ~n24073 ;
  assign n24404 = x88 & n73362 ;
  assign n73363 = ~n24071 ;
  assign n24405 = n73363 & n24404 ;
  assign n24406 = n24075 | n24405 ;
  assign n24408 = n24403 | n24406 ;
  assign n73364 = ~n24075 ;
  assign n24409 = n73364 & n24408 ;
  assign n73365 = ~n24064 ;
  assign n24410 = x89 & n73365 ;
  assign n73366 = ~n24062 ;
  assign n24411 = n73366 & n24410 ;
  assign n24412 = n24066 | n24411 ;
  assign n24413 = n24409 | n24412 ;
  assign n73367 = ~n24066 ;
  assign n24414 = n73367 & n24413 ;
  assign n73368 = ~n24056 ;
  assign n24415 = x90 & n73368 ;
  assign n73369 = ~n24054 ;
  assign n24416 = n73369 & n24415 ;
  assign n24417 = n24058 | n24416 ;
  assign n24419 = n24414 | n24417 ;
  assign n73370 = ~n24058 ;
  assign n24420 = n73370 & n24419 ;
  assign n73371 = ~n24047 ;
  assign n24421 = x91 & n73371 ;
  assign n73372 = ~n24045 ;
  assign n24422 = n73372 & n24421 ;
  assign n24423 = n24049 | n24422 ;
  assign n24424 = n24420 | n24423 ;
  assign n73373 = ~n24049 ;
  assign n24425 = n73373 & n24424 ;
  assign n73374 = ~n24038 ;
  assign n24426 = x92 & n73374 ;
  assign n73375 = ~n24036 ;
  assign n24427 = n73375 & n24426 ;
  assign n24428 = n24040 | n24427 ;
  assign n24430 = n24425 | n24428 ;
  assign n73376 = ~n24040 ;
  assign n24431 = n73376 & n24430 ;
  assign n73377 = ~n24029 ;
  assign n24432 = x93 & n73377 ;
  assign n73378 = ~n24027 ;
  assign n24433 = n73378 & n24432 ;
  assign n24434 = n24031 | n24433 ;
  assign n24435 = n24431 | n24434 ;
  assign n73379 = ~n24031 ;
  assign n24436 = n73379 & n24435 ;
  assign n73380 = ~n24020 ;
  assign n24437 = x94 & n73380 ;
  assign n73381 = ~n24018 ;
  assign n24438 = n73381 & n24437 ;
  assign n24439 = n24022 | n24438 ;
  assign n24441 = n24436 | n24439 ;
  assign n73382 = ~n24022 ;
  assign n24442 = n73382 & n24441 ;
  assign n73383 = ~n24011 ;
  assign n24443 = x95 & n73383 ;
  assign n73384 = ~n24009 ;
  assign n24444 = n73384 & n24443 ;
  assign n24445 = n24013 | n24444 ;
  assign n24446 = n24442 | n24445 ;
  assign n73385 = ~n24013 ;
  assign n24447 = n73385 & n24446 ;
  assign n73386 = ~n24002 ;
  assign n24448 = x96 & n73386 ;
  assign n73387 = ~n24000 ;
  assign n24449 = n73387 & n24448 ;
  assign n24450 = n24004 | n24449 ;
  assign n24452 = n24447 | n24450 ;
  assign n73388 = ~n24004 ;
  assign n24453 = n73388 & n24452 ;
  assign n73389 = ~n23993 ;
  assign n24454 = x97 & n73389 ;
  assign n73390 = ~n23991 ;
  assign n24455 = n73390 & n24454 ;
  assign n24456 = n23995 | n24455 ;
  assign n24457 = n24453 | n24456 ;
  assign n73391 = ~n23995 ;
  assign n24458 = n73391 & n24457 ;
  assign n73392 = ~n23984 ;
  assign n24459 = x98 & n73392 ;
  assign n73393 = ~n23982 ;
  assign n24460 = n73393 & n24459 ;
  assign n24461 = n23986 | n24460 ;
  assign n24463 = n24458 | n24461 ;
  assign n73394 = ~n23986 ;
  assign n24464 = n73394 & n24463 ;
  assign n73395 = ~n23975 ;
  assign n24465 = x99 & n73395 ;
  assign n73396 = ~n23973 ;
  assign n24466 = n73396 & n24465 ;
  assign n24467 = n23977 | n24466 ;
  assign n24468 = n24464 | n24467 ;
  assign n73397 = ~n23977 ;
  assign n24469 = n73397 & n24468 ;
  assign n73398 = ~n23966 ;
  assign n24470 = x100 & n73398 ;
  assign n73399 = ~n23964 ;
  assign n24471 = n73399 & n24470 ;
  assign n24472 = n23968 | n24471 ;
  assign n24474 = n24469 | n24472 ;
  assign n73400 = ~n23968 ;
  assign n24475 = n73400 & n24474 ;
  assign n73401 = ~n23957 ;
  assign n24476 = x101 & n73401 ;
  assign n73402 = ~n23955 ;
  assign n24477 = n73402 & n24476 ;
  assign n24478 = n23959 | n24477 ;
  assign n24479 = n24475 | n24478 ;
  assign n73403 = ~n23959 ;
  assign n24480 = n73403 & n24479 ;
  assign n73404 = ~n23948 ;
  assign n24481 = x102 & n73404 ;
  assign n73405 = ~n23946 ;
  assign n24482 = n73405 & n24481 ;
  assign n24483 = n23950 | n24482 ;
  assign n24485 = n24480 | n24483 ;
  assign n73406 = ~n23950 ;
  assign n24486 = n73406 & n24485 ;
  assign n73407 = ~n23939 ;
  assign n24487 = x103 & n73407 ;
  assign n73408 = ~n23937 ;
  assign n24488 = n73408 & n24487 ;
  assign n24489 = n23941 | n24488 ;
  assign n24490 = n24486 | n24489 ;
  assign n73409 = ~n23941 ;
  assign n24491 = n73409 & n24490 ;
  assign n73410 = ~n23930 ;
  assign n24492 = x104 & n73410 ;
  assign n73411 = ~n23928 ;
  assign n24493 = n73411 & n24492 ;
  assign n24494 = n23932 | n24493 ;
  assign n24496 = n24491 | n24494 ;
  assign n73412 = ~n23932 ;
  assign n24497 = n73412 & n24496 ;
  assign n73413 = ~n23921 ;
  assign n24498 = x105 & n73413 ;
  assign n73414 = ~n23919 ;
  assign n24499 = n73414 & n24498 ;
  assign n24500 = n23923 | n24499 ;
  assign n24501 = n24497 | n24500 ;
  assign n73415 = ~n23923 ;
  assign n24502 = n73415 & n24501 ;
  assign n73416 = ~n23913 ;
  assign n24503 = x106 & n73416 ;
  assign n73417 = ~n23911 ;
  assign n24504 = n73417 & n24503 ;
  assign n24505 = n23915 | n24504 ;
  assign n24507 = n24502 | n24505 ;
  assign n73418 = ~n23915 ;
  assign n24508 = n73418 & n24507 ;
  assign n73419 = ~n23904 ;
  assign n24509 = x107 & n73419 ;
  assign n73420 = ~n23902 ;
  assign n24510 = n73420 & n24509 ;
  assign n24511 = n23906 | n24510 ;
  assign n24512 = n24508 | n24511 ;
  assign n73421 = ~n23906 ;
  assign n24513 = n73421 & n24512 ;
  assign n73422 = ~n23895 ;
  assign n24514 = x108 & n73422 ;
  assign n73423 = ~n23893 ;
  assign n24515 = n73423 & n24514 ;
  assign n24516 = n23897 | n24515 ;
  assign n24518 = n24513 | n24516 ;
  assign n73424 = ~n23897 ;
  assign n24519 = n73424 & n24518 ;
  assign n73425 = ~n23886 ;
  assign n24520 = x109 & n73425 ;
  assign n73426 = ~n23884 ;
  assign n24521 = n73426 & n24520 ;
  assign n24522 = n23888 | n24521 ;
  assign n24523 = n24519 | n24522 ;
  assign n73427 = ~n23888 ;
  assign n24524 = n73427 & n24523 ;
  assign n73428 = ~n23878 ;
  assign n24525 = x110 & n73428 ;
  assign n73429 = ~n23876 ;
  assign n24526 = n73429 & n24525 ;
  assign n24527 = n23880 | n24526 ;
  assign n24529 = n24524 | n24527 ;
  assign n73430 = ~n23880 ;
  assign n24530 = n73430 & n24529 ;
  assign n73431 = ~n23869 ;
  assign n24531 = x111 & n73431 ;
  assign n73432 = ~n23867 ;
  assign n24532 = n73432 & n24531 ;
  assign n24533 = n23871 | n24532 ;
  assign n24534 = n24530 | n24533 ;
  assign n73433 = ~n23871 ;
  assign n24535 = n73433 & n24534 ;
  assign n73434 = ~n23860 ;
  assign n24536 = x112 & n73434 ;
  assign n73435 = ~n23858 ;
  assign n24537 = n73435 & n24536 ;
  assign n24538 = n23862 | n24537 ;
  assign n24540 = n24535 | n24538 ;
  assign n73436 = ~n23862 ;
  assign n24541 = n73436 & n24540 ;
  assign n73437 = ~n23851 ;
  assign n24542 = x113 & n73437 ;
  assign n73438 = ~n23849 ;
  assign n24543 = n73438 & n24542 ;
  assign n24544 = n23853 | n24543 ;
  assign n24545 = n24541 | n24544 ;
  assign n73439 = ~n23853 ;
  assign n24546 = n73439 & n24545 ;
  assign n73440 = ~n23842 ;
  assign n24547 = x114 & n73440 ;
  assign n73441 = ~n23840 ;
  assign n24548 = n73441 & n24547 ;
  assign n24549 = n23844 | n24548 ;
  assign n24551 = n24546 | n24549 ;
  assign n73442 = ~n23844 ;
  assign n24552 = n73442 & n24551 ;
  assign n73443 = ~n23834 ;
  assign n24553 = x115 & n73443 ;
  assign n73444 = ~n23832 ;
  assign n24554 = n73444 & n24553 ;
  assign n24555 = n23836 | n24554 ;
  assign n24556 = n24552 | n24555 ;
  assign n73445 = ~n23836 ;
  assign n24557 = n73445 & n24556 ;
  assign n73446 = ~n23825 ;
  assign n24558 = x116 & n73446 ;
  assign n73447 = ~n23823 ;
  assign n24559 = n73447 & n24558 ;
  assign n24560 = n23827 | n24559 ;
  assign n24562 = n24557 | n24560 ;
  assign n73448 = ~n23827 ;
  assign n24563 = n73448 & n24562 ;
  assign n73449 = ~n23816 ;
  assign n24564 = x117 & n73449 ;
  assign n73450 = ~n23814 ;
  assign n24565 = n73450 & n24564 ;
  assign n24566 = n23818 | n24565 ;
  assign n24567 = n24563 | n24566 ;
  assign n73451 = ~n23818 ;
  assign n24568 = n73451 & n24567 ;
  assign n73452 = ~n23699 ;
  assign n24569 = x118 & n73452 ;
  assign n73453 = ~n23697 ;
  assign n24570 = n73453 & n24569 ;
  assign n24571 = n23701 | n24570 ;
  assign n24573 = n24568 | n24571 ;
  assign n73454 = ~n23701 ;
  assign n24574 = n73454 & n24573 ;
  assign n24575 = n267 | n277 ;
  assign n24576 = n274 | n24575 ;
  assign n24577 = n24574 | n24576 ;
  assign n24578 = n23817 & n24577 ;
  assign n24579 = x65 & n24269 ;
  assign n73455 = ~n24579 ;
  assign n24580 = n24279 & n73455 ;
  assign n24581 = n24281 | n24580 ;
  assign n24582 = n73295 & n24581 ;
  assign n24583 = n24287 | n24582 ;
  assign n24584 = n73298 & n24583 ;
  assign n24585 = n24291 | n24584 ;
  assign n24587 = n73301 & n24585 ;
  assign n24588 = n24250 | n24296 ;
  assign n24590 = n24587 | n24588 ;
  assign n24591 = n73304 & n24590 ;
  assign n24592 = n24300 | n24591 ;
  assign n24594 = n73307 & n24592 ;
  assign n24595 = n24306 | n24594 ;
  assign n24596 = n73310 & n24595 ;
  assign n24597 = n24313 | n24596 ;
  assign n24599 = n73313 & n24597 ;
  assign n24600 = n24318 | n24599 ;
  assign n24601 = n73316 & n24600 ;
  assign n24602 = n24324 | n24601 ;
  assign n24604 = n73319 & n24602 ;
  assign n24605 = n24329 | n24604 ;
  assign n24606 = n73322 & n24605 ;
  assign n24607 = n24335 | n24606 ;
  assign n24609 = n73325 & n24607 ;
  assign n24610 = n24340 | n24609 ;
  assign n24611 = n73328 & n24610 ;
  assign n24612 = n24346 | n24611 ;
  assign n24614 = n73331 & n24612 ;
  assign n24615 = n24351 | n24614 ;
  assign n24616 = n73334 & n24615 ;
  assign n24617 = n24357 | n24616 ;
  assign n24619 = n73337 & n24617 ;
  assign n24620 = n24362 | n24619 ;
  assign n24621 = n73340 & n24620 ;
  assign n24622 = n24368 | n24621 ;
  assign n24624 = n73343 & n24622 ;
  assign n24625 = n24373 | n24624 ;
  assign n24626 = n73346 & n24625 ;
  assign n24627 = n24379 | n24626 ;
  assign n24629 = n73349 & n24627 ;
  assign n24630 = n24384 | n24629 ;
  assign n24631 = n73352 & n24630 ;
  assign n24632 = n24390 | n24631 ;
  assign n24634 = n73355 & n24632 ;
  assign n24635 = n24395 | n24634 ;
  assign n24636 = n73358 & n24635 ;
  assign n24637 = n24401 | n24636 ;
  assign n24639 = n73361 & n24637 ;
  assign n24640 = n24406 | n24639 ;
  assign n24641 = n73364 & n24640 ;
  assign n24642 = n24412 | n24641 ;
  assign n24644 = n73367 & n24642 ;
  assign n24645 = n24417 | n24644 ;
  assign n24646 = n73370 & n24645 ;
  assign n24647 = n24423 | n24646 ;
  assign n24649 = n73373 & n24647 ;
  assign n24650 = n24428 | n24649 ;
  assign n24651 = n73376 & n24650 ;
  assign n24652 = n24434 | n24651 ;
  assign n24654 = n73379 & n24652 ;
  assign n24655 = n24439 | n24654 ;
  assign n24656 = n73382 & n24655 ;
  assign n24657 = n24445 | n24656 ;
  assign n24659 = n73385 & n24657 ;
  assign n24660 = n24450 | n24659 ;
  assign n24661 = n73388 & n24660 ;
  assign n24662 = n24456 | n24661 ;
  assign n24664 = n73391 & n24662 ;
  assign n24665 = n24461 | n24664 ;
  assign n24666 = n73394 & n24665 ;
  assign n24667 = n24467 | n24666 ;
  assign n24669 = n73397 & n24667 ;
  assign n24670 = n24472 | n24669 ;
  assign n24671 = n73400 & n24670 ;
  assign n24672 = n24478 | n24671 ;
  assign n24674 = n73403 & n24672 ;
  assign n24675 = n24483 | n24674 ;
  assign n24676 = n73406 & n24675 ;
  assign n24677 = n24489 | n24676 ;
  assign n24679 = n73409 & n24677 ;
  assign n24680 = n24494 | n24679 ;
  assign n24681 = n73412 & n24680 ;
  assign n24682 = n24500 | n24681 ;
  assign n24684 = n73415 & n24682 ;
  assign n24685 = n24505 | n24684 ;
  assign n24686 = n73418 & n24685 ;
  assign n24687 = n24511 | n24686 ;
  assign n24689 = n73421 & n24687 ;
  assign n24690 = n24516 | n24689 ;
  assign n24691 = n73424 & n24690 ;
  assign n24692 = n24522 | n24691 ;
  assign n24694 = n73427 & n24692 ;
  assign n24695 = n24527 | n24694 ;
  assign n24696 = n73430 & n24695 ;
  assign n24697 = n24533 | n24696 ;
  assign n24699 = n73433 & n24697 ;
  assign n24700 = n24538 | n24699 ;
  assign n24701 = n73436 & n24700 ;
  assign n24702 = n24544 | n24701 ;
  assign n24704 = n73439 & n24702 ;
  assign n24705 = n24549 | n24704 ;
  assign n24706 = n73442 & n24705 ;
  assign n24707 = n24555 | n24706 ;
  assign n24709 = n73445 & n24707 ;
  assign n24710 = n24560 | n24709 ;
  assign n24711 = n73448 & n24710 ;
  assign n73456 = ~n24711 ;
  assign n24712 = n24566 & n73456 ;
  assign n24714 = n23827 | n24566 ;
  assign n73457 = ~n24714 ;
  assign n24715 = n24562 & n73457 ;
  assign n24716 = n24712 | n24715 ;
  assign n73458 = ~n24576 ;
  assign n24717 = n73458 & n24716 ;
  assign n73459 = ~n24574 ;
  assign n24718 = n73459 & n24717 ;
  assign n24719 = n24578 | n24718 ;
  assign n24720 = n73188 & n24719 ;
  assign n73460 = ~n24718 ;
  assign n25426 = x118 & n73460 ;
  assign n73461 = ~n24578 ;
  assign n25427 = n73461 & n25426 ;
  assign n25428 = n24720 | n25427 ;
  assign n24721 = n23826 & n24577 ;
  assign n73462 = ~n24557 ;
  assign n24561 = n73462 & n24560 ;
  assign n24722 = n23836 | n24560 ;
  assign n73463 = ~n24722 ;
  assign n24723 = n24707 & n73463 ;
  assign n24724 = n24561 | n24723 ;
  assign n24725 = n73458 & n24724 ;
  assign n24726 = n73459 & n24725 ;
  assign n24727 = n24721 | n24726 ;
  assign n24728 = n73177 & n24727 ;
  assign n24729 = n23835 & n24577 ;
  assign n73464 = ~n24706 ;
  assign n24708 = n24555 & n73464 ;
  assign n24730 = n23844 | n24555 ;
  assign n73465 = ~n24730 ;
  assign n24731 = n24551 & n73465 ;
  assign n24732 = n24708 | n24731 ;
  assign n24733 = n73458 & n24732 ;
  assign n24734 = n73459 & n24733 ;
  assign n24735 = n24729 | n24734 ;
  assign n24736 = n72752 & n24735 ;
  assign n73466 = ~n24734 ;
  assign n25415 = x116 & n73466 ;
  assign n73467 = ~n24729 ;
  assign n25416 = n73467 & n25415 ;
  assign n25417 = n24736 | n25416 ;
  assign n24737 = n23843 & n24577 ;
  assign n73468 = ~n24546 ;
  assign n24550 = n73468 & n24549 ;
  assign n24738 = n23853 | n24549 ;
  assign n73469 = ~n24738 ;
  assign n24739 = n24702 & n73469 ;
  assign n24740 = n24550 | n24739 ;
  assign n24741 = n73458 & n24740 ;
  assign n24742 = n73459 & n24741 ;
  assign n24743 = n24737 | n24742 ;
  assign n24744 = n72393 & n24743 ;
  assign n24745 = n23852 & n24577 ;
  assign n73470 = ~n24701 ;
  assign n24703 = n24544 & n73470 ;
  assign n24746 = n23862 | n24544 ;
  assign n73471 = ~n24746 ;
  assign n24747 = n24540 & n73471 ;
  assign n24748 = n24703 | n24747 ;
  assign n24749 = n73458 & n24748 ;
  assign n24750 = n73459 & n24749 ;
  assign n24751 = n24745 | n24750 ;
  assign n24752 = n72385 & n24751 ;
  assign n73472 = ~n24750 ;
  assign n25405 = x114 & n73472 ;
  assign n73473 = ~n24745 ;
  assign n25406 = n73473 & n25405 ;
  assign n25407 = n24752 | n25406 ;
  assign n24753 = n23861 & n24577 ;
  assign n73474 = ~n24535 ;
  assign n24539 = n73474 & n24538 ;
  assign n24754 = n23871 | n24538 ;
  assign n73475 = ~n24754 ;
  assign n24755 = n24697 & n73475 ;
  assign n24756 = n24539 | n24755 ;
  assign n24757 = n73458 & n24756 ;
  assign n24758 = n73459 & n24757 ;
  assign n24759 = n24753 | n24758 ;
  assign n24760 = n72025 & n24759 ;
  assign n24761 = n23870 & n24577 ;
  assign n73476 = ~n24696 ;
  assign n24698 = n24533 & n73476 ;
  assign n24762 = n23880 | n24533 ;
  assign n73477 = ~n24762 ;
  assign n24763 = n24529 & n73477 ;
  assign n24764 = n24698 | n24763 ;
  assign n24765 = n73458 & n24764 ;
  assign n24766 = n73459 & n24765 ;
  assign n24767 = n24761 | n24766 ;
  assign n24768 = n71645 & n24767 ;
  assign n73478 = ~n24766 ;
  assign n25394 = x112 & n73478 ;
  assign n73479 = ~n24761 ;
  assign n25395 = n73479 & n25394 ;
  assign n25396 = n24768 | n25395 ;
  assign n24769 = n23879 & n24577 ;
  assign n73480 = ~n24524 ;
  assign n24528 = n73480 & n24527 ;
  assign n24770 = n23888 | n24527 ;
  assign n73481 = ~n24770 ;
  assign n24771 = n24692 & n73481 ;
  assign n24772 = n24528 | n24771 ;
  assign n24773 = n73458 & n24772 ;
  assign n24774 = n73459 & n24773 ;
  assign n24775 = n24769 | n24774 ;
  assign n24776 = n71633 & n24775 ;
  assign n24777 = n23887 & n24577 ;
  assign n73482 = ~n24691 ;
  assign n24693 = n24522 & n73482 ;
  assign n24778 = n23897 | n24522 ;
  assign n73483 = ~n24778 ;
  assign n24779 = n24518 & n73483 ;
  assign n24780 = n24693 | n24779 ;
  assign n24781 = n73458 & n24780 ;
  assign n24782 = n73459 & n24781 ;
  assign n24783 = n24777 | n24782 ;
  assign n24784 = n71253 & n24783 ;
  assign n73484 = ~n24782 ;
  assign n25384 = x110 & n73484 ;
  assign n73485 = ~n24777 ;
  assign n25385 = n73485 & n25384 ;
  assign n25386 = n24784 | n25385 ;
  assign n24785 = n23896 & n24577 ;
  assign n73486 = ~n24513 ;
  assign n24517 = n73486 & n24516 ;
  assign n24786 = n23906 | n24516 ;
  assign n73487 = ~n24786 ;
  assign n24787 = n24687 & n73487 ;
  assign n24788 = n24517 | n24787 ;
  assign n24789 = n73458 & n24788 ;
  assign n24790 = n73459 & n24789 ;
  assign n24791 = n24785 | n24790 ;
  assign n24792 = n70935 & n24791 ;
  assign n24793 = n23905 & n24577 ;
  assign n73488 = ~n24686 ;
  assign n24688 = n24511 & n73488 ;
  assign n24794 = n23915 | n24511 ;
  assign n73489 = ~n24794 ;
  assign n24795 = n24507 & n73489 ;
  assign n24796 = n24688 | n24795 ;
  assign n24797 = n73458 & n24796 ;
  assign n24798 = n73459 & n24797 ;
  assign n24799 = n24793 | n24798 ;
  assign n24800 = n70927 & n24799 ;
  assign n73490 = ~n24798 ;
  assign n25374 = x108 & n73490 ;
  assign n73491 = ~n24793 ;
  assign n25375 = n73491 & n25374 ;
  assign n25376 = n24800 | n25375 ;
  assign n24801 = n23914 & n24577 ;
  assign n73492 = ~n24502 ;
  assign n24506 = n73492 & n24505 ;
  assign n24802 = n23923 | n24505 ;
  assign n73493 = ~n24802 ;
  assign n24803 = n24682 & n73493 ;
  assign n24804 = n24506 | n24803 ;
  assign n24805 = n73458 & n24804 ;
  assign n24806 = n73459 & n24805 ;
  assign n24807 = n24801 | n24806 ;
  assign n24808 = n70609 & n24807 ;
  assign n24809 = n23922 & n24577 ;
  assign n73494 = ~n24681 ;
  assign n24683 = n24500 & n73494 ;
  assign n24810 = n23932 | n24500 ;
  assign n73495 = ~n24810 ;
  assign n24811 = n24496 & n73495 ;
  assign n24812 = n24683 | n24811 ;
  assign n24813 = n73458 & n24812 ;
  assign n24814 = n73459 & n24813 ;
  assign n24815 = n24809 | n24814 ;
  assign n24816 = n70276 & n24815 ;
  assign n73496 = ~n24814 ;
  assign n25363 = x106 & n73496 ;
  assign n73497 = ~n24809 ;
  assign n25364 = n73497 & n25363 ;
  assign n25365 = n24816 | n25364 ;
  assign n24817 = n23931 & n24577 ;
  assign n73498 = ~n24491 ;
  assign n24495 = n73498 & n24494 ;
  assign n24818 = n23941 | n24494 ;
  assign n73499 = ~n24818 ;
  assign n24819 = n24677 & n73499 ;
  assign n24820 = n24495 | n24819 ;
  assign n24821 = n73458 & n24820 ;
  assign n24822 = n73459 & n24821 ;
  assign n24823 = n24817 | n24822 ;
  assign n24824 = n70176 & n24823 ;
  assign n24825 = n23940 & n24577 ;
  assign n73500 = ~n24676 ;
  assign n24678 = n24489 & n73500 ;
  assign n24826 = n23950 | n24489 ;
  assign n73501 = ~n24826 ;
  assign n24827 = n24485 & n73501 ;
  assign n24828 = n24678 | n24827 ;
  assign n24829 = n73458 & n24828 ;
  assign n24830 = n73459 & n24829 ;
  assign n24831 = n24825 | n24830 ;
  assign n24832 = n69857 & n24831 ;
  assign n73502 = ~n24830 ;
  assign n25352 = x104 & n73502 ;
  assign n73503 = ~n24825 ;
  assign n25353 = n73503 & n25352 ;
  assign n25354 = n24832 | n25353 ;
  assign n24833 = n23949 & n24577 ;
  assign n73504 = ~n24480 ;
  assign n24484 = n73504 & n24483 ;
  assign n24834 = n23959 | n24483 ;
  assign n73505 = ~n24834 ;
  assign n24835 = n24672 & n73505 ;
  assign n24836 = n24484 | n24835 ;
  assign n24837 = n73458 & n24836 ;
  assign n24838 = n73459 & n24837 ;
  assign n24839 = n24833 | n24838 ;
  assign n24840 = n69656 & n24839 ;
  assign n24841 = n23958 & n24577 ;
  assign n73506 = ~n24671 ;
  assign n24673 = n24478 & n73506 ;
  assign n24842 = n23968 | n24478 ;
  assign n73507 = ~n24842 ;
  assign n24843 = n24474 & n73507 ;
  assign n24844 = n24673 | n24843 ;
  assign n24845 = n73458 & n24844 ;
  assign n24846 = n73459 & n24845 ;
  assign n24847 = n24841 | n24846 ;
  assign n24848 = n69528 & n24847 ;
  assign n73508 = ~n24846 ;
  assign n25341 = x102 & n73508 ;
  assign n73509 = ~n24841 ;
  assign n25342 = n73509 & n25341 ;
  assign n25343 = n24848 | n25342 ;
  assign n24849 = n23967 & n24577 ;
  assign n73510 = ~n24469 ;
  assign n24473 = n73510 & n24472 ;
  assign n24850 = n23977 | n24472 ;
  assign n73511 = ~n24850 ;
  assign n24851 = n24667 & n73511 ;
  assign n24852 = n24473 | n24851 ;
  assign n24853 = n73458 & n24852 ;
  assign n24854 = n73459 & n24853 ;
  assign n24855 = n24849 | n24854 ;
  assign n24856 = n69261 & n24855 ;
  assign n24857 = n23976 & n24577 ;
  assign n73512 = ~n24666 ;
  assign n24668 = n24467 & n73512 ;
  assign n24858 = n23986 | n24467 ;
  assign n73513 = ~n24858 ;
  assign n24859 = n24463 & n73513 ;
  assign n24860 = n24668 | n24859 ;
  assign n24861 = n73458 & n24860 ;
  assign n24862 = n73459 & n24861 ;
  assign n24863 = n24857 | n24862 ;
  assign n24864 = n69075 & n24863 ;
  assign n73514 = ~n24862 ;
  assign n25331 = x100 & n73514 ;
  assign n73515 = ~n24857 ;
  assign n25332 = n73515 & n25331 ;
  assign n25333 = n24864 | n25332 ;
  assign n24865 = n23985 & n24577 ;
  assign n73516 = ~n24458 ;
  assign n24462 = n73516 & n24461 ;
  assign n24866 = n23995 | n24461 ;
  assign n73517 = ~n24866 ;
  assign n24867 = n24662 & n73517 ;
  assign n24868 = n24462 | n24867 ;
  assign n24869 = n73458 & n24868 ;
  assign n24870 = n73459 & n24869 ;
  assign n24871 = n24865 | n24870 ;
  assign n24872 = n68993 & n24871 ;
  assign n24873 = n23994 & n24577 ;
  assign n73518 = ~n24661 ;
  assign n24663 = n24456 & n73518 ;
  assign n24874 = n24004 | n24456 ;
  assign n73519 = ~n24874 ;
  assign n24875 = n24452 & n73519 ;
  assign n24876 = n24663 | n24875 ;
  assign n24877 = n73458 & n24876 ;
  assign n24878 = n73459 & n24877 ;
  assign n24879 = n24873 | n24878 ;
  assign n24880 = n68716 & n24879 ;
  assign n73520 = ~n24878 ;
  assign n25321 = x98 & n73520 ;
  assign n73521 = ~n24873 ;
  assign n25322 = n73521 & n25321 ;
  assign n25323 = n24880 | n25322 ;
  assign n24881 = n24003 & n24577 ;
  assign n73522 = ~n24447 ;
  assign n24451 = n73522 & n24450 ;
  assign n24882 = n24013 | n24450 ;
  assign n73523 = ~n24882 ;
  assign n24883 = n24657 & n73523 ;
  assign n24884 = n24451 | n24883 ;
  assign n24885 = n73458 & n24884 ;
  assign n24886 = n73459 & n24885 ;
  assign n24887 = n24881 | n24886 ;
  assign n24888 = n68545 & n24887 ;
  assign n24889 = n24012 & n24577 ;
  assign n73524 = ~n24656 ;
  assign n24658 = n24445 & n73524 ;
  assign n24890 = n24022 | n24445 ;
  assign n73525 = ~n24890 ;
  assign n24891 = n24441 & n73525 ;
  assign n24892 = n24658 | n24891 ;
  assign n24893 = n73458 & n24892 ;
  assign n24894 = n73459 & n24893 ;
  assign n24895 = n24889 | n24894 ;
  assign n24896 = n68438 & n24895 ;
  assign n73526 = ~n24894 ;
  assign n25311 = x96 & n73526 ;
  assign n73527 = ~n24889 ;
  assign n25312 = n73527 & n25311 ;
  assign n25313 = n24896 | n25312 ;
  assign n24897 = n24021 & n24577 ;
  assign n73528 = ~n24436 ;
  assign n24440 = n73528 & n24439 ;
  assign n24898 = n24031 | n24439 ;
  assign n73529 = ~n24898 ;
  assign n24899 = n24652 & n73529 ;
  assign n24900 = n24440 | n24899 ;
  assign n24901 = n73458 & n24900 ;
  assign n24902 = n73459 & n24901 ;
  assign n24903 = n24897 | n24902 ;
  assign n24904 = n68214 & n24903 ;
  assign n24905 = n24030 & n24577 ;
  assign n73530 = ~n24651 ;
  assign n24653 = n24434 & n73530 ;
  assign n24906 = n24040 | n24434 ;
  assign n73531 = ~n24906 ;
  assign n24907 = n24430 & n73531 ;
  assign n24908 = n24653 | n24907 ;
  assign n24909 = n73458 & n24908 ;
  assign n24910 = n73459 & n24909 ;
  assign n24911 = n24905 | n24910 ;
  assign n24912 = n68058 & n24911 ;
  assign n73532 = ~n24910 ;
  assign n25301 = x94 & n73532 ;
  assign n73533 = ~n24905 ;
  assign n25302 = n73533 & n25301 ;
  assign n25303 = n24912 | n25302 ;
  assign n24913 = n24039 & n24577 ;
  assign n73534 = ~n24425 ;
  assign n24429 = n73534 & n24428 ;
  assign n24914 = n24049 | n24428 ;
  assign n73535 = ~n24914 ;
  assign n24915 = n24647 & n73535 ;
  assign n24916 = n24429 | n24915 ;
  assign n24917 = n73458 & n24916 ;
  assign n24918 = n73459 & n24917 ;
  assign n24919 = n24913 | n24918 ;
  assign n24920 = n67986 & n24919 ;
  assign n24921 = n24048 & n24577 ;
  assign n73536 = ~n24646 ;
  assign n24648 = n24423 & n73536 ;
  assign n24922 = n24058 | n24423 ;
  assign n73537 = ~n24922 ;
  assign n24923 = n24419 & n73537 ;
  assign n24924 = n24648 | n24923 ;
  assign n24925 = n73458 & n24924 ;
  assign n24926 = n73459 & n24925 ;
  assign n24927 = n24921 | n24926 ;
  assign n24928 = n67763 & n24927 ;
  assign n73538 = ~n24926 ;
  assign n25291 = x92 & n73538 ;
  assign n73539 = ~n24921 ;
  assign n25292 = n73539 & n25291 ;
  assign n25293 = n24928 | n25292 ;
  assign n24929 = n24057 & n24577 ;
  assign n73540 = ~n24414 ;
  assign n24418 = n73540 & n24417 ;
  assign n24930 = n24066 | n24417 ;
  assign n73541 = ~n24930 ;
  assign n24931 = n24642 & n73541 ;
  assign n24932 = n24418 | n24931 ;
  assign n24933 = n73458 & n24932 ;
  assign n24934 = n73459 & n24933 ;
  assign n24935 = n24929 | n24934 ;
  assign n24936 = n67622 & n24935 ;
  assign n24937 = n24065 & n24577 ;
  assign n73542 = ~n24641 ;
  assign n24643 = n24412 & n73542 ;
  assign n24938 = n24075 | n24412 ;
  assign n73543 = ~n24938 ;
  assign n24939 = n24408 & n73543 ;
  assign n24940 = n24643 | n24939 ;
  assign n24941 = n73458 & n24940 ;
  assign n24942 = n73459 & n24941 ;
  assign n24943 = n24937 | n24942 ;
  assign n24944 = n67531 & n24943 ;
  assign n73544 = ~n24942 ;
  assign n25281 = x90 & n73544 ;
  assign n73545 = ~n24937 ;
  assign n25282 = n73545 & n25281 ;
  assign n25283 = n24944 | n25282 ;
  assign n24945 = n24074 & n24577 ;
  assign n73546 = ~n24403 ;
  assign n24407 = n73546 & n24406 ;
  assign n24946 = n24084 | n24406 ;
  assign n73547 = ~n24946 ;
  assign n24947 = n24637 & n73547 ;
  assign n24948 = n24407 | n24947 ;
  assign n24949 = n73458 & n24948 ;
  assign n24950 = n73459 & n24949 ;
  assign n24951 = n24945 | n24950 ;
  assign n24952 = n67348 & n24951 ;
  assign n24953 = n24083 & n24577 ;
  assign n73548 = ~n24636 ;
  assign n24638 = n24401 & n73548 ;
  assign n24954 = n24092 | n24401 ;
  assign n73549 = ~n24954 ;
  assign n24955 = n24397 & n73549 ;
  assign n24956 = n24638 | n24955 ;
  assign n24957 = n73458 & n24956 ;
  assign n24958 = n73459 & n24957 ;
  assign n24959 = n24953 | n24958 ;
  assign n24960 = n67222 & n24959 ;
  assign n73550 = ~n24958 ;
  assign n25271 = x88 & n73550 ;
  assign n73551 = ~n24953 ;
  assign n25272 = n73551 & n25271 ;
  assign n25273 = n24960 | n25272 ;
  assign n24961 = n24091 & n24577 ;
  assign n73552 = ~n24392 ;
  assign n24396 = n73552 & n24395 ;
  assign n24962 = n24100 | n24395 ;
  assign n73553 = ~n24962 ;
  assign n24963 = n24632 & n73553 ;
  assign n24964 = n24396 | n24963 ;
  assign n24965 = n73458 & n24964 ;
  assign n24966 = n73459 & n24965 ;
  assign n24967 = n24961 | n24966 ;
  assign n24968 = n67164 & n24967 ;
  assign n24969 = n24099 & n24577 ;
  assign n73554 = ~n24631 ;
  assign n24633 = n24390 & n73554 ;
  assign n24970 = n24109 | n24390 ;
  assign n73555 = ~n24970 ;
  assign n24971 = n24386 & n73555 ;
  assign n24972 = n24633 | n24971 ;
  assign n24973 = n73458 & n24972 ;
  assign n24974 = n73459 & n24973 ;
  assign n24975 = n24969 | n24974 ;
  assign n24976 = n66979 & n24975 ;
  assign n73556 = ~n24974 ;
  assign n25261 = x86 & n73556 ;
  assign n73557 = ~n24969 ;
  assign n25262 = n73557 & n25261 ;
  assign n25263 = n24976 | n25262 ;
  assign n24977 = n24108 & n24577 ;
  assign n73558 = ~n24381 ;
  assign n24385 = n73558 & n24384 ;
  assign n24978 = n24118 | n24384 ;
  assign n73559 = ~n24978 ;
  assign n24979 = n24627 & n73559 ;
  assign n24980 = n24385 | n24979 ;
  assign n24981 = n73458 & n24980 ;
  assign n24982 = n73459 & n24981 ;
  assign n24983 = n24977 | n24982 ;
  assign n24984 = n66868 & n24983 ;
  assign n24985 = n24117 & n24577 ;
  assign n73560 = ~n24626 ;
  assign n24628 = n24379 & n73560 ;
  assign n24986 = n24127 | n24379 ;
  assign n73561 = ~n24986 ;
  assign n24987 = n24375 & n73561 ;
  assign n24988 = n24628 | n24987 ;
  assign n24989 = n73458 & n24988 ;
  assign n24990 = n73459 & n24989 ;
  assign n24991 = n24985 | n24990 ;
  assign n24992 = n66797 & n24991 ;
  assign n73562 = ~n24990 ;
  assign n25251 = x84 & n73562 ;
  assign n73563 = ~n24985 ;
  assign n25252 = n73563 & n25251 ;
  assign n25253 = n24992 | n25252 ;
  assign n24993 = n24126 & n24577 ;
  assign n73564 = ~n24370 ;
  assign n24374 = n73564 & n24373 ;
  assign n24994 = n24135 | n24373 ;
  assign n73565 = ~n24994 ;
  assign n24995 = n24622 & n73565 ;
  assign n24996 = n24374 | n24995 ;
  assign n24997 = n73458 & n24996 ;
  assign n24998 = n73459 & n24997 ;
  assign n24999 = n24993 | n24998 ;
  assign n25000 = n66654 & n24999 ;
  assign n25001 = n24134 & n24577 ;
  assign n73566 = ~n24621 ;
  assign n24623 = n24368 & n73566 ;
  assign n25002 = n24143 | n24368 ;
  assign n73567 = ~n25002 ;
  assign n25003 = n24364 & n73567 ;
  assign n25004 = n24623 | n25003 ;
  assign n25005 = n73458 & n25004 ;
  assign n25006 = n73459 & n25005 ;
  assign n25007 = n25001 | n25006 ;
  assign n25008 = n66560 & n25007 ;
  assign n73568 = ~n25006 ;
  assign n25241 = x82 & n73568 ;
  assign n73569 = ~n25001 ;
  assign n25242 = n73569 & n25241 ;
  assign n25243 = n25008 | n25242 ;
  assign n25009 = n24142 & n24577 ;
  assign n73570 = ~n24359 ;
  assign n24363 = n73570 & n24362 ;
  assign n25010 = n24152 | n24362 ;
  assign n73571 = ~n25010 ;
  assign n25011 = n24617 & n73571 ;
  assign n25012 = n24363 | n25011 ;
  assign n25013 = n73458 & n25012 ;
  assign n25014 = n73459 & n25013 ;
  assign n25015 = n25009 | n25014 ;
  assign n25016 = n66505 & n25015 ;
  assign n25017 = n24151 & n24577 ;
  assign n73572 = ~n24616 ;
  assign n24618 = n24357 & n73572 ;
  assign n25018 = n24161 | n24357 ;
  assign n73573 = ~n25018 ;
  assign n25019 = n24353 & n73573 ;
  assign n25020 = n24618 | n25019 ;
  assign n25021 = n73458 & n25020 ;
  assign n25022 = n73459 & n25021 ;
  assign n25023 = n25017 | n25022 ;
  assign n25024 = n66379 & n25023 ;
  assign n73574 = ~n25022 ;
  assign n25231 = x80 & n73574 ;
  assign n73575 = ~n25017 ;
  assign n25232 = n73575 & n25231 ;
  assign n25233 = n25024 | n25232 ;
  assign n25025 = n24160 & n24577 ;
  assign n73576 = ~n24348 ;
  assign n24352 = n73576 & n24351 ;
  assign n25026 = n24170 | n24351 ;
  assign n73577 = ~n25026 ;
  assign n25027 = n24612 & n73577 ;
  assign n25028 = n24352 | n25027 ;
  assign n25029 = n73458 & n25028 ;
  assign n25030 = n73459 & n25029 ;
  assign n25031 = n25025 | n25030 ;
  assign n25032 = n66299 & n25031 ;
  assign n25033 = n24169 & n24577 ;
  assign n73578 = ~n24611 ;
  assign n24613 = n24346 & n73578 ;
  assign n25034 = n24179 | n24346 ;
  assign n73579 = ~n25034 ;
  assign n25035 = n24342 & n73579 ;
  assign n25036 = n24613 | n25035 ;
  assign n25037 = n73458 & n25036 ;
  assign n25038 = n73459 & n25037 ;
  assign n25039 = n25033 | n25038 ;
  assign n25040 = n66244 & n25039 ;
  assign n73580 = ~n25038 ;
  assign n25220 = x78 & n73580 ;
  assign n73581 = ~n25033 ;
  assign n25221 = n73581 & n25220 ;
  assign n25222 = n25040 | n25221 ;
  assign n25041 = n24178 & n24577 ;
  assign n73582 = ~n24337 ;
  assign n24341 = n73582 & n24340 ;
  assign n25042 = n24188 | n24340 ;
  assign n73583 = ~n25042 ;
  assign n25043 = n24607 & n73583 ;
  assign n25044 = n24341 | n25043 ;
  assign n25045 = n73458 & n25044 ;
  assign n25046 = n73459 & n25045 ;
  assign n25047 = n25041 | n25046 ;
  assign n25048 = n66145 & n25047 ;
  assign n25049 = n24187 & n24577 ;
  assign n73584 = ~n24606 ;
  assign n24608 = n24335 & n73584 ;
  assign n25050 = n24196 | n24335 ;
  assign n73585 = ~n25050 ;
  assign n25051 = n24331 & n73585 ;
  assign n25052 = n24608 | n25051 ;
  assign n25053 = n73458 & n25052 ;
  assign n25054 = n73459 & n25053 ;
  assign n25055 = n25049 | n25054 ;
  assign n25056 = n66081 & n25055 ;
  assign n73586 = ~n25054 ;
  assign n25210 = x76 & n73586 ;
  assign n73587 = ~n25049 ;
  assign n25211 = n73587 & n25210 ;
  assign n25212 = n25056 | n25211 ;
  assign n25057 = n24195 & n24577 ;
  assign n73588 = ~n24326 ;
  assign n24330 = n73588 & n24329 ;
  assign n25058 = n24205 | n24329 ;
  assign n73589 = ~n25058 ;
  assign n25059 = n24602 & n73589 ;
  assign n25060 = n24330 | n25059 ;
  assign n25061 = n73458 & n25060 ;
  assign n25062 = n73459 & n25061 ;
  assign n25063 = n25057 | n25062 ;
  assign n25064 = n66043 & n25063 ;
  assign n25065 = n24204 & n24577 ;
  assign n73590 = ~n24601 ;
  assign n24603 = n24324 & n73590 ;
  assign n25066 = n24214 | n24324 ;
  assign n73591 = ~n25066 ;
  assign n25067 = n24320 & n73591 ;
  assign n25068 = n24603 | n25067 ;
  assign n25069 = n73458 & n25068 ;
  assign n25070 = n73459 & n25069 ;
  assign n25071 = n25065 | n25070 ;
  assign n25072 = n65960 & n25071 ;
  assign n73592 = ~n25070 ;
  assign n25200 = x74 & n73592 ;
  assign n73593 = ~n25065 ;
  assign n25201 = n73593 & n25200 ;
  assign n25202 = n25072 | n25201 ;
  assign n25073 = n24213 & n24577 ;
  assign n73594 = ~n24315 ;
  assign n24319 = n73594 & n24318 ;
  assign n25074 = n24223 | n24318 ;
  assign n73595 = ~n25074 ;
  assign n25075 = n24597 & n73595 ;
  assign n25076 = n24319 | n25075 ;
  assign n25077 = n73458 & n25076 ;
  assign n25078 = n73459 & n25077 ;
  assign n25079 = n25073 | n25078 ;
  assign n25080 = n65909 & n25079 ;
  assign n25081 = n24222 & n24577 ;
  assign n73596 = ~n24596 ;
  assign n24598 = n24313 & n73596 ;
  assign n25082 = n24232 | n24313 ;
  assign n73597 = ~n25082 ;
  assign n25083 = n24308 & n73597 ;
  assign n25084 = n24598 | n25083 ;
  assign n25085 = n73458 & n25084 ;
  assign n25086 = n73459 & n25085 ;
  assign n25087 = n25081 | n25086 ;
  assign n25088 = n65877 & n25087 ;
  assign n73598 = ~n25086 ;
  assign n25190 = x72 & n73598 ;
  assign n73599 = ~n25081 ;
  assign n25191 = n73599 & n25190 ;
  assign n25192 = n25088 | n25191 ;
  assign n25089 = n24231 & n24577 ;
  assign n73600 = ~n24303 ;
  assign n24307 = n73600 & n24306 ;
  assign n24309 = n24241 | n24306 ;
  assign n25090 = n24301 | n24591 ;
  assign n73601 = ~n24309 ;
  assign n25091 = n73601 & n25090 ;
  assign n25092 = n24307 | n25091 ;
  assign n25093 = n73458 & n25092 ;
  assign n25094 = n73459 & n25093 ;
  assign n25095 = n25089 | n25094 ;
  assign n25096 = n65820 & n25095 ;
  assign n25097 = n24240 & n24577 ;
  assign n73602 = ~n24591 ;
  assign n24593 = n24301 & n73602 ;
  assign n25098 = n24294 | n24588 ;
  assign n25099 = n24250 | n24301 ;
  assign n73603 = ~n25099 ;
  assign n25100 = n25098 & n73603 ;
  assign n25101 = n24593 | n25100 ;
  assign n25102 = n73458 & n25101 ;
  assign n25103 = n73459 & n25102 ;
  assign n25104 = n25097 | n25103 ;
  assign n25105 = n65791 & n25104 ;
  assign n73604 = ~n25103 ;
  assign n25180 = x70 & n73604 ;
  assign n73605 = ~n25097 ;
  assign n25181 = n73605 & n25180 ;
  assign n25182 = n25105 | n25181 ;
  assign n25106 = n24249 & n24577 ;
  assign n73606 = ~n24294 ;
  assign n24589 = n73606 & n24588 ;
  assign n25107 = n24292 | n24584 ;
  assign n25108 = n24258 | n24588 ;
  assign n73607 = ~n25108 ;
  assign n25109 = n25107 & n73607 ;
  assign n25110 = n24589 | n25109 ;
  assign n25111 = n73458 & n25110 ;
  assign n25112 = n73459 & n25111 ;
  assign n25113 = n25106 | n25112 ;
  assign n25114 = n65772 & n25113 ;
  assign n25115 = n24257 & n24577 ;
  assign n73608 = ~n24584 ;
  assign n24586 = n24292 & n73608 ;
  assign n25116 = n24266 | n24292 ;
  assign n73609 = ~n25116 ;
  assign n25117 = n24583 & n73609 ;
  assign n25118 = n24586 | n25117 ;
  assign n25119 = n73458 & n25118 ;
  assign n25120 = n73459 & n25119 ;
  assign n25121 = n25115 | n25120 ;
  assign n25122 = n65746 & n25121 ;
  assign n73610 = ~n25120 ;
  assign n25170 = x68 & n73610 ;
  assign n73611 = ~n25115 ;
  assign n25171 = n73611 & n25170 ;
  assign n25172 = n25122 | n25171 ;
  assign n25123 = n24265 & n24577 ;
  assign n25124 = n24282 | n24287 ;
  assign n73612 = ~n25124 ;
  assign n25125 = n24581 & n73612 ;
  assign n73613 = ~n24284 ;
  assign n25126 = n73613 & n24287 ;
  assign n25127 = n25125 | n25126 ;
  assign n25128 = n73458 & n25127 ;
  assign n25129 = n73459 & n25128 ;
  assign n25130 = n25123 | n25129 ;
  assign n25131 = n65721 & n25130 ;
  assign n25132 = n24276 & n24577 ;
  assign n25133 = n24279 & n24281 ;
  assign n25134 = n73455 & n25133 ;
  assign n25135 = n24576 | n25134 ;
  assign n73614 = ~n25135 ;
  assign n25136 = n24581 & n73614 ;
  assign n25137 = n73459 & n25136 ;
  assign n25138 = n25132 | n25137 ;
  assign n25139 = n65686 & n25138 ;
  assign n73615 = ~n25137 ;
  assign n25160 = x66 & n73615 ;
  assign n73616 = ~n25132 ;
  assign n25161 = n73616 & n25160 ;
  assign n25162 = n25139 | n25161 ;
  assign n24713 = n24566 | n24711 ;
  assign n25140 = n73451 & n24713 ;
  assign n25141 = n24571 | n25140 ;
  assign n25142 = n73454 & n25141 ;
  assign n73617 = ~x119 ;
  assign n25143 = x64 & n73617 ;
  assign n73618 = ~n65392 ;
  assign n25144 = n73618 & n25143 ;
  assign n73619 = ~n65369 ;
  assign n25145 = n73619 & n25144 ;
  assign n73620 = ~n25142 ;
  assign n25146 = n73620 & n25145 ;
  assign n73621 = ~n25146 ;
  assign n25147 = x9 & n73621 ;
  assign n73622 = ~n267 ;
  assign n25148 = n73622 & n24281 ;
  assign n73623 = ~n277 ;
  assign n25149 = n73623 & n25148 ;
  assign n73624 = ~n274 ;
  assign n25150 = n73624 & n25149 ;
  assign n25151 = n73459 & n25150 ;
  assign n25152 = n25147 | n25151 ;
  assign n25153 = x65 & n25152 ;
  assign n25154 = x65 | n25151 ;
  assign n25155 = n25147 | n25154 ;
  assign n73625 = ~n25153 ;
  assign n25156 = n73625 & n25155 ;
  assign n73626 = ~x8 ;
  assign n25157 = n73626 & x64 ;
  assign n25158 = n25156 | n25157 ;
  assign n25159 = n65670 & n25152 ;
  assign n73627 = ~n25159 ;
  assign n25163 = n25158 & n73627 ;
  assign n25164 = n25162 | n25163 ;
  assign n73628 = ~n25139 ;
  assign n25165 = n73628 & n25164 ;
  assign n73629 = ~n25129 ;
  assign n25166 = x67 & n73629 ;
  assign n73630 = ~n25123 ;
  assign n25167 = n73630 & n25166 ;
  assign n25168 = n25131 | n25167 ;
  assign n25169 = n25165 | n25168 ;
  assign n73631 = ~n25131 ;
  assign n25173 = n73631 & n25169 ;
  assign n25174 = n25172 | n25173 ;
  assign n73632 = ~n25122 ;
  assign n25175 = n73632 & n25174 ;
  assign n73633 = ~n25112 ;
  assign n25176 = x69 & n73633 ;
  assign n73634 = ~n25106 ;
  assign n25177 = n73634 & n25176 ;
  assign n25178 = n25114 | n25177 ;
  assign n25179 = n25175 | n25178 ;
  assign n73635 = ~n25114 ;
  assign n25183 = n73635 & n25179 ;
  assign n25184 = n25182 | n25183 ;
  assign n73636 = ~n25105 ;
  assign n25185 = n73636 & n25184 ;
  assign n73637 = ~n25094 ;
  assign n25186 = x71 & n73637 ;
  assign n73638 = ~n25089 ;
  assign n25187 = n73638 & n25186 ;
  assign n25188 = n25096 | n25187 ;
  assign n25189 = n25185 | n25188 ;
  assign n73639 = ~n25096 ;
  assign n25193 = n73639 & n25189 ;
  assign n25194 = n25192 | n25193 ;
  assign n73640 = ~n25088 ;
  assign n25195 = n73640 & n25194 ;
  assign n73641 = ~n25078 ;
  assign n25196 = x73 & n73641 ;
  assign n73642 = ~n25073 ;
  assign n25197 = n73642 & n25196 ;
  assign n25198 = n25080 | n25197 ;
  assign n25199 = n25195 | n25198 ;
  assign n73643 = ~n25080 ;
  assign n25203 = n73643 & n25199 ;
  assign n25204 = n25202 | n25203 ;
  assign n73644 = ~n25072 ;
  assign n25205 = n73644 & n25204 ;
  assign n73645 = ~n25062 ;
  assign n25206 = x75 & n73645 ;
  assign n73646 = ~n25057 ;
  assign n25207 = n73646 & n25206 ;
  assign n25208 = n25064 | n25207 ;
  assign n25209 = n25205 | n25208 ;
  assign n73647 = ~n25064 ;
  assign n25213 = n73647 & n25209 ;
  assign n25214 = n25212 | n25213 ;
  assign n73648 = ~n25056 ;
  assign n25215 = n73648 & n25214 ;
  assign n73649 = ~n25046 ;
  assign n25216 = x77 & n73649 ;
  assign n73650 = ~n25041 ;
  assign n25217 = n73650 & n25216 ;
  assign n25218 = n25048 | n25217 ;
  assign n25219 = n25215 | n25218 ;
  assign n73651 = ~n25048 ;
  assign n25223 = n73651 & n25219 ;
  assign n25224 = n25222 | n25223 ;
  assign n73652 = ~n25040 ;
  assign n25225 = n73652 & n25224 ;
  assign n73653 = ~n25030 ;
  assign n25226 = x79 & n73653 ;
  assign n73654 = ~n25025 ;
  assign n25227 = n73654 & n25226 ;
  assign n25228 = n25032 | n25227 ;
  assign n25230 = n25225 | n25228 ;
  assign n73655 = ~n25032 ;
  assign n25234 = n73655 & n25230 ;
  assign n25235 = n25233 | n25234 ;
  assign n73656 = ~n25024 ;
  assign n25236 = n73656 & n25235 ;
  assign n73657 = ~n25014 ;
  assign n25237 = x81 & n73657 ;
  assign n73658 = ~n25009 ;
  assign n25238 = n73658 & n25237 ;
  assign n25239 = n25016 | n25238 ;
  assign n25240 = n25236 | n25239 ;
  assign n73659 = ~n25016 ;
  assign n25244 = n73659 & n25240 ;
  assign n25245 = n25243 | n25244 ;
  assign n73660 = ~n25008 ;
  assign n25246 = n73660 & n25245 ;
  assign n73661 = ~n24998 ;
  assign n25247 = x83 & n73661 ;
  assign n73662 = ~n24993 ;
  assign n25248 = n73662 & n25247 ;
  assign n25249 = n25000 | n25248 ;
  assign n25250 = n25246 | n25249 ;
  assign n73663 = ~n25000 ;
  assign n25254 = n73663 & n25250 ;
  assign n25255 = n25253 | n25254 ;
  assign n73664 = ~n24992 ;
  assign n25256 = n73664 & n25255 ;
  assign n73665 = ~n24982 ;
  assign n25257 = x85 & n73665 ;
  assign n73666 = ~n24977 ;
  assign n25258 = n73666 & n25257 ;
  assign n25259 = n24984 | n25258 ;
  assign n25260 = n25256 | n25259 ;
  assign n73667 = ~n24984 ;
  assign n25264 = n73667 & n25260 ;
  assign n25265 = n25263 | n25264 ;
  assign n73668 = ~n24976 ;
  assign n25266 = n73668 & n25265 ;
  assign n73669 = ~n24966 ;
  assign n25267 = x87 & n73669 ;
  assign n73670 = ~n24961 ;
  assign n25268 = n73670 & n25267 ;
  assign n25269 = n24968 | n25268 ;
  assign n25270 = n25266 | n25269 ;
  assign n73671 = ~n24968 ;
  assign n25274 = n73671 & n25270 ;
  assign n25275 = n25273 | n25274 ;
  assign n73672 = ~n24960 ;
  assign n25276 = n73672 & n25275 ;
  assign n73673 = ~n24950 ;
  assign n25277 = x89 & n73673 ;
  assign n73674 = ~n24945 ;
  assign n25278 = n73674 & n25277 ;
  assign n25279 = n24952 | n25278 ;
  assign n25280 = n25276 | n25279 ;
  assign n73675 = ~n24952 ;
  assign n25284 = n73675 & n25280 ;
  assign n25285 = n25283 | n25284 ;
  assign n73676 = ~n24944 ;
  assign n25286 = n73676 & n25285 ;
  assign n73677 = ~n24934 ;
  assign n25287 = x91 & n73677 ;
  assign n73678 = ~n24929 ;
  assign n25288 = n73678 & n25287 ;
  assign n25289 = n24936 | n25288 ;
  assign n25290 = n25286 | n25289 ;
  assign n73679 = ~n24936 ;
  assign n25294 = n73679 & n25290 ;
  assign n25295 = n25293 | n25294 ;
  assign n73680 = ~n24928 ;
  assign n25296 = n73680 & n25295 ;
  assign n73681 = ~n24918 ;
  assign n25297 = x93 & n73681 ;
  assign n73682 = ~n24913 ;
  assign n25298 = n73682 & n25297 ;
  assign n25299 = n24920 | n25298 ;
  assign n25300 = n25296 | n25299 ;
  assign n73683 = ~n24920 ;
  assign n25304 = n73683 & n25300 ;
  assign n25305 = n25303 | n25304 ;
  assign n73684 = ~n24912 ;
  assign n25306 = n73684 & n25305 ;
  assign n73685 = ~n24902 ;
  assign n25307 = x95 & n73685 ;
  assign n73686 = ~n24897 ;
  assign n25308 = n73686 & n25307 ;
  assign n25309 = n24904 | n25308 ;
  assign n25310 = n25306 | n25309 ;
  assign n73687 = ~n24904 ;
  assign n25314 = n73687 & n25310 ;
  assign n25315 = n25313 | n25314 ;
  assign n73688 = ~n24896 ;
  assign n25316 = n73688 & n25315 ;
  assign n73689 = ~n24886 ;
  assign n25317 = x97 & n73689 ;
  assign n73690 = ~n24881 ;
  assign n25318 = n73690 & n25317 ;
  assign n25319 = n24888 | n25318 ;
  assign n25320 = n25316 | n25319 ;
  assign n73691 = ~n24888 ;
  assign n25324 = n73691 & n25320 ;
  assign n25325 = n25323 | n25324 ;
  assign n73692 = ~n24880 ;
  assign n25326 = n73692 & n25325 ;
  assign n73693 = ~n24870 ;
  assign n25327 = x99 & n73693 ;
  assign n73694 = ~n24865 ;
  assign n25328 = n73694 & n25327 ;
  assign n25329 = n24872 | n25328 ;
  assign n25330 = n25326 | n25329 ;
  assign n73695 = ~n24872 ;
  assign n25334 = n73695 & n25330 ;
  assign n25335 = n25333 | n25334 ;
  assign n73696 = ~n24864 ;
  assign n25336 = n73696 & n25335 ;
  assign n73697 = ~n24854 ;
  assign n25337 = x101 & n73697 ;
  assign n73698 = ~n24849 ;
  assign n25338 = n73698 & n25337 ;
  assign n25339 = n24856 | n25338 ;
  assign n25340 = n25336 | n25339 ;
  assign n73699 = ~n24856 ;
  assign n25344 = n73699 & n25340 ;
  assign n25345 = n25343 | n25344 ;
  assign n73700 = ~n24848 ;
  assign n25346 = n73700 & n25345 ;
  assign n73701 = ~n24838 ;
  assign n25347 = x103 & n73701 ;
  assign n73702 = ~n24833 ;
  assign n25348 = n73702 & n25347 ;
  assign n25349 = n24840 | n25348 ;
  assign n25351 = n25346 | n25349 ;
  assign n73703 = ~n24840 ;
  assign n25356 = n73703 & n25351 ;
  assign n25357 = n25354 | n25356 ;
  assign n73704 = ~n24832 ;
  assign n25358 = n73704 & n25357 ;
  assign n73705 = ~n24822 ;
  assign n25359 = x105 & n73705 ;
  assign n73706 = ~n24817 ;
  assign n25360 = n73706 & n25359 ;
  assign n25361 = n24824 | n25360 ;
  assign n25362 = n25358 | n25361 ;
  assign n73707 = ~n24824 ;
  assign n25366 = n73707 & n25362 ;
  assign n25367 = n25365 | n25366 ;
  assign n73708 = ~n24816 ;
  assign n25368 = n73708 & n25367 ;
  assign n73709 = ~n24806 ;
  assign n25369 = x107 & n73709 ;
  assign n73710 = ~n24801 ;
  assign n25370 = n73710 & n25369 ;
  assign n25371 = n24808 | n25370 ;
  assign n25373 = n25368 | n25371 ;
  assign n73711 = ~n24808 ;
  assign n25377 = n73711 & n25373 ;
  assign n25378 = n25376 | n25377 ;
  assign n73712 = ~n24800 ;
  assign n25379 = n73712 & n25378 ;
  assign n73713 = ~n24790 ;
  assign n25380 = x109 & n73713 ;
  assign n73714 = ~n24785 ;
  assign n25381 = n73714 & n25380 ;
  assign n25382 = n24792 | n25381 ;
  assign n25383 = n25379 | n25382 ;
  assign n73715 = ~n24792 ;
  assign n25387 = n73715 & n25383 ;
  assign n25388 = n25386 | n25387 ;
  assign n73716 = ~n24784 ;
  assign n25389 = n73716 & n25388 ;
  assign n73717 = ~n24774 ;
  assign n25390 = x111 & n73717 ;
  assign n73718 = ~n24769 ;
  assign n25391 = n73718 & n25390 ;
  assign n25392 = n24776 | n25391 ;
  assign n25393 = n25389 | n25392 ;
  assign n73719 = ~n24776 ;
  assign n25397 = n73719 & n25393 ;
  assign n25398 = n25396 | n25397 ;
  assign n73720 = ~n24768 ;
  assign n25399 = n73720 & n25398 ;
  assign n73721 = ~n24758 ;
  assign n25400 = x113 & n73721 ;
  assign n73722 = ~n24753 ;
  assign n25401 = n73722 & n25400 ;
  assign n25402 = n24760 | n25401 ;
  assign n25404 = n25399 | n25402 ;
  assign n73723 = ~n24760 ;
  assign n25408 = n73723 & n25404 ;
  assign n25409 = n25407 | n25408 ;
  assign n73724 = ~n24752 ;
  assign n25410 = n73724 & n25409 ;
  assign n73725 = ~n24742 ;
  assign n25411 = x115 & n73725 ;
  assign n73726 = ~n24737 ;
  assign n25412 = n73726 & n25411 ;
  assign n25413 = n24744 | n25412 ;
  assign n25414 = n25410 | n25413 ;
  assign n73727 = ~n24744 ;
  assign n25419 = n73727 & n25414 ;
  assign n25420 = n25417 | n25419 ;
  assign n73728 = ~n24736 ;
  assign n25421 = n73728 & n25420 ;
  assign n73729 = ~n24726 ;
  assign n25422 = x117 & n73729 ;
  assign n73730 = ~n24721 ;
  assign n25423 = n73730 & n25422 ;
  assign n25424 = n24728 | n25423 ;
  assign n25425 = n25421 | n25424 ;
  assign n73731 = ~n24728 ;
  assign n25430 = n73731 & n25425 ;
  assign n25431 = n25428 | n25430 ;
  assign n73732 = ~n24720 ;
  assign n25432 = n73732 & n25431 ;
  assign n73733 = ~n24568 ;
  assign n24572 = n73733 & n24571 ;
  assign n25433 = n23818 | n24571 ;
  assign n73734 = ~n25433 ;
  assign n25434 = n24713 & n73734 ;
  assign n25435 = n24572 | n25434 ;
  assign n25436 = n24577 | n25435 ;
  assign n73735 = ~n23700 ;
  assign n25437 = n73735 & n24577 ;
  assign n73736 = ~n25437 ;
  assign n25438 = n25436 & n73736 ;
  assign n25439 = n73617 & n25438 ;
  assign n138 = ~n24577 ;
  assign n25440 = n138 & n25435 ;
  assign n25441 = n23700 & n24577 ;
  assign n73738 = ~n25441 ;
  assign n25442 = x119 & n73738 ;
  assign n73739 = ~n25440 ;
  assign n25443 = n73739 & n25442 ;
  assign n25444 = n66655 | n25443 ;
  assign n25445 = n25439 | n25444 ;
  assign n25446 = n25432 | n25445 ;
  assign n25447 = n73458 & n25438 ;
  assign n73740 = ~n25447 ;
  assign n25448 = n25446 & n73740 ;
  assign n26352 = n24720 | n25443 ;
  assign n26353 = n25439 | n26352 ;
  assign n73741 = ~n26353 ;
  assign n26354 = n25431 & n73741 ;
  assign n25458 = n73459 & n25145 ;
  assign n73742 = ~n25458 ;
  assign n25459 = x9 & n73742 ;
  assign n25460 = n25151 | n25459 ;
  assign n25461 = x65 & n25460 ;
  assign n73743 = ~n25461 ;
  assign n25462 = n25155 & n73743 ;
  assign n25463 = n25157 | n25462 ;
  assign n25464 = n73627 & n25463 ;
  assign n25465 = n25162 | n25464 ;
  assign n25466 = n73628 & n25465 ;
  assign n25467 = n25168 | n25466 ;
  assign n25468 = n73631 & n25467 ;
  assign n25469 = n25172 | n25468 ;
  assign n25470 = n73632 & n25469 ;
  assign n25471 = n25178 | n25470 ;
  assign n25472 = n73635 & n25471 ;
  assign n25473 = n25182 | n25472 ;
  assign n25474 = n73636 & n25473 ;
  assign n25475 = n25188 | n25474 ;
  assign n25476 = n73639 & n25475 ;
  assign n25477 = n25192 | n25476 ;
  assign n25478 = n73640 & n25477 ;
  assign n25479 = n25198 | n25478 ;
  assign n25480 = n73643 & n25479 ;
  assign n25481 = n25202 | n25480 ;
  assign n25482 = n73644 & n25481 ;
  assign n25483 = n25208 | n25482 ;
  assign n25484 = n73647 & n25483 ;
  assign n25485 = n25212 | n25484 ;
  assign n25486 = n73648 & n25485 ;
  assign n25487 = n25218 | n25486 ;
  assign n25488 = n73651 & n25487 ;
  assign n25489 = n25222 | n25488 ;
  assign n25490 = n73652 & n25489 ;
  assign n25491 = n25228 | n25490 ;
  assign n25492 = n73655 & n25491 ;
  assign n25493 = n25233 | n25492 ;
  assign n25494 = n73656 & n25493 ;
  assign n25495 = n25239 | n25494 ;
  assign n25496 = n73659 & n25495 ;
  assign n25497 = n25243 | n25496 ;
  assign n25498 = n73660 & n25497 ;
  assign n25499 = n25249 | n25498 ;
  assign n25500 = n73663 & n25499 ;
  assign n25501 = n25253 | n25500 ;
  assign n25502 = n73664 & n25501 ;
  assign n25503 = n25259 | n25502 ;
  assign n25504 = n73667 & n25503 ;
  assign n25505 = n25263 | n25504 ;
  assign n25506 = n73668 & n25505 ;
  assign n25507 = n25269 | n25506 ;
  assign n25508 = n73671 & n25507 ;
  assign n25509 = n25273 | n25508 ;
  assign n25510 = n73672 & n25509 ;
  assign n25511 = n25279 | n25510 ;
  assign n25512 = n73675 & n25511 ;
  assign n25513 = n25283 | n25512 ;
  assign n25514 = n73676 & n25513 ;
  assign n25515 = n25289 | n25514 ;
  assign n25516 = n73679 & n25515 ;
  assign n25517 = n25293 | n25516 ;
  assign n25518 = n73680 & n25517 ;
  assign n25519 = n25299 | n25518 ;
  assign n25520 = n73683 & n25519 ;
  assign n25521 = n25303 | n25520 ;
  assign n25522 = n73684 & n25521 ;
  assign n25523 = n25309 | n25522 ;
  assign n25524 = n73687 & n25523 ;
  assign n25525 = n25313 | n25524 ;
  assign n25526 = n73688 & n25525 ;
  assign n25527 = n25319 | n25526 ;
  assign n25528 = n73691 & n25527 ;
  assign n25529 = n25323 | n25528 ;
  assign n25530 = n73692 & n25529 ;
  assign n25531 = n25329 | n25530 ;
  assign n25532 = n73695 & n25531 ;
  assign n25533 = n25333 | n25532 ;
  assign n25534 = n73696 & n25533 ;
  assign n25535 = n25339 | n25534 ;
  assign n25536 = n73699 & n25535 ;
  assign n25537 = n25343 | n25536 ;
  assign n25538 = n73700 & n25537 ;
  assign n25539 = n25349 | n25538 ;
  assign n25540 = n73703 & n25539 ;
  assign n25541 = n25354 | n25540 ;
  assign n25542 = n73704 & n25541 ;
  assign n25543 = n25361 | n25542 ;
  assign n25544 = n73707 & n25543 ;
  assign n25545 = n25365 | n25544 ;
  assign n25546 = n73708 & n25545 ;
  assign n25547 = n25371 | n25546 ;
  assign n25548 = n73711 & n25547 ;
  assign n25549 = n25376 | n25548 ;
  assign n25550 = n73712 & n25549 ;
  assign n25551 = n25382 | n25550 ;
  assign n25552 = n73715 & n25551 ;
  assign n25553 = n25386 | n25552 ;
  assign n25554 = n73716 & n25553 ;
  assign n25555 = n25392 | n25554 ;
  assign n25556 = n73719 & n25555 ;
  assign n25557 = n25396 | n25556 ;
  assign n25558 = n73720 & n25557 ;
  assign n25559 = n25402 | n25558 ;
  assign n25560 = n73723 & n25559 ;
  assign n25561 = n25407 | n25560 ;
  assign n25562 = n73724 & n25561 ;
  assign n25563 = n25413 | n25562 ;
  assign n25564 = n73727 & n25563 ;
  assign n25565 = n25417 | n25564 ;
  assign n25566 = n73728 & n25565 ;
  assign n26037 = n25424 | n25566 ;
  assign n26038 = n73731 & n26037 ;
  assign n26039 = n25428 | n26038 ;
  assign n26040 = n73732 & n26039 ;
  assign n26355 = n25439 | n25443 ;
  assign n73744 = ~n26040 ;
  assign n26356 = n73744 & n26355 ;
  assign n26357 = n26354 | n26356 ;
  assign n137 = ~n25448 ;
  assign n26358 = n137 & n26357 ;
  assign n26359 = n24576 & n25438 ;
  assign n26360 = n25446 & n26359 ;
  assign n26361 = n26358 | n26360 ;
  assign n26367 = n65681 & n26361 ;
  assign n73746 = ~n25430 ;
  assign n25450 = n25428 & n73746 ;
  assign n25429 = n24728 | n25428 ;
  assign n73747 = ~n25429 ;
  assign n25451 = n25425 & n73747 ;
  assign n25452 = n25450 | n25451 ;
  assign n25453 = n137 & n25452 ;
  assign n25454 = n24719 & n73740 ;
  assign n25455 = n25446 & n25454 ;
  assign n25456 = n25453 | n25455 ;
  assign n25457 = n73617 & n25456 ;
  assign n73748 = ~n25566 ;
  assign n25567 = n25424 & n73748 ;
  assign n25568 = n24736 | n25424 ;
  assign n73749 = ~n25568 ;
  assign n25569 = n25420 & n73749 ;
  assign n25570 = n25567 | n25569 ;
  assign n25571 = n137 & n25570 ;
  assign n25572 = n24727 & n73740 ;
  assign n25573 = n25446 & n25572 ;
  assign n25574 = n25571 | n25573 ;
  assign n25575 = n73188 & n25574 ;
  assign n73750 = ~n25419 ;
  assign n25576 = n25417 & n73750 ;
  assign n25418 = n24744 | n25417 ;
  assign n73751 = ~n25418 ;
  assign n25577 = n25414 & n73751 ;
  assign n25578 = n25576 | n25577 ;
  assign n25579 = n137 & n25578 ;
  assign n25580 = n24735 & n73740 ;
  assign n25581 = n25446 & n25580 ;
  assign n25582 = n25579 | n25581 ;
  assign n25583 = n73177 & n25582 ;
  assign n73752 = ~n25562 ;
  assign n25584 = n25413 & n73752 ;
  assign n25585 = n24752 | n25413 ;
  assign n73753 = ~n25585 ;
  assign n25586 = n25409 & n73753 ;
  assign n25587 = n25584 | n25586 ;
  assign n25588 = n137 & n25587 ;
  assign n25589 = n24743 & n73740 ;
  assign n25590 = n25446 & n25589 ;
  assign n25591 = n25588 | n25590 ;
  assign n25592 = n72752 & n25591 ;
  assign n73754 = ~n25408 ;
  assign n25593 = n25407 & n73754 ;
  assign n25594 = n24760 | n25407 ;
  assign n73755 = ~n25594 ;
  assign n25595 = n25559 & n73755 ;
  assign n25596 = n25593 | n25595 ;
  assign n25597 = n137 & n25596 ;
  assign n25598 = n24751 & n73740 ;
  assign n25599 = n25446 & n25598 ;
  assign n25600 = n25597 | n25599 ;
  assign n25601 = n72393 & n25600 ;
  assign n73756 = ~n25558 ;
  assign n25602 = n25402 & n73756 ;
  assign n25403 = n24768 | n25402 ;
  assign n73757 = ~n25403 ;
  assign n25603 = n73757 & n25557 ;
  assign n25604 = n25602 | n25603 ;
  assign n25605 = n137 & n25604 ;
  assign n25606 = n24759 & n73740 ;
  assign n25607 = n25446 & n25606 ;
  assign n25608 = n25605 | n25607 ;
  assign n25609 = n72385 & n25608 ;
  assign n73758 = ~n25397 ;
  assign n25610 = n25396 & n73758 ;
  assign n25611 = n24776 | n25396 ;
  assign n73759 = ~n25611 ;
  assign n25612 = n25555 & n73759 ;
  assign n25613 = n25610 | n25612 ;
  assign n25614 = n137 & n25613 ;
  assign n25615 = n24767 & n73740 ;
  assign n25616 = n25446 & n25615 ;
  assign n25617 = n25614 | n25616 ;
  assign n25618 = n72025 & n25617 ;
  assign n73760 = ~n25554 ;
  assign n25619 = n25392 & n73760 ;
  assign n25620 = n24784 | n25392 ;
  assign n73761 = ~n25620 ;
  assign n25621 = n25388 & n73761 ;
  assign n25622 = n25619 | n25621 ;
  assign n25623 = n137 & n25622 ;
  assign n25624 = n24775 & n73740 ;
  assign n25625 = n25446 & n25624 ;
  assign n25626 = n25623 | n25625 ;
  assign n25627 = n71645 & n25626 ;
  assign n73762 = ~n25387 ;
  assign n25628 = n25386 & n73762 ;
  assign n25629 = n24792 | n25386 ;
  assign n73763 = ~n25629 ;
  assign n25630 = n25551 & n73763 ;
  assign n25631 = n25628 | n25630 ;
  assign n25632 = n137 & n25631 ;
  assign n25633 = n24783 & n73740 ;
  assign n25634 = n25446 & n25633 ;
  assign n25635 = n25632 | n25634 ;
  assign n25636 = n71633 & n25635 ;
  assign n73764 = ~n25550 ;
  assign n25637 = n25382 & n73764 ;
  assign n25638 = n24800 | n25382 ;
  assign n73765 = ~n25638 ;
  assign n25639 = n25378 & n73765 ;
  assign n25640 = n25637 | n25639 ;
  assign n25641 = n137 & n25640 ;
  assign n25642 = n24791 & n73740 ;
  assign n25643 = n25446 & n25642 ;
  assign n25644 = n25641 | n25643 ;
  assign n25645 = n71253 & n25644 ;
  assign n73766 = ~n25377 ;
  assign n25646 = n25376 & n73766 ;
  assign n25647 = n24808 | n25376 ;
  assign n73767 = ~n25647 ;
  assign n25648 = n25547 & n73767 ;
  assign n25649 = n25646 | n25648 ;
  assign n25650 = n137 & n25649 ;
  assign n25651 = n24799 & n73740 ;
  assign n25652 = n25446 & n25651 ;
  assign n25653 = n25650 | n25652 ;
  assign n25654 = n70935 & n25653 ;
  assign n73768 = ~n25546 ;
  assign n25655 = n25371 & n73768 ;
  assign n25372 = n24816 | n25371 ;
  assign n73769 = ~n25372 ;
  assign n25656 = n73769 & n25545 ;
  assign n25657 = n25655 | n25656 ;
  assign n25658 = n137 & n25657 ;
  assign n25659 = n24807 & n73740 ;
  assign n25660 = n25446 & n25659 ;
  assign n25661 = n25658 | n25660 ;
  assign n25662 = n70927 & n25661 ;
  assign n73770 = ~n25366 ;
  assign n25663 = n25365 & n73770 ;
  assign n25664 = n24824 | n25365 ;
  assign n73771 = ~n25664 ;
  assign n25665 = n25543 & n73771 ;
  assign n25666 = n25663 | n25665 ;
  assign n25667 = n137 & n25666 ;
  assign n25668 = n24815 & n73740 ;
  assign n25669 = n25446 & n25668 ;
  assign n25670 = n25667 | n25669 ;
  assign n25671 = n70609 & n25670 ;
  assign n73772 = ~n25542 ;
  assign n25672 = n25361 & n73772 ;
  assign n25673 = n24832 | n25361 ;
  assign n73773 = ~n25673 ;
  assign n25674 = n25357 & n73773 ;
  assign n25675 = n25672 | n25674 ;
  assign n25676 = n137 & n25675 ;
  assign n25677 = n24823 & n73740 ;
  assign n25678 = n25446 & n25677 ;
  assign n25679 = n25676 | n25678 ;
  assign n25680 = n70276 & n25679 ;
  assign n73774 = ~n25356 ;
  assign n25681 = n25354 & n73774 ;
  assign n25355 = n24840 | n25354 ;
  assign n73775 = ~n25355 ;
  assign n25682 = n25351 & n73775 ;
  assign n25683 = n25681 | n25682 ;
  assign n25684 = n137 & n25683 ;
  assign n25685 = n24831 & n73740 ;
  assign n25686 = n25446 & n25685 ;
  assign n25687 = n25684 | n25686 ;
  assign n25688 = n70176 & n25687 ;
  assign n73776 = ~n25538 ;
  assign n25689 = n25349 & n73776 ;
  assign n25350 = n24848 | n25349 ;
  assign n73777 = ~n25350 ;
  assign n25690 = n73777 & n25537 ;
  assign n25691 = n25689 | n25690 ;
  assign n25692 = n137 & n25691 ;
  assign n25693 = n24839 & n73740 ;
  assign n25694 = n25446 & n25693 ;
  assign n25695 = n25692 | n25694 ;
  assign n25696 = n69857 & n25695 ;
  assign n73778 = ~n25344 ;
  assign n25697 = n25343 & n73778 ;
  assign n25698 = n24856 | n25343 ;
  assign n73779 = ~n25698 ;
  assign n25699 = n25535 & n73779 ;
  assign n25700 = n25697 | n25699 ;
  assign n25701 = n137 & n25700 ;
  assign n25702 = n24847 & n73740 ;
  assign n25703 = n25446 & n25702 ;
  assign n25704 = n25701 | n25703 ;
  assign n25705 = n69656 & n25704 ;
  assign n73780 = ~n25534 ;
  assign n25706 = n25339 & n73780 ;
  assign n25707 = n24864 | n25339 ;
  assign n73781 = ~n25707 ;
  assign n25708 = n25335 & n73781 ;
  assign n25709 = n25706 | n25708 ;
  assign n25710 = n137 & n25709 ;
  assign n25711 = n24855 & n73740 ;
  assign n25712 = n25446 & n25711 ;
  assign n25713 = n25710 | n25712 ;
  assign n25714 = n69528 & n25713 ;
  assign n73782 = ~n25334 ;
  assign n25715 = n25333 & n73782 ;
  assign n25716 = n24872 | n25333 ;
  assign n73783 = ~n25716 ;
  assign n25717 = n25531 & n73783 ;
  assign n25718 = n25715 | n25717 ;
  assign n25719 = n137 & n25718 ;
  assign n25720 = n24863 & n73740 ;
  assign n25721 = n25446 & n25720 ;
  assign n25722 = n25719 | n25721 ;
  assign n25723 = n69261 & n25722 ;
  assign n73784 = ~n25530 ;
  assign n25724 = n25329 & n73784 ;
  assign n25725 = n24880 | n25329 ;
  assign n73785 = ~n25725 ;
  assign n25726 = n25325 & n73785 ;
  assign n25727 = n25724 | n25726 ;
  assign n25728 = n137 & n25727 ;
  assign n25729 = n24871 & n73740 ;
  assign n25730 = n25446 & n25729 ;
  assign n25731 = n25728 | n25730 ;
  assign n25732 = n69075 & n25731 ;
  assign n73786 = ~n25324 ;
  assign n25733 = n25323 & n73786 ;
  assign n25734 = n24888 | n25323 ;
  assign n73787 = ~n25734 ;
  assign n25735 = n25527 & n73787 ;
  assign n25736 = n25733 | n25735 ;
  assign n25737 = n137 & n25736 ;
  assign n25738 = n24879 & n73740 ;
  assign n25739 = n25446 & n25738 ;
  assign n25740 = n25737 | n25739 ;
  assign n25741 = n68993 & n25740 ;
  assign n73788 = ~n25526 ;
  assign n25742 = n25319 & n73788 ;
  assign n25743 = n24896 | n25319 ;
  assign n73789 = ~n25743 ;
  assign n25744 = n25315 & n73789 ;
  assign n25745 = n25742 | n25744 ;
  assign n25746 = n137 & n25745 ;
  assign n25747 = n24887 & n73740 ;
  assign n25748 = n25446 & n25747 ;
  assign n25749 = n25746 | n25748 ;
  assign n25750 = n68716 & n25749 ;
  assign n73790 = ~n25314 ;
  assign n25751 = n25313 & n73790 ;
  assign n25752 = n24904 | n25313 ;
  assign n73791 = ~n25752 ;
  assign n25753 = n25523 & n73791 ;
  assign n25754 = n25751 | n25753 ;
  assign n25755 = n137 & n25754 ;
  assign n25756 = n24895 & n73740 ;
  assign n25757 = n25446 & n25756 ;
  assign n25758 = n25755 | n25757 ;
  assign n25759 = n68545 & n25758 ;
  assign n73792 = ~n25522 ;
  assign n25760 = n25309 & n73792 ;
  assign n25761 = n24912 | n25309 ;
  assign n73793 = ~n25761 ;
  assign n25762 = n25305 & n73793 ;
  assign n25763 = n25760 | n25762 ;
  assign n25764 = n137 & n25763 ;
  assign n25765 = n24903 & n73740 ;
  assign n25766 = n25446 & n25765 ;
  assign n25767 = n25764 | n25766 ;
  assign n25768 = n68438 & n25767 ;
  assign n73794 = ~n25304 ;
  assign n25769 = n25303 & n73794 ;
  assign n25770 = n24920 | n25303 ;
  assign n73795 = ~n25770 ;
  assign n25771 = n25519 & n73795 ;
  assign n25772 = n25769 | n25771 ;
  assign n25773 = n137 & n25772 ;
  assign n25774 = n24911 & n73740 ;
  assign n25775 = n25446 & n25774 ;
  assign n25776 = n25773 | n25775 ;
  assign n25777 = n68214 & n25776 ;
  assign n73796 = ~n25518 ;
  assign n25778 = n25299 & n73796 ;
  assign n25779 = n24928 | n25299 ;
  assign n73797 = ~n25779 ;
  assign n25780 = n25295 & n73797 ;
  assign n25781 = n25778 | n25780 ;
  assign n25782 = n137 & n25781 ;
  assign n25783 = n24919 & n73740 ;
  assign n25784 = n25446 & n25783 ;
  assign n25785 = n25782 | n25784 ;
  assign n25786 = n68058 & n25785 ;
  assign n73798 = ~n25294 ;
  assign n25787 = n25293 & n73798 ;
  assign n25788 = n24936 | n25293 ;
  assign n73799 = ~n25788 ;
  assign n25789 = n25515 & n73799 ;
  assign n25790 = n25787 | n25789 ;
  assign n25791 = n137 & n25790 ;
  assign n25792 = n24927 & n73740 ;
  assign n25793 = n25446 & n25792 ;
  assign n25794 = n25791 | n25793 ;
  assign n25795 = n67986 & n25794 ;
  assign n73800 = ~n25514 ;
  assign n25796 = n25289 & n73800 ;
  assign n25797 = n24944 | n25289 ;
  assign n73801 = ~n25797 ;
  assign n25798 = n25285 & n73801 ;
  assign n25799 = n25796 | n25798 ;
  assign n25800 = n137 & n25799 ;
  assign n25801 = n24935 & n73740 ;
  assign n25802 = n25446 & n25801 ;
  assign n25803 = n25800 | n25802 ;
  assign n25804 = n67763 & n25803 ;
  assign n73802 = ~n25284 ;
  assign n25805 = n25283 & n73802 ;
  assign n25806 = n24952 | n25283 ;
  assign n73803 = ~n25806 ;
  assign n25807 = n25511 & n73803 ;
  assign n25808 = n25805 | n25807 ;
  assign n25809 = n137 & n25808 ;
  assign n25810 = n24943 & n73740 ;
  assign n25811 = n25446 & n25810 ;
  assign n25812 = n25809 | n25811 ;
  assign n25813 = n67622 & n25812 ;
  assign n73804 = ~n25510 ;
  assign n25814 = n25279 & n73804 ;
  assign n25815 = n24960 | n25279 ;
  assign n73805 = ~n25815 ;
  assign n25816 = n25275 & n73805 ;
  assign n25817 = n25814 | n25816 ;
  assign n25818 = n137 & n25817 ;
  assign n25819 = n24951 & n73740 ;
  assign n25820 = n25446 & n25819 ;
  assign n25821 = n25818 | n25820 ;
  assign n25822 = n67531 & n25821 ;
  assign n73806 = ~n25274 ;
  assign n25823 = n25273 & n73806 ;
  assign n25824 = n24968 | n25273 ;
  assign n73807 = ~n25824 ;
  assign n25825 = n25507 & n73807 ;
  assign n25826 = n25823 | n25825 ;
  assign n25827 = n137 & n25826 ;
  assign n25828 = n24959 & n73740 ;
  assign n25829 = n25446 & n25828 ;
  assign n25830 = n25827 | n25829 ;
  assign n25831 = n67348 & n25830 ;
  assign n73808 = ~n25506 ;
  assign n25832 = n25269 & n73808 ;
  assign n25833 = n24976 | n25269 ;
  assign n73809 = ~n25833 ;
  assign n25834 = n25265 & n73809 ;
  assign n25835 = n25832 | n25834 ;
  assign n25836 = n137 & n25835 ;
  assign n25837 = n24967 & n73740 ;
  assign n25838 = n25446 & n25837 ;
  assign n25839 = n25836 | n25838 ;
  assign n25840 = n67222 & n25839 ;
  assign n73810 = ~n25264 ;
  assign n25841 = n25263 & n73810 ;
  assign n25842 = n24984 | n25263 ;
  assign n73811 = ~n25842 ;
  assign n25843 = n25503 & n73811 ;
  assign n25844 = n25841 | n25843 ;
  assign n25845 = n137 & n25844 ;
  assign n25846 = n24975 & n73740 ;
  assign n25847 = n25446 & n25846 ;
  assign n25848 = n25845 | n25847 ;
  assign n25849 = n67164 & n25848 ;
  assign n73812 = ~n25502 ;
  assign n25850 = n25259 & n73812 ;
  assign n25851 = n24992 | n25259 ;
  assign n73813 = ~n25851 ;
  assign n25852 = n25255 & n73813 ;
  assign n25853 = n25850 | n25852 ;
  assign n25854 = n137 & n25853 ;
  assign n25855 = n24983 & n73740 ;
  assign n25856 = n25446 & n25855 ;
  assign n25857 = n25854 | n25856 ;
  assign n25858 = n66979 & n25857 ;
  assign n73814 = ~n25254 ;
  assign n25859 = n25253 & n73814 ;
  assign n25860 = n25000 | n25253 ;
  assign n73815 = ~n25860 ;
  assign n25861 = n25499 & n73815 ;
  assign n25862 = n25859 | n25861 ;
  assign n25863 = n137 & n25862 ;
  assign n25864 = n24991 & n73740 ;
  assign n25865 = n25446 & n25864 ;
  assign n25866 = n25863 | n25865 ;
  assign n25867 = n66868 & n25866 ;
  assign n73816 = ~n25498 ;
  assign n25868 = n25249 & n73816 ;
  assign n25869 = n25008 | n25249 ;
  assign n73817 = ~n25869 ;
  assign n25870 = n25245 & n73817 ;
  assign n25871 = n25868 | n25870 ;
  assign n25872 = n137 & n25871 ;
  assign n25873 = n24999 & n73740 ;
  assign n25874 = n25446 & n25873 ;
  assign n25875 = n25872 | n25874 ;
  assign n25876 = n66797 & n25875 ;
  assign n73818 = ~n25244 ;
  assign n25877 = n25243 & n73818 ;
  assign n25878 = n25016 | n25243 ;
  assign n73819 = ~n25878 ;
  assign n25879 = n25495 & n73819 ;
  assign n25880 = n25877 | n25879 ;
  assign n25881 = n137 & n25880 ;
  assign n25882 = n25007 & n73740 ;
  assign n25883 = n25446 & n25882 ;
  assign n25884 = n25881 | n25883 ;
  assign n25885 = n66654 & n25884 ;
  assign n73820 = ~n25494 ;
  assign n25886 = n25239 & n73820 ;
  assign n25887 = n25024 | n25239 ;
  assign n73821 = ~n25887 ;
  assign n25888 = n25235 & n73821 ;
  assign n25889 = n25886 | n25888 ;
  assign n25890 = n137 & n25889 ;
  assign n25891 = n25015 & n73740 ;
  assign n25892 = n25446 & n25891 ;
  assign n25893 = n25890 | n25892 ;
  assign n25894 = n66560 & n25893 ;
  assign n73822 = ~n25234 ;
  assign n25895 = n25233 & n73822 ;
  assign n25896 = n25032 | n25233 ;
  assign n73823 = ~n25896 ;
  assign n25897 = n25491 & n73823 ;
  assign n25898 = n25895 | n25897 ;
  assign n25899 = n137 & n25898 ;
  assign n25900 = n25023 & n73740 ;
  assign n25901 = n25446 & n25900 ;
  assign n25902 = n25899 | n25901 ;
  assign n25903 = n66505 & n25902 ;
  assign n73824 = ~n25490 ;
  assign n25904 = n25228 & n73824 ;
  assign n25229 = n25040 | n25228 ;
  assign n73825 = ~n25229 ;
  assign n25905 = n73825 & n25489 ;
  assign n25906 = n25904 | n25905 ;
  assign n25907 = n137 & n25906 ;
  assign n25908 = n25031 & n73740 ;
  assign n25909 = n25446 & n25908 ;
  assign n25910 = n25907 | n25909 ;
  assign n25911 = n66379 & n25910 ;
  assign n73826 = ~n25223 ;
  assign n25912 = n25222 & n73826 ;
  assign n25913 = n25048 | n25222 ;
  assign n73827 = ~n25913 ;
  assign n25914 = n25487 & n73827 ;
  assign n25915 = n25912 | n25914 ;
  assign n25916 = n137 & n25915 ;
  assign n25917 = n25039 & n73740 ;
  assign n25918 = n25446 & n25917 ;
  assign n25919 = n25916 | n25918 ;
  assign n25920 = n66299 & n25919 ;
  assign n73828 = ~n25486 ;
  assign n25921 = n25218 & n73828 ;
  assign n25922 = n25056 | n25218 ;
  assign n73829 = ~n25922 ;
  assign n25923 = n25214 & n73829 ;
  assign n25924 = n25921 | n25923 ;
  assign n25925 = n137 & n25924 ;
  assign n25926 = n25047 & n73740 ;
  assign n25927 = n25446 & n25926 ;
  assign n25928 = n25925 | n25927 ;
  assign n25929 = n66244 & n25928 ;
  assign n73830 = ~n25213 ;
  assign n25930 = n25212 & n73830 ;
  assign n25931 = n25064 | n25212 ;
  assign n73831 = ~n25931 ;
  assign n25932 = n25483 & n73831 ;
  assign n25933 = n25930 | n25932 ;
  assign n25934 = n137 & n25933 ;
  assign n25935 = n25055 & n73740 ;
  assign n25936 = n25446 & n25935 ;
  assign n25937 = n25934 | n25936 ;
  assign n25938 = n66145 & n25937 ;
  assign n73832 = ~n25482 ;
  assign n25939 = n25208 & n73832 ;
  assign n25940 = n25072 | n25208 ;
  assign n73833 = ~n25940 ;
  assign n25941 = n25204 & n73833 ;
  assign n25942 = n25939 | n25941 ;
  assign n25943 = n137 & n25942 ;
  assign n25944 = n25063 & n73740 ;
  assign n25945 = n25446 & n25944 ;
  assign n25946 = n25943 | n25945 ;
  assign n25947 = n66081 & n25946 ;
  assign n73834 = ~n25203 ;
  assign n25948 = n25202 & n73834 ;
  assign n25949 = n25080 | n25202 ;
  assign n73835 = ~n25949 ;
  assign n25950 = n25479 & n73835 ;
  assign n25951 = n25948 | n25950 ;
  assign n25952 = n137 & n25951 ;
  assign n25953 = n25071 & n73740 ;
  assign n25954 = n25446 & n25953 ;
  assign n25955 = n25952 | n25954 ;
  assign n25956 = n66043 & n25955 ;
  assign n73836 = ~n25478 ;
  assign n25957 = n25198 & n73836 ;
  assign n25958 = n25088 | n25198 ;
  assign n73837 = ~n25958 ;
  assign n25959 = n25194 & n73837 ;
  assign n25960 = n25957 | n25959 ;
  assign n25961 = n137 & n25960 ;
  assign n25962 = n25079 & n73740 ;
  assign n25963 = n25446 & n25962 ;
  assign n25964 = n25961 | n25963 ;
  assign n25965 = n65960 & n25964 ;
  assign n73838 = ~n25193 ;
  assign n25966 = n25192 & n73838 ;
  assign n25967 = n25096 | n25192 ;
  assign n73839 = ~n25967 ;
  assign n25968 = n25475 & n73839 ;
  assign n25969 = n25966 | n25968 ;
  assign n25970 = n137 & n25969 ;
  assign n25971 = n25087 & n73740 ;
  assign n25972 = n25446 & n25971 ;
  assign n25973 = n25970 | n25972 ;
  assign n25974 = n65909 & n25973 ;
  assign n73840 = ~n25474 ;
  assign n25975 = n25188 & n73840 ;
  assign n25976 = n25105 | n25188 ;
  assign n73841 = ~n25976 ;
  assign n25977 = n25184 & n73841 ;
  assign n25978 = n25975 | n25977 ;
  assign n25979 = n137 & n25978 ;
  assign n25980 = n25095 & n73740 ;
  assign n25981 = n25446 & n25980 ;
  assign n25982 = n25979 | n25981 ;
  assign n25983 = n65877 & n25982 ;
  assign n73842 = ~n25183 ;
  assign n25984 = n25182 & n73842 ;
  assign n25985 = n25114 | n25182 ;
  assign n73843 = ~n25985 ;
  assign n25986 = n25471 & n73843 ;
  assign n25987 = n25984 | n25986 ;
  assign n25988 = n137 & n25987 ;
  assign n25989 = n25104 & n73740 ;
  assign n25990 = n25446 & n25989 ;
  assign n25991 = n25988 | n25990 ;
  assign n25992 = n65820 & n25991 ;
  assign n73844 = ~n25470 ;
  assign n25993 = n25178 & n73844 ;
  assign n25994 = n25122 | n25178 ;
  assign n73845 = ~n25994 ;
  assign n25995 = n25174 & n73845 ;
  assign n25996 = n25993 | n25995 ;
  assign n25997 = n137 & n25996 ;
  assign n25998 = n25113 & n73740 ;
  assign n25999 = n25446 & n25998 ;
  assign n26000 = n25997 | n25999 ;
  assign n26001 = n65791 & n26000 ;
  assign n73846 = ~n25173 ;
  assign n26003 = n25172 & n73846 ;
  assign n26002 = n25131 | n25172 ;
  assign n73847 = ~n26002 ;
  assign n26004 = n25169 & n73847 ;
  assign n26005 = n26003 | n26004 ;
  assign n26006 = n137 & n26005 ;
  assign n26007 = n25121 & n73740 ;
  assign n26008 = n25446 & n26007 ;
  assign n26009 = n26006 | n26008 ;
  assign n26010 = n65772 & n26009 ;
  assign n73848 = ~n25466 ;
  assign n26012 = n25168 & n73848 ;
  assign n26011 = n25139 | n25168 ;
  assign n73849 = ~n26011 ;
  assign n26013 = n25465 & n73849 ;
  assign n26014 = n26012 | n26013 ;
  assign n26015 = n137 & n26014 ;
  assign n26016 = n25130 & n73740 ;
  assign n26017 = n25446 & n26016 ;
  assign n26018 = n26015 | n26017 ;
  assign n26019 = n65746 & n26018 ;
  assign n73850 = ~n25163 ;
  assign n26021 = n25162 & n73850 ;
  assign n26020 = n25159 | n25162 ;
  assign n73851 = ~n26020 ;
  assign n26022 = n25158 & n73851 ;
  assign n26023 = n26021 | n26022 ;
  assign n26024 = n137 & n26023 ;
  assign n26025 = n25138 & n73740 ;
  assign n26026 = n25446 & n26025 ;
  assign n26027 = n26024 | n26026 ;
  assign n26028 = n65721 & n26027 ;
  assign n26029 = n25155 & n25157 ;
  assign n26030 = n73625 & n26029 ;
  assign n73852 = ~n26030 ;
  assign n26031 = n25158 & n73852 ;
  assign n26032 = n137 & n26031 ;
  assign n26033 = n25152 & n73740 ;
  assign n26034 = n25446 & n26033 ;
  assign n26035 = n26032 | n26034 ;
  assign n26036 = n65686 & n26035 ;
  assign n25449 = n25157 & n137 ;
  assign n26045 = x64 & n137 ;
  assign n73853 = ~n26045 ;
  assign n26046 = x8 & n73853 ;
  assign n26047 = n25449 | n26046 ;
  assign n26049 = x65 & n26047 ;
  assign n26041 = n25445 | n26040 ;
  assign n26042 = n73740 & n26041 ;
  assign n73854 = ~n26042 ;
  assign n26043 = x64 & n73854 ;
  assign n73855 = ~n26043 ;
  assign n26044 = x8 & n73855 ;
  assign n26048 = x65 | n25449 ;
  assign n26050 = n26044 | n26048 ;
  assign n73856 = ~n26049 ;
  assign n26051 = n73856 & n26050 ;
  assign n73857 = ~x7 ;
  assign n26052 = n73857 & x64 ;
  assign n26053 = n26051 | n26052 ;
  assign n26054 = n65670 & n26047 ;
  assign n73858 = ~n26054 ;
  assign n26055 = n26053 & n73858 ;
  assign n73859 = ~n26034 ;
  assign n26056 = x66 & n73859 ;
  assign n73860 = ~n26032 ;
  assign n26057 = n73860 & n26056 ;
  assign n26058 = n26036 | n26057 ;
  assign n26059 = n26055 | n26058 ;
  assign n73861 = ~n26036 ;
  assign n26060 = n73861 & n26059 ;
  assign n73862 = ~n26026 ;
  assign n26061 = x67 & n73862 ;
  assign n73863 = ~n26024 ;
  assign n26062 = n73863 & n26061 ;
  assign n26063 = n26028 | n26062 ;
  assign n26064 = n26060 | n26063 ;
  assign n73864 = ~n26028 ;
  assign n26065 = n73864 & n26064 ;
  assign n73865 = ~n26017 ;
  assign n26066 = x68 & n73865 ;
  assign n73866 = ~n26015 ;
  assign n26067 = n73866 & n26066 ;
  assign n26068 = n26019 | n26067 ;
  assign n26069 = n26065 | n26068 ;
  assign n73867 = ~n26019 ;
  assign n26070 = n73867 & n26069 ;
  assign n73868 = ~n26008 ;
  assign n26071 = x69 & n73868 ;
  assign n73869 = ~n26006 ;
  assign n26072 = n73869 & n26071 ;
  assign n26073 = n26010 | n26072 ;
  assign n26075 = n26070 | n26073 ;
  assign n73870 = ~n26010 ;
  assign n26076 = n73870 & n26075 ;
  assign n73871 = ~n25999 ;
  assign n26077 = x70 & n73871 ;
  assign n73872 = ~n25997 ;
  assign n26078 = n73872 & n26077 ;
  assign n26079 = n26001 | n26078 ;
  assign n26080 = n26076 | n26079 ;
  assign n73873 = ~n26001 ;
  assign n26081 = n73873 & n26080 ;
  assign n73874 = ~n25990 ;
  assign n26082 = x71 & n73874 ;
  assign n73875 = ~n25988 ;
  assign n26083 = n73875 & n26082 ;
  assign n26084 = n25992 | n26083 ;
  assign n26086 = n26081 | n26084 ;
  assign n73876 = ~n25992 ;
  assign n26087 = n73876 & n26086 ;
  assign n73877 = ~n25981 ;
  assign n26088 = x72 & n73877 ;
  assign n73878 = ~n25979 ;
  assign n26089 = n73878 & n26088 ;
  assign n26090 = n25983 | n26089 ;
  assign n26091 = n26087 | n26090 ;
  assign n73879 = ~n25983 ;
  assign n26092 = n73879 & n26091 ;
  assign n73880 = ~n25972 ;
  assign n26093 = x73 & n73880 ;
  assign n73881 = ~n25970 ;
  assign n26094 = n73881 & n26093 ;
  assign n26095 = n25974 | n26094 ;
  assign n26097 = n26092 | n26095 ;
  assign n73882 = ~n25974 ;
  assign n26098 = n73882 & n26097 ;
  assign n73883 = ~n25963 ;
  assign n26099 = x74 & n73883 ;
  assign n73884 = ~n25961 ;
  assign n26100 = n73884 & n26099 ;
  assign n26101 = n25965 | n26100 ;
  assign n26102 = n26098 | n26101 ;
  assign n73885 = ~n25965 ;
  assign n26103 = n73885 & n26102 ;
  assign n73886 = ~n25954 ;
  assign n26104 = x75 & n73886 ;
  assign n73887 = ~n25952 ;
  assign n26105 = n73887 & n26104 ;
  assign n26106 = n25956 | n26105 ;
  assign n26108 = n26103 | n26106 ;
  assign n73888 = ~n25956 ;
  assign n26109 = n73888 & n26108 ;
  assign n73889 = ~n25945 ;
  assign n26110 = x76 & n73889 ;
  assign n73890 = ~n25943 ;
  assign n26111 = n73890 & n26110 ;
  assign n26112 = n25947 | n26111 ;
  assign n26113 = n26109 | n26112 ;
  assign n73891 = ~n25947 ;
  assign n26114 = n73891 & n26113 ;
  assign n73892 = ~n25936 ;
  assign n26115 = x77 & n73892 ;
  assign n73893 = ~n25934 ;
  assign n26116 = n73893 & n26115 ;
  assign n26117 = n25938 | n26116 ;
  assign n26119 = n26114 | n26117 ;
  assign n73894 = ~n25938 ;
  assign n26120 = n73894 & n26119 ;
  assign n73895 = ~n25927 ;
  assign n26121 = x78 & n73895 ;
  assign n73896 = ~n25925 ;
  assign n26122 = n73896 & n26121 ;
  assign n26123 = n25929 | n26122 ;
  assign n26124 = n26120 | n26123 ;
  assign n73897 = ~n25929 ;
  assign n26125 = n73897 & n26124 ;
  assign n73898 = ~n25918 ;
  assign n26126 = x79 & n73898 ;
  assign n73899 = ~n25916 ;
  assign n26127 = n73899 & n26126 ;
  assign n26128 = n25920 | n26127 ;
  assign n26130 = n26125 | n26128 ;
  assign n73900 = ~n25920 ;
  assign n26131 = n73900 & n26130 ;
  assign n73901 = ~n25909 ;
  assign n26132 = x80 & n73901 ;
  assign n73902 = ~n25907 ;
  assign n26133 = n73902 & n26132 ;
  assign n26134 = n25911 | n26133 ;
  assign n26135 = n26131 | n26134 ;
  assign n73903 = ~n25911 ;
  assign n26136 = n73903 & n26135 ;
  assign n73904 = ~n25901 ;
  assign n26137 = x81 & n73904 ;
  assign n73905 = ~n25899 ;
  assign n26138 = n73905 & n26137 ;
  assign n26139 = n25903 | n26138 ;
  assign n26141 = n26136 | n26139 ;
  assign n73906 = ~n25903 ;
  assign n26142 = n73906 & n26141 ;
  assign n73907 = ~n25892 ;
  assign n26143 = x82 & n73907 ;
  assign n73908 = ~n25890 ;
  assign n26144 = n73908 & n26143 ;
  assign n26145 = n25894 | n26144 ;
  assign n26146 = n26142 | n26145 ;
  assign n73909 = ~n25894 ;
  assign n26147 = n73909 & n26146 ;
  assign n73910 = ~n25883 ;
  assign n26148 = x83 & n73910 ;
  assign n73911 = ~n25881 ;
  assign n26149 = n73911 & n26148 ;
  assign n26150 = n25885 | n26149 ;
  assign n26152 = n26147 | n26150 ;
  assign n73912 = ~n25885 ;
  assign n26153 = n73912 & n26152 ;
  assign n73913 = ~n25874 ;
  assign n26154 = x84 & n73913 ;
  assign n73914 = ~n25872 ;
  assign n26155 = n73914 & n26154 ;
  assign n26156 = n25876 | n26155 ;
  assign n26157 = n26153 | n26156 ;
  assign n73915 = ~n25876 ;
  assign n26158 = n73915 & n26157 ;
  assign n73916 = ~n25865 ;
  assign n26159 = x85 & n73916 ;
  assign n73917 = ~n25863 ;
  assign n26160 = n73917 & n26159 ;
  assign n26161 = n25867 | n26160 ;
  assign n26163 = n26158 | n26161 ;
  assign n73918 = ~n25867 ;
  assign n26164 = n73918 & n26163 ;
  assign n73919 = ~n25856 ;
  assign n26165 = x86 & n73919 ;
  assign n73920 = ~n25854 ;
  assign n26166 = n73920 & n26165 ;
  assign n26167 = n25858 | n26166 ;
  assign n26168 = n26164 | n26167 ;
  assign n73921 = ~n25858 ;
  assign n26169 = n73921 & n26168 ;
  assign n73922 = ~n25847 ;
  assign n26170 = x87 & n73922 ;
  assign n73923 = ~n25845 ;
  assign n26171 = n73923 & n26170 ;
  assign n26172 = n25849 | n26171 ;
  assign n26174 = n26169 | n26172 ;
  assign n73924 = ~n25849 ;
  assign n26175 = n73924 & n26174 ;
  assign n73925 = ~n25838 ;
  assign n26176 = x88 & n73925 ;
  assign n73926 = ~n25836 ;
  assign n26177 = n73926 & n26176 ;
  assign n26178 = n25840 | n26177 ;
  assign n26179 = n26175 | n26178 ;
  assign n73927 = ~n25840 ;
  assign n26180 = n73927 & n26179 ;
  assign n73928 = ~n25829 ;
  assign n26181 = x89 & n73928 ;
  assign n73929 = ~n25827 ;
  assign n26182 = n73929 & n26181 ;
  assign n26183 = n25831 | n26182 ;
  assign n26185 = n26180 | n26183 ;
  assign n73930 = ~n25831 ;
  assign n26186 = n73930 & n26185 ;
  assign n73931 = ~n25820 ;
  assign n26187 = x90 & n73931 ;
  assign n73932 = ~n25818 ;
  assign n26188 = n73932 & n26187 ;
  assign n26189 = n25822 | n26188 ;
  assign n26190 = n26186 | n26189 ;
  assign n73933 = ~n25822 ;
  assign n26191 = n73933 & n26190 ;
  assign n73934 = ~n25811 ;
  assign n26192 = x91 & n73934 ;
  assign n73935 = ~n25809 ;
  assign n26193 = n73935 & n26192 ;
  assign n26194 = n25813 | n26193 ;
  assign n26196 = n26191 | n26194 ;
  assign n73936 = ~n25813 ;
  assign n26197 = n73936 & n26196 ;
  assign n73937 = ~n25802 ;
  assign n26198 = x92 & n73937 ;
  assign n73938 = ~n25800 ;
  assign n26199 = n73938 & n26198 ;
  assign n26200 = n25804 | n26199 ;
  assign n26201 = n26197 | n26200 ;
  assign n73939 = ~n25804 ;
  assign n26202 = n73939 & n26201 ;
  assign n73940 = ~n25793 ;
  assign n26203 = x93 & n73940 ;
  assign n73941 = ~n25791 ;
  assign n26204 = n73941 & n26203 ;
  assign n26205 = n25795 | n26204 ;
  assign n26207 = n26202 | n26205 ;
  assign n73942 = ~n25795 ;
  assign n26208 = n73942 & n26207 ;
  assign n73943 = ~n25784 ;
  assign n26209 = x94 & n73943 ;
  assign n73944 = ~n25782 ;
  assign n26210 = n73944 & n26209 ;
  assign n26211 = n25786 | n26210 ;
  assign n26212 = n26208 | n26211 ;
  assign n73945 = ~n25786 ;
  assign n26213 = n73945 & n26212 ;
  assign n73946 = ~n25775 ;
  assign n26214 = x95 & n73946 ;
  assign n73947 = ~n25773 ;
  assign n26215 = n73947 & n26214 ;
  assign n26216 = n25777 | n26215 ;
  assign n26218 = n26213 | n26216 ;
  assign n73948 = ~n25777 ;
  assign n26219 = n73948 & n26218 ;
  assign n73949 = ~n25766 ;
  assign n26220 = x96 & n73949 ;
  assign n73950 = ~n25764 ;
  assign n26221 = n73950 & n26220 ;
  assign n26222 = n25768 | n26221 ;
  assign n26223 = n26219 | n26222 ;
  assign n73951 = ~n25768 ;
  assign n26224 = n73951 & n26223 ;
  assign n73952 = ~n25757 ;
  assign n26225 = x97 & n73952 ;
  assign n73953 = ~n25755 ;
  assign n26226 = n73953 & n26225 ;
  assign n26227 = n25759 | n26226 ;
  assign n26229 = n26224 | n26227 ;
  assign n73954 = ~n25759 ;
  assign n26230 = n73954 & n26229 ;
  assign n73955 = ~n25748 ;
  assign n26231 = x98 & n73955 ;
  assign n73956 = ~n25746 ;
  assign n26232 = n73956 & n26231 ;
  assign n26233 = n25750 | n26232 ;
  assign n26234 = n26230 | n26233 ;
  assign n73957 = ~n25750 ;
  assign n26235 = n73957 & n26234 ;
  assign n73958 = ~n25739 ;
  assign n26236 = x99 & n73958 ;
  assign n73959 = ~n25737 ;
  assign n26237 = n73959 & n26236 ;
  assign n26238 = n25741 | n26237 ;
  assign n26240 = n26235 | n26238 ;
  assign n73960 = ~n25741 ;
  assign n26241 = n73960 & n26240 ;
  assign n73961 = ~n25730 ;
  assign n26242 = x100 & n73961 ;
  assign n73962 = ~n25728 ;
  assign n26243 = n73962 & n26242 ;
  assign n26244 = n25732 | n26243 ;
  assign n26245 = n26241 | n26244 ;
  assign n73963 = ~n25732 ;
  assign n26246 = n73963 & n26245 ;
  assign n73964 = ~n25721 ;
  assign n26247 = x101 & n73964 ;
  assign n73965 = ~n25719 ;
  assign n26248 = n73965 & n26247 ;
  assign n26249 = n25723 | n26248 ;
  assign n26251 = n26246 | n26249 ;
  assign n73966 = ~n25723 ;
  assign n26252 = n73966 & n26251 ;
  assign n73967 = ~n25712 ;
  assign n26253 = x102 & n73967 ;
  assign n73968 = ~n25710 ;
  assign n26254 = n73968 & n26253 ;
  assign n26255 = n25714 | n26254 ;
  assign n26256 = n26252 | n26255 ;
  assign n73969 = ~n25714 ;
  assign n26257 = n73969 & n26256 ;
  assign n73970 = ~n25703 ;
  assign n26258 = x103 & n73970 ;
  assign n73971 = ~n25701 ;
  assign n26259 = n73971 & n26258 ;
  assign n26260 = n25705 | n26259 ;
  assign n26262 = n26257 | n26260 ;
  assign n73972 = ~n25705 ;
  assign n26263 = n73972 & n26262 ;
  assign n73973 = ~n25694 ;
  assign n26264 = x104 & n73973 ;
  assign n73974 = ~n25692 ;
  assign n26265 = n73974 & n26264 ;
  assign n26266 = n25696 | n26265 ;
  assign n26267 = n26263 | n26266 ;
  assign n73975 = ~n25696 ;
  assign n26268 = n73975 & n26267 ;
  assign n73976 = ~n25686 ;
  assign n26269 = x105 & n73976 ;
  assign n73977 = ~n25684 ;
  assign n26270 = n73977 & n26269 ;
  assign n26271 = n25688 | n26270 ;
  assign n26273 = n26268 | n26271 ;
  assign n73978 = ~n25688 ;
  assign n26274 = n73978 & n26273 ;
  assign n73979 = ~n25678 ;
  assign n26275 = x106 & n73979 ;
  assign n73980 = ~n25676 ;
  assign n26276 = n73980 & n26275 ;
  assign n26277 = n25680 | n26276 ;
  assign n26278 = n26274 | n26277 ;
  assign n73981 = ~n25680 ;
  assign n26279 = n73981 & n26278 ;
  assign n73982 = ~n25669 ;
  assign n26280 = x107 & n73982 ;
  assign n73983 = ~n25667 ;
  assign n26281 = n73983 & n26280 ;
  assign n26282 = n25671 | n26281 ;
  assign n26284 = n26279 | n26282 ;
  assign n73984 = ~n25671 ;
  assign n26285 = n73984 & n26284 ;
  assign n73985 = ~n25660 ;
  assign n26286 = x108 & n73985 ;
  assign n73986 = ~n25658 ;
  assign n26287 = n73986 & n26286 ;
  assign n26288 = n25662 | n26287 ;
  assign n26289 = n26285 | n26288 ;
  assign n73987 = ~n25662 ;
  assign n26290 = n73987 & n26289 ;
  assign n73988 = ~n25652 ;
  assign n26291 = x109 & n73988 ;
  assign n73989 = ~n25650 ;
  assign n26292 = n73989 & n26291 ;
  assign n26293 = n25654 | n26292 ;
  assign n26295 = n26290 | n26293 ;
  assign n73990 = ~n25654 ;
  assign n26296 = n73990 & n26295 ;
  assign n73991 = ~n25643 ;
  assign n26297 = x110 & n73991 ;
  assign n73992 = ~n25641 ;
  assign n26298 = n73992 & n26297 ;
  assign n26299 = n25645 | n26298 ;
  assign n26300 = n26296 | n26299 ;
  assign n73993 = ~n25645 ;
  assign n26301 = n73993 & n26300 ;
  assign n73994 = ~n25634 ;
  assign n26302 = x111 & n73994 ;
  assign n73995 = ~n25632 ;
  assign n26303 = n73995 & n26302 ;
  assign n26304 = n25636 | n26303 ;
  assign n26306 = n26301 | n26304 ;
  assign n73996 = ~n25636 ;
  assign n26307 = n73996 & n26306 ;
  assign n73997 = ~n25625 ;
  assign n26308 = x112 & n73997 ;
  assign n73998 = ~n25623 ;
  assign n26309 = n73998 & n26308 ;
  assign n26310 = n25627 | n26309 ;
  assign n26311 = n26307 | n26310 ;
  assign n73999 = ~n25627 ;
  assign n26312 = n73999 & n26311 ;
  assign n74000 = ~n25616 ;
  assign n26313 = x113 & n74000 ;
  assign n74001 = ~n25614 ;
  assign n26314 = n74001 & n26313 ;
  assign n26315 = n25618 | n26314 ;
  assign n26317 = n26312 | n26315 ;
  assign n74002 = ~n25618 ;
  assign n26318 = n74002 & n26317 ;
  assign n74003 = ~n25607 ;
  assign n26319 = x114 & n74003 ;
  assign n74004 = ~n25605 ;
  assign n26320 = n74004 & n26319 ;
  assign n26321 = n25609 | n26320 ;
  assign n26322 = n26318 | n26321 ;
  assign n74005 = ~n25609 ;
  assign n26323 = n74005 & n26322 ;
  assign n74006 = ~n25599 ;
  assign n26324 = x115 & n74006 ;
  assign n74007 = ~n25597 ;
  assign n26325 = n74007 & n26324 ;
  assign n26326 = n25601 | n26325 ;
  assign n26328 = n26323 | n26326 ;
  assign n74008 = ~n25601 ;
  assign n26329 = n74008 & n26328 ;
  assign n74009 = ~n25590 ;
  assign n26330 = x116 & n74009 ;
  assign n74010 = ~n25588 ;
  assign n26331 = n74010 & n26330 ;
  assign n26332 = n25592 | n26331 ;
  assign n26333 = n26329 | n26332 ;
  assign n74011 = ~n25592 ;
  assign n26334 = n74011 & n26333 ;
  assign n74012 = ~n25581 ;
  assign n26335 = x117 & n74012 ;
  assign n74013 = ~n25579 ;
  assign n26336 = n74013 & n26335 ;
  assign n26337 = n25583 | n26336 ;
  assign n26339 = n26334 | n26337 ;
  assign n74014 = ~n25583 ;
  assign n26340 = n74014 & n26339 ;
  assign n74015 = ~n25573 ;
  assign n26341 = x118 & n74015 ;
  assign n74016 = ~n25571 ;
  assign n26342 = n74016 & n26341 ;
  assign n26343 = n25575 | n26342 ;
  assign n26344 = n26340 | n26343 ;
  assign n74017 = ~n25575 ;
  assign n26345 = n74017 & n26344 ;
  assign n74018 = ~n25455 ;
  assign n26346 = x119 & n74018 ;
  assign n74019 = ~n25453 ;
  assign n26347 = n74019 & n26346 ;
  assign n26348 = n25457 | n26347 ;
  assign n26350 = n26345 | n26348 ;
  assign n74020 = ~n25457 ;
  assign n26351 = n74020 & n26350 ;
  assign n74021 = ~x120 ;
  assign n26362 = n74021 & n26361 ;
  assign n74022 = ~n26360 ;
  assign n26363 = x120 & n74022 ;
  assign n74023 = ~n26358 ;
  assign n26364 = n74023 & n26363 ;
  assign n26365 = n278 | n26364 ;
  assign n26366 = n26362 | n26365 ;
  assign n26368 = n26351 | n26366 ;
  assign n74024 = ~n26367 ;
  assign n26369 = n74024 & n26368 ;
  assign n26513 = n25457 | n26364 ;
  assign n26514 = n26362 | n26513 ;
  assign n74025 = ~n26514 ;
  assign n26515 = n26350 & n74025 ;
  assign n26372 = n25449 | n26044 ;
  assign n26373 = x65 & n26372 ;
  assign n74026 = ~n26373 ;
  assign n26374 = n26050 & n74026 ;
  assign n26375 = n26052 | n26374 ;
  assign n26376 = n73858 & n26375 ;
  assign n26377 = n26058 | n26376 ;
  assign n26378 = n73861 & n26377 ;
  assign n26380 = n26063 | n26378 ;
  assign n26381 = n73864 & n26380 ;
  assign n26383 = n26068 | n26381 ;
  assign n26384 = n73867 & n26383 ;
  assign n26385 = n26073 | n26384 ;
  assign n26386 = n73870 & n26385 ;
  assign n26387 = n26079 | n26386 ;
  assign n26389 = n73873 & n26387 ;
  assign n26390 = n26084 | n26389 ;
  assign n26391 = n73876 & n26390 ;
  assign n26392 = n26090 | n26391 ;
  assign n26394 = n73879 & n26392 ;
  assign n26395 = n26095 | n26394 ;
  assign n26396 = n73882 & n26395 ;
  assign n26397 = n26101 | n26396 ;
  assign n26399 = n73885 & n26397 ;
  assign n26400 = n26106 | n26399 ;
  assign n26401 = n73888 & n26400 ;
  assign n26402 = n26112 | n26401 ;
  assign n26404 = n73891 & n26402 ;
  assign n26405 = n26117 | n26404 ;
  assign n26406 = n73894 & n26405 ;
  assign n26407 = n26123 | n26406 ;
  assign n26409 = n73897 & n26407 ;
  assign n26410 = n26128 | n26409 ;
  assign n26411 = n73900 & n26410 ;
  assign n26412 = n26134 | n26411 ;
  assign n26414 = n73903 & n26412 ;
  assign n26415 = n26139 | n26414 ;
  assign n26416 = n73906 & n26415 ;
  assign n26417 = n26145 | n26416 ;
  assign n26419 = n73909 & n26417 ;
  assign n26420 = n26150 | n26419 ;
  assign n26421 = n73912 & n26420 ;
  assign n26422 = n26156 | n26421 ;
  assign n26424 = n73915 & n26422 ;
  assign n26425 = n26161 | n26424 ;
  assign n26426 = n73918 & n26425 ;
  assign n26427 = n26167 | n26426 ;
  assign n26429 = n73921 & n26427 ;
  assign n26430 = n26172 | n26429 ;
  assign n26431 = n73924 & n26430 ;
  assign n26432 = n26178 | n26431 ;
  assign n26434 = n73927 & n26432 ;
  assign n26435 = n26183 | n26434 ;
  assign n26436 = n73930 & n26435 ;
  assign n26437 = n26189 | n26436 ;
  assign n26439 = n73933 & n26437 ;
  assign n26440 = n26194 | n26439 ;
  assign n26441 = n73936 & n26440 ;
  assign n26442 = n26200 | n26441 ;
  assign n26444 = n73939 & n26442 ;
  assign n26445 = n26205 | n26444 ;
  assign n26446 = n73942 & n26445 ;
  assign n26447 = n26211 | n26446 ;
  assign n26449 = n73945 & n26447 ;
  assign n26450 = n26216 | n26449 ;
  assign n26451 = n73948 & n26450 ;
  assign n26452 = n26222 | n26451 ;
  assign n26454 = n73951 & n26452 ;
  assign n26455 = n26227 | n26454 ;
  assign n26456 = n73954 & n26455 ;
  assign n26457 = n26233 | n26456 ;
  assign n26459 = n73957 & n26457 ;
  assign n26460 = n26238 | n26459 ;
  assign n26461 = n73960 & n26460 ;
  assign n26462 = n26244 | n26461 ;
  assign n26464 = n73963 & n26462 ;
  assign n26465 = n26249 | n26464 ;
  assign n26466 = n73966 & n26465 ;
  assign n26467 = n26255 | n26466 ;
  assign n26469 = n73969 & n26467 ;
  assign n26470 = n26260 | n26469 ;
  assign n26471 = n73972 & n26470 ;
  assign n26472 = n26266 | n26471 ;
  assign n26474 = n73975 & n26472 ;
  assign n26475 = n26271 | n26474 ;
  assign n26476 = n73978 & n26475 ;
  assign n26477 = n26277 | n26476 ;
  assign n26479 = n73981 & n26477 ;
  assign n26480 = n26282 | n26479 ;
  assign n26481 = n73984 & n26480 ;
  assign n26482 = n26288 | n26481 ;
  assign n26484 = n73987 & n26482 ;
  assign n26485 = n26293 | n26484 ;
  assign n26486 = n73990 & n26485 ;
  assign n26487 = n26299 | n26486 ;
  assign n26489 = n73993 & n26487 ;
  assign n26490 = n26304 | n26489 ;
  assign n26491 = n73996 & n26490 ;
  assign n26492 = n26310 | n26491 ;
  assign n26494 = n73999 & n26492 ;
  assign n26495 = n26315 | n26494 ;
  assign n26496 = n74002 & n26495 ;
  assign n26497 = n26321 | n26496 ;
  assign n26499 = n74005 & n26497 ;
  assign n26500 = n26326 | n26499 ;
  assign n26501 = n74008 & n26500 ;
  assign n26502 = n26332 | n26501 ;
  assign n26504 = n74011 & n26502 ;
  assign n26505 = n26337 | n26504 ;
  assign n26506 = n74014 & n26505 ;
  assign n26507 = n26343 | n26506 ;
  assign n26509 = n74017 & n26507 ;
  assign n26510 = n26348 | n26509 ;
  assign n26511 = n74020 & n26510 ;
  assign n26516 = n26362 | n26364 ;
  assign n74027 = ~n26511 ;
  assign n26517 = n74027 & n26516 ;
  assign n26518 = n26515 | n26517 ;
  assign n136 = ~n26369 ;
  assign n26519 = n136 & n26518 ;
  assign n26512 = n26366 | n26511 ;
  assign n26520 = n66655 & n26361 ;
  assign n26521 = n26512 & n26520 ;
  assign n26522 = n26519 | n26521 ;
  assign n74029 = ~x121 ;
  assign n26523 = n74029 & n26522 ;
  assign n74030 = ~n26521 ;
  assign n27305 = x121 & n74030 ;
  assign n74031 = ~n26519 ;
  assign n27306 = n74031 & n27305 ;
  assign n27307 = n26523 | n27306 ;
  assign n74032 = ~n26345 ;
  assign n26349 = n74032 & n26348 ;
  assign n26524 = n25575 | n26348 ;
  assign n74033 = ~n26524 ;
  assign n26525 = n26507 & n74033 ;
  assign n26526 = n26349 | n26525 ;
  assign n26527 = n136 & n26526 ;
  assign n26528 = n25456 & n74024 ;
  assign n26529 = n26512 & n26528 ;
  assign n26530 = n26527 | n26529 ;
  assign n26531 = n74021 & n26530 ;
  assign n74034 = ~n26506 ;
  assign n26508 = n26343 & n74034 ;
  assign n26532 = n25583 | n26343 ;
  assign n74035 = ~n26532 ;
  assign n26533 = n26339 & n74035 ;
  assign n26534 = n26508 | n26533 ;
  assign n26535 = n136 & n26534 ;
  assign n26536 = n25574 & n74024 ;
  assign n26537 = n26512 & n26536 ;
  assign n26538 = n26535 | n26537 ;
  assign n26539 = n73617 & n26538 ;
  assign n74036 = ~n26537 ;
  assign n27293 = x119 & n74036 ;
  assign n74037 = ~n26535 ;
  assign n27294 = n74037 & n27293 ;
  assign n27295 = n26539 | n27294 ;
  assign n74038 = ~n26334 ;
  assign n26338 = n74038 & n26337 ;
  assign n26540 = n25592 | n26337 ;
  assign n74039 = ~n26540 ;
  assign n26541 = n26502 & n74039 ;
  assign n26542 = n26338 | n26541 ;
  assign n26543 = n136 & n26542 ;
  assign n26544 = n25582 & n74024 ;
  assign n26545 = n26512 & n26544 ;
  assign n26546 = n26543 | n26545 ;
  assign n26547 = n73188 & n26546 ;
  assign n74040 = ~n26501 ;
  assign n26503 = n26332 & n74040 ;
  assign n26548 = n25601 | n26332 ;
  assign n74041 = ~n26548 ;
  assign n26549 = n26328 & n74041 ;
  assign n26550 = n26503 | n26549 ;
  assign n26551 = n136 & n26550 ;
  assign n26552 = n25591 & n74024 ;
  assign n26553 = n26512 & n26552 ;
  assign n26554 = n26551 | n26553 ;
  assign n26555 = n73177 & n26554 ;
  assign n74042 = ~n26553 ;
  assign n27281 = x117 & n74042 ;
  assign n74043 = ~n26551 ;
  assign n27282 = n74043 & n27281 ;
  assign n27283 = n26555 | n27282 ;
  assign n74044 = ~n26323 ;
  assign n26327 = n74044 & n26326 ;
  assign n26556 = n25609 | n26326 ;
  assign n74045 = ~n26556 ;
  assign n26557 = n26497 & n74045 ;
  assign n26558 = n26327 | n26557 ;
  assign n26559 = n136 & n26558 ;
  assign n26560 = n25600 & n74024 ;
  assign n26561 = n26512 & n26560 ;
  assign n26562 = n26559 | n26561 ;
  assign n26563 = n72752 & n26562 ;
  assign n74046 = ~n26496 ;
  assign n26498 = n26321 & n74046 ;
  assign n26564 = n25618 | n26321 ;
  assign n74047 = ~n26564 ;
  assign n26565 = n26317 & n74047 ;
  assign n26566 = n26498 | n26565 ;
  assign n26567 = n136 & n26566 ;
  assign n26568 = n25608 & n74024 ;
  assign n26569 = n26512 & n26568 ;
  assign n26570 = n26567 | n26569 ;
  assign n26571 = n72393 & n26570 ;
  assign n74048 = ~n26569 ;
  assign n27269 = x115 & n74048 ;
  assign n74049 = ~n26567 ;
  assign n27270 = n74049 & n27269 ;
  assign n27271 = n26571 | n27270 ;
  assign n74050 = ~n26312 ;
  assign n26316 = n74050 & n26315 ;
  assign n26572 = n25627 | n26315 ;
  assign n74051 = ~n26572 ;
  assign n26573 = n26492 & n74051 ;
  assign n26574 = n26316 | n26573 ;
  assign n26575 = n136 & n26574 ;
  assign n26576 = n25617 & n74024 ;
  assign n26577 = n26512 & n26576 ;
  assign n26578 = n26575 | n26577 ;
  assign n26579 = n72385 & n26578 ;
  assign n74052 = ~n26491 ;
  assign n26493 = n26310 & n74052 ;
  assign n26580 = n25636 | n26310 ;
  assign n74053 = ~n26580 ;
  assign n26581 = n26306 & n74053 ;
  assign n26582 = n26493 | n26581 ;
  assign n26583 = n136 & n26582 ;
  assign n26584 = n25626 & n74024 ;
  assign n26585 = n26512 & n26584 ;
  assign n26586 = n26583 | n26585 ;
  assign n26587 = n72025 & n26586 ;
  assign n74054 = ~n26585 ;
  assign n27257 = x113 & n74054 ;
  assign n74055 = ~n26583 ;
  assign n27258 = n74055 & n27257 ;
  assign n27259 = n26587 | n27258 ;
  assign n74056 = ~n26301 ;
  assign n26305 = n74056 & n26304 ;
  assign n26588 = n25645 | n26304 ;
  assign n74057 = ~n26588 ;
  assign n26589 = n26487 & n74057 ;
  assign n26590 = n26305 | n26589 ;
  assign n26591 = n136 & n26590 ;
  assign n26592 = n25635 & n74024 ;
  assign n26593 = n26512 & n26592 ;
  assign n26594 = n26591 | n26593 ;
  assign n26595 = n71645 & n26594 ;
  assign n74058 = ~n26486 ;
  assign n26488 = n26299 & n74058 ;
  assign n26596 = n25654 | n26299 ;
  assign n74059 = ~n26596 ;
  assign n26597 = n26295 & n74059 ;
  assign n26598 = n26488 | n26597 ;
  assign n26599 = n136 & n26598 ;
  assign n26600 = n25644 & n74024 ;
  assign n26601 = n26512 & n26600 ;
  assign n26602 = n26599 | n26601 ;
  assign n26603 = n71633 & n26602 ;
  assign n74060 = ~n26601 ;
  assign n27245 = x111 & n74060 ;
  assign n74061 = ~n26599 ;
  assign n27246 = n74061 & n27245 ;
  assign n27247 = n26603 | n27246 ;
  assign n74062 = ~n26290 ;
  assign n26294 = n74062 & n26293 ;
  assign n26604 = n25662 | n26293 ;
  assign n74063 = ~n26604 ;
  assign n26605 = n26482 & n74063 ;
  assign n26606 = n26294 | n26605 ;
  assign n26607 = n136 & n26606 ;
  assign n26608 = n25653 & n74024 ;
  assign n26609 = n26512 & n26608 ;
  assign n26610 = n26607 | n26609 ;
  assign n26611 = n71253 & n26610 ;
  assign n74064 = ~n26481 ;
  assign n26483 = n26288 & n74064 ;
  assign n26612 = n25671 | n26288 ;
  assign n74065 = ~n26612 ;
  assign n26613 = n26284 & n74065 ;
  assign n26614 = n26483 | n26613 ;
  assign n26615 = n136 & n26614 ;
  assign n26616 = n25661 & n74024 ;
  assign n26617 = n26512 & n26616 ;
  assign n26618 = n26615 | n26617 ;
  assign n26619 = n70935 & n26618 ;
  assign n74066 = ~n26617 ;
  assign n27233 = x109 & n74066 ;
  assign n74067 = ~n26615 ;
  assign n27234 = n74067 & n27233 ;
  assign n27235 = n26619 | n27234 ;
  assign n74068 = ~n26279 ;
  assign n26283 = n74068 & n26282 ;
  assign n26620 = n25680 | n26282 ;
  assign n74069 = ~n26620 ;
  assign n26621 = n26477 & n74069 ;
  assign n26622 = n26283 | n26621 ;
  assign n26623 = n136 & n26622 ;
  assign n26624 = n25670 & n74024 ;
  assign n26625 = n26512 & n26624 ;
  assign n26626 = n26623 | n26625 ;
  assign n26627 = n70927 & n26626 ;
  assign n74070 = ~n26476 ;
  assign n26478 = n26277 & n74070 ;
  assign n26628 = n25688 | n26277 ;
  assign n74071 = ~n26628 ;
  assign n26629 = n26273 & n74071 ;
  assign n26630 = n26478 | n26629 ;
  assign n26631 = n136 & n26630 ;
  assign n26632 = n25679 & n74024 ;
  assign n26633 = n26512 & n26632 ;
  assign n26634 = n26631 | n26633 ;
  assign n26635 = n70609 & n26634 ;
  assign n74072 = ~n26633 ;
  assign n27221 = x107 & n74072 ;
  assign n74073 = ~n26631 ;
  assign n27222 = n74073 & n27221 ;
  assign n27223 = n26635 | n27222 ;
  assign n74074 = ~n26268 ;
  assign n26272 = n74074 & n26271 ;
  assign n26636 = n25696 | n26271 ;
  assign n74075 = ~n26636 ;
  assign n26637 = n26472 & n74075 ;
  assign n26638 = n26272 | n26637 ;
  assign n26639 = n136 & n26638 ;
  assign n26640 = n25687 & n74024 ;
  assign n26641 = n26512 & n26640 ;
  assign n26642 = n26639 | n26641 ;
  assign n26643 = n70276 & n26642 ;
  assign n74076 = ~n26471 ;
  assign n26473 = n26266 & n74076 ;
  assign n26644 = n25705 | n26266 ;
  assign n74077 = ~n26644 ;
  assign n26645 = n26262 & n74077 ;
  assign n26646 = n26473 | n26645 ;
  assign n26647 = n136 & n26646 ;
  assign n26648 = n25695 & n74024 ;
  assign n26649 = n26512 & n26648 ;
  assign n26650 = n26647 | n26649 ;
  assign n26651 = n70176 & n26650 ;
  assign n74078 = ~n26649 ;
  assign n27209 = x105 & n74078 ;
  assign n74079 = ~n26647 ;
  assign n27210 = n74079 & n27209 ;
  assign n27211 = n26651 | n27210 ;
  assign n74080 = ~n26257 ;
  assign n26261 = n74080 & n26260 ;
  assign n26652 = n25714 | n26260 ;
  assign n74081 = ~n26652 ;
  assign n26653 = n26467 & n74081 ;
  assign n26654 = n26261 | n26653 ;
  assign n26655 = n136 & n26654 ;
  assign n26656 = n25704 & n74024 ;
  assign n26657 = n26512 & n26656 ;
  assign n26658 = n26655 | n26657 ;
  assign n26659 = n69857 & n26658 ;
  assign n74082 = ~n26466 ;
  assign n26468 = n26255 & n74082 ;
  assign n26660 = n25723 | n26255 ;
  assign n74083 = ~n26660 ;
  assign n26661 = n26251 & n74083 ;
  assign n26662 = n26468 | n26661 ;
  assign n26663 = n136 & n26662 ;
  assign n26664 = n25713 & n74024 ;
  assign n26665 = n26512 & n26664 ;
  assign n26666 = n26663 | n26665 ;
  assign n26667 = n69656 & n26666 ;
  assign n74084 = ~n26665 ;
  assign n27197 = x103 & n74084 ;
  assign n74085 = ~n26663 ;
  assign n27198 = n74085 & n27197 ;
  assign n27199 = n26667 | n27198 ;
  assign n74086 = ~n26246 ;
  assign n26250 = n74086 & n26249 ;
  assign n26668 = n25732 | n26249 ;
  assign n74087 = ~n26668 ;
  assign n26669 = n26462 & n74087 ;
  assign n26670 = n26250 | n26669 ;
  assign n26671 = n136 & n26670 ;
  assign n26672 = n25722 & n74024 ;
  assign n26673 = n26512 & n26672 ;
  assign n26674 = n26671 | n26673 ;
  assign n26675 = n69528 & n26674 ;
  assign n74088 = ~n26461 ;
  assign n26463 = n26244 & n74088 ;
  assign n26676 = n25741 | n26244 ;
  assign n74089 = ~n26676 ;
  assign n26677 = n26240 & n74089 ;
  assign n26678 = n26463 | n26677 ;
  assign n26679 = n136 & n26678 ;
  assign n26680 = n25731 & n74024 ;
  assign n26681 = n26512 & n26680 ;
  assign n26682 = n26679 | n26681 ;
  assign n26683 = n69261 & n26682 ;
  assign n74090 = ~n26681 ;
  assign n27185 = x101 & n74090 ;
  assign n74091 = ~n26679 ;
  assign n27186 = n74091 & n27185 ;
  assign n27187 = n26683 | n27186 ;
  assign n74092 = ~n26235 ;
  assign n26239 = n74092 & n26238 ;
  assign n26684 = n25750 | n26238 ;
  assign n74093 = ~n26684 ;
  assign n26685 = n26457 & n74093 ;
  assign n26686 = n26239 | n26685 ;
  assign n26687 = n136 & n26686 ;
  assign n26688 = n25740 & n74024 ;
  assign n26689 = n26512 & n26688 ;
  assign n26690 = n26687 | n26689 ;
  assign n26691 = n69075 & n26690 ;
  assign n74094 = ~n26456 ;
  assign n26458 = n26233 & n74094 ;
  assign n26692 = n25759 | n26233 ;
  assign n74095 = ~n26692 ;
  assign n26693 = n26229 & n74095 ;
  assign n26694 = n26458 | n26693 ;
  assign n26695 = n136 & n26694 ;
  assign n26696 = n25749 & n74024 ;
  assign n26697 = n26512 & n26696 ;
  assign n26698 = n26695 | n26697 ;
  assign n26699 = n68993 & n26698 ;
  assign n74096 = ~n26697 ;
  assign n27173 = x99 & n74096 ;
  assign n74097 = ~n26695 ;
  assign n27174 = n74097 & n27173 ;
  assign n27175 = n26699 | n27174 ;
  assign n74098 = ~n26224 ;
  assign n26228 = n74098 & n26227 ;
  assign n26700 = n25768 | n26227 ;
  assign n74099 = ~n26700 ;
  assign n26701 = n26452 & n74099 ;
  assign n26702 = n26228 | n26701 ;
  assign n26703 = n136 & n26702 ;
  assign n26704 = n25758 & n74024 ;
  assign n26705 = n26512 & n26704 ;
  assign n26706 = n26703 | n26705 ;
  assign n26707 = n68716 & n26706 ;
  assign n74100 = ~n26451 ;
  assign n26453 = n26222 & n74100 ;
  assign n26708 = n25777 | n26222 ;
  assign n74101 = ~n26708 ;
  assign n26709 = n26218 & n74101 ;
  assign n26710 = n26453 | n26709 ;
  assign n26711 = n136 & n26710 ;
  assign n26712 = n25767 & n74024 ;
  assign n26713 = n26512 & n26712 ;
  assign n26714 = n26711 | n26713 ;
  assign n26715 = n68545 & n26714 ;
  assign n74102 = ~n26713 ;
  assign n27161 = x97 & n74102 ;
  assign n74103 = ~n26711 ;
  assign n27162 = n74103 & n27161 ;
  assign n27163 = n26715 | n27162 ;
  assign n74104 = ~n26213 ;
  assign n26217 = n74104 & n26216 ;
  assign n26716 = n25786 | n26216 ;
  assign n74105 = ~n26716 ;
  assign n26717 = n26447 & n74105 ;
  assign n26718 = n26217 | n26717 ;
  assign n26719 = n136 & n26718 ;
  assign n26720 = n25776 & n74024 ;
  assign n26721 = n26512 & n26720 ;
  assign n26722 = n26719 | n26721 ;
  assign n26723 = n68438 & n26722 ;
  assign n74106 = ~n26446 ;
  assign n26448 = n26211 & n74106 ;
  assign n26724 = n25795 | n26211 ;
  assign n74107 = ~n26724 ;
  assign n26725 = n26207 & n74107 ;
  assign n26726 = n26448 | n26725 ;
  assign n26727 = n136 & n26726 ;
  assign n26728 = n25785 & n74024 ;
  assign n26729 = n26512 & n26728 ;
  assign n26730 = n26727 | n26729 ;
  assign n26731 = n68214 & n26730 ;
  assign n74108 = ~n26729 ;
  assign n27149 = x95 & n74108 ;
  assign n74109 = ~n26727 ;
  assign n27150 = n74109 & n27149 ;
  assign n27151 = n26731 | n27150 ;
  assign n74110 = ~n26202 ;
  assign n26206 = n74110 & n26205 ;
  assign n26732 = n25804 | n26205 ;
  assign n74111 = ~n26732 ;
  assign n26733 = n26442 & n74111 ;
  assign n26734 = n26206 | n26733 ;
  assign n26735 = n136 & n26734 ;
  assign n26736 = n25794 & n74024 ;
  assign n26737 = n26512 & n26736 ;
  assign n26738 = n26735 | n26737 ;
  assign n26739 = n68058 & n26738 ;
  assign n74112 = ~n26441 ;
  assign n26443 = n26200 & n74112 ;
  assign n26740 = n25813 | n26200 ;
  assign n74113 = ~n26740 ;
  assign n26741 = n26196 & n74113 ;
  assign n26742 = n26443 | n26741 ;
  assign n26743 = n136 & n26742 ;
  assign n26744 = n25803 & n74024 ;
  assign n26745 = n26512 & n26744 ;
  assign n26746 = n26743 | n26745 ;
  assign n26747 = n67986 & n26746 ;
  assign n74114 = ~n26745 ;
  assign n27137 = x93 & n74114 ;
  assign n74115 = ~n26743 ;
  assign n27138 = n74115 & n27137 ;
  assign n27139 = n26747 | n27138 ;
  assign n74116 = ~n26191 ;
  assign n26195 = n74116 & n26194 ;
  assign n26748 = n25822 | n26194 ;
  assign n74117 = ~n26748 ;
  assign n26749 = n26437 & n74117 ;
  assign n26750 = n26195 | n26749 ;
  assign n26751 = n136 & n26750 ;
  assign n26752 = n25812 & n74024 ;
  assign n26753 = n26512 & n26752 ;
  assign n26754 = n26751 | n26753 ;
  assign n26755 = n67763 & n26754 ;
  assign n74118 = ~n26436 ;
  assign n26438 = n26189 & n74118 ;
  assign n26756 = n25831 | n26189 ;
  assign n74119 = ~n26756 ;
  assign n26757 = n26185 & n74119 ;
  assign n26758 = n26438 | n26757 ;
  assign n26759 = n136 & n26758 ;
  assign n26760 = n25821 & n74024 ;
  assign n26761 = n26512 & n26760 ;
  assign n26762 = n26759 | n26761 ;
  assign n26763 = n67622 & n26762 ;
  assign n74120 = ~n26761 ;
  assign n27125 = x91 & n74120 ;
  assign n74121 = ~n26759 ;
  assign n27126 = n74121 & n27125 ;
  assign n27127 = n26763 | n27126 ;
  assign n74122 = ~n26180 ;
  assign n26184 = n74122 & n26183 ;
  assign n26764 = n25840 | n26183 ;
  assign n74123 = ~n26764 ;
  assign n26765 = n26432 & n74123 ;
  assign n26766 = n26184 | n26765 ;
  assign n26767 = n136 & n26766 ;
  assign n26768 = n25830 & n74024 ;
  assign n26769 = n26512 & n26768 ;
  assign n26770 = n26767 | n26769 ;
  assign n26771 = n67531 & n26770 ;
  assign n74124 = ~n26431 ;
  assign n26433 = n26178 & n74124 ;
  assign n26772 = n25849 | n26178 ;
  assign n74125 = ~n26772 ;
  assign n26773 = n26174 & n74125 ;
  assign n26774 = n26433 | n26773 ;
  assign n26775 = n136 & n26774 ;
  assign n26776 = n25839 & n74024 ;
  assign n26777 = n26512 & n26776 ;
  assign n26778 = n26775 | n26777 ;
  assign n26779 = n67348 & n26778 ;
  assign n74126 = ~n26777 ;
  assign n27113 = x89 & n74126 ;
  assign n74127 = ~n26775 ;
  assign n27114 = n74127 & n27113 ;
  assign n27115 = n26779 | n27114 ;
  assign n74128 = ~n26169 ;
  assign n26173 = n74128 & n26172 ;
  assign n26780 = n25858 | n26172 ;
  assign n74129 = ~n26780 ;
  assign n26781 = n26427 & n74129 ;
  assign n26782 = n26173 | n26781 ;
  assign n26783 = n136 & n26782 ;
  assign n26784 = n25848 & n74024 ;
  assign n26785 = n26512 & n26784 ;
  assign n26786 = n26783 | n26785 ;
  assign n26787 = n67222 & n26786 ;
  assign n74130 = ~n26426 ;
  assign n26428 = n26167 & n74130 ;
  assign n26788 = n25867 | n26167 ;
  assign n74131 = ~n26788 ;
  assign n26789 = n26163 & n74131 ;
  assign n26790 = n26428 | n26789 ;
  assign n26791 = n136 & n26790 ;
  assign n26792 = n25857 & n74024 ;
  assign n26793 = n26512 & n26792 ;
  assign n26794 = n26791 | n26793 ;
  assign n26795 = n67164 & n26794 ;
  assign n74132 = ~n26793 ;
  assign n27101 = x87 & n74132 ;
  assign n74133 = ~n26791 ;
  assign n27102 = n74133 & n27101 ;
  assign n27103 = n26795 | n27102 ;
  assign n74134 = ~n26158 ;
  assign n26162 = n74134 & n26161 ;
  assign n26796 = n25876 | n26161 ;
  assign n74135 = ~n26796 ;
  assign n26797 = n26422 & n74135 ;
  assign n26798 = n26162 | n26797 ;
  assign n26799 = n136 & n26798 ;
  assign n26800 = n25866 & n74024 ;
  assign n26801 = n26512 & n26800 ;
  assign n26802 = n26799 | n26801 ;
  assign n26803 = n66979 & n26802 ;
  assign n74136 = ~n26421 ;
  assign n26423 = n26156 & n74136 ;
  assign n26804 = n25885 | n26156 ;
  assign n74137 = ~n26804 ;
  assign n26805 = n26152 & n74137 ;
  assign n26806 = n26423 | n26805 ;
  assign n26807 = n136 & n26806 ;
  assign n26808 = n25875 & n74024 ;
  assign n26809 = n26512 & n26808 ;
  assign n26810 = n26807 | n26809 ;
  assign n26811 = n66868 & n26810 ;
  assign n74138 = ~n26809 ;
  assign n27089 = x85 & n74138 ;
  assign n74139 = ~n26807 ;
  assign n27090 = n74139 & n27089 ;
  assign n27091 = n26811 | n27090 ;
  assign n74140 = ~n26147 ;
  assign n26151 = n74140 & n26150 ;
  assign n26812 = n25894 | n26150 ;
  assign n74141 = ~n26812 ;
  assign n26813 = n26417 & n74141 ;
  assign n26814 = n26151 | n26813 ;
  assign n26815 = n136 & n26814 ;
  assign n26816 = n25884 & n74024 ;
  assign n26817 = n26512 & n26816 ;
  assign n26818 = n26815 | n26817 ;
  assign n26819 = n66797 & n26818 ;
  assign n74142 = ~n26416 ;
  assign n26418 = n26145 & n74142 ;
  assign n26820 = n25903 | n26145 ;
  assign n74143 = ~n26820 ;
  assign n26821 = n26141 & n74143 ;
  assign n26822 = n26418 | n26821 ;
  assign n26823 = n136 & n26822 ;
  assign n26824 = n25893 & n74024 ;
  assign n26825 = n26512 & n26824 ;
  assign n26826 = n26823 | n26825 ;
  assign n26827 = n66654 & n26826 ;
  assign n74144 = ~n26825 ;
  assign n27077 = x83 & n74144 ;
  assign n74145 = ~n26823 ;
  assign n27078 = n74145 & n27077 ;
  assign n27079 = n26827 | n27078 ;
  assign n74146 = ~n26136 ;
  assign n26140 = n74146 & n26139 ;
  assign n26828 = n25911 | n26139 ;
  assign n74147 = ~n26828 ;
  assign n26829 = n26412 & n74147 ;
  assign n26830 = n26140 | n26829 ;
  assign n26831 = n136 & n26830 ;
  assign n26832 = n25902 & n74024 ;
  assign n26833 = n26512 & n26832 ;
  assign n26834 = n26831 | n26833 ;
  assign n26835 = n66560 & n26834 ;
  assign n74148 = ~n26411 ;
  assign n26413 = n26134 & n74148 ;
  assign n26836 = n25920 | n26134 ;
  assign n74149 = ~n26836 ;
  assign n26837 = n26130 & n74149 ;
  assign n26838 = n26413 | n26837 ;
  assign n26839 = n136 & n26838 ;
  assign n26840 = n25910 & n74024 ;
  assign n26841 = n26512 & n26840 ;
  assign n26842 = n26839 | n26841 ;
  assign n26843 = n66505 & n26842 ;
  assign n74150 = ~n26841 ;
  assign n27065 = x81 & n74150 ;
  assign n74151 = ~n26839 ;
  assign n27066 = n74151 & n27065 ;
  assign n27067 = n26843 | n27066 ;
  assign n74152 = ~n26125 ;
  assign n26129 = n74152 & n26128 ;
  assign n26844 = n25929 | n26128 ;
  assign n74153 = ~n26844 ;
  assign n26845 = n26407 & n74153 ;
  assign n26846 = n26129 | n26845 ;
  assign n26847 = n136 & n26846 ;
  assign n26848 = n25919 & n74024 ;
  assign n26849 = n26512 & n26848 ;
  assign n26850 = n26847 | n26849 ;
  assign n26851 = n66379 & n26850 ;
  assign n74154 = ~n26406 ;
  assign n26408 = n26123 & n74154 ;
  assign n26852 = n25938 | n26123 ;
  assign n74155 = ~n26852 ;
  assign n26853 = n26119 & n74155 ;
  assign n26854 = n26408 | n26853 ;
  assign n26855 = n136 & n26854 ;
  assign n26856 = n25928 & n74024 ;
  assign n26857 = n26512 & n26856 ;
  assign n26858 = n26855 | n26857 ;
  assign n26859 = n66299 & n26858 ;
  assign n74156 = ~n26857 ;
  assign n27053 = x79 & n74156 ;
  assign n74157 = ~n26855 ;
  assign n27054 = n74157 & n27053 ;
  assign n27055 = n26859 | n27054 ;
  assign n74158 = ~n26114 ;
  assign n26118 = n74158 & n26117 ;
  assign n26860 = n25947 | n26117 ;
  assign n74159 = ~n26860 ;
  assign n26861 = n26402 & n74159 ;
  assign n26862 = n26118 | n26861 ;
  assign n26863 = n136 & n26862 ;
  assign n26864 = n25937 & n74024 ;
  assign n26865 = n26512 & n26864 ;
  assign n26866 = n26863 | n26865 ;
  assign n26867 = n66244 & n26866 ;
  assign n74160 = ~n26401 ;
  assign n26403 = n26112 & n74160 ;
  assign n26868 = n25956 | n26112 ;
  assign n74161 = ~n26868 ;
  assign n26869 = n26108 & n74161 ;
  assign n26870 = n26403 | n26869 ;
  assign n26871 = n136 & n26870 ;
  assign n26872 = n25946 & n74024 ;
  assign n26873 = n26512 & n26872 ;
  assign n26874 = n26871 | n26873 ;
  assign n26875 = n66145 & n26874 ;
  assign n74162 = ~n26873 ;
  assign n27041 = x77 & n74162 ;
  assign n74163 = ~n26871 ;
  assign n27042 = n74163 & n27041 ;
  assign n27043 = n26875 | n27042 ;
  assign n74164 = ~n26103 ;
  assign n26107 = n74164 & n26106 ;
  assign n26876 = n25965 | n26106 ;
  assign n74165 = ~n26876 ;
  assign n26877 = n26397 & n74165 ;
  assign n26878 = n26107 | n26877 ;
  assign n26879 = n136 & n26878 ;
  assign n26880 = n25955 & n74024 ;
  assign n26881 = n26512 & n26880 ;
  assign n26882 = n26879 | n26881 ;
  assign n26883 = n66081 & n26882 ;
  assign n74166 = ~n26396 ;
  assign n26398 = n26101 & n74166 ;
  assign n26884 = n25974 | n26101 ;
  assign n74167 = ~n26884 ;
  assign n26885 = n26097 & n74167 ;
  assign n26886 = n26398 | n26885 ;
  assign n26887 = n136 & n26886 ;
  assign n26888 = n25964 & n74024 ;
  assign n26889 = n26512 & n26888 ;
  assign n26890 = n26887 | n26889 ;
  assign n26891 = n66043 & n26890 ;
  assign n74168 = ~n26889 ;
  assign n27029 = x75 & n74168 ;
  assign n74169 = ~n26887 ;
  assign n27030 = n74169 & n27029 ;
  assign n27031 = n26891 | n27030 ;
  assign n74170 = ~n26092 ;
  assign n26096 = n74170 & n26095 ;
  assign n26892 = n25983 | n26095 ;
  assign n74171 = ~n26892 ;
  assign n26893 = n26392 & n74171 ;
  assign n26894 = n26096 | n26893 ;
  assign n26895 = n136 & n26894 ;
  assign n26896 = n25973 & n74024 ;
  assign n26897 = n26512 & n26896 ;
  assign n26898 = n26895 | n26897 ;
  assign n26899 = n65960 & n26898 ;
  assign n74172 = ~n26391 ;
  assign n26393 = n26090 & n74172 ;
  assign n26900 = n25992 | n26090 ;
  assign n74173 = ~n26900 ;
  assign n26901 = n26086 & n74173 ;
  assign n26902 = n26393 | n26901 ;
  assign n26903 = n136 & n26902 ;
  assign n26904 = n25982 & n74024 ;
  assign n26905 = n26512 & n26904 ;
  assign n26906 = n26903 | n26905 ;
  assign n26907 = n65909 & n26906 ;
  assign n74174 = ~n26905 ;
  assign n27017 = x73 & n74174 ;
  assign n74175 = ~n26903 ;
  assign n27018 = n74175 & n27017 ;
  assign n27019 = n26907 | n27018 ;
  assign n74176 = ~n26081 ;
  assign n26085 = n74176 & n26084 ;
  assign n26908 = n26001 | n26084 ;
  assign n74177 = ~n26908 ;
  assign n26909 = n26387 & n74177 ;
  assign n26910 = n26085 | n26909 ;
  assign n26911 = n136 & n26910 ;
  assign n26912 = n25991 & n74024 ;
  assign n26913 = n26512 & n26912 ;
  assign n26914 = n26911 | n26913 ;
  assign n26915 = n65877 & n26914 ;
  assign n74178 = ~n26386 ;
  assign n26388 = n26079 & n74178 ;
  assign n26916 = n26010 | n26079 ;
  assign n74179 = ~n26916 ;
  assign n26917 = n26075 & n74179 ;
  assign n26918 = n26388 | n26917 ;
  assign n26919 = n136 & n26918 ;
  assign n26920 = n26000 & n74024 ;
  assign n26921 = n26512 & n26920 ;
  assign n26922 = n26919 | n26921 ;
  assign n26923 = n65820 & n26922 ;
  assign n74180 = ~n26921 ;
  assign n27005 = x71 & n74180 ;
  assign n74181 = ~n26919 ;
  assign n27006 = n74181 & n27005 ;
  assign n27007 = n26923 | n27006 ;
  assign n74182 = ~n26070 ;
  assign n26074 = n74182 & n26073 ;
  assign n26924 = n26019 | n26073 ;
  assign n74183 = ~n26924 ;
  assign n26925 = n26383 & n74183 ;
  assign n26926 = n26074 | n26925 ;
  assign n26927 = n136 & n26926 ;
  assign n26928 = n26009 & n74024 ;
  assign n26929 = n26512 & n26928 ;
  assign n26930 = n26927 | n26929 ;
  assign n26931 = n65791 & n26930 ;
  assign n74184 = ~n26381 ;
  assign n26382 = n26068 & n74184 ;
  assign n26932 = n26028 | n26068 ;
  assign n74185 = ~n26932 ;
  assign n26933 = n26064 & n74185 ;
  assign n26934 = n26382 | n26933 ;
  assign n26935 = n136 & n26934 ;
  assign n26936 = n26018 & n74024 ;
  assign n26937 = n26512 & n26936 ;
  assign n26938 = n26935 | n26937 ;
  assign n26939 = n65772 & n26938 ;
  assign n74186 = ~n26937 ;
  assign n26994 = x69 & n74186 ;
  assign n74187 = ~n26935 ;
  assign n26995 = n74187 & n26994 ;
  assign n26996 = n26939 | n26995 ;
  assign n74188 = ~n26060 ;
  assign n26379 = n74188 & n26063 ;
  assign n26940 = n26036 | n26063 ;
  assign n74189 = ~n26940 ;
  assign n26941 = n26059 & n74189 ;
  assign n26942 = n26379 | n26941 ;
  assign n26943 = n136 & n26942 ;
  assign n26944 = n26027 & n74024 ;
  assign n26945 = n26512 & n26944 ;
  assign n26946 = n26943 | n26945 ;
  assign n26947 = n65746 & n26946 ;
  assign n74190 = ~n26055 ;
  assign n26949 = n74190 & n26058 ;
  assign n26948 = n26054 | n26058 ;
  assign n74191 = ~n26948 ;
  assign n26950 = n26053 & n74191 ;
  assign n26951 = n26949 | n26950 ;
  assign n26952 = n136 & n26951 ;
  assign n26953 = n26035 & n74024 ;
  assign n26954 = n26512 & n26953 ;
  assign n26955 = n26952 | n26954 ;
  assign n26956 = n65721 & n26955 ;
  assign n74192 = ~n26954 ;
  assign n26984 = x67 & n74192 ;
  assign n74193 = ~n26952 ;
  assign n26985 = n74193 & n26984 ;
  assign n26986 = n26956 | n26985 ;
  assign n26957 = n26050 & n26052 ;
  assign n26958 = n73856 & n26957 ;
  assign n74194 = ~n26958 ;
  assign n26959 = n26375 & n74194 ;
  assign n26960 = n136 & n26959 ;
  assign n26961 = n26047 & n74024 ;
  assign n26962 = n26512 & n26961 ;
  assign n26963 = n26960 | n26962 ;
  assign n26964 = n65686 & n26963 ;
  assign n74195 = ~x6 ;
  assign n26974 = n74195 & x64 ;
  assign n26370 = n26052 & n136 ;
  assign n26965 = n74024 & n26512 ;
  assign n74196 = ~n26965 ;
  assign n26966 = x64 & n74196 ;
  assign n74197 = ~n26966 ;
  assign n26967 = x7 & n74197 ;
  assign n26968 = n26370 | n26967 ;
  assign n26969 = x65 & n26968 ;
  assign n26371 = x64 & n136 ;
  assign n74198 = ~n26371 ;
  assign n26970 = x7 & n74198 ;
  assign n26971 = n26052 & n74196 ;
  assign n26972 = x65 | n26971 ;
  assign n26973 = n26970 | n26972 ;
  assign n74199 = ~n26969 ;
  assign n26975 = n74199 & n26973 ;
  assign n26976 = n26974 | n26975 ;
  assign n26977 = n26370 | n26970 ;
  assign n26978 = n65670 & n26977 ;
  assign n74200 = ~n26978 ;
  assign n26979 = n26976 & n74200 ;
  assign n74201 = ~n26962 ;
  assign n26980 = x66 & n74201 ;
  assign n74202 = ~n26960 ;
  assign n26981 = n74202 & n26980 ;
  assign n26982 = n26964 | n26981 ;
  assign n26983 = n26979 | n26982 ;
  assign n74203 = ~n26964 ;
  assign n26987 = n74203 & n26983 ;
  assign n26988 = n26986 | n26987 ;
  assign n74204 = ~n26956 ;
  assign n26989 = n74204 & n26988 ;
  assign n74205 = ~n26945 ;
  assign n26990 = x68 & n74205 ;
  assign n74206 = ~n26943 ;
  assign n26991 = n74206 & n26990 ;
  assign n26992 = n26947 | n26991 ;
  assign n26993 = n26989 | n26992 ;
  assign n74207 = ~n26947 ;
  assign n26997 = n74207 & n26993 ;
  assign n26998 = n26996 | n26997 ;
  assign n74208 = ~n26939 ;
  assign n26999 = n74208 & n26998 ;
  assign n74209 = ~n26929 ;
  assign n27000 = x70 & n74209 ;
  assign n74210 = ~n26927 ;
  assign n27001 = n74210 & n27000 ;
  assign n27002 = n26931 | n27001 ;
  assign n27004 = n26999 | n27002 ;
  assign n74211 = ~n26931 ;
  assign n27009 = n74211 & n27004 ;
  assign n27010 = n27007 | n27009 ;
  assign n74212 = ~n26923 ;
  assign n27011 = n74212 & n27010 ;
  assign n74213 = ~n26913 ;
  assign n27012 = x72 & n74213 ;
  assign n74214 = ~n26911 ;
  assign n27013 = n74214 & n27012 ;
  assign n27014 = n26915 | n27013 ;
  assign n27016 = n27011 | n27014 ;
  assign n74215 = ~n26915 ;
  assign n27021 = n74215 & n27016 ;
  assign n27022 = n27019 | n27021 ;
  assign n74216 = ~n26907 ;
  assign n27023 = n74216 & n27022 ;
  assign n74217 = ~n26897 ;
  assign n27024 = x74 & n74217 ;
  assign n74218 = ~n26895 ;
  assign n27025 = n74218 & n27024 ;
  assign n27026 = n26899 | n27025 ;
  assign n27028 = n27023 | n27026 ;
  assign n74219 = ~n26899 ;
  assign n27033 = n74219 & n27028 ;
  assign n27034 = n27031 | n27033 ;
  assign n74220 = ~n26891 ;
  assign n27035 = n74220 & n27034 ;
  assign n74221 = ~n26881 ;
  assign n27036 = x76 & n74221 ;
  assign n74222 = ~n26879 ;
  assign n27037 = n74222 & n27036 ;
  assign n27038 = n26883 | n27037 ;
  assign n27040 = n27035 | n27038 ;
  assign n74223 = ~n26883 ;
  assign n27045 = n74223 & n27040 ;
  assign n27046 = n27043 | n27045 ;
  assign n74224 = ~n26875 ;
  assign n27047 = n74224 & n27046 ;
  assign n74225 = ~n26865 ;
  assign n27048 = x78 & n74225 ;
  assign n74226 = ~n26863 ;
  assign n27049 = n74226 & n27048 ;
  assign n27050 = n26867 | n27049 ;
  assign n27052 = n27047 | n27050 ;
  assign n74227 = ~n26867 ;
  assign n27057 = n74227 & n27052 ;
  assign n27058 = n27055 | n27057 ;
  assign n74228 = ~n26859 ;
  assign n27059 = n74228 & n27058 ;
  assign n74229 = ~n26849 ;
  assign n27060 = x80 & n74229 ;
  assign n74230 = ~n26847 ;
  assign n27061 = n74230 & n27060 ;
  assign n27062 = n26851 | n27061 ;
  assign n27064 = n27059 | n27062 ;
  assign n74231 = ~n26851 ;
  assign n27069 = n74231 & n27064 ;
  assign n27070 = n27067 | n27069 ;
  assign n74232 = ~n26843 ;
  assign n27071 = n74232 & n27070 ;
  assign n74233 = ~n26833 ;
  assign n27072 = x82 & n74233 ;
  assign n74234 = ~n26831 ;
  assign n27073 = n74234 & n27072 ;
  assign n27074 = n26835 | n27073 ;
  assign n27076 = n27071 | n27074 ;
  assign n74235 = ~n26835 ;
  assign n27081 = n74235 & n27076 ;
  assign n27082 = n27079 | n27081 ;
  assign n74236 = ~n26827 ;
  assign n27083 = n74236 & n27082 ;
  assign n74237 = ~n26817 ;
  assign n27084 = x84 & n74237 ;
  assign n74238 = ~n26815 ;
  assign n27085 = n74238 & n27084 ;
  assign n27086 = n26819 | n27085 ;
  assign n27088 = n27083 | n27086 ;
  assign n74239 = ~n26819 ;
  assign n27093 = n74239 & n27088 ;
  assign n27094 = n27091 | n27093 ;
  assign n74240 = ~n26811 ;
  assign n27095 = n74240 & n27094 ;
  assign n74241 = ~n26801 ;
  assign n27096 = x86 & n74241 ;
  assign n74242 = ~n26799 ;
  assign n27097 = n74242 & n27096 ;
  assign n27098 = n26803 | n27097 ;
  assign n27100 = n27095 | n27098 ;
  assign n74243 = ~n26803 ;
  assign n27105 = n74243 & n27100 ;
  assign n27106 = n27103 | n27105 ;
  assign n74244 = ~n26795 ;
  assign n27107 = n74244 & n27106 ;
  assign n74245 = ~n26785 ;
  assign n27108 = x88 & n74245 ;
  assign n74246 = ~n26783 ;
  assign n27109 = n74246 & n27108 ;
  assign n27110 = n26787 | n27109 ;
  assign n27112 = n27107 | n27110 ;
  assign n74247 = ~n26787 ;
  assign n27117 = n74247 & n27112 ;
  assign n27118 = n27115 | n27117 ;
  assign n74248 = ~n26779 ;
  assign n27119 = n74248 & n27118 ;
  assign n74249 = ~n26769 ;
  assign n27120 = x90 & n74249 ;
  assign n74250 = ~n26767 ;
  assign n27121 = n74250 & n27120 ;
  assign n27122 = n26771 | n27121 ;
  assign n27124 = n27119 | n27122 ;
  assign n74251 = ~n26771 ;
  assign n27129 = n74251 & n27124 ;
  assign n27130 = n27127 | n27129 ;
  assign n74252 = ~n26763 ;
  assign n27131 = n74252 & n27130 ;
  assign n74253 = ~n26753 ;
  assign n27132 = x92 & n74253 ;
  assign n74254 = ~n26751 ;
  assign n27133 = n74254 & n27132 ;
  assign n27134 = n26755 | n27133 ;
  assign n27136 = n27131 | n27134 ;
  assign n74255 = ~n26755 ;
  assign n27141 = n74255 & n27136 ;
  assign n27142 = n27139 | n27141 ;
  assign n74256 = ~n26747 ;
  assign n27143 = n74256 & n27142 ;
  assign n74257 = ~n26737 ;
  assign n27144 = x94 & n74257 ;
  assign n74258 = ~n26735 ;
  assign n27145 = n74258 & n27144 ;
  assign n27146 = n26739 | n27145 ;
  assign n27148 = n27143 | n27146 ;
  assign n74259 = ~n26739 ;
  assign n27153 = n74259 & n27148 ;
  assign n27154 = n27151 | n27153 ;
  assign n74260 = ~n26731 ;
  assign n27155 = n74260 & n27154 ;
  assign n74261 = ~n26721 ;
  assign n27156 = x96 & n74261 ;
  assign n74262 = ~n26719 ;
  assign n27157 = n74262 & n27156 ;
  assign n27158 = n26723 | n27157 ;
  assign n27160 = n27155 | n27158 ;
  assign n74263 = ~n26723 ;
  assign n27165 = n74263 & n27160 ;
  assign n27166 = n27163 | n27165 ;
  assign n74264 = ~n26715 ;
  assign n27167 = n74264 & n27166 ;
  assign n74265 = ~n26705 ;
  assign n27168 = x98 & n74265 ;
  assign n74266 = ~n26703 ;
  assign n27169 = n74266 & n27168 ;
  assign n27170 = n26707 | n27169 ;
  assign n27172 = n27167 | n27170 ;
  assign n74267 = ~n26707 ;
  assign n27177 = n74267 & n27172 ;
  assign n27178 = n27175 | n27177 ;
  assign n74268 = ~n26699 ;
  assign n27179 = n74268 & n27178 ;
  assign n74269 = ~n26689 ;
  assign n27180 = x100 & n74269 ;
  assign n74270 = ~n26687 ;
  assign n27181 = n74270 & n27180 ;
  assign n27182 = n26691 | n27181 ;
  assign n27184 = n27179 | n27182 ;
  assign n74271 = ~n26691 ;
  assign n27189 = n74271 & n27184 ;
  assign n27190 = n27187 | n27189 ;
  assign n74272 = ~n26683 ;
  assign n27191 = n74272 & n27190 ;
  assign n74273 = ~n26673 ;
  assign n27192 = x102 & n74273 ;
  assign n74274 = ~n26671 ;
  assign n27193 = n74274 & n27192 ;
  assign n27194 = n26675 | n27193 ;
  assign n27196 = n27191 | n27194 ;
  assign n74275 = ~n26675 ;
  assign n27201 = n74275 & n27196 ;
  assign n27202 = n27199 | n27201 ;
  assign n74276 = ~n26667 ;
  assign n27203 = n74276 & n27202 ;
  assign n74277 = ~n26657 ;
  assign n27204 = x104 & n74277 ;
  assign n74278 = ~n26655 ;
  assign n27205 = n74278 & n27204 ;
  assign n27206 = n26659 | n27205 ;
  assign n27208 = n27203 | n27206 ;
  assign n74279 = ~n26659 ;
  assign n27213 = n74279 & n27208 ;
  assign n27214 = n27211 | n27213 ;
  assign n74280 = ~n26651 ;
  assign n27215 = n74280 & n27214 ;
  assign n74281 = ~n26641 ;
  assign n27216 = x106 & n74281 ;
  assign n74282 = ~n26639 ;
  assign n27217 = n74282 & n27216 ;
  assign n27218 = n26643 | n27217 ;
  assign n27220 = n27215 | n27218 ;
  assign n74283 = ~n26643 ;
  assign n27225 = n74283 & n27220 ;
  assign n27226 = n27223 | n27225 ;
  assign n74284 = ~n26635 ;
  assign n27227 = n74284 & n27226 ;
  assign n74285 = ~n26625 ;
  assign n27228 = x108 & n74285 ;
  assign n74286 = ~n26623 ;
  assign n27229 = n74286 & n27228 ;
  assign n27230 = n26627 | n27229 ;
  assign n27232 = n27227 | n27230 ;
  assign n74287 = ~n26627 ;
  assign n27237 = n74287 & n27232 ;
  assign n27238 = n27235 | n27237 ;
  assign n74288 = ~n26619 ;
  assign n27239 = n74288 & n27238 ;
  assign n74289 = ~n26609 ;
  assign n27240 = x110 & n74289 ;
  assign n74290 = ~n26607 ;
  assign n27241 = n74290 & n27240 ;
  assign n27242 = n26611 | n27241 ;
  assign n27244 = n27239 | n27242 ;
  assign n74291 = ~n26611 ;
  assign n27249 = n74291 & n27244 ;
  assign n27250 = n27247 | n27249 ;
  assign n74292 = ~n26603 ;
  assign n27251 = n74292 & n27250 ;
  assign n74293 = ~n26593 ;
  assign n27252 = x112 & n74293 ;
  assign n74294 = ~n26591 ;
  assign n27253 = n74294 & n27252 ;
  assign n27254 = n26595 | n27253 ;
  assign n27256 = n27251 | n27254 ;
  assign n74295 = ~n26595 ;
  assign n27261 = n74295 & n27256 ;
  assign n27262 = n27259 | n27261 ;
  assign n74296 = ~n26587 ;
  assign n27263 = n74296 & n27262 ;
  assign n74297 = ~n26577 ;
  assign n27264 = x114 & n74297 ;
  assign n74298 = ~n26575 ;
  assign n27265 = n74298 & n27264 ;
  assign n27266 = n26579 | n27265 ;
  assign n27268 = n27263 | n27266 ;
  assign n74299 = ~n26579 ;
  assign n27273 = n74299 & n27268 ;
  assign n27274 = n27271 | n27273 ;
  assign n74300 = ~n26571 ;
  assign n27275 = n74300 & n27274 ;
  assign n74301 = ~n26561 ;
  assign n27276 = x116 & n74301 ;
  assign n74302 = ~n26559 ;
  assign n27277 = n74302 & n27276 ;
  assign n27278 = n26563 | n27277 ;
  assign n27280 = n27275 | n27278 ;
  assign n74303 = ~n26563 ;
  assign n27285 = n74303 & n27280 ;
  assign n27286 = n27283 | n27285 ;
  assign n74304 = ~n26555 ;
  assign n27287 = n74304 & n27286 ;
  assign n74305 = ~n26545 ;
  assign n27288 = x118 & n74305 ;
  assign n74306 = ~n26543 ;
  assign n27289 = n74306 & n27288 ;
  assign n27290 = n26547 | n27289 ;
  assign n27292 = n27287 | n27290 ;
  assign n74307 = ~n26547 ;
  assign n27297 = n74307 & n27292 ;
  assign n27298 = n27295 | n27297 ;
  assign n74308 = ~n26539 ;
  assign n27299 = n74308 & n27298 ;
  assign n74309 = ~n26529 ;
  assign n27300 = x120 & n74309 ;
  assign n74310 = ~n26527 ;
  assign n27301 = n74310 & n27300 ;
  assign n27302 = n26531 | n27301 ;
  assign n27304 = n27299 | n27302 ;
  assign n74311 = ~n26531 ;
  assign n27308 = n74311 & n27304 ;
  assign n27309 = n27307 | n27308 ;
  assign n74312 = ~n26523 ;
  assign n27310 = n74312 & n27309 ;
  assign n27312 = n27310 | n27311 ;
  assign n74313 = ~n26522 ;
  assign n27313 = n74313 & n27312 ;
  assign n74314 = ~n27308 ;
  assign n28206 = n27307 & n74314 ;
  assign n27317 = x65 & n26977 ;
  assign n74315 = ~n27317 ;
  assign n27318 = n26973 & n74315 ;
  assign n27320 = n26974 | n27318 ;
  assign n27322 = n74200 & n27320 ;
  assign n27323 = n26982 | n27322 ;
  assign n27324 = n74203 & n27323 ;
  assign n27325 = n26986 | n27324 ;
  assign n27326 = n74204 & n27325 ;
  assign n27327 = n26992 | n27326 ;
  assign n27328 = n74207 & n27327 ;
  assign n27329 = n26996 | n27328 ;
  assign n27330 = n74208 & n27329 ;
  assign n27331 = n27002 | n27330 ;
  assign n27332 = n74211 & n27331 ;
  assign n27333 = n27007 | n27332 ;
  assign n27334 = n74212 & n27333 ;
  assign n27335 = n27014 | n27334 ;
  assign n27336 = n74215 & n27335 ;
  assign n27337 = n27019 | n27336 ;
  assign n27338 = n74216 & n27337 ;
  assign n27339 = n27026 | n27338 ;
  assign n27340 = n74219 & n27339 ;
  assign n27341 = n27031 | n27340 ;
  assign n27342 = n74220 & n27341 ;
  assign n27343 = n27038 | n27342 ;
  assign n27344 = n74223 & n27343 ;
  assign n27345 = n27043 | n27344 ;
  assign n27346 = n74224 & n27345 ;
  assign n27347 = n27050 | n27346 ;
  assign n27348 = n74227 & n27347 ;
  assign n27349 = n27055 | n27348 ;
  assign n27350 = n74228 & n27349 ;
  assign n27351 = n27062 | n27350 ;
  assign n27352 = n74231 & n27351 ;
  assign n27353 = n27067 | n27352 ;
  assign n27354 = n74232 & n27353 ;
  assign n27355 = n27074 | n27354 ;
  assign n27356 = n74235 & n27355 ;
  assign n27357 = n27079 | n27356 ;
  assign n27358 = n74236 & n27357 ;
  assign n27359 = n27086 | n27358 ;
  assign n27360 = n74239 & n27359 ;
  assign n27361 = n27091 | n27360 ;
  assign n27362 = n74240 & n27361 ;
  assign n27363 = n27098 | n27362 ;
  assign n27364 = n74243 & n27363 ;
  assign n27365 = n27103 | n27364 ;
  assign n27366 = n74244 & n27365 ;
  assign n27367 = n27110 | n27366 ;
  assign n27368 = n74247 & n27367 ;
  assign n27369 = n27115 | n27368 ;
  assign n27370 = n74248 & n27369 ;
  assign n27371 = n27122 | n27370 ;
  assign n27372 = n74251 & n27371 ;
  assign n27373 = n27127 | n27372 ;
  assign n27374 = n74252 & n27373 ;
  assign n27375 = n27134 | n27374 ;
  assign n27376 = n74255 & n27375 ;
  assign n27377 = n27139 | n27376 ;
  assign n27378 = n74256 & n27377 ;
  assign n27379 = n27146 | n27378 ;
  assign n27380 = n74259 & n27379 ;
  assign n27381 = n27151 | n27380 ;
  assign n27382 = n74260 & n27381 ;
  assign n27383 = n27158 | n27382 ;
  assign n27384 = n74263 & n27383 ;
  assign n27385 = n27163 | n27384 ;
  assign n27386 = n74264 & n27385 ;
  assign n27387 = n27170 | n27386 ;
  assign n27388 = n74267 & n27387 ;
  assign n27389 = n27175 | n27388 ;
  assign n27390 = n74268 & n27389 ;
  assign n27391 = n27182 | n27390 ;
  assign n27392 = n74271 & n27391 ;
  assign n27393 = n27187 | n27392 ;
  assign n27394 = n74272 & n27393 ;
  assign n27395 = n27194 | n27394 ;
  assign n27396 = n74275 & n27395 ;
  assign n27397 = n27199 | n27396 ;
  assign n27398 = n74276 & n27397 ;
  assign n27399 = n27206 | n27398 ;
  assign n27400 = n74279 & n27399 ;
  assign n27401 = n27211 | n27400 ;
  assign n27402 = n74280 & n27401 ;
  assign n27403 = n27218 | n27402 ;
  assign n27404 = n74283 & n27403 ;
  assign n27405 = n27223 | n27404 ;
  assign n27406 = n74284 & n27405 ;
  assign n27407 = n27230 | n27406 ;
  assign n27408 = n74287 & n27407 ;
  assign n27409 = n27235 | n27408 ;
  assign n27410 = n74288 & n27409 ;
  assign n27411 = n27242 | n27410 ;
  assign n27412 = n74291 & n27411 ;
  assign n27413 = n27247 | n27412 ;
  assign n27414 = n74292 & n27413 ;
  assign n27415 = n27254 | n27414 ;
  assign n27416 = n74295 & n27415 ;
  assign n27417 = n27259 | n27416 ;
  assign n27418 = n74296 & n27417 ;
  assign n27419 = n27266 | n27418 ;
  assign n27420 = n74299 & n27419 ;
  assign n27421 = n27271 | n27420 ;
  assign n27422 = n74300 & n27421 ;
  assign n27423 = n27278 | n27422 ;
  assign n27424 = n74303 & n27423 ;
  assign n27425 = n27283 | n27424 ;
  assign n27426 = n74304 & n27425 ;
  assign n27427 = n27290 | n27426 ;
  assign n27428 = n74307 & n27427 ;
  assign n27429 = n27295 | n27428 ;
  assign n27431 = n74308 & n27429 ;
  assign n27883 = n27302 | n27431 ;
  assign n28207 = n26531 | n27307 ;
  assign n74316 = ~n28207 ;
  assign n28208 = n27883 & n74316 ;
  assign n28209 = n28206 | n28208 ;
  assign n28210 = n27312 | n28209 ;
  assign n74317 = ~n27313 ;
  assign n28211 = n74317 & n28210 ;
  assign n74318 = ~n27311 ;
  assign n28220 = n74318 & n28211 ;
  assign n27315 = n26530 & n27312 ;
  assign n27303 = n26539 | n27302 ;
  assign n74319 = ~n27303 ;
  assign n27430 = n74319 & n27429 ;
  assign n74320 = ~n27431 ;
  assign n27432 = n27302 & n74320 ;
  assign n27433 = n27430 | n27432 ;
  assign n27434 = n74318 & n27433 ;
  assign n74321 = ~n27310 ;
  assign n27435 = n74321 & n27434 ;
  assign n27436 = n27315 | n27435 ;
  assign n27437 = n74029 & n27436 ;
  assign n27438 = n26538 & n27312 ;
  assign n27296 = n26547 | n27295 ;
  assign n74322 = ~n27296 ;
  assign n27439 = n27292 & n74322 ;
  assign n74323 = ~n27297 ;
  assign n27440 = n27295 & n74323 ;
  assign n27441 = n27439 | n27440 ;
  assign n27442 = n74318 & n27441 ;
  assign n27443 = n74321 & n27442 ;
  assign n27444 = n27438 | n27443 ;
  assign n27445 = n74021 & n27444 ;
  assign n27446 = n26546 & n27312 ;
  assign n27291 = n26555 | n27290 ;
  assign n74324 = ~n27291 ;
  assign n27447 = n74324 & n27425 ;
  assign n74325 = ~n27426 ;
  assign n27448 = n27290 & n74325 ;
  assign n27449 = n27447 | n27448 ;
  assign n27450 = n74318 & n27449 ;
  assign n27451 = n74321 & n27450 ;
  assign n27452 = n27446 | n27451 ;
  assign n27453 = n73617 & n27452 ;
  assign n27454 = n26554 & n27312 ;
  assign n27284 = n26563 | n27283 ;
  assign n74326 = ~n27284 ;
  assign n27455 = n27280 & n74326 ;
  assign n74327 = ~n27285 ;
  assign n27456 = n27283 & n74327 ;
  assign n27457 = n27455 | n27456 ;
  assign n27458 = n74318 & n27457 ;
  assign n27459 = n74321 & n27458 ;
  assign n27460 = n27454 | n27459 ;
  assign n27461 = n73188 & n27460 ;
  assign n27462 = n26562 & n27312 ;
  assign n27279 = n26571 | n27278 ;
  assign n74328 = ~n27279 ;
  assign n27463 = n74328 & n27421 ;
  assign n74329 = ~n27422 ;
  assign n27464 = n27278 & n74329 ;
  assign n27465 = n27463 | n27464 ;
  assign n27466 = n74318 & n27465 ;
  assign n27467 = n74321 & n27466 ;
  assign n27468 = n27462 | n27467 ;
  assign n27469 = n73177 & n27468 ;
  assign n27470 = n26570 & n27312 ;
  assign n27272 = n26579 | n27271 ;
  assign n74330 = ~n27272 ;
  assign n27471 = n27268 & n74330 ;
  assign n74331 = ~n27273 ;
  assign n27472 = n27271 & n74331 ;
  assign n27473 = n27471 | n27472 ;
  assign n27474 = n74318 & n27473 ;
  assign n27475 = n74321 & n27474 ;
  assign n27476 = n27470 | n27475 ;
  assign n27477 = n72752 & n27476 ;
  assign n27478 = n26578 & n27312 ;
  assign n27267 = n26587 | n27266 ;
  assign n74332 = ~n27267 ;
  assign n27479 = n74332 & n27417 ;
  assign n74333 = ~n27418 ;
  assign n27480 = n27266 & n74333 ;
  assign n27481 = n27479 | n27480 ;
  assign n27482 = n74318 & n27481 ;
  assign n27483 = n74321 & n27482 ;
  assign n27484 = n27478 | n27483 ;
  assign n27485 = n72393 & n27484 ;
  assign n27486 = n26586 & n27312 ;
  assign n27260 = n26595 | n27259 ;
  assign n74334 = ~n27260 ;
  assign n27487 = n27256 & n74334 ;
  assign n74335 = ~n27261 ;
  assign n27488 = n27259 & n74335 ;
  assign n27489 = n27487 | n27488 ;
  assign n27490 = n74318 & n27489 ;
  assign n27491 = n74321 & n27490 ;
  assign n27492 = n27486 | n27491 ;
  assign n27493 = n72385 & n27492 ;
  assign n27494 = n26594 & n27312 ;
  assign n27255 = n26603 | n27254 ;
  assign n74336 = ~n27255 ;
  assign n27495 = n74336 & n27413 ;
  assign n74337 = ~n27414 ;
  assign n27496 = n27254 & n74337 ;
  assign n27497 = n27495 | n27496 ;
  assign n27498 = n74318 & n27497 ;
  assign n27499 = n74321 & n27498 ;
  assign n27500 = n27494 | n27499 ;
  assign n27501 = n72025 & n27500 ;
  assign n27502 = n26602 & n27312 ;
  assign n27248 = n26611 | n27247 ;
  assign n74338 = ~n27248 ;
  assign n27503 = n27244 & n74338 ;
  assign n74339 = ~n27249 ;
  assign n27504 = n27247 & n74339 ;
  assign n27505 = n27503 | n27504 ;
  assign n27506 = n74318 & n27505 ;
  assign n27507 = n74321 & n27506 ;
  assign n27508 = n27502 | n27507 ;
  assign n27509 = n71645 & n27508 ;
  assign n27510 = n26610 & n27312 ;
  assign n27243 = n26619 | n27242 ;
  assign n74340 = ~n27243 ;
  assign n27511 = n74340 & n27409 ;
  assign n74341 = ~n27410 ;
  assign n27512 = n27242 & n74341 ;
  assign n27513 = n27511 | n27512 ;
  assign n27514 = n74318 & n27513 ;
  assign n27515 = n74321 & n27514 ;
  assign n27516 = n27510 | n27515 ;
  assign n27517 = n71633 & n27516 ;
  assign n27518 = n26618 & n27312 ;
  assign n27236 = n26627 | n27235 ;
  assign n74342 = ~n27236 ;
  assign n27519 = n27232 & n74342 ;
  assign n74343 = ~n27237 ;
  assign n27520 = n27235 & n74343 ;
  assign n27521 = n27519 | n27520 ;
  assign n27522 = n74318 & n27521 ;
  assign n27523 = n74321 & n27522 ;
  assign n27524 = n27518 | n27523 ;
  assign n27525 = n71253 & n27524 ;
  assign n27526 = n26626 & n27312 ;
  assign n27231 = n26635 | n27230 ;
  assign n74344 = ~n27231 ;
  assign n27527 = n74344 & n27405 ;
  assign n74345 = ~n27406 ;
  assign n27528 = n27230 & n74345 ;
  assign n27529 = n27527 | n27528 ;
  assign n27530 = n74318 & n27529 ;
  assign n27531 = n74321 & n27530 ;
  assign n27532 = n27526 | n27531 ;
  assign n27533 = n70935 & n27532 ;
  assign n27534 = n26634 & n27312 ;
  assign n27224 = n26643 | n27223 ;
  assign n74346 = ~n27224 ;
  assign n27535 = n27220 & n74346 ;
  assign n74347 = ~n27225 ;
  assign n27536 = n27223 & n74347 ;
  assign n27537 = n27535 | n27536 ;
  assign n27538 = n74318 & n27537 ;
  assign n27539 = n74321 & n27538 ;
  assign n27540 = n27534 | n27539 ;
  assign n27541 = n70927 & n27540 ;
  assign n27542 = n26642 & n27312 ;
  assign n27219 = n26651 | n27218 ;
  assign n74348 = ~n27219 ;
  assign n27543 = n74348 & n27401 ;
  assign n74349 = ~n27402 ;
  assign n27544 = n27218 & n74349 ;
  assign n27545 = n27543 | n27544 ;
  assign n27546 = n74318 & n27545 ;
  assign n27547 = n74321 & n27546 ;
  assign n27548 = n27542 | n27547 ;
  assign n27549 = n70609 & n27548 ;
  assign n27550 = n26650 & n27312 ;
  assign n27212 = n26659 | n27211 ;
  assign n74350 = ~n27212 ;
  assign n27551 = n27208 & n74350 ;
  assign n74351 = ~n27213 ;
  assign n27552 = n27211 & n74351 ;
  assign n27553 = n27551 | n27552 ;
  assign n27554 = n74318 & n27553 ;
  assign n27555 = n74321 & n27554 ;
  assign n27556 = n27550 | n27555 ;
  assign n27557 = n70276 & n27556 ;
  assign n27558 = n26658 & n27312 ;
  assign n27207 = n26667 | n27206 ;
  assign n74352 = ~n27207 ;
  assign n27559 = n74352 & n27397 ;
  assign n74353 = ~n27398 ;
  assign n27560 = n27206 & n74353 ;
  assign n27561 = n27559 | n27560 ;
  assign n27562 = n74318 & n27561 ;
  assign n27563 = n74321 & n27562 ;
  assign n27564 = n27558 | n27563 ;
  assign n27565 = n70176 & n27564 ;
  assign n27566 = n26666 & n27312 ;
  assign n27200 = n26675 | n27199 ;
  assign n74354 = ~n27200 ;
  assign n27567 = n27196 & n74354 ;
  assign n74355 = ~n27201 ;
  assign n27568 = n27199 & n74355 ;
  assign n27569 = n27567 | n27568 ;
  assign n27570 = n74318 & n27569 ;
  assign n27571 = n74321 & n27570 ;
  assign n27572 = n27566 | n27571 ;
  assign n27573 = n69857 & n27572 ;
  assign n27574 = n26674 & n27312 ;
  assign n27195 = n26683 | n27194 ;
  assign n74356 = ~n27195 ;
  assign n27575 = n74356 & n27393 ;
  assign n74357 = ~n27394 ;
  assign n27576 = n27194 & n74357 ;
  assign n27577 = n27575 | n27576 ;
  assign n27578 = n74318 & n27577 ;
  assign n27579 = n74321 & n27578 ;
  assign n27580 = n27574 | n27579 ;
  assign n27581 = n69656 & n27580 ;
  assign n27582 = n26682 & n27312 ;
  assign n27188 = n26691 | n27187 ;
  assign n74358 = ~n27188 ;
  assign n27583 = n27184 & n74358 ;
  assign n74359 = ~n27189 ;
  assign n27584 = n27187 & n74359 ;
  assign n27585 = n27583 | n27584 ;
  assign n27586 = n74318 & n27585 ;
  assign n27587 = n74321 & n27586 ;
  assign n27588 = n27582 | n27587 ;
  assign n27589 = n69528 & n27588 ;
  assign n27590 = n26690 & n27312 ;
  assign n27183 = n26699 | n27182 ;
  assign n74360 = ~n27183 ;
  assign n27591 = n74360 & n27389 ;
  assign n74361 = ~n27390 ;
  assign n27592 = n27182 & n74361 ;
  assign n27593 = n27591 | n27592 ;
  assign n27594 = n74318 & n27593 ;
  assign n27595 = n74321 & n27594 ;
  assign n27596 = n27590 | n27595 ;
  assign n27597 = n69261 & n27596 ;
  assign n27598 = n26698 & n27312 ;
  assign n27176 = n26707 | n27175 ;
  assign n74362 = ~n27176 ;
  assign n27599 = n27172 & n74362 ;
  assign n74363 = ~n27177 ;
  assign n27600 = n27175 & n74363 ;
  assign n27601 = n27599 | n27600 ;
  assign n27602 = n74318 & n27601 ;
  assign n27603 = n74321 & n27602 ;
  assign n27604 = n27598 | n27603 ;
  assign n27605 = n69075 & n27604 ;
  assign n27606 = n26706 & n27312 ;
  assign n27171 = n26715 | n27170 ;
  assign n74364 = ~n27171 ;
  assign n27607 = n74364 & n27385 ;
  assign n74365 = ~n27386 ;
  assign n27608 = n27170 & n74365 ;
  assign n27609 = n27607 | n27608 ;
  assign n27610 = n74318 & n27609 ;
  assign n27611 = n74321 & n27610 ;
  assign n27612 = n27606 | n27611 ;
  assign n27613 = n68993 & n27612 ;
  assign n27614 = n26714 & n27312 ;
  assign n27164 = n26723 | n27163 ;
  assign n74366 = ~n27164 ;
  assign n27615 = n27160 & n74366 ;
  assign n74367 = ~n27165 ;
  assign n27616 = n27163 & n74367 ;
  assign n27617 = n27615 | n27616 ;
  assign n27618 = n74318 & n27617 ;
  assign n27619 = n74321 & n27618 ;
  assign n27620 = n27614 | n27619 ;
  assign n27621 = n68716 & n27620 ;
  assign n27622 = n26722 & n27312 ;
  assign n27159 = n26731 | n27158 ;
  assign n74368 = ~n27159 ;
  assign n27623 = n74368 & n27381 ;
  assign n74369 = ~n27382 ;
  assign n27624 = n27158 & n74369 ;
  assign n27625 = n27623 | n27624 ;
  assign n27626 = n74318 & n27625 ;
  assign n27627 = n74321 & n27626 ;
  assign n27628 = n27622 | n27627 ;
  assign n27629 = n68545 & n27628 ;
  assign n27630 = n26730 & n27312 ;
  assign n27152 = n26739 | n27151 ;
  assign n74370 = ~n27152 ;
  assign n27631 = n27148 & n74370 ;
  assign n74371 = ~n27153 ;
  assign n27632 = n27151 & n74371 ;
  assign n27633 = n27631 | n27632 ;
  assign n27634 = n74318 & n27633 ;
  assign n27635 = n74321 & n27634 ;
  assign n27636 = n27630 | n27635 ;
  assign n27637 = n68438 & n27636 ;
  assign n27638 = n26738 & n27312 ;
  assign n27147 = n26747 | n27146 ;
  assign n74372 = ~n27147 ;
  assign n27639 = n74372 & n27377 ;
  assign n74373 = ~n27378 ;
  assign n27640 = n27146 & n74373 ;
  assign n27641 = n27639 | n27640 ;
  assign n27642 = n74318 & n27641 ;
  assign n27643 = n74321 & n27642 ;
  assign n27644 = n27638 | n27643 ;
  assign n27645 = n68214 & n27644 ;
  assign n27646 = n26746 & n27312 ;
  assign n27140 = n26755 | n27139 ;
  assign n74374 = ~n27140 ;
  assign n27647 = n27136 & n74374 ;
  assign n74375 = ~n27141 ;
  assign n27648 = n27139 & n74375 ;
  assign n27649 = n27647 | n27648 ;
  assign n27650 = n74318 & n27649 ;
  assign n27651 = n74321 & n27650 ;
  assign n27652 = n27646 | n27651 ;
  assign n27653 = n68058 & n27652 ;
  assign n27654 = n26754 & n27312 ;
  assign n27135 = n26763 | n27134 ;
  assign n74376 = ~n27135 ;
  assign n27655 = n74376 & n27373 ;
  assign n74377 = ~n27374 ;
  assign n27656 = n27134 & n74377 ;
  assign n27657 = n27655 | n27656 ;
  assign n27658 = n74318 & n27657 ;
  assign n27659 = n74321 & n27658 ;
  assign n27660 = n27654 | n27659 ;
  assign n27661 = n67986 & n27660 ;
  assign n27662 = n26762 & n27312 ;
  assign n27128 = n26771 | n27127 ;
  assign n74378 = ~n27128 ;
  assign n27663 = n27124 & n74378 ;
  assign n74379 = ~n27129 ;
  assign n27664 = n27127 & n74379 ;
  assign n27665 = n27663 | n27664 ;
  assign n27666 = n74318 & n27665 ;
  assign n27667 = n74321 & n27666 ;
  assign n27668 = n27662 | n27667 ;
  assign n27669 = n67763 & n27668 ;
  assign n27670 = n26770 & n27312 ;
  assign n27123 = n26779 | n27122 ;
  assign n74380 = ~n27123 ;
  assign n27671 = n74380 & n27369 ;
  assign n74381 = ~n27370 ;
  assign n27672 = n27122 & n74381 ;
  assign n27673 = n27671 | n27672 ;
  assign n27674 = n74318 & n27673 ;
  assign n27675 = n74321 & n27674 ;
  assign n27676 = n27670 | n27675 ;
  assign n27677 = n67622 & n27676 ;
  assign n27678 = n26778 & n27312 ;
  assign n27116 = n26787 | n27115 ;
  assign n74382 = ~n27116 ;
  assign n27679 = n27112 & n74382 ;
  assign n74383 = ~n27117 ;
  assign n27680 = n27115 & n74383 ;
  assign n27681 = n27679 | n27680 ;
  assign n27682 = n74318 & n27681 ;
  assign n27683 = n74321 & n27682 ;
  assign n27684 = n27678 | n27683 ;
  assign n27685 = n67531 & n27684 ;
  assign n27686 = n26786 & n27312 ;
  assign n27111 = n26795 | n27110 ;
  assign n74384 = ~n27111 ;
  assign n27687 = n74384 & n27365 ;
  assign n74385 = ~n27366 ;
  assign n27688 = n27110 & n74385 ;
  assign n27689 = n27687 | n27688 ;
  assign n27690 = n74318 & n27689 ;
  assign n27691 = n74321 & n27690 ;
  assign n27692 = n27686 | n27691 ;
  assign n27693 = n67348 & n27692 ;
  assign n27694 = n26794 & n27312 ;
  assign n27104 = n26803 | n27103 ;
  assign n74386 = ~n27104 ;
  assign n27695 = n27100 & n74386 ;
  assign n74387 = ~n27105 ;
  assign n27696 = n27103 & n74387 ;
  assign n27697 = n27695 | n27696 ;
  assign n27698 = n74318 & n27697 ;
  assign n27699 = n74321 & n27698 ;
  assign n27700 = n27694 | n27699 ;
  assign n27701 = n67222 & n27700 ;
  assign n27702 = n26802 & n27312 ;
  assign n27099 = n26811 | n27098 ;
  assign n74388 = ~n27099 ;
  assign n27703 = n74388 & n27361 ;
  assign n74389 = ~n27362 ;
  assign n27704 = n27098 & n74389 ;
  assign n27705 = n27703 | n27704 ;
  assign n27706 = n74318 & n27705 ;
  assign n27707 = n74321 & n27706 ;
  assign n27708 = n27702 | n27707 ;
  assign n27709 = n67164 & n27708 ;
  assign n27710 = n26810 & n27312 ;
  assign n27092 = n26819 | n27091 ;
  assign n74390 = ~n27092 ;
  assign n27711 = n27088 & n74390 ;
  assign n74391 = ~n27093 ;
  assign n27712 = n27091 & n74391 ;
  assign n27713 = n27711 | n27712 ;
  assign n27714 = n74318 & n27713 ;
  assign n27715 = n74321 & n27714 ;
  assign n27716 = n27710 | n27715 ;
  assign n27717 = n66979 & n27716 ;
  assign n27718 = n26818 & n27312 ;
  assign n27087 = n26827 | n27086 ;
  assign n74392 = ~n27087 ;
  assign n27719 = n74392 & n27357 ;
  assign n74393 = ~n27358 ;
  assign n27720 = n27086 & n74393 ;
  assign n27721 = n27719 | n27720 ;
  assign n27722 = n74318 & n27721 ;
  assign n27723 = n74321 & n27722 ;
  assign n27724 = n27718 | n27723 ;
  assign n27725 = n66868 & n27724 ;
  assign n27726 = n26826 & n27312 ;
  assign n27080 = n26835 | n27079 ;
  assign n74394 = ~n27080 ;
  assign n27727 = n27076 & n74394 ;
  assign n74395 = ~n27081 ;
  assign n27728 = n27079 & n74395 ;
  assign n27729 = n27727 | n27728 ;
  assign n27730 = n74318 & n27729 ;
  assign n27731 = n74321 & n27730 ;
  assign n27732 = n27726 | n27731 ;
  assign n27733 = n66797 & n27732 ;
  assign n27734 = n26834 & n27312 ;
  assign n27075 = n26843 | n27074 ;
  assign n74396 = ~n27075 ;
  assign n27735 = n74396 & n27353 ;
  assign n74397 = ~n27354 ;
  assign n27736 = n27074 & n74397 ;
  assign n27737 = n27735 | n27736 ;
  assign n27738 = n74318 & n27737 ;
  assign n27739 = n74321 & n27738 ;
  assign n27740 = n27734 | n27739 ;
  assign n27741 = n66654 & n27740 ;
  assign n27742 = n26842 & n27312 ;
  assign n27068 = n26851 | n27067 ;
  assign n74398 = ~n27068 ;
  assign n27743 = n27064 & n74398 ;
  assign n74399 = ~n27069 ;
  assign n27744 = n27067 & n74399 ;
  assign n27745 = n27743 | n27744 ;
  assign n27746 = n74318 & n27745 ;
  assign n27747 = n74321 & n27746 ;
  assign n27748 = n27742 | n27747 ;
  assign n27749 = n66560 & n27748 ;
  assign n27750 = n26850 & n27312 ;
  assign n27063 = n26859 | n27062 ;
  assign n74400 = ~n27063 ;
  assign n27751 = n74400 & n27349 ;
  assign n74401 = ~n27350 ;
  assign n27752 = n27062 & n74401 ;
  assign n27753 = n27751 | n27752 ;
  assign n27754 = n74318 & n27753 ;
  assign n27755 = n74321 & n27754 ;
  assign n27756 = n27750 | n27755 ;
  assign n27757 = n66505 & n27756 ;
  assign n27758 = n26858 & n27312 ;
  assign n27056 = n26867 | n27055 ;
  assign n74402 = ~n27056 ;
  assign n27759 = n27052 & n74402 ;
  assign n74403 = ~n27057 ;
  assign n27760 = n27055 & n74403 ;
  assign n27761 = n27759 | n27760 ;
  assign n27762 = n74318 & n27761 ;
  assign n27763 = n74321 & n27762 ;
  assign n27764 = n27758 | n27763 ;
  assign n27765 = n66379 & n27764 ;
  assign n27766 = n26866 & n27312 ;
  assign n27051 = n26875 | n27050 ;
  assign n74404 = ~n27051 ;
  assign n27767 = n74404 & n27345 ;
  assign n74405 = ~n27346 ;
  assign n27768 = n27050 & n74405 ;
  assign n27769 = n27767 | n27768 ;
  assign n27770 = n74318 & n27769 ;
  assign n27771 = n74321 & n27770 ;
  assign n27772 = n27766 | n27771 ;
  assign n27773 = n66299 & n27772 ;
  assign n27774 = n26874 & n27312 ;
  assign n27044 = n26883 | n27043 ;
  assign n74406 = ~n27044 ;
  assign n27775 = n27040 & n74406 ;
  assign n74407 = ~n27045 ;
  assign n27776 = n27043 & n74407 ;
  assign n27777 = n27775 | n27776 ;
  assign n27778 = n74318 & n27777 ;
  assign n27779 = n74321 & n27778 ;
  assign n27780 = n27774 | n27779 ;
  assign n27781 = n66244 & n27780 ;
  assign n27782 = n26882 & n27312 ;
  assign n27039 = n26891 | n27038 ;
  assign n74408 = ~n27039 ;
  assign n27783 = n74408 & n27341 ;
  assign n74409 = ~n27342 ;
  assign n27784 = n27038 & n74409 ;
  assign n27785 = n27783 | n27784 ;
  assign n27786 = n74318 & n27785 ;
  assign n27787 = n74321 & n27786 ;
  assign n27788 = n27782 | n27787 ;
  assign n27789 = n66145 & n27788 ;
  assign n27790 = n26890 & n27312 ;
  assign n27032 = n26899 | n27031 ;
  assign n74410 = ~n27032 ;
  assign n27791 = n27028 & n74410 ;
  assign n74411 = ~n27033 ;
  assign n27792 = n27031 & n74411 ;
  assign n27793 = n27791 | n27792 ;
  assign n27794 = n74318 & n27793 ;
  assign n27795 = n74321 & n27794 ;
  assign n27796 = n27790 | n27795 ;
  assign n27797 = n66081 & n27796 ;
  assign n27798 = n26898 & n27312 ;
  assign n27027 = n26907 | n27026 ;
  assign n74412 = ~n27027 ;
  assign n27799 = n74412 & n27337 ;
  assign n74413 = ~n27338 ;
  assign n27800 = n27026 & n74413 ;
  assign n27801 = n27799 | n27800 ;
  assign n27802 = n74318 & n27801 ;
  assign n27803 = n74321 & n27802 ;
  assign n27804 = n27798 | n27803 ;
  assign n27805 = n66043 & n27804 ;
  assign n27806 = n26906 & n27312 ;
  assign n27020 = n26915 | n27019 ;
  assign n74414 = ~n27020 ;
  assign n27807 = n27016 & n74414 ;
  assign n74415 = ~n27021 ;
  assign n27808 = n27019 & n74415 ;
  assign n27809 = n27807 | n27808 ;
  assign n27810 = n74318 & n27809 ;
  assign n27811 = n74321 & n27810 ;
  assign n27812 = n27806 | n27811 ;
  assign n27813 = n65960 & n27812 ;
  assign n27814 = n26914 & n27312 ;
  assign n27015 = n26923 | n27014 ;
  assign n74416 = ~n27015 ;
  assign n27815 = n74416 & n27333 ;
  assign n74417 = ~n27334 ;
  assign n27816 = n27014 & n74417 ;
  assign n27817 = n27815 | n27816 ;
  assign n27818 = n74318 & n27817 ;
  assign n27819 = n74321 & n27818 ;
  assign n27820 = n27814 | n27819 ;
  assign n27821 = n65909 & n27820 ;
  assign n27822 = n26922 & n27312 ;
  assign n27008 = n26931 | n27007 ;
  assign n74418 = ~n27008 ;
  assign n27823 = n27004 & n74418 ;
  assign n74419 = ~n27009 ;
  assign n27824 = n27007 & n74419 ;
  assign n27825 = n27823 | n27824 ;
  assign n27826 = n74318 & n27825 ;
  assign n27827 = n74321 & n27826 ;
  assign n27828 = n27822 | n27827 ;
  assign n27829 = n65877 & n27828 ;
  assign n27830 = n26930 & n27312 ;
  assign n27003 = n26939 | n27002 ;
  assign n74420 = ~n27003 ;
  assign n27831 = n74420 & n27329 ;
  assign n74421 = ~n27330 ;
  assign n27832 = n27002 & n74421 ;
  assign n27833 = n27831 | n27832 ;
  assign n27834 = n74318 & n27833 ;
  assign n27835 = n74321 & n27834 ;
  assign n27836 = n27830 | n27835 ;
  assign n27837 = n65820 & n27836 ;
  assign n27838 = n26938 & n27312 ;
  assign n27316 = n26947 | n26996 ;
  assign n74422 = ~n27316 ;
  assign n27839 = n26993 & n74422 ;
  assign n74423 = ~n26997 ;
  assign n27840 = n26996 & n74423 ;
  assign n27841 = n27839 | n27840 ;
  assign n27842 = n74318 & n27841 ;
  assign n27843 = n74321 & n27842 ;
  assign n27844 = n27838 | n27843 ;
  assign n27845 = n65791 & n27844 ;
  assign n27846 = n26946 & n27312 ;
  assign n27847 = n26956 | n26992 ;
  assign n74424 = ~n27847 ;
  assign n27848 = n27325 & n74424 ;
  assign n74425 = ~n27326 ;
  assign n27849 = n26992 & n74425 ;
  assign n27850 = n27848 | n27849 ;
  assign n27851 = n74318 & n27850 ;
  assign n27852 = n74321 & n27851 ;
  assign n27853 = n27846 | n27852 ;
  assign n27854 = n65772 & n27853 ;
  assign n27855 = n26955 & n27312 ;
  assign n27856 = n26964 | n26986 ;
  assign n74426 = ~n27856 ;
  assign n27857 = n27323 & n74426 ;
  assign n74427 = ~n26987 ;
  assign n27858 = n26986 & n74427 ;
  assign n27859 = n27857 | n27858 ;
  assign n27860 = n74318 & n27859 ;
  assign n27861 = n74321 & n27860 ;
  assign n27862 = n27855 | n27861 ;
  assign n27863 = n65746 & n27862 ;
  assign n27864 = n26963 & n27312 ;
  assign n27321 = n26978 | n26982 ;
  assign n74428 = ~n27321 ;
  assign n27865 = n26976 & n74428 ;
  assign n74429 = ~n27322 ;
  assign n27866 = n26982 & n74429 ;
  assign n27867 = n27865 | n27866 ;
  assign n27868 = n74318 & n27867 ;
  assign n27869 = n74321 & n27868 ;
  assign n27870 = n27864 | n27869 ;
  assign n27871 = n65721 & n27870 ;
  assign n27314 = n26977 & n27312 ;
  assign n27319 = n26973 & n26974 ;
  assign n27872 = n74199 & n27319 ;
  assign n27873 = n27311 | n27872 ;
  assign n74430 = ~n27873 ;
  assign n27874 = n26976 & n74430 ;
  assign n27875 = n74321 & n27874 ;
  assign n27876 = n27314 | n27875 ;
  assign n27877 = n65686 & n27876 ;
  assign n74431 = ~x122 ;
  assign n27878 = x64 & n74431 ;
  assign n74432 = ~n276 ;
  assign n27879 = n74432 & n27878 ;
  assign n27880 = n73624 & n27879 ;
  assign n27884 = n74311 & n27883 ;
  assign n27885 = n27307 | n27884 ;
  assign n27886 = n74312 & n27885 ;
  assign n74433 = ~n27886 ;
  assign n27887 = n27880 & n74433 ;
  assign n74434 = ~n27887 ;
  assign n27888 = x6 & n74434 ;
  assign n74435 = ~n65384 ;
  assign n27889 = n74435 & n26974 ;
  assign n27890 = n73619 & n27889 ;
  assign n27891 = n74321 & n27890 ;
  assign n27892 = n27888 | n27891 ;
  assign n27894 = x65 & n27892 ;
  assign n27881 = n74321 & n27880 ;
  assign n74436 = ~n27881 ;
  assign n27882 = x6 & n74436 ;
  assign n27893 = x65 | n27891 ;
  assign n27895 = n27882 | n27893 ;
  assign n74437 = ~n27894 ;
  assign n27896 = n74437 & n27895 ;
  assign n74438 = ~x5 ;
  assign n27897 = n74438 & x64 ;
  assign n27898 = n27896 | n27897 ;
  assign n27899 = n65670 & n27892 ;
  assign n74439 = ~n27899 ;
  assign n27900 = n27898 & n74439 ;
  assign n74440 = ~n27875 ;
  assign n27901 = x66 & n74440 ;
  assign n74441 = ~n27314 ;
  assign n27902 = n74441 & n27901 ;
  assign n27903 = n27877 | n27902 ;
  assign n27904 = n27900 | n27903 ;
  assign n74442 = ~n27877 ;
  assign n27905 = n74442 & n27904 ;
  assign n74443 = ~n27869 ;
  assign n27906 = x67 & n74443 ;
  assign n74444 = ~n27864 ;
  assign n27907 = n74444 & n27906 ;
  assign n27908 = n27905 | n27907 ;
  assign n74445 = ~n27871 ;
  assign n27909 = n74445 & n27908 ;
  assign n74446 = ~n27861 ;
  assign n27910 = x68 & n74446 ;
  assign n74447 = ~n27855 ;
  assign n27911 = n74447 & n27910 ;
  assign n27912 = n27863 | n27911 ;
  assign n27913 = n27909 | n27912 ;
  assign n74448 = ~n27863 ;
  assign n27914 = n74448 & n27913 ;
  assign n74449 = ~n27852 ;
  assign n27915 = x69 & n74449 ;
  assign n74450 = ~n27846 ;
  assign n27916 = n74450 & n27915 ;
  assign n27917 = n27854 | n27916 ;
  assign n27918 = n27914 | n27917 ;
  assign n74451 = ~n27854 ;
  assign n27919 = n74451 & n27918 ;
  assign n74452 = ~n27843 ;
  assign n27920 = x70 & n74452 ;
  assign n74453 = ~n27838 ;
  assign n27921 = n74453 & n27920 ;
  assign n27922 = n27845 | n27921 ;
  assign n27923 = n27919 | n27922 ;
  assign n74454 = ~n27845 ;
  assign n27924 = n74454 & n27923 ;
  assign n74455 = ~n27835 ;
  assign n27925 = x71 & n74455 ;
  assign n74456 = ~n27830 ;
  assign n27926 = n74456 & n27925 ;
  assign n27927 = n27837 | n27926 ;
  assign n27929 = n27924 | n27927 ;
  assign n74457 = ~n27837 ;
  assign n27930 = n74457 & n27929 ;
  assign n74458 = ~n27827 ;
  assign n27931 = x72 & n74458 ;
  assign n74459 = ~n27822 ;
  assign n27932 = n74459 & n27931 ;
  assign n27933 = n27829 | n27932 ;
  assign n27934 = n27930 | n27933 ;
  assign n74460 = ~n27829 ;
  assign n27935 = n74460 & n27934 ;
  assign n74461 = ~n27819 ;
  assign n27936 = x73 & n74461 ;
  assign n74462 = ~n27814 ;
  assign n27937 = n74462 & n27936 ;
  assign n27938 = n27821 | n27937 ;
  assign n27940 = n27935 | n27938 ;
  assign n74463 = ~n27821 ;
  assign n27941 = n74463 & n27940 ;
  assign n74464 = ~n27811 ;
  assign n27942 = x74 & n74464 ;
  assign n74465 = ~n27806 ;
  assign n27943 = n74465 & n27942 ;
  assign n27944 = n27813 | n27943 ;
  assign n27945 = n27941 | n27944 ;
  assign n74466 = ~n27813 ;
  assign n27946 = n74466 & n27945 ;
  assign n74467 = ~n27803 ;
  assign n27947 = x75 & n74467 ;
  assign n74468 = ~n27798 ;
  assign n27948 = n74468 & n27947 ;
  assign n27949 = n27805 | n27948 ;
  assign n27951 = n27946 | n27949 ;
  assign n74469 = ~n27805 ;
  assign n27952 = n74469 & n27951 ;
  assign n74470 = ~n27795 ;
  assign n27953 = x76 & n74470 ;
  assign n74471 = ~n27790 ;
  assign n27954 = n74471 & n27953 ;
  assign n27955 = n27797 | n27954 ;
  assign n27956 = n27952 | n27955 ;
  assign n74472 = ~n27797 ;
  assign n27957 = n74472 & n27956 ;
  assign n74473 = ~n27787 ;
  assign n27958 = x77 & n74473 ;
  assign n74474 = ~n27782 ;
  assign n27959 = n74474 & n27958 ;
  assign n27960 = n27789 | n27959 ;
  assign n27962 = n27957 | n27960 ;
  assign n74475 = ~n27789 ;
  assign n27963 = n74475 & n27962 ;
  assign n74476 = ~n27779 ;
  assign n27964 = x78 & n74476 ;
  assign n74477 = ~n27774 ;
  assign n27965 = n74477 & n27964 ;
  assign n27966 = n27781 | n27965 ;
  assign n27967 = n27963 | n27966 ;
  assign n74478 = ~n27781 ;
  assign n27968 = n74478 & n27967 ;
  assign n74479 = ~n27771 ;
  assign n27969 = x79 & n74479 ;
  assign n74480 = ~n27766 ;
  assign n27970 = n74480 & n27969 ;
  assign n27971 = n27773 | n27970 ;
  assign n27973 = n27968 | n27971 ;
  assign n74481 = ~n27773 ;
  assign n27974 = n74481 & n27973 ;
  assign n74482 = ~n27763 ;
  assign n27975 = x80 & n74482 ;
  assign n74483 = ~n27758 ;
  assign n27976 = n74483 & n27975 ;
  assign n27977 = n27765 | n27976 ;
  assign n27978 = n27974 | n27977 ;
  assign n74484 = ~n27765 ;
  assign n27979 = n74484 & n27978 ;
  assign n74485 = ~n27755 ;
  assign n27980 = x81 & n74485 ;
  assign n74486 = ~n27750 ;
  assign n27981 = n74486 & n27980 ;
  assign n27982 = n27757 | n27981 ;
  assign n27984 = n27979 | n27982 ;
  assign n74487 = ~n27757 ;
  assign n27985 = n74487 & n27984 ;
  assign n74488 = ~n27747 ;
  assign n27986 = x82 & n74488 ;
  assign n74489 = ~n27742 ;
  assign n27987 = n74489 & n27986 ;
  assign n27988 = n27749 | n27987 ;
  assign n27989 = n27985 | n27988 ;
  assign n74490 = ~n27749 ;
  assign n27990 = n74490 & n27989 ;
  assign n74491 = ~n27739 ;
  assign n27991 = x83 & n74491 ;
  assign n74492 = ~n27734 ;
  assign n27992 = n74492 & n27991 ;
  assign n27993 = n27741 | n27992 ;
  assign n27995 = n27990 | n27993 ;
  assign n74493 = ~n27741 ;
  assign n27996 = n74493 & n27995 ;
  assign n74494 = ~n27731 ;
  assign n27997 = x84 & n74494 ;
  assign n74495 = ~n27726 ;
  assign n27998 = n74495 & n27997 ;
  assign n27999 = n27733 | n27998 ;
  assign n28000 = n27996 | n27999 ;
  assign n74496 = ~n27733 ;
  assign n28001 = n74496 & n28000 ;
  assign n74497 = ~n27723 ;
  assign n28002 = x85 & n74497 ;
  assign n74498 = ~n27718 ;
  assign n28003 = n74498 & n28002 ;
  assign n28004 = n27725 | n28003 ;
  assign n28006 = n28001 | n28004 ;
  assign n74499 = ~n27725 ;
  assign n28007 = n74499 & n28006 ;
  assign n74500 = ~n27715 ;
  assign n28008 = x86 & n74500 ;
  assign n74501 = ~n27710 ;
  assign n28009 = n74501 & n28008 ;
  assign n28010 = n27717 | n28009 ;
  assign n28011 = n28007 | n28010 ;
  assign n74502 = ~n27717 ;
  assign n28012 = n74502 & n28011 ;
  assign n74503 = ~n27707 ;
  assign n28013 = x87 & n74503 ;
  assign n74504 = ~n27702 ;
  assign n28014 = n74504 & n28013 ;
  assign n28015 = n27709 | n28014 ;
  assign n28017 = n28012 | n28015 ;
  assign n74505 = ~n27709 ;
  assign n28018 = n74505 & n28017 ;
  assign n74506 = ~n27699 ;
  assign n28019 = x88 & n74506 ;
  assign n74507 = ~n27694 ;
  assign n28020 = n74507 & n28019 ;
  assign n28021 = n27701 | n28020 ;
  assign n28022 = n28018 | n28021 ;
  assign n74508 = ~n27701 ;
  assign n28023 = n74508 & n28022 ;
  assign n74509 = ~n27691 ;
  assign n28024 = x89 & n74509 ;
  assign n74510 = ~n27686 ;
  assign n28025 = n74510 & n28024 ;
  assign n28026 = n27693 | n28025 ;
  assign n28028 = n28023 | n28026 ;
  assign n74511 = ~n27693 ;
  assign n28029 = n74511 & n28028 ;
  assign n74512 = ~n27683 ;
  assign n28030 = x90 & n74512 ;
  assign n74513 = ~n27678 ;
  assign n28031 = n74513 & n28030 ;
  assign n28032 = n27685 | n28031 ;
  assign n28033 = n28029 | n28032 ;
  assign n74514 = ~n27685 ;
  assign n28034 = n74514 & n28033 ;
  assign n74515 = ~n27675 ;
  assign n28035 = x91 & n74515 ;
  assign n74516 = ~n27670 ;
  assign n28036 = n74516 & n28035 ;
  assign n28037 = n27677 | n28036 ;
  assign n28039 = n28034 | n28037 ;
  assign n74517 = ~n27677 ;
  assign n28040 = n74517 & n28039 ;
  assign n74518 = ~n27667 ;
  assign n28041 = x92 & n74518 ;
  assign n74519 = ~n27662 ;
  assign n28042 = n74519 & n28041 ;
  assign n28043 = n27669 | n28042 ;
  assign n28044 = n28040 | n28043 ;
  assign n74520 = ~n27669 ;
  assign n28045 = n74520 & n28044 ;
  assign n74521 = ~n27659 ;
  assign n28046 = x93 & n74521 ;
  assign n74522 = ~n27654 ;
  assign n28047 = n74522 & n28046 ;
  assign n28048 = n27661 | n28047 ;
  assign n28050 = n28045 | n28048 ;
  assign n74523 = ~n27661 ;
  assign n28051 = n74523 & n28050 ;
  assign n74524 = ~n27651 ;
  assign n28052 = x94 & n74524 ;
  assign n74525 = ~n27646 ;
  assign n28053 = n74525 & n28052 ;
  assign n28054 = n27653 | n28053 ;
  assign n28055 = n28051 | n28054 ;
  assign n74526 = ~n27653 ;
  assign n28056 = n74526 & n28055 ;
  assign n74527 = ~n27643 ;
  assign n28057 = x95 & n74527 ;
  assign n74528 = ~n27638 ;
  assign n28058 = n74528 & n28057 ;
  assign n28059 = n27645 | n28058 ;
  assign n28061 = n28056 | n28059 ;
  assign n74529 = ~n27645 ;
  assign n28062 = n74529 & n28061 ;
  assign n74530 = ~n27635 ;
  assign n28063 = x96 & n74530 ;
  assign n74531 = ~n27630 ;
  assign n28064 = n74531 & n28063 ;
  assign n28065 = n27637 | n28064 ;
  assign n28066 = n28062 | n28065 ;
  assign n74532 = ~n27637 ;
  assign n28067 = n74532 & n28066 ;
  assign n74533 = ~n27627 ;
  assign n28068 = x97 & n74533 ;
  assign n74534 = ~n27622 ;
  assign n28069 = n74534 & n28068 ;
  assign n28070 = n27629 | n28069 ;
  assign n28072 = n28067 | n28070 ;
  assign n74535 = ~n27629 ;
  assign n28073 = n74535 & n28072 ;
  assign n74536 = ~n27619 ;
  assign n28074 = x98 & n74536 ;
  assign n74537 = ~n27614 ;
  assign n28075 = n74537 & n28074 ;
  assign n28076 = n27621 | n28075 ;
  assign n28077 = n28073 | n28076 ;
  assign n74538 = ~n27621 ;
  assign n28078 = n74538 & n28077 ;
  assign n74539 = ~n27611 ;
  assign n28079 = x99 & n74539 ;
  assign n74540 = ~n27606 ;
  assign n28080 = n74540 & n28079 ;
  assign n28081 = n27613 | n28080 ;
  assign n28083 = n28078 | n28081 ;
  assign n74541 = ~n27613 ;
  assign n28084 = n74541 & n28083 ;
  assign n74542 = ~n27603 ;
  assign n28085 = x100 & n74542 ;
  assign n74543 = ~n27598 ;
  assign n28086 = n74543 & n28085 ;
  assign n28087 = n27605 | n28086 ;
  assign n28088 = n28084 | n28087 ;
  assign n74544 = ~n27605 ;
  assign n28089 = n74544 & n28088 ;
  assign n74545 = ~n27595 ;
  assign n28090 = x101 & n74545 ;
  assign n74546 = ~n27590 ;
  assign n28091 = n74546 & n28090 ;
  assign n28092 = n27597 | n28091 ;
  assign n28094 = n28089 | n28092 ;
  assign n74547 = ~n27597 ;
  assign n28095 = n74547 & n28094 ;
  assign n74548 = ~n27587 ;
  assign n28096 = x102 & n74548 ;
  assign n74549 = ~n27582 ;
  assign n28097 = n74549 & n28096 ;
  assign n28098 = n27589 | n28097 ;
  assign n28099 = n28095 | n28098 ;
  assign n74550 = ~n27589 ;
  assign n28100 = n74550 & n28099 ;
  assign n74551 = ~n27579 ;
  assign n28101 = x103 & n74551 ;
  assign n74552 = ~n27574 ;
  assign n28102 = n74552 & n28101 ;
  assign n28103 = n27581 | n28102 ;
  assign n28105 = n28100 | n28103 ;
  assign n74553 = ~n27581 ;
  assign n28106 = n74553 & n28105 ;
  assign n74554 = ~n27571 ;
  assign n28107 = x104 & n74554 ;
  assign n74555 = ~n27566 ;
  assign n28108 = n74555 & n28107 ;
  assign n28109 = n27573 | n28108 ;
  assign n28110 = n28106 | n28109 ;
  assign n74556 = ~n27573 ;
  assign n28111 = n74556 & n28110 ;
  assign n74557 = ~n27563 ;
  assign n28112 = x105 & n74557 ;
  assign n74558 = ~n27558 ;
  assign n28113 = n74558 & n28112 ;
  assign n28114 = n27565 | n28113 ;
  assign n28116 = n28111 | n28114 ;
  assign n74559 = ~n27565 ;
  assign n28117 = n74559 & n28116 ;
  assign n74560 = ~n27555 ;
  assign n28118 = x106 & n74560 ;
  assign n74561 = ~n27550 ;
  assign n28119 = n74561 & n28118 ;
  assign n28120 = n27557 | n28119 ;
  assign n28121 = n28117 | n28120 ;
  assign n74562 = ~n27557 ;
  assign n28122 = n74562 & n28121 ;
  assign n74563 = ~n27547 ;
  assign n28123 = x107 & n74563 ;
  assign n74564 = ~n27542 ;
  assign n28124 = n74564 & n28123 ;
  assign n28125 = n27549 | n28124 ;
  assign n28127 = n28122 | n28125 ;
  assign n74565 = ~n27549 ;
  assign n28128 = n74565 & n28127 ;
  assign n74566 = ~n27539 ;
  assign n28129 = x108 & n74566 ;
  assign n74567 = ~n27534 ;
  assign n28130 = n74567 & n28129 ;
  assign n28131 = n27541 | n28130 ;
  assign n28132 = n28128 | n28131 ;
  assign n74568 = ~n27541 ;
  assign n28133 = n74568 & n28132 ;
  assign n74569 = ~n27531 ;
  assign n28134 = x109 & n74569 ;
  assign n74570 = ~n27526 ;
  assign n28135 = n74570 & n28134 ;
  assign n28136 = n27533 | n28135 ;
  assign n28138 = n28133 | n28136 ;
  assign n74571 = ~n27533 ;
  assign n28139 = n74571 & n28138 ;
  assign n74572 = ~n27523 ;
  assign n28140 = x110 & n74572 ;
  assign n74573 = ~n27518 ;
  assign n28141 = n74573 & n28140 ;
  assign n28142 = n27525 | n28141 ;
  assign n28143 = n28139 | n28142 ;
  assign n74574 = ~n27525 ;
  assign n28144 = n74574 & n28143 ;
  assign n74575 = ~n27515 ;
  assign n28145 = x111 & n74575 ;
  assign n74576 = ~n27510 ;
  assign n28146 = n74576 & n28145 ;
  assign n28147 = n27517 | n28146 ;
  assign n28149 = n28144 | n28147 ;
  assign n74577 = ~n27517 ;
  assign n28150 = n74577 & n28149 ;
  assign n74578 = ~n27507 ;
  assign n28151 = x112 & n74578 ;
  assign n74579 = ~n27502 ;
  assign n28152 = n74579 & n28151 ;
  assign n28153 = n27509 | n28152 ;
  assign n28154 = n28150 | n28153 ;
  assign n74580 = ~n27509 ;
  assign n28155 = n74580 & n28154 ;
  assign n74581 = ~n27499 ;
  assign n28156 = x113 & n74581 ;
  assign n74582 = ~n27494 ;
  assign n28157 = n74582 & n28156 ;
  assign n28158 = n27501 | n28157 ;
  assign n28160 = n28155 | n28158 ;
  assign n74583 = ~n27501 ;
  assign n28161 = n74583 & n28160 ;
  assign n74584 = ~n27491 ;
  assign n28162 = x114 & n74584 ;
  assign n74585 = ~n27486 ;
  assign n28163 = n74585 & n28162 ;
  assign n28164 = n27493 | n28163 ;
  assign n28165 = n28161 | n28164 ;
  assign n74586 = ~n27493 ;
  assign n28166 = n74586 & n28165 ;
  assign n74587 = ~n27483 ;
  assign n28167 = x115 & n74587 ;
  assign n74588 = ~n27478 ;
  assign n28168 = n74588 & n28167 ;
  assign n28169 = n27485 | n28168 ;
  assign n28171 = n28166 | n28169 ;
  assign n74589 = ~n27485 ;
  assign n28172 = n74589 & n28171 ;
  assign n74590 = ~n27475 ;
  assign n28173 = x116 & n74590 ;
  assign n74591 = ~n27470 ;
  assign n28174 = n74591 & n28173 ;
  assign n28175 = n27477 | n28174 ;
  assign n28176 = n28172 | n28175 ;
  assign n74592 = ~n27477 ;
  assign n28177 = n74592 & n28176 ;
  assign n74593 = ~n27467 ;
  assign n28178 = x117 & n74593 ;
  assign n74594 = ~n27462 ;
  assign n28179 = n74594 & n28178 ;
  assign n28180 = n27469 | n28179 ;
  assign n28182 = n28177 | n28180 ;
  assign n74595 = ~n27469 ;
  assign n28183 = n74595 & n28182 ;
  assign n74596 = ~n27459 ;
  assign n28184 = x118 & n74596 ;
  assign n74597 = ~n27454 ;
  assign n28185 = n74597 & n28184 ;
  assign n28186 = n27461 | n28185 ;
  assign n28187 = n28183 | n28186 ;
  assign n74598 = ~n27461 ;
  assign n28188 = n74598 & n28187 ;
  assign n74599 = ~n27451 ;
  assign n28189 = x119 & n74599 ;
  assign n74600 = ~n27446 ;
  assign n28190 = n74600 & n28189 ;
  assign n28191 = n27453 | n28190 ;
  assign n28193 = n28188 | n28191 ;
  assign n74601 = ~n27453 ;
  assign n28194 = n74601 & n28193 ;
  assign n74602 = ~n27443 ;
  assign n28195 = x120 & n74602 ;
  assign n74603 = ~n27438 ;
  assign n28196 = n74603 & n28195 ;
  assign n28197 = n27445 | n28196 ;
  assign n28198 = n28194 | n28197 ;
  assign n74604 = ~n27445 ;
  assign n28199 = n74604 & n28198 ;
  assign n74605 = ~n27435 ;
  assign n28200 = x121 & n74605 ;
  assign n74606 = ~n27315 ;
  assign n28201 = n74606 & n28200 ;
  assign n28202 = n27437 | n28201 ;
  assign n28204 = n28199 | n28202 ;
  assign n74607 = ~n27437 ;
  assign n28205 = n74607 & n28204 ;
  assign n28212 = n74431 & n28211 ;
  assign n135 = ~n27312 ;
  assign n28213 = n135 & n28209 ;
  assign n28214 = n26522 & n27312 ;
  assign n74609 = ~n28214 ;
  assign n28215 = x122 & n74609 ;
  assign n74610 = ~n28213 ;
  assign n28216 = n74610 & n28215 ;
  assign n28217 = n274 | n276 ;
  assign n28218 = n28216 | n28217 ;
  assign n28219 = n28212 | n28218 ;
  assign n28221 = n28205 | n28219 ;
  assign n74611 = ~n28220 ;
  assign n28222 = n74611 & n28221 ;
  assign n74612 = ~n28199 ;
  assign n28203 = n74612 & n28202 ;
  assign n28225 = n27882 | n27891 ;
  assign n28226 = x65 & n28225 ;
  assign n74613 = ~n28226 ;
  assign n28227 = n27895 & n74613 ;
  assign n28228 = n27897 | n28227 ;
  assign n28229 = n74439 & n28228 ;
  assign n28231 = n27902 | n28229 ;
  assign n28232 = n74442 & n28231 ;
  assign n28233 = n27871 | n27907 ;
  assign n28235 = n28232 | n28233 ;
  assign n28236 = n74445 & n28235 ;
  assign n28238 = n27912 | n28236 ;
  assign n28239 = n74448 & n28238 ;
  assign n28241 = n27917 | n28239 ;
  assign n28242 = n74451 & n28241 ;
  assign n28243 = n27922 | n28242 ;
  assign n28245 = n74454 & n28243 ;
  assign n28246 = n27927 | n28245 ;
  assign n28247 = n74457 & n28246 ;
  assign n28248 = n27933 | n28247 ;
  assign n28250 = n74460 & n28248 ;
  assign n28251 = n27938 | n28250 ;
  assign n28252 = n74463 & n28251 ;
  assign n28253 = n27944 | n28252 ;
  assign n28255 = n74466 & n28253 ;
  assign n28256 = n27949 | n28255 ;
  assign n28257 = n74469 & n28256 ;
  assign n28258 = n27955 | n28257 ;
  assign n28260 = n74472 & n28258 ;
  assign n28261 = n27960 | n28260 ;
  assign n28262 = n74475 & n28261 ;
  assign n28263 = n27966 | n28262 ;
  assign n28265 = n74478 & n28263 ;
  assign n28266 = n27971 | n28265 ;
  assign n28267 = n74481 & n28266 ;
  assign n28268 = n27977 | n28267 ;
  assign n28270 = n74484 & n28268 ;
  assign n28271 = n27982 | n28270 ;
  assign n28272 = n74487 & n28271 ;
  assign n28273 = n27988 | n28272 ;
  assign n28275 = n74490 & n28273 ;
  assign n28276 = n27993 | n28275 ;
  assign n28277 = n74493 & n28276 ;
  assign n28278 = n27999 | n28277 ;
  assign n28280 = n74496 & n28278 ;
  assign n28281 = n28004 | n28280 ;
  assign n28282 = n74499 & n28281 ;
  assign n28283 = n28010 | n28282 ;
  assign n28285 = n74502 & n28283 ;
  assign n28286 = n28015 | n28285 ;
  assign n28287 = n74505 & n28286 ;
  assign n28288 = n28021 | n28287 ;
  assign n28290 = n74508 & n28288 ;
  assign n28291 = n28026 | n28290 ;
  assign n28292 = n74511 & n28291 ;
  assign n28293 = n28032 | n28292 ;
  assign n28295 = n74514 & n28293 ;
  assign n28296 = n28037 | n28295 ;
  assign n28297 = n74517 & n28296 ;
  assign n28298 = n28043 | n28297 ;
  assign n28300 = n74520 & n28298 ;
  assign n28301 = n28048 | n28300 ;
  assign n28302 = n74523 & n28301 ;
  assign n28303 = n28054 | n28302 ;
  assign n28305 = n74526 & n28303 ;
  assign n28306 = n28059 | n28305 ;
  assign n28307 = n74529 & n28306 ;
  assign n28308 = n28065 | n28307 ;
  assign n28310 = n74532 & n28308 ;
  assign n28311 = n28070 | n28310 ;
  assign n28312 = n74535 & n28311 ;
  assign n28313 = n28076 | n28312 ;
  assign n28315 = n74538 & n28313 ;
  assign n28316 = n28081 | n28315 ;
  assign n28317 = n74541 & n28316 ;
  assign n28318 = n28087 | n28317 ;
  assign n28320 = n74544 & n28318 ;
  assign n28321 = n28092 | n28320 ;
  assign n28322 = n74547 & n28321 ;
  assign n28323 = n28098 | n28322 ;
  assign n28325 = n74550 & n28323 ;
  assign n28326 = n28103 | n28325 ;
  assign n28327 = n74553 & n28326 ;
  assign n28328 = n28109 | n28327 ;
  assign n28330 = n74556 & n28328 ;
  assign n28331 = n28114 | n28330 ;
  assign n28332 = n74559 & n28331 ;
  assign n28333 = n28120 | n28332 ;
  assign n28335 = n74562 & n28333 ;
  assign n28336 = n28125 | n28335 ;
  assign n28337 = n74565 & n28336 ;
  assign n28338 = n28131 | n28337 ;
  assign n28340 = n74568 & n28338 ;
  assign n28341 = n28136 | n28340 ;
  assign n28342 = n74571 & n28341 ;
  assign n28343 = n28142 | n28342 ;
  assign n28345 = n74574 & n28343 ;
  assign n28346 = n28147 | n28345 ;
  assign n28347 = n74577 & n28346 ;
  assign n28348 = n28153 | n28347 ;
  assign n28350 = n74580 & n28348 ;
  assign n28351 = n28158 | n28350 ;
  assign n28352 = n74583 & n28351 ;
  assign n28353 = n28164 | n28352 ;
  assign n28355 = n74586 & n28353 ;
  assign n28356 = n28169 | n28355 ;
  assign n28357 = n74589 & n28356 ;
  assign n28358 = n28175 | n28357 ;
  assign n28360 = n74592 & n28358 ;
  assign n28361 = n28180 | n28360 ;
  assign n28362 = n74595 & n28361 ;
  assign n28363 = n28186 | n28362 ;
  assign n28365 = n74598 & n28363 ;
  assign n28366 = n28191 | n28365 ;
  assign n28367 = n74601 & n28366 ;
  assign n28368 = n28197 | n28367 ;
  assign n28370 = n27445 | n28202 ;
  assign n74614 = ~n28370 ;
  assign n28371 = n28368 & n74614 ;
  assign n28372 = n28203 | n28371 ;
  assign n134 = ~n28222 ;
  assign n28373 = n134 & n28372 ;
  assign n28374 = n74604 & n28368 ;
  assign n28375 = n28202 | n28374 ;
  assign n28376 = n74607 & n28375 ;
  assign n28377 = n28219 | n28376 ;
  assign n28378 = n27436 & n74611 ;
  assign n28379 = n28377 & n28378 ;
  assign n28380 = n28373 | n28379 ;
  assign n28381 = n74431 & n28380 ;
  assign n74616 = ~n28379 ;
  assign n29129 = x122 & n74616 ;
  assign n74617 = ~n28373 ;
  assign n29130 = n74617 & n29129 ;
  assign n29131 = n28381 | n29130 ;
  assign n74618 = ~n28367 ;
  assign n28369 = n28197 & n74618 ;
  assign n28382 = n27453 | n28197 ;
  assign n74619 = ~n28382 ;
  assign n28383 = n28193 & n74619 ;
  assign n28384 = n28369 | n28383 ;
  assign n28385 = n134 & n28384 ;
  assign n28386 = n27444 & n74611 ;
  assign n28387 = n28377 & n28386 ;
  assign n28388 = n28385 | n28387 ;
  assign n28389 = n74029 & n28388 ;
  assign n74620 = ~n28188 ;
  assign n28192 = n74620 & n28191 ;
  assign n28390 = n27461 | n28191 ;
  assign n74621 = ~n28390 ;
  assign n28391 = n28363 & n74621 ;
  assign n28392 = n28192 | n28391 ;
  assign n28393 = n134 & n28392 ;
  assign n28394 = n27452 & n74611 ;
  assign n28395 = n28377 & n28394 ;
  assign n28396 = n28393 | n28395 ;
  assign n28397 = n74021 & n28396 ;
  assign n74622 = ~n28395 ;
  assign n29119 = x120 & n74622 ;
  assign n74623 = ~n28393 ;
  assign n29120 = n74623 & n29119 ;
  assign n29121 = n28397 | n29120 ;
  assign n74624 = ~n28362 ;
  assign n28364 = n28186 & n74624 ;
  assign n28398 = n27469 | n28186 ;
  assign n74625 = ~n28398 ;
  assign n28399 = n28182 & n74625 ;
  assign n28400 = n28364 | n28399 ;
  assign n28401 = n134 & n28400 ;
  assign n28402 = n27460 & n74611 ;
  assign n28403 = n28377 & n28402 ;
  assign n28404 = n28401 | n28403 ;
  assign n28405 = n73617 & n28404 ;
  assign n74626 = ~n28177 ;
  assign n28181 = n74626 & n28180 ;
  assign n28406 = n27477 | n28180 ;
  assign n74627 = ~n28406 ;
  assign n28407 = n28358 & n74627 ;
  assign n28408 = n28181 | n28407 ;
  assign n28409 = n134 & n28408 ;
  assign n28410 = n27468 & n74611 ;
  assign n28411 = n28377 & n28410 ;
  assign n28412 = n28409 | n28411 ;
  assign n28413 = n73188 & n28412 ;
  assign n74628 = ~n28411 ;
  assign n29109 = x118 & n74628 ;
  assign n74629 = ~n28409 ;
  assign n29110 = n74629 & n29109 ;
  assign n29111 = n28413 | n29110 ;
  assign n74630 = ~n28357 ;
  assign n28359 = n28175 & n74630 ;
  assign n28414 = n27485 | n28175 ;
  assign n74631 = ~n28414 ;
  assign n28415 = n28171 & n74631 ;
  assign n28416 = n28359 | n28415 ;
  assign n28417 = n134 & n28416 ;
  assign n28418 = n27476 & n74611 ;
  assign n28419 = n28377 & n28418 ;
  assign n28420 = n28417 | n28419 ;
  assign n28421 = n73177 & n28420 ;
  assign n74632 = ~n28166 ;
  assign n28170 = n74632 & n28169 ;
  assign n28422 = n27493 | n28169 ;
  assign n74633 = ~n28422 ;
  assign n28423 = n28353 & n74633 ;
  assign n28424 = n28170 | n28423 ;
  assign n28425 = n134 & n28424 ;
  assign n28426 = n27484 & n74611 ;
  assign n28427 = n28377 & n28426 ;
  assign n28428 = n28425 | n28427 ;
  assign n28429 = n72752 & n28428 ;
  assign n74634 = ~n28427 ;
  assign n29098 = x116 & n74634 ;
  assign n74635 = ~n28425 ;
  assign n29099 = n74635 & n29098 ;
  assign n29100 = n28429 | n29099 ;
  assign n74636 = ~n28352 ;
  assign n28354 = n28164 & n74636 ;
  assign n28430 = n27501 | n28164 ;
  assign n74637 = ~n28430 ;
  assign n28431 = n28160 & n74637 ;
  assign n28432 = n28354 | n28431 ;
  assign n28433 = n134 & n28432 ;
  assign n28434 = n27492 & n74611 ;
  assign n28435 = n28377 & n28434 ;
  assign n28436 = n28433 | n28435 ;
  assign n28437 = n72393 & n28436 ;
  assign n74638 = ~n28155 ;
  assign n28159 = n74638 & n28158 ;
  assign n28438 = n27509 | n28158 ;
  assign n74639 = ~n28438 ;
  assign n28439 = n28348 & n74639 ;
  assign n28440 = n28159 | n28439 ;
  assign n28441 = n134 & n28440 ;
  assign n28442 = n27500 & n74611 ;
  assign n28443 = n28377 & n28442 ;
  assign n28444 = n28441 | n28443 ;
  assign n28445 = n72385 & n28444 ;
  assign n74640 = ~n28443 ;
  assign n29088 = x114 & n74640 ;
  assign n74641 = ~n28441 ;
  assign n29089 = n74641 & n29088 ;
  assign n29090 = n28445 | n29089 ;
  assign n74642 = ~n28347 ;
  assign n28349 = n28153 & n74642 ;
  assign n28446 = n27517 | n28153 ;
  assign n74643 = ~n28446 ;
  assign n28447 = n28149 & n74643 ;
  assign n28448 = n28349 | n28447 ;
  assign n28449 = n134 & n28448 ;
  assign n28450 = n27508 & n74611 ;
  assign n28451 = n28377 & n28450 ;
  assign n28452 = n28449 | n28451 ;
  assign n28453 = n72025 & n28452 ;
  assign n74644 = ~n28144 ;
  assign n28148 = n74644 & n28147 ;
  assign n28454 = n27525 | n28147 ;
  assign n74645 = ~n28454 ;
  assign n28455 = n28343 & n74645 ;
  assign n28456 = n28148 | n28455 ;
  assign n28457 = n134 & n28456 ;
  assign n28458 = n27516 & n74611 ;
  assign n28459 = n28377 & n28458 ;
  assign n28460 = n28457 | n28459 ;
  assign n28461 = n71645 & n28460 ;
  assign n74646 = ~n28459 ;
  assign n29078 = x112 & n74646 ;
  assign n74647 = ~n28457 ;
  assign n29079 = n74647 & n29078 ;
  assign n29080 = n28461 | n29079 ;
  assign n74648 = ~n28342 ;
  assign n28344 = n28142 & n74648 ;
  assign n28462 = n27533 | n28142 ;
  assign n74649 = ~n28462 ;
  assign n28463 = n28138 & n74649 ;
  assign n28464 = n28344 | n28463 ;
  assign n28465 = n134 & n28464 ;
  assign n28466 = n27524 & n74611 ;
  assign n28467 = n28377 & n28466 ;
  assign n28468 = n28465 | n28467 ;
  assign n28469 = n71633 & n28468 ;
  assign n74650 = ~n28133 ;
  assign n28137 = n74650 & n28136 ;
  assign n28470 = n27541 | n28136 ;
  assign n74651 = ~n28470 ;
  assign n28471 = n28338 & n74651 ;
  assign n28472 = n28137 | n28471 ;
  assign n28473 = n134 & n28472 ;
  assign n28474 = n27532 & n74611 ;
  assign n28475 = n28377 & n28474 ;
  assign n28476 = n28473 | n28475 ;
  assign n28477 = n71253 & n28476 ;
  assign n74652 = ~n28475 ;
  assign n29068 = x110 & n74652 ;
  assign n74653 = ~n28473 ;
  assign n29069 = n74653 & n29068 ;
  assign n29070 = n28477 | n29069 ;
  assign n74654 = ~n28337 ;
  assign n28339 = n28131 & n74654 ;
  assign n28478 = n27549 | n28131 ;
  assign n74655 = ~n28478 ;
  assign n28479 = n28127 & n74655 ;
  assign n28480 = n28339 | n28479 ;
  assign n28481 = n134 & n28480 ;
  assign n28482 = n27540 & n74611 ;
  assign n28483 = n28377 & n28482 ;
  assign n28484 = n28481 | n28483 ;
  assign n28485 = n70935 & n28484 ;
  assign n74656 = ~n28122 ;
  assign n28126 = n74656 & n28125 ;
  assign n28486 = n27557 | n28125 ;
  assign n74657 = ~n28486 ;
  assign n28487 = n28333 & n74657 ;
  assign n28488 = n28126 | n28487 ;
  assign n28489 = n134 & n28488 ;
  assign n28490 = n27548 & n74611 ;
  assign n28491 = n28377 & n28490 ;
  assign n28492 = n28489 | n28491 ;
  assign n28493 = n70927 & n28492 ;
  assign n74658 = ~n28491 ;
  assign n29057 = x108 & n74658 ;
  assign n74659 = ~n28489 ;
  assign n29058 = n74659 & n29057 ;
  assign n29059 = n28493 | n29058 ;
  assign n74660 = ~n28332 ;
  assign n28334 = n28120 & n74660 ;
  assign n28494 = n27565 | n28120 ;
  assign n74661 = ~n28494 ;
  assign n28495 = n28116 & n74661 ;
  assign n28496 = n28334 | n28495 ;
  assign n28497 = n134 & n28496 ;
  assign n28498 = n27556 & n74611 ;
  assign n28499 = n28377 & n28498 ;
  assign n28500 = n28497 | n28499 ;
  assign n28501 = n70609 & n28500 ;
  assign n74662 = ~n28111 ;
  assign n28115 = n74662 & n28114 ;
  assign n28502 = n27573 | n28114 ;
  assign n74663 = ~n28502 ;
  assign n28503 = n28328 & n74663 ;
  assign n28504 = n28115 | n28503 ;
  assign n28505 = n134 & n28504 ;
  assign n28506 = n27564 & n74611 ;
  assign n28507 = n28377 & n28506 ;
  assign n28508 = n28505 | n28507 ;
  assign n28509 = n70276 & n28508 ;
  assign n74664 = ~n28507 ;
  assign n29046 = x106 & n74664 ;
  assign n74665 = ~n28505 ;
  assign n29047 = n74665 & n29046 ;
  assign n29048 = n28509 | n29047 ;
  assign n74666 = ~n28327 ;
  assign n28329 = n28109 & n74666 ;
  assign n28510 = n27581 | n28109 ;
  assign n74667 = ~n28510 ;
  assign n28511 = n28105 & n74667 ;
  assign n28512 = n28329 | n28511 ;
  assign n28513 = n134 & n28512 ;
  assign n28514 = n27572 & n74611 ;
  assign n28515 = n28377 & n28514 ;
  assign n28516 = n28513 | n28515 ;
  assign n28517 = n70176 & n28516 ;
  assign n74668 = ~n28100 ;
  assign n28104 = n74668 & n28103 ;
  assign n28518 = n27589 | n28103 ;
  assign n74669 = ~n28518 ;
  assign n28519 = n28323 & n74669 ;
  assign n28520 = n28104 | n28519 ;
  assign n28521 = n134 & n28520 ;
  assign n28522 = n27580 & n74611 ;
  assign n28523 = n28377 & n28522 ;
  assign n28524 = n28521 | n28523 ;
  assign n28525 = n69857 & n28524 ;
  assign n74670 = ~n28523 ;
  assign n29035 = x104 & n74670 ;
  assign n74671 = ~n28521 ;
  assign n29036 = n74671 & n29035 ;
  assign n29037 = n28525 | n29036 ;
  assign n74672 = ~n28322 ;
  assign n28324 = n28098 & n74672 ;
  assign n28526 = n27597 | n28098 ;
  assign n74673 = ~n28526 ;
  assign n28527 = n28094 & n74673 ;
  assign n28528 = n28324 | n28527 ;
  assign n28529 = n134 & n28528 ;
  assign n28530 = n27588 & n74611 ;
  assign n28531 = n28377 & n28530 ;
  assign n28532 = n28529 | n28531 ;
  assign n28533 = n69656 & n28532 ;
  assign n74674 = ~n28089 ;
  assign n28093 = n74674 & n28092 ;
  assign n28534 = n27605 | n28092 ;
  assign n74675 = ~n28534 ;
  assign n28535 = n28318 & n74675 ;
  assign n28536 = n28093 | n28535 ;
  assign n28537 = n134 & n28536 ;
  assign n28538 = n27596 & n74611 ;
  assign n28539 = n28377 & n28538 ;
  assign n28540 = n28537 | n28539 ;
  assign n28541 = n69528 & n28540 ;
  assign n74676 = ~n28539 ;
  assign n29024 = x102 & n74676 ;
  assign n74677 = ~n28537 ;
  assign n29025 = n74677 & n29024 ;
  assign n29026 = n28541 | n29025 ;
  assign n74678 = ~n28317 ;
  assign n28319 = n28087 & n74678 ;
  assign n28542 = n27613 | n28087 ;
  assign n74679 = ~n28542 ;
  assign n28543 = n28083 & n74679 ;
  assign n28544 = n28319 | n28543 ;
  assign n28545 = n134 & n28544 ;
  assign n28546 = n27604 & n74611 ;
  assign n28547 = n28377 & n28546 ;
  assign n28548 = n28545 | n28547 ;
  assign n28549 = n69261 & n28548 ;
  assign n74680 = ~n28078 ;
  assign n28082 = n74680 & n28081 ;
  assign n28550 = n27621 | n28081 ;
  assign n74681 = ~n28550 ;
  assign n28551 = n28313 & n74681 ;
  assign n28552 = n28082 | n28551 ;
  assign n28553 = n134 & n28552 ;
  assign n28554 = n27612 & n74611 ;
  assign n28555 = n28377 & n28554 ;
  assign n28556 = n28553 | n28555 ;
  assign n28557 = n69075 & n28556 ;
  assign n74682 = ~n28555 ;
  assign n29014 = x100 & n74682 ;
  assign n74683 = ~n28553 ;
  assign n29015 = n74683 & n29014 ;
  assign n29016 = n28557 | n29015 ;
  assign n74684 = ~n28312 ;
  assign n28314 = n28076 & n74684 ;
  assign n28558 = n27629 | n28076 ;
  assign n74685 = ~n28558 ;
  assign n28559 = n28072 & n74685 ;
  assign n28560 = n28314 | n28559 ;
  assign n28561 = n134 & n28560 ;
  assign n28562 = n27620 & n74611 ;
  assign n28563 = n28377 & n28562 ;
  assign n28564 = n28561 | n28563 ;
  assign n28565 = n68993 & n28564 ;
  assign n74686 = ~n28067 ;
  assign n28071 = n74686 & n28070 ;
  assign n28566 = n27637 | n28070 ;
  assign n74687 = ~n28566 ;
  assign n28567 = n28308 & n74687 ;
  assign n28568 = n28071 | n28567 ;
  assign n28569 = n134 & n28568 ;
  assign n28570 = n27628 & n74611 ;
  assign n28571 = n28377 & n28570 ;
  assign n28572 = n28569 | n28571 ;
  assign n28573 = n68716 & n28572 ;
  assign n74688 = ~n28571 ;
  assign n29004 = x98 & n74688 ;
  assign n74689 = ~n28569 ;
  assign n29005 = n74689 & n29004 ;
  assign n29006 = n28573 | n29005 ;
  assign n74690 = ~n28307 ;
  assign n28309 = n28065 & n74690 ;
  assign n28574 = n27645 | n28065 ;
  assign n74691 = ~n28574 ;
  assign n28575 = n28061 & n74691 ;
  assign n28576 = n28309 | n28575 ;
  assign n28577 = n134 & n28576 ;
  assign n28578 = n27636 & n74611 ;
  assign n28579 = n28377 & n28578 ;
  assign n28580 = n28577 | n28579 ;
  assign n28581 = n68545 & n28580 ;
  assign n74692 = ~n28056 ;
  assign n28060 = n74692 & n28059 ;
  assign n28582 = n27653 | n28059 ;
  assign n74693 = ~n28582 ;
  assign n28583 = n28303 & n74693 ;
  assign n28584 = n28060 | n28583 ;
  assign n28585 = n134 & n28584 ;
  assign n28586 = n27644 & n74611 ;
  assign n28587 = n28377 & n28586 ;
  assign n28588 = n28585 | n28587 ;
  assign n28589 = n68438 & n28588 ;
  assign n74694 = ~n28587 ;
  assign n28994 = x96 & n74694 ;
  assign n74695 = ~n28585 ;
  assign n28995 = n74695 & n28994 ;
  assign n28996 = n28589 | n28995 ;
  assign n74696 = ~n28302 ;
  assign n28304 = n28054 & n74696 ;
  assign n28590 = n27661 | n28054 ;
  assign n74697 = ~n28590 ;
  assign n28591 = n28050 & n74697 ;
  assign n28592 = n28304 | n28591 ;
  assign n28593 = n134 & n28592 ;
  assign n28594 = n27652 & n74611 ;
  assign n28595 = n28377 & n28594 ;
  assign n28596 = n28593 | n28595 ;
  assign n28597 = n68214 & n28596 ;
  assign n74698 = ~n28045 ;
  assign n28049 = n74698 & n28048 ;
  assign n28598 = n27669 | n28048 ;
  assign n74699 = ~n28598 ;
  assign n28599 = n28298 & n74699 ;
  assign n28600 = n28049 | n28599 ;
  assign n28601 = n134 & n28600 ;
  assign n28602 = n27660 & n74611 ;
  assign n28603 = n28377 & n28602 ;
  assign n28604 = n28601 | n28603 ;
  assign n28605 = n68058 & n28604 ;
  assign n74700 = ~n28603 ;
  assign n28983 = x94 & n74700 ;
  assign n74701 = ~n28601 ;
  assign n28984 = n74701 & n28983 ;
  assign n28985 = n28605 | n28984 ;
  assign n74702 = ~n28297 ;
  assign n28299 = n28043 & n74702 ;
  assign n28606 = n27677 | n28043 ;
  assign n74703 = ~n28606 ;
  assign n28607 = n28039 & n74703 ;
  assign n28608 = n28299 | n28607 ;
  assign n28609 = n134 & n28608 ;
  assign n28610 = n27668 & n74611 ;
  assign n28611 = n28377 & n28610 ;
  assign n28612 = n28609 | n28611 ;
  assign n28613 = n67986 & n28612 ;
  assign n74704 = ~n28034 ;
  assign n28038 = n74704 & n28037 ;
  assign n28614 = n27685 | n28037 ;
  assign n74705 = ~n28614 ;
  assign n28615 = n28293 & n74705 ;
  assign n28616 = n28038 | n28615 ;
  assign n28617 = n134 & n28616 ;
  assign n28618 = n27676 & n74611 ;
  assign n28619 = n28377 & n28618 ;
  assign n28620 = n28617 | n28619 ;
  assign n28621 = n67763 & n28620 ;
  assign n74706 = ~n28619 ;
  assign n28973 = x92 & n74706 ;
  assign n74707 = ~n28617 ;
  assign n28974 = n74707 & n28973 ;
  assign n28975 = n28621 | n28974 ;
  assign n74708 = ~n28292 ;
  assign n28294 = n28032 & n74708 ;
  assign n28622 = n27693 | n28032 ;
  assign n74709 = ~n28622 ;
  assign n28623 = n28028 & n74709 ;
  assign n28624 = n28294 | n28623 ;
  assign n28625 = n134 & n28624 ;
  assign n28626 = n27684 & n74611 ;
  assign n28627 = n28377 & n28626 ;
  assign n28628 = n28625 | n28627 ;
  assign n28629 = n67622 & n28628 ;
  assign n74710 = ~n28023 ;
  assign n28027 = n74710 & n28026 ;
  assign n28630 = n27701 | n28026 ;
  assign n74711 = ~n28630 ;
  assign n28631 = n28288 & n74711 ;
  assign n28632 = n28027 | n28631 ;
  assign n28633 = n134 & n28632 ;
  assign n28634 = n27692 & n74611 ;
  assign n28635 = n28377 & n28634 ;
  assign n28636 = n28633 | n28635 ;
  assign n28637 = n67531 & n28636 ;
  assign n74712 = ~n28635 ;
  assign n28963 = x90 & n74712 ;
  assign n74713 = ~n28633 ;
  assign n28964 = n74713 & n28963 ;
  assign n28965 = n28637 | n28964 ;
  assign n74714 = ~n28287 ;
  assign n28289 = n28021 & n74714 ;
  assign n28638 = n27709 | n28021 ;
  assign n74715 = ~n28638 ;
  assign n28639 = n28017 & n74715 ;
  assign n28640 = n28289 | n28639 ;
  assign n28641 = n134 & n28640 ;
  assign n28642 = n27700 & n74611 ;
  assign n28643 = n28377 & n28642 ;
  assign n28644 = n28641 | n28643 ;
  assign n28645 = n67348 & n28644 ;
  assign n74716 = ~n28012 ;
  assign n28016 = n74716 & n28015 ;
  assign n28646 = n27717 | n28015 ;
  assign n74717 = ~n28646 ;
  assign n28647 = n28283 & n74717 ;
  assign n28648 = n28016 | n28647 ;
  assign n28649 = n134 & n28648 ;
  assign n28650 = n27708 & n74611 ;
  assign n28651 = n28377 & n28650 ;
  assign n28652 = n28649 | n28651 ;
  assign n28653 = n67222 & n28652 ;
  assign n74718 = ~n28651 ;
  assign n28953 = x88 & n74718 ;
  assign n74719 = ~n28649 ;
  assign n28954 = n74719 & n28953 ;
  assign n28955 = n28653 | n28954 ;
  assign n74720 = ~n28282 ;
  assign n28284 = n28010 & n74720 ;
  assign n28654 = n27725 | n28010 ;
  assign n74721 = ~n28654 ;
  assign n28655 = n28006 & n74721 ;
  assign n28656 = n28284 | n28655 ;
  assign n28657 = n134 & n28656 ;
  assign n28658 = n27716 & n74611 ;
  assign n28659 = n28377 & n28658 ;
  assign n28660 = n28657 | n28659 ;
  assign n28661 = n67164 & n28660 ;
  assign n74722 = ~n28001 ;
  assign n28005 = n74722 & n28004 ;
  assign n28662 = n27733 | n28004 ;
  assign n74723 = ~n28662 ;
  assign n28663 = n28278 & n74723 ;
  assign n28664 = n28005 | n28663 ;
  assign n28665 = n134 & n28664 ;
  assign n28666 = n27724 & n74611 ;
  assign n28667 = n28377 & n28666 ;
  assign n28668 = n28665 | n28667 ;
  assign n28669 = n66979 & n28668 ;
  assign n74724 = ~n28667 ;
  assign n28943 = x86 & n74724 ;
  assign n74725 = ~n28665 ;
  assign n28944 = n74725 & n28943 ;
  assign n28945 = n28669 | n28944 ;
  assign n74726 = ~n28277 ;
  assign n28279 = n27999 & n74726 ;
  assign n28670 = n27741 | n27999 ;
  assign n74727 = ~n28670 ;
  assign n28671 = n27995 & n74727 ;
  assign n28672 = n28279 | n28671 ;
  assign n28673 = n134 & n28672 ;
  assign n28674 = n27732 & n74611 ;
  assign n28675 = n28377 & n28674 ;
  assign n28676 = n28673 | n28675 ;
  assign n28677 = n66868 & n28676 ;
  assign n74728 = ~n27990 ;
  assign n27994 = n74728 & n27993 ;
  assign n28678 = n27749 | n27993 ;
  assign n74729 = ~n28678 ;
  assign n28679 = n28273 & n74729 ;
  assign n28680 = n27994 | n28679 ;
  assign n28681 = n134 & n28680 ;
  assign n28682 = n27740 & n74611 ;
  assign n28683 = n28377 & n28682 ;
  assign n28684 = n28681 | n28683 ;
  assign n28685 = n66797 & n28684 ;
  assign n74730 = ~n28683 ;
  assign n28933 = x84 & n74730 ;
  assign n74731 = ~n28681 ;
  assign n28934 = n74731 & n28933 ;
  assign n28935 = n28685 | n28934 ;
  assign n74732 = ~n28272 ;
  assign n28274 = n27988 & n74732 ;
  assign n28686 = n27757 | n27988 ;
  assign n74733 = ~n28686 ;
  assign n28687 = n27984 & n74733 ;
  assign n28688 = n28274 | n28687 ;
  assign n28689 = n134 & n28688 ;
  assign n28690 = n27748 & n74611 ;
  assign n28691 = n28377 & n28690 ;
  assign n28692 = n28689 | n28691 ;
  assign n28693 = n66654 & n28692 ;
  assign n74734 = ~n27979 ;
  assign n27983 = n74734 & n27982 ;
  assign n28694 = n27765 | n27982 ;
  assign n74735 = ~n28694 ;
  assign n28695 = n28268 & n74735 ;
  assign n28696 = n27983 | n28695 ;
  assign n28697 = n134 & n28696 ;
  assign n28698 = n27756 & n74611 ;
  assign n28699 = n28377 & n28698 ;
  assign n28700 = n28697 | n28699 ;
  assign n28701 = n66560 & n28700 ;
  assign n74736 = ~n28699 ;
  assign n28923 = x82 & n74736 ;
  assign n74737 = ~n28697 ;
  assign n28924 = n74737 & n28923 ;
  assign n28925 = n28701 | n28924 ;
  assign n74738 = ~n28267 ;
  assign n28269 = n27977 & n74738 ;
  assign n28702 = n27773 | n27977 ;
  assign n74739 = ~n28702 ;
  assign n28703 = n27973 & n74739 ;
  assign n28704 = n28269 | n28703 ;
  assign n28705 = n134 & n28704 ;
  assign n28706 = n27764 & n74611 ;
  assign n28707 = n28377 & n28706 ;
  assign n28708 = n28705 | n28707 ;
  assign n28709 = n66505 & n28708 ;
  assign n74740 = ~n27968 ;
  assign n27972 = n74740 & n27971 ;
  assign n28710 = n27781 | n27971 ;
  assign n74741 = ~n28710 ;
  assign n28711 = n28263 & n74741 ;
  assign n28712 = n27972 | n28711 ;
  assign n28713 = n134 & n28712 ;
  assign n28714 = n27772 & n74611 ;
  assign n28715 = n28377 & n28714 ;
  assign n28716 = n28713 | n28715 ;
  assign n28717 = n66379 & n28716 ;
  assign n74742 = ~n28715 ;
  assign n28913 = x80 & n74742 ;
  assign n74743 = ~n28713 ;
  assign n28914 = n74743 & n28913 ;
  assign n28915 = n28717 | n28914 ;
  assign n74744 = ~n28262 ;
  assign n28264 = n27966 & n74744 ;
  assign n28718 = n27789 | n27966 ;
  assign n74745 = ~n28718 ;
  assign n28719 = n27962 & n74745 ;
  assign n28720 = n28264 | n28719 ;
  assign n28721 = n134 & n28720 ;
  assign n28722 = n27780 & n74611 ;
  assign n28723 = n28377 & n28722 ;
  assign n28724 = n28721 | n28723 ;
  assign n28725 = n66299 & n28724 ;
  assign n74746 = ~n27957 ;
  assign n27961 = n74746 & n27960 ;
  assign n28726 = n27797 | n27960 ;
  assign n74747 = ~n28726 ;
  assign n28727 = n28258 & n74747 ;
  assign n28728 = n27961 | n28727 ;
  assign n28729 = n134 & n28728 ;
  assign n28730 = n27788 & n74611 ;
  assign n28731 = n28377 & n28730 ;
  assign n28732 = n28729 | n28731 ;
  assign n28733 = n66244 & n28732 ;
  assign n74748 = ~n28731 ;
  assign n28903 = x78 & n74748 ;
  assign n74749 = ~n28729 ;
  assign n28904 = n74749 & n28903 ;
  assign n28905 = n28733 | n28904 ;
  assign n74750 = ~n28257 ;
  assign n28259 = n27955 & n74750 ;
  assign n28734 = n27805 | n27955 ;
  assign n74751 = ~n28734 ;
  assign n28735 = n27951 & n74751 ;
  assign n28736 = n28259 | n28735 ;
  assign n28737 = n134 & n28736 ;
  assign n28738 = n27796 & n74611 ;
  assign n28739 = n28377 & n28738 ;
  assign n28740 = n28737 | n28739 ;
  assign n28741 = n66145 & n28740 ;
  assign n74752 = ~n27946 ;
  assign n27950 = n74752 & n27949 ;
  assign n28742 = n27813 | n27949 ;
  assign n74753 = ~n28742 ;
  assign n28743 = n28253 & n74753 ;
  assign n28744 = n27950 | n28743 ;
  assign n28745 = n134 & n28744 ;
  assign n28746 = n27804 & n74611 ;
  assign n28747 = n28377 & n28746 ;
  assign n28748 = n28745 | n28747 ;
  assign n28749 = n66081 & n28748 ;
  assign n74754 = ~n28747 ;
  assign n28893 = x76 & n74754 ;
  assign n74755 = ~n28745 ;
  assign n28894 = n74755 & n28893 ;
  assign n28895 = n28749 | n28894 ;
  assign n74756 = ~n28252 ;
  assign n28254 = n27944 & n74756 ;
  assign n28750 = n27821 | n27944 ;
  assign n74757 = ~n28750 ;
  assign n28751 = n27940 & n74757 ;
  assign n28752 = n28254 | n28751 ;
  assign n28753 = n134 & n28752 ;
  assign n28754 = n27812 & n74611 ;
  assign n28755 = n28377 & n28754 ;
  assign n28756 = n28753 | n28755 ;
  assign n28757 = n66043 & n28756 ;
  assign n74758 = ~n27935 ;
  assign n27939 = n74758 & n27938 ;
  assign n28758 = n27829 | n27938 ;
  assign n74759 = ~n28758 ;
  assign n28759 = n28248 & n74759 ;
  assign n28760 = n27939 | n28759 ;
  assign n28761 = n134 & n28760 ;
  assign n28762 = n27820 & n74611 ;
  assign n28763 = n28377 & n28762 ;
  assign n28764 = n28761 | n28763 ;
  assign n28765 = n65960 & n28764 ;
  assign n74760 = ~n28763 ;
  assign n28883 = x74 & n74760 ;
  assign n74761 = ~n28761 ;
  assign n28884 = n74761 & n28883 ;
  assign n28885 = n28765 | n28884 ;
  assign n74762 = ~n28247 ;
  assign n28249 = n27933 & n74762 ;
  assign n28766 = n27837 | n27933 ;
  assign n74763 = ~n28766 ;
  assign n28767 = n27929 & n74763 ;
  assign n28768 = n28249 | n28767 ;
  assign n28769 = n134 & n28768 ;
  assign n28770 = n27828 & n74611 ;
  assign n28771 = n28377 & n28770 ;
  assign n28772 = n28769 | n28771 ;
  assign n28773 = n65909 & n28772 ;
  assign n74764 = ~n27924 ;
  assign n27928 = n74764 & n27927 ;
  assign n28774 = n27845 | n27927 ;
  assign n74765 = ~n28774 ;
  assign n28775 = n28243 & n74765 ;
  assign n28776 = n27928 | n28775 ;
  assign n28777 = n134 & n28776 ;
  assign n28778 = n27836 & n74611 ;
  assign n28779 = n28377 & n28778 ;
  assign n28780 = n28777 | n28779 ;
  assign n28781 = n65877 & n28780 ;
  assign n74766 = ~n28779 ;
  assign n28873 = x72 & n74766 ;
  assign n74767 = ~n28777 ;
  assign n28874 = n74767 & n28873 ;
  assign n28875 = n28781 | n28874 ;
  assign n74768 = ~n28242 ;
  assign n28244 = n27922 & n74768 ;
  assign n28782 = n27854 | n27922 ;
  assign n74769 = ~n28782 ;
  assign n28783 = n27918 & n74769 ;
  assign n28784 = n28244 | n28783 ;
  assign n28785 = n134 & n28784 ;
  assign n28786 = n27844 & n74611 ;
  assign n28787 = n28377 & n28786 ;
  assign n28788 = n28785 | n28787 ;
  assign n28789 = n65820 & n28788 ;
  assign n74770 = ~n27914 ;
  assign n28240 = n74770 & n27917 ;
  assign n28790 = n27863 | n27917 ;
  assign n74771 = ~n28790 ;
  assign n28791 = n28238 & n74771 ;
  assign n28792 = n28240 | n28791 ;
  assign n28793 = n134 & n28792 ;
  assign n28794 = n27853 & n74611 ;
  assign n28795 = n28377 & n28794 ;
  assign n28796 = n28793 | n28795 ;
  assign n28797 = n65791 & n28796 ;
  assign n74772 = ~n28795 ;
  assign n28863 = x70 & n74772 ;
  assign n74773 = ~n28793 ;
  assign n28864 = n74773 & n28863 ;
  assign n28865 = n28797 | n28864 ;
  assign n74774 = ~n28236 ;
  assign n28237 = n27912 & n74774 ;
  assign n28798 = n27905 | n28233 ;
  assign n28799 = n27871 | n27912 ;
  assign n74775 = ~n28799 ;
  assign n28800 = n28798 & n74775 ;
  assign n28801 = n28237 | n28800 ;
  assign n28802 = n134 & n28801 ;
  assign n28803 = n27862 & n74611 ;
  assign n28804 = n28377 & n28803 ;
  assign n28805 = n28802 | n28804 ;
  assign n28806 = n65772 & n28805 ;
  assign n74776 = ~n27905 ;
  assign n28234 = n74776 & n28233 ;
  assign n28807 = n27877 | n28233 ;
  assign n74777 = ~n28807 ;
  assign n28808 = n27904 & n74777 ;
  assign n28809 = n28234 | n28808 ;
  assign n28810 = n134 & n28809 ;
  assign n28811 = n27870 & n74611 ;
  assign n28812 = n28377 & n28811 ;
  assign n28813 = n28810 | n28812 ;
  assign n28814 = n65746 & n28813 ;
  assign n74778 = ~n28812 ;
  assign n28852 = x68 & n74778 ;
  assign n74779 = ~n28810 ;
  assign n28853 = n74779 & n28852 ;
  assign n28854 = n28814 | n28853 ;
  assign n74780 = ~n28229 ;
  assign n28230 = n27903 & n74780 ;
  assign n28815 = n27899 | n27903 ;
  assign n74781 = ~n28815 ;
  assign n28816 = n27898 & n74781 ;
  assign n28817 = n28230 | n28816 ;
  assign n28818 = n134 & n28817 ;
  assign n28819 = n27876 & n74611 ;
  assign n28820 = n28377 & n28819 ;
  assign n28821 = n28818 | n28820 ;
  assign n28822 = n65721 & n28821 ;
  assign n28823 = n27895 & n27897 ;
  assign n28824 = n74437 & n28823 ;
  assign n74782 = ~n28824 ;
  assign n28825 = n28228 & n74782 ;
  assign n28826 = n134 & n28825 ;
  assign n28827 = n74611 & n28225 ;
  assign n28828 = n28377 & n28827 ;
  assign n28829 = n28826 | n28828 ;
  assign n28830 = n65686 & n28829 ;
  assign n74783 = ~n28828 ;
  assign n28842 = x66 & n74783 ;
  assign n74784 = ~n28826 ;
  assign n28843 = n74784 & n28842 ;
  assign n28844 = n28830 | n28843 ;
  assign n28223 = n27897 & n134 ;
  assign n28224 = x64 & n134 ;
  assign n74785 = ~n28224 ;
  assign n28831 = x5 & n74785 ;
  assign n28832 = n28223 | n28831 ;
  assign n28833 = x65 & n28832 ;
  assign n28834 = n74611 & n28377 ;
  assign n74786 = ~n28834 ;
  assign n28835 = n27897 & n74786 ;
  assign n28836 = x65 | n28835 ;
  assign n28837 = n28831 | n28836 ;
  assign n74787 = ~n28833 ;
  assign n28838 = n74787 & n28837 ;
  assign n74788 = ~x4 ;
  assign n28839 = n74788 & x64 ;
  assign n28840 = n28838 | n28839 ;
  assign n28841 = n65670 & n28832 ;
  assign n74789 = ~n28841 ;
  assign n28845 = n28840 & n74789 ;
  assign n28846 = n28844 | n28845 ;
  assign n74790 = ~n28830 ;
  assign n28847 = n74790 & n28846 ;
  assign n74791 = ~n28820 ;
  assign n28848 = x67 & n74791 ;
  assign n74792 = ~n28818 ;
  assign n28849 = n74792 & n28848 ;
  assign n28850 = n28822 | n28849 ;
  assign n28851 = n28847 | n28850 ;
  assign n74793 = ~n28822 ;
  assign n28855 = n74793 & n28851 ;
  assign n28856 = n28854 | n28855 ;
  assign n74794 = ~n28814 ;
  assign n28857 = n74794 & n28856 ;
  assign n74795 = ~n28804 ;
  assign n28858 = x69 & n74795 ;
  assign n74796 = ~n28802 ;
  assign n28859 = n74796 & n28858 ;
  assign n28860 = n28806 | n28859 ;
  assign n28862 = n28857 | n28860 ;
  assign n74797 = ~n28806 ;
  assign n28866 = n74797 & n28862 ;
  assign n28867 = n28865 | n28866 ;
  assign n74798 = ~n28797 ;
  assign n28868 = n74798 & n28867 ;
  assign n74799 = ~n28787 ;
  assign n28869 = x71 & n74799 ;
  assign n74800 = ~n28785 ;
  assign n28870 = n74800 & n28869 ;
  assign n28871 = n28789 | n28870 ;
  assign n28872 = n28868 | n28871 ;
  assign n74801 = ~n28789 ;
  assign n28876 = n74801 & n28872 ;
  assign n28877 = n28875 | n28876 ;
  assign n74802 = ~n28781 ;
  assign n28878 = n74802 & n28877 ;
  assign n74803 = ~n28771 ;
  assign n28879 = x73 & n74803 ;
  assign n74804 = ~n28769 ;
  assign n28880 = n74804 & n28879 ;
  assign n28881 = n28773 | n28880 ;
  assign n28882 = n28878 | n28881 ;
  assign n74805 = ~n28773 ;
  assign n28886 = n74805 & n28882 ;
  assign n28887 = n28885 | n28886 ;
  assign n74806 = ~n28765 ;
  assign n28888 = n74806 & n28887 ;
  assign n74807 = ~n28755 ;
  assign n28889 = x75 & n74807 ;
  assign n74808 = ~n28753 ;
  assign n28890 = n74808 & n28889 ;
  assign n28891 = n28757 | n28890 ;
  assign n28892 = n28888 | n28891 ;
  assign n74809 = ~n28757 ;
  assign n28896 = n74809 & n28892 ;
  assign n28897 = n28895 | n28896 ;
  assign n74810 = ~n28749 ;
  assign n28898 = n74810 & n28897 ;
  assign n74811 = ~n28739 ;
  assign n28899 = x77 & n74811 ;
  assign n74812 = ~n28737 ;
  assign n28900 = n74812 & n28899 ;
  assign n28901 = n28741 | n28900 ;
  assign n28902 = n28898 | n28901 ;
  assign n74813 = ~n28741 ;
  assign n28906 = n74813 & n28902 ;
  assign n28907 = n28905 | n28906 ;
  assign n74814 = ~n28733 ;
  assign n28908 = n74814 & n28907 ;
  assign n74815 = ~n28723 ;
  assign n28909 = x79 & n74815 ;
  assign n74816 = ~n28721 ;
  assign n28910 = n74816 & n28909 ;
  assign n28911 = n28725 | n28910 ;
  assign n28912 = n28908 | n28911 ;
  assign n74817 = ~n28725 ;
  assign n28916 = n74817 & n28912 ;
  assign n28917 = n28915 | n28916 ;
  assign n74818 = ~n28717 ;
  assign n28918 = n74818 & n28917 ;
  assign n74819 = ~n28707 ;
  assign n28919 = x81 & n74819 ;
  assign n74820 = ~n28705 ;
  assign n28920 = n74820 & n28919 ;
  assign n28921 = n28709 | n28920 ;
  assign n28922 = n28918 | n28921 ;
  assign n74821 = ~n28709 ;
  assign n28926 = n74821 & n28922 ;
  assign n28927 = n28925 | n28926 ;
  assign n74822 = ~n28701 ;
  assign n28928 = n74822 & n28927 ;
  assign n74823 = ~n28691 ;
  assign n28929 = x83 & n74823 ;
  assign n74824 = ~n28689 ;
  assign n28930 = n74824 & n28929 ;
  assign n28931 = n28693 | n28930 ;
  assign n28932 = n28928 | n28931 ;
  assign n74825 = ~n28693 ;
  assign n28936 = n74825 & n28932 ;
  assign n28937 = n28935 | n28936 ;
  assign n74826 = ~n28685 ;
  assign n28938 = n74826 & n28937 ;
  assign n74827 = ~n28675 ;
  assign n28939 = x85 & n74827 ;
  assign n74828 = ~n28673 ;
  assign n28940 = n74828 & n28939 ;
  assign n28941 = n28677 | n28940 ;
  assign n28942 = n28938 | n28941 ;
  assign n74829 = ~n28677 ;
  assign n28946 = n74829 & n28942 ;
  assign n28947 = n28945 | n28946 ;
  assign n74830 = ~n28669 ;
  assign n28948 = n74830 & n28947 ;
  assign n74831 = ~n28659 ;
  assign n28949 = x87 & n74831 ;
  assign n74832 = ~n28657 ;
  assign n28950 = n74832 & n28949 ;
  assign n28951 = n28661 | n28950 ;
  assign n28952 = n28948 | n28951 ;
  assign n74833 = ~n28661 ;
  assign n28956 = n74833 & n28952 ;
  assign n28957 = n28955 | n28956 ;
  assign n74834 = ~n28653 ;
  assign n28958 = n74834 & n28957 ;
  assign n74835 = ~n28643 ;
  assign n28959 = x89 & n74835 ;
  assign n74836 = ~n28641 ;
  assign n28960 = n74836 & n28959 ;
  assign n28961 = n28645 | n28960 ;
  assign n28962 = n28958 | n28961 ;
  assign n74837 = ~n28645 ;
  assign n28966 = n74837 & n28962 ;
  assign n28967 = n28965 | n28966 ;
  assign n74838 = ~n28637 ;
  assign n28968 = n74838 & n28967 ;
  assign n74839 = ~n28627 ;
  assign n28969 = x91 & n74839 ;
  assign n74840 = ~n28625 ;
  assign n28970 = n74840 & n28969 ;
  assign n28971 = n28629 | n28970 ;
  assign n28972 = n28968 | n28971 ;
  assign n74841 = ~n28629 ;
  assign n28976 = n74841 & n28972 ;
  assign n28977 = n28975 | n28976 ;
  assign n74842 = ~n28621 ;
  assign n28978 = n74842 & n28977 ;
  assign n74843 = ~n28611 ;
  assign n28979 = x93 & n74843 ;
  assign n74844 = ~n28609 ;
  assign n28980 = n74844 & n28979 ;
  assign n28981 = n28613 | n28980 ;
  assign n28982 = n28978 | n28981 ;
  assign n74845 = ~n28613 ;
  assign n28986 = n74845 & n28982 ;
  assign n28987 = n28985 | n28986 ;
  assign n74846 = ~n28605 ;
  assign n28988 = n74846 & n28987 ;
  assign n74847 = ~n28595 ;
  assign n28989 = x95 & n74847 ;
  assign n74848 = ~n28593 ;
  assign n28990 = n74848 & n28989 ;
  assign n28991 = n28597 | n28990 ;
  assign n28993 = n28988 | n28991 ;
  assign n74849 = ~n28597 ;
  assign n28997 = n74849 & n28993 ;
  assign n28998 = n28996 | n28997 ;
  assign n74850 = ~n28589 ;
  assign n28999 = n74850 & n28998 ;
  assign n74851 = ~n28579 ;
  assign n29000 = x97 & n74851 ;
  assign n74852 = ~n28577 ;
  assign n29001 = n74852 & n29000 ;
  assign n29002 = n28581 | n29001 ;
  assign n29003 = n28999 | n29002 ;
  assign n74853 = ~n28581 ;
  assign n29007 = n74853 & n29003 ;
  assign n29008 = n29006 | n29007 ;
  assign n74854 = ~n28573 ;
  assign n29009 = n74854 & n29008 ;
  assign n74855 = ~n28563 ;
  assign n29010 = x99 & n74855 ;
  assign n74856 = ~n28561 ;
  assign n29011 = n74856 & n29010 ;
  assign n29012 = n28565 | n29011 ;
  assign n29013 = n29009 | n29012 ;
  assign n74857 = ~n28565 ;
  assign n29017 = n74857 & n29013 ;
  assign n29018 = n29016 | n29017 ;
  assign n74858 = ~n28557 ;
  assign n29019 = n74858 & n29018 ;
  assign n74859 = ~n28547 ;
  assign n29020 = x101 & n74859 ;
  assign n74860 = ~n28545 ;
  assign n29021 = n74860 & n29020 ;
  assign n29022 = n28549 | n29021 ;
  assign n29023 = n29019 | n29022 ;
  assign n74861 = ~n28549 ;
  assign n29027 = n74861 & n29023 ;
  assign n29028 = n29026 | n29027 ;
  assign n74862 = ~n28541 ;
  assign n29029 = n74862 & n29028 ;
  assign n74863 = ~n28531 ;
  assign n29030 = x103 & n74863 ;
  assign n74864 = ~n28529 ;
  assign n29031 = n74864 & n29030 ;
  assign n29032 = n28533 | n29031 ;
  assign n29034 = n29029 | n29032 ;
  assign n74865 = ~n28533 ;
  assign n29038 = n74865 & n29034 ;
  assign n29039 = n29037 | n29038 ;
  assign n74866 = ~n28525 ;
  assign n29040 = n74866 & n29039 ;
  assign n74867 = ~n28515 ;
  assign n29041 = x105 & n74867 ;
  assign n74868 = ~n28513 ;
  assign n29042 = n74868 & n29041 ;
  assign n29043 = n28517 | n29042 ;
  assign n29045 = n29040 | n29043 ;
  assign n74869 = ~n28517 ;
  assign n29049 = n74869 & n29045 ;
  assign n29050 = n29048 | n29049 ;
  assign n74870 = ~n28509 ;
  assign n29051 = n74870 & n29050 ;
  assign n74871 = ~n28499 ;
  assign n29052 = x107 & n74871 ;
  assign n74872 = ~n28497 ;
  assign n29053 = n74872 & n29052 ;
  assign n29054 = n28501 | n29053 ;
  assign n29056 = n29051 | n29054 ;
  assign n74873 = ~n28501 ;
  assign n29061 = n74873 & n29056 ;
  assign n29062 = n29059 | n29061 ;
  assign n74874 = ~n28493 ;
  assign n29063 = n74874 & n29062 ;
  assign n74875 = ~n28483 ;
  assign n29064 = x109 & n74875 ;
  assign n74876 = ~n28481 ;
  assign n29065 = n74876 & n29064 ;
  assign n29066 = n28485 | n29065 ;
  assign n29067 = n29063 | n29066 ;
  assign n74877 = ~n28485 ;
  assign n29071 = n74877 & n29067 ;
  assign n29072 = n29070 | n29071 ;
  assign n74878 = ~n28477 ;
  assign n29073 = n74878 & n29072 ;
  assign n74879 = ~n28467 ;
  assign n29074 = x111 & n74879 ;
  assign n74880 = ~n28465 ;
  assign n29075 = n74880 & n29074 ;
  assign n29076 = n28469 | n29075 ;
  assign n29077 = n29073 | n29076 ;
  assign n74881 = ~n28469 ;
  assign n29081 = n74881 & n29077 ;
  assign n29082 = n29080 | n29081 ;
  assign n74882 = ~n28461 ;
  assign n29083 = n74882 & n29082 ;
  assign n74883 = ~n28451 ;
  assign n29084 = x113 & n74883 ;
  assign n74884 = ~n28449 ;
  assign n29085 = n74884 & n29084 ;
  assign n29086 = n28453 | n29085 ;
  assign n29087 = n29083 | n29086 ;
  assign n74885 = ~n28453 ;
  assign n29091 = n74885 & n29087 ;
  assign n29092 = n29090 | n29091 ;
  assign n74886 = ~n28445 ;
  assign n29093 = n74886 & n29092 ;
  assign n74887 = ~n28435 ;
  assign n29094 = x115 & n74887 ;
  assign n74888 = ~n28433 ;
  assign n29095 = n74888 & n29094 ;
  assign n29096 = n28437 | n29095 ;
  assign n29097 = n29093 | n29096 ;
  assign n74889 = ~n28437 ;
  assign n29102 = n74889 & n29097 ;
  assign n29103 = n29100 | n29102 ;
  assign n74890 = ~n28429 ;
  assign n29104 = n74890 & n29103 ;
  assign n74891 = ~n28419 ;
  assign n29105 = x117 & n74891 ;
  assign n74892 = ~n28417 ;
  assign n29106 = n74892 & n29105 ;
  assign n29107 = n28421 | n29106 ;
  assign n29108 = n29104 | n29107 ;
  assign n74893 = ~n28421 ;
  assign n29112 = n74893 & n29108 ;
  assign n29113 = n29111 | n29112 ;
  assign n74894 = ~n28413 ;
  assign n29114 = n74894 & n29113 ;
  assign n74895 = ~n28403 ;
  assign n29115 = x119 & n74895 ;
  assign n74896 = ~n28401 ;
  assign n29116 = n74896 & n29115 ;
  assign n29117 = n28405 | n29116 ;
  assign n29118 = n29114 | n29117 ;
  assign n74897 = ~n28405 ;
  assign n29122 = n74897 & n29118 ;
  assign n29123 = n29121 | n29122 ;
  assign n74898 = ~n28397 ;
  assign n29124 = n74898 & n29123 ;
  assign n74899 = ~n28387 ;
  assign n29125 = x121 & n74899 ;
  assign n74900 = ~n28385 ;
  assign n29126 = n74900 & n29125 ;
  assign n29127 = n28389 | n29126 ;
  assign n29128 = n29124 | n29127 ;
  assign n74901 = ~n28389 ;
  assign n29132 = n74901 & n29128 ;
  assign n29133 = n29131 | n29132 ;
  assign n74902 = ~n28381 ;
  assign n29134 = n74902 & n29133 ;
  assign n29135 = n27437 | n28216 ;
  assign n29136 = n28212 | n29135 ;
  assign n74903 = ~n29136 ;
  assign n29137 = n28204 & n74903 ;
  assign n29138 = n28212 | n28216 ;
  assign n74904 = ~n28376 ;
  assign n29139 = n74904 & n29138 ;
  assign n29140 = n29137 | n29139 ;
  assign n29141 = n134 & n29140 ;
  assign n29142 = n27311 & n28211 ;
  assign n29143 = n28377 & n29142 ;
  assign n29144 = n29141 | n29143 ;
  assign n74905 = ~x123 ;
  assign n29145 = n74905 & n29144 ;
  assign n74906 = ~n29143 ;
  assign n29146 = x123 & n74906 ;
  assign n74907 = ~n29141 ;
  assign n29147 = n74907 & n29146 ;
  assign n29148 = n65369 | n29147 ;
  assign n29149 = n29145 | n29148 ;
  assign n29150 = n29134 | n29149 ;
  assign n74908 = ~n28217 ;
  assign n29151 = n74908 & n29144 ;
  assign n74909 = ~n29151 ;
  assign n29152 = n29150 & n74909 ;
  assign n30122 = n28381 | n29147 ;
  assign n30123 = n29145 | n30122 ;
  assign n74910 = ~n30123 ;
  assign n30124 = n29133 & n74910 ;
  assign n29154 = x64 & n74786 ;
  assign n74911 = ~n29154 ;
  assign n29155 = x5 & n74911 ;
  assign n29156 = n28223 | n29155 ;
  assign n29157 = x65 & n29156 ;
  assign n74912 = ~n29157 ;
  assign n29158 = n28837 & n74912 ;
  assign n29159 = n28839 | n29158 ;
  assign n29160 = n74789 & n29159 ;
  assign n29162 = n28844 | n29160 ;
  assign n29163 = n74790 & n29162 ;
  assign n29164 = n28850 | n29163 ;
  assign n29165 = n74793 & n29164 ;
  assign n29166 = n28854 | n29165 ;
  assign n29167 = n74794 & n29166 ;
  assign n29168 = n28860 | n29167 ;
  assign n29169 = n74797 & n29168 ;
  assign n29170 = n28865 | n29169 ;
  assign n29171 = n74798 & n29170 ;
  assign n29172 = n28871 | n29171 ;
  assign n29173 = n74801 & n29172 ;
  assign n29174 = n28875 | n29173 ;
  assign n29175 = n74802 & n29174 ;
  assign n29176 = n28881 | n29175 ;
  assign n29177 = n74805 & n29176 ;
  assign n29178 = n28885 | n29177 ;
  assign n29179 = n74806 & n29178 ;
  assign n29180 = n28891 | n29179 ;
  assign n29181 = n74809 & n29180 ;
  assign n29182 = n28895 | n29181 ;
  assign n29183 = n74810 & n29182 ;
  assign n29184 = n28901 | n29183 ;
  assign n29185 = n74813 & n29184 ;
  assign n29186 = n28905 | n29185 ;
  assign n29187 = n74814 & n29186 ;
  assign n29188 = n28911 | n29187 ;
  assign n29189 = n74817 & n29188 ;
  assign n29190 = n28915 | n29189 ;
  assign n29191 = n74818 & n29190 ;
  assign n29192 = n28921 | n29191 ;
  assign n29193 = n74821 & n29192 ;
  assign n29194 = n28925 | n29193 ;
  assign n29195 = n74822 & n29194 ;
  assign n29196 = n28931 | n29195 ;
  assign n29197 = n74825 & n29196 ;
  assign n29198 = n28935 | n29197 ;
  assign n29199 = n74826 & n29198 ;
  assign n29200 = n28941 | n29199 ;
  assign n29201 = n74829 & n29200 ;
  assign n29202 = n28945 | n29201 ;
  assign n29203 = n74830 & n29202 ;
  assign n29204 = n28951 | n29203 ;
  assign n29205 = n74833 & n29204 ;
  assign n29206 = n28955 | n29205 ;
  assign n29207 = n74834 & n29206 ;
  assign n29208 = n28961 | n29207 ;
  assign n29209 = n74837 & n29208 ;
  assign n29210 = n28965 | n29209 ;
  assign n29211 = n74838 & n29210 ;
  assign n29212 = n28971 | n29211 ;
  assign n29213 = n74841 & n29212 ;
  assign n29214 = n28975 | n29213 ;
  assign n29215 = n74842 & n29214 ;
  assign n29216 = n28981 | n29215 ;
  assign n29217 = n74845 & n29216 ;
  assign n29218 = n28985 | n29217 ;
  assign n29219 = n74846 & n29218 ;
  assign n29220 = n28991 | n29219 ;
  assign n29221 = n74849 & n29220 ;
  assign n29222 = n28996 | n29221 ;
  assign n29223 = n74850 & n29222 ;
  assign n29224 = n29002 | n29223 ;
  assign n29225 = n74853 & n29224 ;
  assign n29226 = n29006 | n29225 ;
  assign n29227 = n74854 & n29226 ;
  assign n29228 = n29012 | n29227 ;
  assign n29229 = n74857 & n29228 ;
  assign n29230 = n29016 | n29229 ;
  assign n29231 = n74858 & n29230 ;
  assign n29232 = n29022 | n29231 ;
  assign n29233 = n74861 & n29232 ;
  assign n29234 = n29026 | n29233 ;
  assign n29235 = n74862 & n29234 ;
  assign n29236 = n29032 | n29235 ;
  assign n29237 = n74865 & n29236 ;
  assign n29238 = n29037 | n29237 ;
  assign n29239 = n74866 & n29238 ;
  assign n29240 = n29043 | n29239 ;
  assign n29241 = n74869 & n29240 ;
  assign n29242 = n29048 | n29241 ;
  assign n29243 = n74870 & n29242 ;
  assign n29244 = n29054 | n29243 ;
  assign n29245 = n74873 & n29244 ;
  assign n29246 = n29059 | n29245 ;
  assign n29247 = n74874 & n29246 ;
  assign n29248 = n29066 | n29247 ;
  assign n29249 = n74877 & n29248 ;
  assign n29250 = n29070 | n29249 ;
  assign n29251 = n74878 & n29250 ;
  assign n29252 = n29076 | n29251 ;
  assign n29253 = n74881 & n29252 ;
  assign n29254 = n29080 | n29253 ;
  assign n29255 = n74882 & n29254 ;
  assign n29256 = n29086 | n29255 ;
  assign n29257 = n74885 & n29256 ;
  assign n29258 = n29090 | n29257 ;
  assign n29259 = n74886 & n29258 ;
  assign n29260 = n29096 | n29259 ;
  assign n29261 = n74889 & n29260 ;
  assign n29262 = n29100 | n29261 ;
  assign n29263 = n74890 & n29262 ;
  assign n29264 = n29107 | n29263 ;
  assign n29265 = n74893 & n29264 ;
  assign n29266 = n29111 | n29265 ;
  assign n29267 = n74894 & n29266 ;
  assign n29268 = n29117 | n29267 ;
  assign n29269 = n74897 & n29268 ;
  assign n29270 = n29121 | n29269 ;
  assign n29271 = n74898 & n29270 ;
  assign n29272 = n29127 | n29271 ;
  assign n29273 = n74901 & n29272 ;
  assign n29787 = n29131 | n29273 ;
  assign n29788 = n74902 & n29787 ;
  assign n30125 = n29145 | n29147 ;
  assign n74913 = ~n29788 ;
  assign n30126 = n74913 & n30125 ;
  assign n30127 = n30124 | n30126 ;
  assign n133 = ~n29152 ;
  assign n30128 = n133 & n30127 ;
  assign n30129 = n28217 & n29144 ;
  assign n30130 = n29150 & n30129 ;
  assign n30131 = n30128 | n30130 ;
  assign n30137 = n73619 & n30131 ;
  assign n74915 = ~n29132 ;
  assign n29274 = n29131 & n74915 ;
  assign n29275 = n28389 | n29131 ;
  assign n74916 = ~n29275 ;
  assign n29276 = n29272 & n74916 ;
  assign n29277 = n29274 | n29276 ;
  assign n29278 = n133 & n29277 ;
  assign n29279 = n28380 & n74909 ;
  assign n29280 = n29150 & n29279 ;
  assign n29281 = n29278 | n29280 ;
  assign n29282 = n74905 & n29281 ;
  assign n74917 = ~n29271 ;
  assign n29283 = n29127 & n74917 ;
  assign n29284 = n28397 | n29127 ;
  assign n74918 = ~n29284 ;
  assign n29285 = n29123 & n74918 ;
  assign n29286 = n29283 | n29285 ;
  assign n29287 = n133 & n29286 ;
  assign n29288 = n28388 & n74909 ;
  assign n29289 = n29150 & n29288 ;
  assign n29290 = n29287 | n29289 ;
  assign n29291 = n74431 & n29290 ;
  assign n74919 = ~n29122 ;
  assign n29292 = n29121 & n74919 ;
  assign n29293 = n28405 | n29121 ;
  assign n74920 = ~n29293 ;
  assign n29294 = n29268 & n74920 ;
  assign n29295 = n29292 | n29294 ;
  assign n29296 = n133 & n29295 ;
  assign n29297 = n28396 & n74909 ;
  assign n29298 = n29150 & n29297 ;
  assign n29299 = n29296 | n29298 ;
  assign n29300 = n74029 & n29299 ;
  assign n74921 = ~n29267 ;
  assign n29301 = n29117 & n74921 ;
  assign n29302 = n28413 | n29117 ;
  assign n74922 = ~n29302 ;
  assign n29303 = n29113 & n74922 ;
  assign n29304 = n29301 | n29303 ;
  assign n29305 = n133 & n29304 ;
  assign n29306 = n28404 & n74909 ;
  assign n29307 = n29150 & n29306 ;
  assign n29308 = n29305 | n29307 ;
  assign n29309 = n74021 & n29308 ;
  assign n74923 = ~n29112 ;
  assign n29310 = n29111 & n74923 ;
  assign n29311 = n28421 | n29111 ;
  assign n74924 = ~n29311 ;
  assign n29312 = n29264 & n74924 ;
  assign n29313 = n29310 | n29312 ;
  assign n29314 = n133 & n29313 ;
  assign n29315 = n28412 & n74909 ;
  assign n29316 = n29150 & n29315 ;
  assign n29317 = n29314 | n29316 ;
  assign n29318 = n73617 & n29317 ;
  assign n74925 = ~n29263 ;
  assign n29319 = n29107 & n74925 ;
  assign n29320 = n28429 | n29107 ;
  assign n74926 = ~n29320 ;
  assign n29321 = n29103 & n74926 ;
  assign n29322 = n29319 | n29321 ;
  assign n29323 = n133 & n29322 ;
  assign n29324 = n28420 & n74909 ;
  assign n29325 = n29150 & n29324 ;
  assign n29326 = n29323 | n29325 ;
  assign n29327 = n73188 & n29326 ;
  assign n74927 = ~n29102 ;
  assign n29328 = n29100 & n74927 ;
  assign n29101 = n28437 | n29100 ;
  assign n74928 = ~n29101 ;
  assign n29329 = n29097 & n74928 ;
  assign n29330 = n29328 | n29329 ;
  assign n29331 = n133 & n29330 ;
  assign n29332 = n28428 & n74909 ;
  assign n29333 = n29150 & n29332 ;
  assign n29334 = n29331 | n29333 ;
  assign n29335 = n73177 & n29334 ;
  assign n74929 = ~n29259 ;
  assign n29336 = n29096 & n74929 ;
  assign n29337 = n28445 | n29096 ;
  assign n74930 = ~n29337 ;
  assign n29338 = n29092 & n74930 ;
  assign n29339 = n29336 | n29338 ;
  assign n29340 = n133 & n29339 ;
  assign n29341 = n28436 & n74909 ;
  assign n29342 = n29150 & n29341 ;
  assign n29343 = n29340 | n29342 ;
  assign n29344 = n72752 & n29343 ;
  assign n74931 = ~n29091 ;
  assign n29345 = n29090 & n74931 ;
  assign n29346 = n28453 | n29090 ;
  assign n74932 = ~n29346 ;
  assign n29347 = n29256 & n74932 ;
  assign n29348 = n29345 | n29347 ;
  assign n29349 = n133 & n29348 ;
  assign n29350 = n28444 & n74909 ;
  assign n29351 = n29150 & n29350 ;
  assign n29352 = n29349 | n29351 ;
  assign n29353 = n72393 & n29352 ;
  assign n74933 = ~n29255 ;
  assign n29354 = n29086 & n74933 ;
  assign n29355 = n28461 | n29086 ;
  assign n74934 = ~n29355 ;
  assign n29356 = n29082 & n74934 ;
  assign n29357 = n29354 | n29356 ;
  assign n29358 = n133 & n29357 ;
  assign n29359 = n28452 & n74909 ;
  assign n29360 = n29150 & n29359 ;
  assign n29361 = n29358 | n29360 ;
  assign n29362 = n72385 & n29361 ;
  assign n74935 = ~n29081 ;
  assign n29363 = n29080 & n74935 ;
  assign n29364 = n28469 | n29080 ;
  assign n74936 = ~n29364 ;
  assign n29365 = n29252 & n74936 ;
  assign n29366 = n29363 | n29365 ;
  assign n29367 = n133 & n29366 ;
  assign n29368 = n28460 & n74909 ;
  assign n29369 = n29150 & n29368 ;
  assign n29370 = n29367 | n29369 ;
  assign n29371 = n72025 & n29370 ;
  assign n74937 = ~n29251 ;
  assign n29372 = n29076 & n74937 ;
  assign n29373 = n28477 | n29076 ;
  assign n74938 = ~n29373 ;
  assign n29374 = n29072 & n74938 ;
  assign n29375 = n29372 | n29374 ;
  assign n29376 = n133 & n29375 ;
  assign n29377 = n28468 & n74909 ;
  assign n29378 = n29150 & n29377 ;
  assign n29379 = n29376 | n29378 ;
  assign n29380 = n71645 & n29379 ;
  assign n74939 = ~n29071 ;
  assign n29381 = n29070 & n74939 ;
  assign n29382 = n28485 | n29070 ;
  assign n74940 = ~n29382 ;
  assign n29383 = n29248 & n74940 ;
  assign n29384 = n29381 | n29383 ;
  assign n29385 = n133 & n29384 ;
  assign n29386 = n28476 & n74909 ;
  assign n29387 = n29150 & n29386 ;
  assign n29388 = n29385 | n29387 ;
  assign n29389 = n71633 & n29388 ;
  assign n74941 = ~n29247 ;
  assign n29390 = n29066 & n74941 ;
  assign n29391 = n28493 | n29066 ;
  assign n74942 = ~n29391 ;
  assign n29392 = n29062 & n74942 ;
  assign n29393 = n29390 | n29392 ;
  assign n29394 = n133 & n29393 ;
  assign n29395 = n28484 & n74909 ;
  assign n29396 = n29150 & n29395 ;
  assign n29397 = n29394 | n29396 ;
  assign n29398 = n71253 & n29397 ;
  assign n74943 = ~n29061 ;
  assign n29399 = n29059 & n74943 ;
  assign n29060 = n28501 | n29059 ;
  assign n74944 = ~n29060 ;
  assign n29400 = n29056 & n74944 ;
  assign n29401 = n29399 | n29400 ;
  assign n29402 = n133 & n29401 ;
  assign n29403 = n28492 & n74909 ;
  assign n29404 = n29150 & n29403 ;
  assign n29405 = n29402 | n29404 ;
  assign n29406 = n70935 & n29405 ;
  assign n74945 = ~n29243 ;
  assign n29407 = n29054 & n74945 ;
  assign n29055 = n28509 | n29054 ;
  assign n74946 = ~n29055 ;
  assign n29408 = n74946 & n29242 ;
  assign n29409 = n29407 | n29408 ;
  assign n29410 = n133 & n29409 ;
  assign n29411 = n28500 & n74909 ;
  assign n29412 = n29150 & n29411 ;
  assign n29413 = n29410 | n29412 ;
  assign n29414 = n70927 & n29413 ;
  assign n74947 = ~n29049 ;
  assign n29415 = n29048 & n74947 ;
  assign n29416 = n28517 | n29048 ;
  assign n74948 = ~n29416 ;
  assign n29417 = n29240 & n74948 ;
  assign n29418 = n29415 | n29417 ;
  assign n29419 = n133 & n29418 ;
  assign n29420 = n28508 & n74909 ;
  assign n29421 = n29150 & n29420 ;
  assign n29422 = n29419 | n29421 ;
  assign n29423 = n70609 & n29422 ;
  assign n74949 = ~n29239 ;
  assign n29424 = n29043 & n74949 ;
  assign n29044 = n28525 | n29043 ;
  assign n74950 = ~n29044 ;
  assign n29425 = n74950 & n29238 ;
  assign n29426 = n29424 | n29425 ;
  assign n29427 = n133 & n29426 ;
  assign n29428 = n28516 & n74909 ;
  assign n29429 = n29150 & n29428 ;
  assign n29430 = n29427 | n29429 ;
  assign n29431 = n70276 & n29430 ;
  assign n74951 = ~n29038 ;
  assign n29432 = n29037 & n74951 ;
  assign n29433 = n28533 | n29037 ;
  assign n74952 = ~n29433 ;
  assign n29434 = n29236 & n74952 ;
  assign n29435 = n29432 | n29434 ;
  assign n29436 = n133 & n29435 ;
  assign n29437 = n28524 & n74909 ;
  assign n29438 = n29150 & n29437 ;
  assign n29439 = n29436 | n29438 ;
  assign n29440 = n70176 & n29439 ;
  assign n74953 = ~n29235 ;
  assign n29441 = n29032 & n74953 ;
  assign n29033 = n28541 | n29032 ;
  assign n74954 = ~n29033 ;
  assign n29442 = n74954 & n29234 ;
  assign n29443 = n29441 | n29442 ;
  assign n29444 = n133 & n29443 ;
  assign n29445 = n28532 & n74909 ;
  assign n29446 = n29150 & n29445 ;
  assign n29447 = n29444 | n29446 ;
  assign n29448 = n69857 & n29447 ;
  assign n74955 = ~n29027 ;
  assign n29449 = n29026 & n74955 ;
  assign n29450 = n28549 | n29026 ;
  assign n74956 = ~n29450 ;
  assign n29451 = n29232 & n74956 ;
  assign n29452 = n29449 | n29451 ;
  assign n29453 = n133 & n29452 ;
  assign n29454 = n28540 & n74909 ;
  assign n29455 = n29150 & n29454 ;
  assign n29456 = n29453 | n29455 ;
  assign n29457 = n69656 & n29456 ;
  assign n74957 = ~n29231 ;
  assign n29458 = n29022 & n74957 ;
  assign n29459 = n28557 | n29022 ;
  assign n74958 = ~n29459 ;
  assign n29460 = n29018 & n74958 ;
  assign n29461 = n29458 | n29460 ;
  assign n29462 = n133 & n29461 ;
  assign n29463 = n28548 & n74909 ;
  assign n29464 = n29150 & n29463 ;
  assign n29465 = n29462 | n29464 ;
  assign n29466 = n69528 & n29465 ;
  assign n74959 = ~n29017 ;
  assign n29467 = n29016 & n74959 ;
  assign n29468 = n28565 | n29016 ;
  assign n74960 = ~n29468 ;
  assign n29469 = n29228 & n74960 ;
  assign n29470 = n29467 | n29469 ;
  assign n29471 = n133 & n29470 ;
  assign n29472 = n28556 & n74909 ;
  assign n29473 = n29150 & n29472 ;
  assign n29474 = n29471 | n29473 ;
  assign n29475 = n69261 & n29474 ;
  assign n74961 = ~n29227 ;
  assign n29476 = n29012 & n74961 ;
  assign n29477 = n28573 | n29012 ;
  assign n74962 = ~n29477 ;
  assign n29478 = n29008 & n74962 ;
  assign n29479 = n29476 | n29478 ;
  assign n29480 = n133 & n29479 ;
  assign n29481 = n28564 & n74909 ;
  assign n29482 = n29150 & n29481 ;
  assign n29483 = n29480 | n29482 ;
  assign n29484 = n69075 & n29483 ;
  assign n74963 = ~n29007 ;
  assign n29485 = n29006 & n74963 ;
  assign n29486 = n28581 | n29006 ;
  assign n74964 = ~n29486 ;
  assign n29487 = n29224 & n74964 ;
  assign n29488 = n29485 | n29487 ;
  assign n29489 = n133 & n29488 ;
  assign n29490 = n28572 & n74909 ;
  assign n29491 = n29150 & n29490 ;
  assign n29492 = n29489 | n29491 ;
  assign n29493 = n68993 & n29492 ;
  assign n74965 = ~n29223 ;
  assign n29494 = n29002 & n74965 ;
  assign n29495 = n28589 | n29002 ;
  assign n74966 = ~n29495 ;
  assign n29496 = n28998 & n74966 ;
  assign n29497 = n29494 | n29496 ;
  assign n29498 = n133 & n29497 ;
  assign n29499 = n28580 & n74909 ;
  assign n29500 = n29150 & n29499 ;
  assign n29501 = n29498 | n29500 ;
  assign n29502 = n68716 & n29501 ;
  assign n74967 = ~n28997 ;
  assign n29503 = n28996 & n74967 ;
  assign n29504 = n28597 | n28996 ;
  assign n74968 = ~n29504 ;
  assign n29505 = n29220 & n74968 ;
  assign n29506 = n29503 | n29505 ;
  assign n29507 = n133 & n29506 ;
  assign n29508 = n28588 & n74909 ;
  assign n29509 = n29150 & n29508 ;
  assign n29510 = n29507 | n29509 ;
  assign n29511 = n68545 & n29510 ;
  assign n74969 = ~n29219 ;
  assign n29512 = n28991 & n74969 ;
  assign n28992 = n28605 | n28991 ;
  assign n74970 = ~n28992 ;
  assign n29513 = n74970 & n29218 ;
  assign n29514 = n29512 | n29513 ;
  assign n29515 = n133 & n29514 ;
  assign n29516 = n28596 & n74909 ;
  assign n29517 = n29150 & n29516 ;
  assign n29518 = n29515 | n29517 ;
  assign n29519 = n68438 & n29518 ;
  assign n74971 = ~n28986 ;
  assign n29520 = n28985 & n74971 ;
  assign n29521 = n28613 | n28985 ;
  assign n74972 = ~n29521 ;
  assign n29522 = n29216 & n74972 ;
  assign n29523 = n29520 | n29522 ;
  assign n29524 = n133 & n29523 ;
  assign n29525 = n28604 & n74909 ;
  assign n29526 = n29150 & n29525 ;
  assign n29527 = n29524 | n29526 ;
  assign n29528 = n68214 & n29527 ;
  assign n74973 = ~n29215 ;
  assign n29529 = n28981 & n74973 ;
  assign n29530 = n28621 | n28981 ;
  assign n74974 = ~n29530 ;
  assign n29531 = n28977 & n74974 ;
  assign n29532 = n29529 | n29531 ;
  assign n29533 = n133 & n29532 ;
  assign n29534 = n28612 & n74909 ;
  assign n29535 = n29150 & n29534 ;
  assign n29536 = n29533 | n29535 ;
  assign n29537 = n68058 & n29536 ;
  assign n74975 = ~n28976 ;
  assign n29538 = n28975 & n74975 ;
  assign n29539 = n28629 | n28975 ;
  assign n74976 = ~n29539 ;
  assign n29540 = n29212 & n74976 ;
  assign n29541 = n29538 | n29540 ;
  assign n29542 = n133 & n29541 ;
  assign n29543 = n28620 & n74909 ;
  assign n29544 = n29150 & n29543 ;
  assign n29545 = n29542 | n29544 ;
  assign n29546 = n67986 & n29545 ;
  assign n74977 = ~n29211 ;
  assign n29547 = n28971 & n74977 ;
  assign n29548 = n28637 | n28971 ;
  assign n74978 = ~n29548 ;
  assign n29549 = n28967 & n74978 ;
  assign n29550 = n29547 | n29549 ;
  assign n29551 = n133 & n29550 ;
  assign n29552 = n28628 & n74909 ;
  assign n29553 = n29150 & n29552 ;
  assign n29554 = n29551 | n29553 ;
  assign n29555 = n67763 & n29554 ;
  assign n74979 = ~n28966 ;
  assign n29556 = n28965 & n74979 ;
  assign n29557 = n28645 | n28965 ;
  assign n74980 = ~n29557 ;
  assign n29558 = n29208 & n74980 ;
  assign n29559 = n29556 | n29558 ;
  assign n29560 = n133 & n29559 ;
  assign n29561 = n28636 & n74909 ;
  assign n29562 = n29150 & n29561 ;
  assign n29563 = n29560 | n29562 ;
  assign n29564 = n67622 & n29563 ;
  assign n74981 = ~n29207 ;
  assign n29565 = n28961 & n74981 ;
  assign n29566 = n28653 | n28961 ;
  assign n74982 = ~n29566 ;
  assign n29567 = n28957 & n74982 ;
  assign n29568 = n29565 | n29567 ;
  assign n29569 = n133 & n29568 ;
  assign n29570 = n28644 & n74909 ;
  assign n29571 = n29150 & n29570 ;
  assign n29572 = n29569 | n29571 ;
  assign n29573 = n67531 & n29572 ;
  assign n74983 = ~n28956 ;
  assign n29574 = n28955 & n74983 ;
  assign n29575 = n28661 | n28955 ;
  assign n74984 = ~n29575 ;
  assign n29576 = n29204 & n74984 ;
  assign n29577 = n29574 | n29576 ;
  assign n29578 = n133 & n29577 ;
  assign n29579 = n28652 & n74909 ;
  assign n29580 = n29150 & n29579 ;
  assign n29581 = n29578 | n29580 ;
  assign n29582 = n67348 & n29581 ;
  assign n74985 = ~n29203 ;
  assign n29583 = n28951 & n74985 ;
  assign n29584 = n28669 | n28951 ;
  assign n74986 = ~n29584 ;
  assign n29585 = n28947 & n74986 ;
  assign n29586 = n29583 | n29585 ;
  assign n29587 = n133 & n29586 ;
  assign n29588 = n28660 & n74909 ;
  assign n29589 = n29150 & n29588 ;
  assign n29590 = n29587 | n29589 ;
  assign n29591 = n67222 & n29590 ;
  assign n74987 = ~n28946 ;
  assign n29592 = n28945 & n74987 ;
  assign n29593 = n28677 | n28945 ;
  assign n74988 = ~n29593 ;
  assign n29594 = n29200 & n74988 ;
  assign n29595 = n29592 | n29594 ;
  assign n29596 = n133 & n29595 ;
  assign n29597 = n28668 & n74909 ;
  assign n29598 = n29150 & n29597 ;
  assign n29599 = n29596 | n29598 ;
  assign n29600 = n67164 & n29599 ;
  assign n74989 = ~n29199 ;
  assign n29601 = n28941 & n74989 ;
  assign n29602 = n28685 | n28941 ;
  assign n74990 = ~n29602 ;
  assign n29603 = n28937 & n74990 ;
  assign n29604 = n29601 | n29603 ;
  assign n29605 = n133 & n29604 ;
  assign n29606 = n28676 & n74909 ;
  assign n29607 = n29150 & n29606 ;
  assign n29608 = n29605 | n29607 ;
  assign n29609 = n66979 & n29608 ;
  assign n74991 = ~n28936 ;
  assign n29610 = n28935 & n74991 ;
  assign n29611 = n28693 | n28935 ;
  assign n74992 = ~n29611 ;
  assign n29612 = n29196 & n74992 ;
  assign n29613 = n29610 | n29612 ;
  assign n29614 = n133 & n29613 ;
  assign n29615 = n28684 & n74909 ;
  assign n29616 = n29150 & n29615 ;
  assign n29617 = n29614 | n29616 ;
  assign n29618 = n66868 & n29617 ;
  assign n74993 = ~n29195 ;
  assign n29619 = n28931 & n74993 ;
  assign n29620 = n28701 | n28931 ;
  assign n74994 = ~n29620 ;
  assign n29621 = n28927 & n74994 ;
  assign n29622 = n29619 | n29621 ;
  assign n29623 = n133 & n29622 ;
  assign n29624 = n28692 & n74909 ;
  assign n29625 = n29150 & n29624 ;
  assign n29626 = n29623 | n29625 ;
  assign n29627 = n66797 & n29626 ;
  assign n74995 = ~n28926 ;
  assign n29628 = n28925 & n74995 ;
  assign n29629 = n28709 | n28925 ;
  assign n74996 = ~n29629 ;
  assign n29630 = n29192 & n74996 ;
  assign n29631 = n29628 | n29630 ;
  assign n29632 = n133 & n29631 ;
  assign n29633 = n28700 & n74909 ;
  assign n29634 = n29150 & n29633 ;
  assign n29635 = n29632 | n29634 ;
  assign n29636 = n66654 & n29635 ;
  assign n74997 = ~n29191 ;
  assign n29637 = n28921 & n74997 ;
  assign n29638 = n28717 | n28921 ;
  assign n74998 = ~n29638 ;
  assign n29639 = n28917 & n74998 ;
  assign n29640 = n29637 | n29639 ;
  assign n29641 = n133 & n29640 ;
  assign n29642 = n28708 & n74909 ;
  assign n29643 = n29150 & n29642 ;
  assign n29644 = n29641 | n29643 ;
  assign n29645 = n66560 & n29644 ;
  assign n74999 = ~n28916 ;
  assign n29646 = n28915 & n74999 ;
  assign n29647 = n28725 | n28915 ;
  assign n75000 = ~n29647 ;
  assign n29648 = n29188 & n75000 ;
  assign n29649 = n29646 | n29648 ;
  assign n29650 = n133 & n29649 ;
  assign n29651 = n28716 & n74909 ;
  assign n29652 = n29150 & n29651 ;
  assign n29653 = n29650 | n29652 ;
  assign n29654 = n66505 & n29653 ;
  assign n75001 = ~n29187 ;
  assign n29655 = n28911 & n75001 ;
  assign n29656 = n28733 | n28911 ;
  assign n75002 = ~n29656 ;
  assign n29657 = n28907 & n75002 ;
  assign n29658 = n29655 | n29657 ;
  assign n29659 = n133 & n29658 ;
  assign n29660 = n28724 & n74909 ;
  assign n29661 = n29150 & n29660 ;
  assign n29662 = n29659 | n29661 ;
  assign n29663 = n66379 & n29662 ;
  assign n75003 = ~n28906 ;
  assign n29664 = n28905 & n75003 ;
  assign n29665 = n28741 | n28905 ;
  assign n75004 = ~n29665 ;
  assign n29666 = n29184 & n75004 ;
  assign n29667 = n29664 | n29666 ;
  assign n29668 = n133 & n29667 ;
  assign n29669 = n28732 & n74909 ;
  assign n29670 = n29150 & n29669 ;
  assign n29671 = n29668 | n29670 ;
  assign n29672 = n66299 & n29671 ;
  assign n75005 = ~n29183 ;
  assign n29673 = n28901 & n75005 ;
  assign n29674 = n28749 | n28901 ;
  assign n75006 = ~n29674 ;
  assign n29675 = n28897 & n75006 ;
  assign n29676 = n29673 | n29675 ;
  assign n29677 = n133 & n29676 ;
  assign n29678 = n28740 & n74909 ;
  assign n29679 = n29150 & n29678 ;
  assign n29680 = n29677 | n29679 ;
  assign n29681 = n66244 & n29680 ;
  assign n75007 = ~n28896 ;
  assign n29682 = n28895 & n75007 ;
  assign n29683 = n28757 | n28895 ;
  assign n75008 = ~n29683 ;
  assign n29684 = n29180 & n75008 ;
  assign n29685 = n29682 | n29684 ;
  assign n29686 = n133 & n29685 ;
  assign n29687 = n28748 & n74909 ;
  assign n29688 = n29150 & n29687 ;
  assign n29689 = n29686 | n29688 ;
  assign n29690 = n66145 & n29689 ;
  assign n75009 = ~n29179 ;
  assign n29691 = n28891 & n75009 ;
  assign n29692 = n28765 | n28891 ;
  assign n75010 = ~n29692 ;
  assign n29693 = n28887 & n75010 ;
  assign n29694 = n29691 | n29693 ;
  assign n29695 = n133 & n29694 ;
  assign n29696 = n28756 & n74909 ;
  assign n29697 = n29150 & n29696 ;
  assign n29698 = n29695 | n29697 ;
  assign n29699 = n66081 & n29698 ;
  assign n75011 = ~n28886 ;
  assign n29700 = n28885 & n75011 ;
  assign n29701 = n28773 | n28885 ;
  assign n75012 = ~n29701 ;
  assign n29702 = n29176 & n75012 ;
  assign n29703 = n29700 | n29702 ;
  assign n29704 = n133 & n29703 ;
  assign n29705 = n28764 & n74909 ;
  assign n29706 = n29150 & n29705 ;
  assign n29707 = n29704 | n29706 ;
  assign n29708 = n66043 & n29707 ;
  assign n75013 = ~n29175 ;
  assign n29709 = n28881 & n75013 ;
  assign n29710 = n28781 | n28881 ;
  assign n75014 = ~n29710 ;
  assign n29711 = n28877 & n75014 ;
  assign n29712 = n29709 | n29711 ;
  assign n29713 = n133 & n29712 ;
  assign n29714 = n28772 & n74909 ;
  assign n29715 = n29150 & n29714 ;
  assign n29716 = n29713 | n29715 ;
  assign n29717 = n65960 & n29716 ;
  assign n75015 = ~n28876 ;
  assign n29718 = n28875 & n75015 ;
  assign n29719 = n28789 | n28875 ;
  assign n75016 = ~n29719 ;
  assign n29720 = n29172 & n75016 ;
  assign n29721 = n29718 | n29720 ;
  assign n29722 = n133 & n29721 ;
  assign n29723 = n28780 & n74909 ;
  assign n29724 = n29150 & n29723 ;
  assign n29725 = n29722 | n29724 ;
  assign n29726 = n65909 & n29725 ;
  assign n75017 = ~n29171 ;
  assign n29727 = n28871 & n75017 ;
  assign n29728 = n28797 | n28871 ;
  assign n75018 = ~n29728 ;
  assign n29729 = n28867 & n75018 ;
  assign n29730 = n29727 | n29729 ;
  assign n29731 = n133 & n29730 ;
  assign n29732 = n28788 & n74909 ;
  assign n29733 = n29150 & n29732 ;
  assign n29734 = n29731 | n29733 ;
  assign n29735 = n65877 & n29734 ;
  assign n75019 = ~n28866 ;
  assign n29736 = n28865 & n75019 ;
  assign n29737 = n28806 | n28865 ;
  assign n75020 = ~n29737 ;
  assign n29738 = n29168 & n75020 ;
  assign n29739 = n29736 | n29738 ;
  assign n29740 = n133 & n29739 ;
  assign n29741 = n28796 & n74909 ;
  assign n29742 = n29150 & n29741 ;
  assign n29743 = n29740 | n29742 ;
  assign n29744 = n65820 & n29743 ;
  assign n75021 = ~n29167 ;
  assign n29745 = n28860 & n75021 ;
  assign n28861 = n28814 | n28860 ;
  assign n75022 = ~n28861 ;
  assign n29746 = n75022 & n29166 ;
  assign n29747 = n29745 | n29746 ;
  assign n29748 = n133 & n29747 ;
  assign n29749 = n28805 & n74909 ;
  assign n29750 = n29150 & n29749 ;
  assign n29751 = n29748 | n29750 ;
  assign n29752 = n65791 & n29751 ;
  assign n75023 = ~n28855 ;
  assign n29753 = n28854 & n75023 ;
  assign n29754 = n28822 | n28854 ;
  assign n75024 = ~n29754 ;
  assign n29755 = n29164 & n75024 ;
  assign n29756 = n29753 | n29755 ;
  assign n29757 = n133 & n29756 ;
  assign n29758 = n28813 & n74909 ;
  assign n29759 = n29150 & n29758 ;
  assign n29760 = n29757 | n29759 ;
  assign n29761 = n65772 & n29760 ;
  assign n75025 = ~n29163 ;
  assign n29763 = n28850 & n75025 ;
  assign n29762 = n28830 | n28850 ;
  assign n75026 = ~n29762 ;
  assign n29764 = n29162 & n75026 ;
  assign n29765 = n29763 | n29764 ;
  assign n29766 = n133 & n29765 ;
  assign n29767 = n28821 & n74909 ;
  assign n29768 = n29150 & n29767 ;
  assign n29769 = n29766 | n29768 ;
  assign n29770 = n65746 & n29769 ;
  assign n75027 = ~n28845 ;
  assign n29771 = n28844 & n75027 ;
  assign n29161 = n28841 | n28844 ;
  assign n75028 = ~n29161 ;
  assign n29772 = n28840 & n75028 ;
  assign n29773 = n29771 | n29772 ;
  assign n29774 = n133 & n29773 ;
  assign n29775 = n28829 & n74909 ;
  assign n29776 = n29150 & n29775 ;
  assign n29777 = n29774 | n29776 ;
  assign n29778 = n65721 & n29777 ;
  assign n29779 = n28837 & n28839 ;
  assign n29780 = n74787 & n29779 ;
  assign n75029 = ~n29780 ;
  assign n29781 = n28840 & n75029 ;
  assign n29782 = n133 & n29781 ;
  assign n29783 = n28832 & n74909 ;
  assign n29784 = n29150 & n29783 ;
  assign n29785 = n29782 | n29784 ;
  assign n29786 = n65686 & n29785 ;
  assign n29153 = n28839 & n133 ;
  assign n29793 = x64 & n133 ;
  assign n75030 = ~n29793 ;
  assign n29794 = x4 & n75030 ;
  assign n29795 = n29153 | n29794 ;
  assign n29797 = x65 & n29795 ;
  assign n29789 = n29149 | n29788 ;
  assign n29790 = n74909 & n29789 ;
  assign n75031 = ~n29790 ;
  assign n29791 = x64 & n75031 ;
  assign n75032 = ~n29791 ;
  assign n29792 = x4 & n75032 ;
  assign n29796 = x65 | n29153 ;
  assign n29798 = n29792 | n29796 ;
  assign n75033 = ~n29797 ;
  assign n29799 = n75033 & n29798 ;
  assign n75034 = ~x3 ;
  assign n29800 = n75034 & x64 ;
  assign n29801 = n29799 | n29800 ;
  assign n29802 = n65670 & n29795 ;
  assign n75035 = ~n29802 ;
  assign n29803 = n29801 & n75035 ;
  assign n75036 = ~n29784 ;
  assign n29804 = x66 & n75036 ;
  assign n75037 = ~n29782 ;
  assign n29805 = n75037 & n29804 ;
  assign n29806 = n29786 | n29805 ;
  assign n29807 = n29803 | n29806 ;
  assign n75038 = ~n29786 ;
  assign n29808 = n75038 & n29807 ;
  assign n75039 = ~n29776 ;
  assign n29809 = x67 & n75039 ;
  assign n75040 = ~n29774 ;
  assign n29810 = n75040 & n29809 ;
  assign n29811 = n29778 | n29810 ;
  assign n29812 = n29808 | n29811 ;
  assign n75041 = ~n29778 ;
  assign n29813 = n75041 & n29812 ;
  assign n75042 = ~n29768 ;
  assign n29814 = x68 & n75042 ;
  assign n75043 = ~n29766 ;
  assign n29815 = n75043 & n29814 ;
  assign n29816 = n29770 | n29815 ;
  assign n29817 = n29813 | n29816 ;
  assign n75044 = ~n29770 ;
  assign n29818 = n75044 & n29817 ;
  assign n75045 = ~n29759 ;
  assign n29819 = x69 & n75045 ;
  assign n75046 = ~n29757 ;
  assign n29820 = n75046 & n29819 ;
  assign n29821 = n29761 | n29820 ;
  assign n29823 = n29818 | n29821 ;
  assign n75047 = ~n29761 ;
  assign n29824 = n75047 & n29823 ;
  assign n75048 = ~n29750 ;
  assign n29825 = x70 & n75048 ;
  assign n75049 = ~n29748 ;
  assign n29826 = n75049 & n29825 ;
  assign n29827 = n29752 | n29826 ;
  assign n29828 = n29824 | n29827 ;
  assign n75050 = ~n29752 ;
  assign n29829 = n75050 & n29828 ;
  assign n75051 = ~n29742 ;
  assign n29830 = x71 & n75051 ;
  assign n75052 = ~n29740 ;
  assign n29831 = n75052 & n29830 ;
  assign n29832 = n29744 | n29831 ;
  assign n29834 = n29829 | n29832 ;
  assign n75053 = ~n29744 ;
  assign n29835 = n75053 & n29834 ;
  assign n75054 = ~n29733 ;
  assign n29836 = x72 & n75054 ;
  assign n75055 = ~n29731 ;
  assign n29837 = n75055 & n29836 ;
  assign n29838 = n29735 | n29837 ;
  assign n29839 = n29835 | n29838 ;
  assign n75056 = ~n29735 ;
  assign n29840 = n75056 & n29839 ;
  assign n75057 = ~n29724 ;
  assign n29841 = x73 & n75057 ;
  assign n75058 = ~n29722 ;
  assign n29842 = n75058 & n29841 ;
  assign n29843 = n29726 | n29842 ;
  assign n29845 = n29840 | n29843 ;
  assign n75059 = ~n29726 ;
  assign n29846 = n75059 & n29845 ;
  assign n75060 = ~n29715 ;
  assign n29847 = x74 & n75060 ;
  assign n75061 = ~n29713 ;
  assign n29848 = n75061 & n29847 ;
  assign n29849 = n29717 | n29848 ;
  assign n29850 = n29846 | n29849 ;
  assign n75062 = ~n29717 ;
  assign n29851 = n75062 & n29850 ;
  assign n75063 = ~n29706 ;
  assign n29852 = x75 & n75063 ;
  assign n75064 = ~n29704 ;
  assign n29853 = n75064 & n29852 ;
  assign n29854 = n29708 | n29853 ;
  assign n29856 = n29851 | n29854 ;
  assign n75065 = ~n29708 ;
  assign n29857 = n75065 & n29856 ;
  assign n75066 = ~n29697 ;
  assign n29858 = x76 & n75066 ;
  assign n75067 = ~n29695 ;
  assign n29859 = n75067 & n29858 ;
  assign n29860 = n29699 | n29859 ;
  assign n29861 = n29857 | n29860 ;
  assign n75068 = ~n29699 ;
  assign n29862 = n75068 & n29861 ;
  assign n75069 = ~n29688 ;
  assign n29863 = x77 & n75069 ;
  assign n75070 = ~n29686 ;
  assign n29864 = n75070 & n29863 ;
  assign n29865 = n29690 | n29864 ;
  assign n29867 = n29862 | n29865 ;
  assign n75071 = ~n29690 ;
  assign n29868 = n75071 & n29867 ;
  assign n75072 = ~n29679 ;
  assign n29869 = x78 & n75072 ;
  assign n75073 = ~n29677 ;
  assign n29870 = n75073 & n29869 ;
  assign n29871 = n29681 | n29870 ;
  assign n29872 = n29868 | n29871 ;
  assign n75074 = ~n29681 ;
  assign n29873 = n75074 & n29872 ;
  assign n75075 = ~n29670 ;
  assign n29874 = x79 & n75075 ;
  assign n75076 = ~n29668 ;
  assign n29875 = n75076 & n29874 ;
  assign n29876 = n29672 | n29875 ;
  assign n29878 = n29873 | n29876 ;
  assign n75077 = ~n29672 ;
  assign n29879 = n75077 & n29878 ;
  assign n75078 = ~n29661 ;
  assign n29880 = x80 & n75078 ;
  assign n75079 = ~n29659 ;
  assign n29881 = n75079 & n29880 ;
  assign n29882 = n29663 | n29881 ;
  assign n29883 = n29879 | n29882 ;
  assign n75080 = ~n29663 ;
  assign n29884 = n75080 & n29883 ;
  assign n75081 = ~n29652 ;
  assign n29885 = x81 & n75081 ;
  assign n75082 = ~n29650 ;
  assign n29886 = n75082 & n29885 ;
  assign n29887 = n29654 | n29886 ;
  assign n29889 = n29884 | n29887 ;
  assign n75083 = ~n29654 ;
  assign n29890 = n75083 & n29889 ;
  assign n75084 = ~n29643 ;
  assign n29891 = x82 & n75084 ;
  assign n75085 = ~n29641 ;
  assign n29892 = n75085 & n29891 ;
  assign n29893 = n29645 | n29892 ;
  assign n29894 = n29890 | n29893 ;
  assign n75086 = ~n29645 ;
  assign n29895 = n75086 & n29894 ;
  assign n75087 = ~n29634 ;
  assign n29896 = x83 & n75087 ;
  assign n75088 = ~n29632 ;
  assign n29897 = n75088 & n29896 ;
  assign n29898 = n29636 | n29897 ;
  assign n29900 = n29895 | n29898 ;
  assign n75089 = ~n29636 ;
  assign n29901 = n75089 & n29900 ;
  assign n75090 = ~n29625 ;
  assign n29902 = x84 & n75090 ;
  assign n75091 = ~n29623 ;
  assign n29903 = n75091 & n29902 ;
  assign n29904 = n29627 | n29903 ;
  assign n29905 = n29901 | n29904 ;
  assign n75092 = ~n29627 ;
  assign n29906 = n75092 & n29905 ;
  assign n75093 = ~n29616 ;
  assign n29907 = x85 & n75093 ;
  assign n75094 = ~n29614 ;
  assign n29908 = n75094 & n29907 ;
  assign n29909 = n29618 | n29908 ;
  assign n29911 = n29906 | n29909 ;
  assign n75095 = ~n29618 ;
  assign n29912 = n75095 & n29911 ;
  assign n75096 = ~n29607 ;
  assign n29913 = x86 & n75096 ;
  assign n75097 = ~n29605 ;
  assign n29914 = n75097 & n29913 ;
  assign n29915 = n29609 | n29914 ;
  assign n29916 = n29912 | n29915 ;
  assign n75098 = ~n29609 ;
  assign n29917 = n75098 & n29916 ;
  assign n75099 = ~n29598 ;
  assign n29918 = x87 & n75099 ;
  assign n75100 = ~n29596 ;
  assign n29919 = n75100 & n29918 ;
  assign n29920 = n29600 | n29919 ;
  assign n29922 = n29917 | n29920 ;
  assign n75101 = ~n29600 ;
  assign n29923 = n75101 & n29922 ;
  assign n75102 = ~n29589 ;
  assign n29924 = x88 & n75102 ;
  assign n75103 = ~n29587 ;
  assign n29925 = n75103 & n29924 ;
  assign n29926 = n29591 | n29925 ;
  assign n29927 = n29923 | n29926 ;
  assign n75104 = ~n29591 ;
  assign n29928 = n75104 & n29927 ;
  assign n75105 = ~n29580 ;
  assign n29929 = x89 & n75105 ;
  assign n75106 = ~n29578 ;
  assign n29930 = n75106 & n29929 ;
  assign n29931 = n29582 | n29930 ;
  assign n29933 = n29928 | n29931 ;
  assign n75107 = ~n29582 ;
  assign n29934 = n75107 & n29933 ;
  assign n75108 = ~n29571 ;
  assign n29935 = x90 & n75108 ;
  assign n75109 = ~n29569 ;
  assign n29936 = n75109 & n29935 ;
  assign n29937 = n29573 | n29936 ;
  assign n29938 = n29934 | n29937 ;
  assign n75110 = ~n29573 ;
  assign n29939 = n75110 & n29938 ;
  assign n75111 = ~n29562 ;
  assign n29940 = x91 & n75111 ;
  assign n75112 = ~n29560 ;
  assign n29941 = n75112 & n29940 ;
  assign n29942 = n29564 | n29941 ;
  assign n29944 = n29939 | n29942 ;
  assign n75113 = ~n29564 ;
  assign n29945 = n75113 & n29944 ;
  assign n75114 = ~n29553 ;
  assign n29946 = x92 & n75114 ;
  assign n75115 = ~n29551 ;
  assign n29947 = n75115 & n29946 ;
  assign n29948 = n29555 | n29947 ;
  assign n29949 = n29945 | n29948 ;
  assign n75116 = ~n29555 ;
  assign n29950 = n75116 & n29949 ;
  assign n75117 = ~n29544 ;
  assign n29951 = x93 & n75117 ;
  assign n75118 = ~n29542 ;
  assign n29952 = n75118 & n29951 ;
  assign n29953 = n29546 | n29952 ;
  assign n29955 = n29950 | n29953 ;
  assign n75119 = ~n29546 ;
  assign n29956 = n75119 & n29955 ;
  assign n75120 = ~n29535 ;
  assign n29957 = x94 & n75120 ;
  assign n75121 = ~n29533 ;
  assign n29958 = n75121 & n29957 ;
  assign n29959 = n29537 | n29958 ;
  assign n29960 = n29956 | n29959 ;
  assign n75122 = ~n29537 ;
  assign n29961 = n75122 & n29960 ;
  assign n75123 = ~n29526 ;
  assign n29962 = x95 & n75123 ;
  assign n75124 = ~n29524 ;
  assign n29963 = n75124 & n29962 ;
  assign n29964 = n29528 | n29963 ;
  assign n29966 = n29961 | n29964 ;
  assign n75125 = ~n29528 ;
  assign n29967 = n75125 & n29966 ;
  assign n75126 = ~n29517 ;
  assign n29968 = x96 & n75126 ;
  assign n75127 = ~n29515 ;
  assign n29969 = n75127 & n29968 ;
  assign n29970 = n29519 | n29969 ;
  assign n29971 = n29967 | n29970 ;
  assign n75128 = ~n29519 ;
  assign n29972 = n75128 & n29971 ;
  assign n75129 = ~n29509 ;
  assign n29973 = x97 & n75129 ;
  assign n75130 = ~n29507 ;
  assign n29974 = n75130 & n29973 ;
  assign n29975 = n29511 | n29974 ;
  assign n29977 = n29972 | n29975 ;
  assign n75131 = ~n29511 ;
  assign n29978 = n75131 & n29977 ;
  assign n75132 = ~n29500 ;
  assign n29979 = x98 & n75132 ;
  assign n75133 = ~n29498 ;
  assign n29980 = n75133 & n29979 ;
  assign n29981 = n29502 | n29980 ;
  assign n29982 = n29978 | n29981 ;
  assign n75134 = ~n29502 ;
  assign n29983 = n75134 & n29982 ;
  assign n75135 = ~n29491 ;
  assign n29984 = x99 & n75135 ;
  assign n75136 = ~n29489 ;
  assign n29985 = n75136 & n29984 ;
  assign n29986 = n29493 | n29985 ;
  assign n29988 = n29983 | n29986 ;
  assign n75137 = ~n29493 ;
  assign n29989 = n75137 & n29988 ;
  assign n75138 = ~n29482 ;
  assign n29990 = x100 & n75138 ;
  assign n75139 = ~n29480 ;
  assign n29991 = n75139 & n29990 ;
  assign n29992 = n29484 | n29991 ;
  assign n29993 = n29989 | n29992 ;
  assign n75140 = ~n29484 ;
  assign n29994 = n75140 & n29993 ;
  assign n75141 = ~n29473 ;
  assign n29995 = x101 & n75141 ;
  assign n75142 = ~n29471 ;
  assign n29996 = n75142 & n29995 ;
  assign n29997 = n29475 | n29996 ;
  assign n29999 = n29994 | n29997 ;
  assign n75143 = ~n29475 ;
  assign n30000 = n75143 & n29999 ;
  assign n75144 = ~n29464 ;
  assign n30001 = x102 & n75144 ;
  assign n75145 = ~n29462 ;
  assign n30002 = n75145 & n30001 ;
  assign n30003 = n29466 | n30002 ;
  assign n30004 = n30000 | n30003 ;
  assign n75146 = ~n29466 ;
  assign n30005 = n75146 & n30004 ;
  assign n75147 = ~n29455 ;
  assign n30006 = x103 & n75147 ;
  assign n75148 = ~n29453 ;
  assign n30007 = n75148 & n30006 ;
  assign n30008 = n29457 | n30007 ;
  assign n30010 = n30005 | n30008 ;
  assign n75149 = ~n29457 ;
  assign n30011 = n75149 & n30010 ;
  assign n75150 = ~n29446 ;
  assign n30012 = x104 & n75150 ;
  assign n75151 = ~n29444 ;
  assign n30013 = n75151 & n30012 ;
  assign n30014 = n29448 | n30013 ;
  assign n30015 = n30011 | n30014 ;
  assign n75152 = ~n29448 ;
  assign n30016 = n75152 & n30015 ;
  assign n75153 = ~n29438 ;
  assign n30017 = x105 & n75153 ;
  assign n75154 = ~n29436 ;
  assign n30018 = n75154 & n30017 ;
  assign n30019 = n29440 | n30018 ;
  assign n30021 = n30016 | n30019 ;
  assign n75155 = ~n29440 ;
  assign n30022 = n75155 & n30021 ;
  assign n75156 = ~n29429 ;
  assign n30023 = x106 & n75156 ;
  assign n75157 = ~n29427 ;
  assign n30024 = n75157 & n30023 ;
  assign n30025 = n29431 | n30024 ;
  assign n30026 = n30022 | n30025 ;
  assign n75158 = ~n29431 ;
  assign n30027 = n75158 & n30026 ;
  assign n75159 = ~n29421 ;
  assign n30028 = x107 & n75159 ;
  assign n75160 = ~n29419 ;
  assign n30029 = n75160 & n30028 ;
  assign n30030 = n29423 | n30029 ;
  assign n30032 = n30027 | n30030 ;
  assign n75161 = ~n29423 ;
  assign n30033 = n75161 & n30032 ;
  assign n75162 = ~n29412 ;
  assign n30034 = x108 & n75162 ;
  assign n75163 = ~n29410 ;
  assign n30035 = n75163 & n30034 ;
  assign n30036 = n29414 | n30035 ;
  assign n30037 = n30033 | n30036 ;
  assign n75164 = ~n29414 ;
  assign n30038 = n75164 & n30037 ;
  assign n75165 = ~n29404 ;
  assign n30039 = x109 & n75165 ;
  assign n75166 = ~n29402 ;
  assign n30040 = n75166 & n30039 ;
  assign n30041 = n29406 | n30040 ;
  assign n30043 = n30038 | n30041 ;
  assign n75167 = ~n29406 ;
  assign n30044 = n75167 & n30043 ;
  assign n75168 = ~n29396 ;
  assign n30045 = x110 & n75168 ;
  assign n75169 = ~n29394 ;
  assign n30046 = n75169 & n30045 ;
  assign n30047 = n29398 | n30046 ;
  assign n30048 = n30044 | n30047 ;
  assign n75170 = ~n29398 ;
  assign n30049 = n75170 & n30048 ;
  assign n75171 = ~n29387 ;
  assign n30050 = x111 & n75171 ;
  assign n75172 = ~n29385 ;
  assign n30051 = n75172 & n30050 ;
  assign n30052 = n29389 | n30051 ;
  assign n30054 = n30049 | n30052 ;
  assign n75173 = ~n29389 ;
  assign n30055 = n75173 & n30054 ;
  assign n75174 = ~n29378 ;
  assign n30056 = x112 & n75174 ;
  assign n75175 = ~n29376 ;
  assign n30057 = n75175 & n30056 ;
  assign n30058 = n29380 | n30057 ;
  assign n30059 = n30055 | n30058 ;
  assign n75176 = ~n29380 ;
  assign n30060 = n75176 & n30059 ;
  assign n75177 = ~n29369 ;
  assign n30061 = x113 & n75177 ;
  assign n75178 = ~n29367 ;
  assign n30062 = n75178 & n30061 ;
  assign n30063 = n29371 | n30062 ;
  assign n30065 = n30060 | n30063 ;
  assign n75179 = ~n29371 ;
  assign n30066 = n75179 & n30065 ;
  assign n75180 = ~n29360 ;
  assign n30067 = x114 & n75180 ;
  assign n75181 = ~n29358 ;
  assign n30068 = n75181 & n30067 ;
  assign n30069 = n29362 | n30068 ;
  assign n30070 = n30066 | n30069 ;
  assign n75182 = ~n29362 ;
  assign n30071 = n75182 & n30070 ;
  assign n75183 = ~n29351 ;
  assign n30072 = x115 & n75183 ;
  assign n75184 = ~n29349 ;
  assign n30073 = n75184 & n30072 ;
  assign n30074 = n29353 | n30073 ;
  assign n30076 = n30071 | n30074 ;
  assign n75185 = ~n29353 ;
  assign n30077 = n75185 & n30076 ;
  assign n75186 = ~n29342 ;
  assign n30078 = x116 & n75186 ;
  assign n75187 = ~n29340 ;
  assign n30079 = n75187 & n30078 ;
  assign n30080 = n29344 | n30079 ;
  assign n30081 = n30077 | n30080 ;
  assign n75188 = ~n29344 ;
  assign n30082 = n75188 & n30081 ;
  assign n75189 = ~n29333 ;
  assign n30083 = x117 & n75189 ;
  assign n75190 = ~n29331 ;
  assign n30084 = n75190 & n30083 ;
  assign n30085 = n29335 | n30084 ;
  assign n30087 = n30082 | n30085 ;
  assign n75191 = ~n29335 ;
  assign n30088 = n75191 & n30087 ;
  assign n75192 = ~n29325 ;
  assign n30089 = x118 & n75192 ;
  assign n75193 = ~n29323 ;
  assign n30090 = n75193 & n30089 ;
  assign n30091 = n29327 | n30090 ;
  assign n30092 = n30088 | n30091 ;
  assign n75194 = ~n29327 ;
  assign n30093 = n75194 & n30092 ;
  assign n75195 = ~n29316 ;
  assign n30094 = x119 & n75195 ;
  assign n75196 = ~n29314 ;
  assign n30095 = n75196 & n30094 ;
  assign n30096 = n29318 | n30095 ;
  assign n30098 = n30093 | n30096 ;
  assign n75197 = ~n29318 ;
  assign n30099 = n75197 & n30098 ;
  assign n75198 = ~n29307 ;
  assign n30100 = x120 & n75198 ;
  assign n75199 = ~n29305 ;
  assign n30101 = n75199 & n30100 ;
  assign n30102 = n29309 | n30101 ;
  assign n30103 = n30099 | n30102 ;
  assign n75200 = ~n29309 ;
  assign n30104 = n75200 & n30103 ;
  assign n75201 = ~n29298 ;
  assign n30105 = x121 & n75201 ;
  assign n75202 = ~n29296 ;
  assign n30106 = n75202 & n30105 ;
  assign n30107 = n29300 | n30106 ;
  assign n30109 = n30104 | n30107 ;
  assign n75203 = ~n29300 ;
  assign n30110 = n75203 & n30109 ;
  assign n75204 = ~n29289 ;
  assign n30111 = x122 & n75204 ;
  assign n75205 = ~n29287 ;
  assign n30112 = n75205 & n30111 ;
  assign n30113 = n29291 | n30112 ;
  assign n30114 = n30110 | n30113 ;
  assign n75206 = ~n29291 ;
  assign n30115 = n75206 & n30114 ;
  assign n75207 = ~n29280 ;
  assign n30116 = x123 & n75207 ;
  assign n75208 = ~n29278 ;
  assign n30117 = n75208 & n30116 ;
  assign n30118 = n29282 | n30117 ;
  assign n30120 = n30115 | n30118 ;
  assign n75209 = ~n29282 ;
  assign n30121 = n75209 & n30120 ;
  assign n75210 = ~x124 ;
  assign n30132 = n75210 & n30131 ;
  assign n75211 = ~n30130 ;
  assign n30133 = x124 & n75211 ;
  assign n75212 = ~n30128 ;
  assign n30134 = n75212 & n30133 ;
  assign n30135 = n274 | n30134 ;
  assign n30136 = n30132 | n30135 ;
  assign n30138 = n30121 | n30136 ;
  assign n75213 = ~n30137 ;
  assign n30139 = n75213 & n30138 ;
  assign n75214 = ~n30115 ;
  assign n30119 = n75214 & n30118 ;
  assign n30142 = n29153 | n29792 ;
  assign n30143 = x65 & n30142 ;
  assign n75215 = ~n30143 ;
  assign n30144 = n29798 & n75215 ;
  assign n30145 = n29800 | n30144 ;
  assign n30146 = n75035 & n30145 ;
  assign n30147 = n29806 | n30146 ;
  assign n30148 = n75038 & n30147 ;
  assign n30150 = n29811 | n30148 ;
  assign n30151 = n75041 & n30150 ;
  assign n30153 = n29816 | n30151 ;
  assign n30154 = n75044 & n30153 ;
  assign n30155 = n29821 | n30154 ;
  assign n30156 = n75047 & n30155 ;
  assign n30157 = n29827 | n30156 ;
  assign n30159 = n75050 & n30157 ;
  assign n30160 = n29832 | n30159 ;
  assign n30161 = n75053 & n30160 ;
  assign n30162 = n29838 | n30161 ;
  assign n30164 = n75056 & n30162 ;
  assign n30165 = n29843 | n30164 ;
  assign n30166 = n75059 & n30165 ;
  assign n30167 = n29849 | n30166 ;
  assign n30169 = n75062 & n30167 ;
  assign n30170 = n29854 | n30169 ;
  assign n30171 = n75065 & n30170 ;
  assign n30172 = n29860 | n30171 ;
  assign n30174 = n75068 & n30172 ;
  assign n30175 = n29865 | n30174 ;
  assign n30176 = n75071 & n30175 ;
  assign n30177 = n29871 | n30176 ;
  assign n30179 = n75074 & n30177 ;
  assign n30180 = n29876 | n30179 ;
  assign n30181 = n75077 & n30180 ;
  assign n30182 = n29882 | n30181 ;
  assign n30184 = n75080 & n30182 ;
  assign n30185 = n29887 | n30184 ;
  assign n30186 = n75083 & n30185 ;
  assign n30187 = n29893 | n30186 ;
  assign n30189 = n75086 & n30187 ;
  assign n30190 = n29898 | n30189 ;
  assign n30191 = n75089 & n30190 ;
  assign n30192 = n29904 | n30191 ;
  assign n30194 = n75092 & n30192 ;
  assign n30195 = n29909 | n30194 ;
  assign n30196 = n75095 & n30195 ;
  assign n30197 = n29915 | n30196 ;
  assign n30199 = n75098 & n30197 ;
  assign n30200 = n29920 | n30199 ;
  assign n30201 = n75101 & n30200 ;
  assign n30202 = n29926 | n30201 ;
  assign n30204 = n75104 & n30202 ;
  assign n30205 = n29931 | n30204 ;
  assign n30206 = n75107 & n30205 ;
  assign n30207 = n29937 | n30206 ;
  assign n30209 = n75110 & n30207 ;
  assign n30210 = n29942 | n30209 ;
  assign n30211 = n75113 & n30210 ;
  assign n30212 = n29948 | n30211 ;
  assign n30214 = n75116 & n30212 ;
  assign n30215 = n29953 | n30214 ;
  assign n30216 = n75119 & n30215 ;
  assign n30217 = n29959 | n30216 ;
  assign n30219 = n75122 & n30217 ;
  assign n30220 = n29964 | n30219 ;
  assign n30221 = n75125 & n30220 ;
  assign n30222 = n29970 | n30221 ;
  assign n30224 = n75128 & n30222 ;
  assign n30225 = n29975 | n30224 ;
  assign n30226 = n75131 & n30225 ;
  assign n30227 = n29981 | n30226 ;
  assign n30229 = n75134 & n30227 ;
  assign n30230 = n29986 | n30229 ;
  assign n30231 = n75137 & n30230 ;
  assign n30232 = n29992 | n30231 ;
  assign n30234 = n75140 & n30232 ;
  assign n30235 = n29997 | n30234 ;
  assign n30236 = n75143 & n30235 ;
  assign n30237 = n30003 | n30236 ;
  assign n30239 = n75146 & n30237 ;
  assign n30240 = n30008 | n30239 ;
  assign n30241 = n75149 & n30240 ;
  assign n30242 = n30014 | n30241 ;
  assign n30244 = n75152 & n30242 ;
  assign n30245 = n30019 | n30244 ;
  assign n30246 = n75155 & n30245 ;
  assign n30247 = n30025 | n30246 ;
  assign n30249 = n75158 & n30247 ;
  assign n30250 = n30030 | n30249 ;
  assign n30251 = n75161 & n30250 ;
  assign n30252 = n30036 | n30251 ;
  assign n30254 = n75164 & n30252 ;
  assign n30255 = n30041 | n30254 ;
  assign n30256 = n75167 & n30255 ;
  assign n30257 = n30047 | n30256 ;
  assign n30259 = n75170 & n30257 ;
  assign n30260 = n30052 | n30259 ;
  assign n30261 = n75173 & n30260 ;
  assign n30262 = n30058 | n30261 ;
  assign n30264 = n75176 & n30262 ;
  assign n30265 = n30063 | n30264 ;
  assign n30266 = n75179 & n30265 ;
  assign n30267 = n30069 | n30266 ;
  assign n30269 = n75182 & n30267 ;
  assign n30270 = n30074 | n30269 ;
  assign n30271 = n75185 & n30270 ;
  assign n30272 = n30080 | n30271 ;
  assign n30274 = n75188 & n30272 ;
  assign n30275 = n30085 | n30274 ;
  assign n30276 = n75191 & n30275 ;
  assign n30277 = n30091 | n30276 ;
  assign n30279 = n75194 & n30277 ;
  assign n30280 = n30096 | n30279 ;
  assign n30281 = n75197 & n30280 ;
  assign n30282 = n30102 | n30281 ;
  assign n30284 = n75200 & n30282 ;
  assign n30285 = n30107 | n30284 ;
  assign n30286 = n75203 & n30285 ;
  assign n30287 = n30113 | n30286 ;
  assign n30289 = n29291 | n30118 ;
  assign n75216 = ~n30289 ;
  assign n30290 = n30287 & n75216 ;
  assign n30291 = n30119 | n30290 ;
  assign n132 = ~n30139 ;
  assign n30292 = n132 & n30291 ;
  assign n30293 = n75206 & n30287 ;
  assign n30294 = n30118 | n30293 ;
  assign n30295 = n75209 & n30294 ;
  assign n30296 = n30136 | n30295 ;
  assign n30297 = n29281 & n75213 ;
  assign n30298 = n30296 & n30297 ;
  assign n30299 = n30292 | n30298 ;
  assign n30300 = n75210 & n30299 ;
  assign n75218 = ~n30298 ;
  assign n31071 = x124 & n75218 ;
  assign n75219 = ~n30292 ;
  assign n31072 = n75219 & n31071 ;
  assign n31073 = n30300 | n31072 ;
  assign n75220 = ~n30286 ;
  assign n30288 = n30113 & n75220 ;
  assign n30301 = n29300 | n30113 ;
  assign n75221 = ~n30301 ;
  assign n30302 = n30109 & n75221 ;
  assign n30303 = n30288 | n30302 ;
  assign n30304 = n132 & n30303 ;
  assign n30305 = n29290 & n75213 ;
  assign n30306 = n30296 & n30305 ;
  assign n30307 = n30304 | n30306 ;
  assign n30308 = n74905 & n30307 ;
  assign n75222 = ~n30104 ;
  assign n30108 = n75222 & n30107 ;
  assign n30309 = n29309 | n30107 ;
  assign n75223 = ~n30309 ;
  assign n30310 = n30282 & n75223 ;
  assign n30311 = n30108 | n30310 ;
  assign n30312 = n132 & n30311 ;
  assign n30313 = n29299 & n75213 ;
  assign n30314 = n30296 & n30313 ;
  assign n30315 = n30312 | n30314 ;
  assign n30316 = n74431 & n30315 ;
  assign n75224 = ~n30314 ;
  assign n31061 = x122 & n75224 ;
  assign n75225 = ~n30312 ;
  assign n31062 = n75225 & n31061 ;
  assign n31063 = n30316 | n31062 ;
  assign n75226 = ~n30281 ;
  assign n30283 = n30102 & n75226 ;
  assign n30317 = n29318 | n30102 ;
  assign n75227 = ~n30317 ;
  assign n30318 = n30098 & n75227 ;
  assign n30319 = n30283 | n30318 ;
  assign n30320 = n132 & n30319 ;
  assign n30321 = n29308 & n75213 ;
  assign n30322 = n30296 & n30321 ;
  assign n30323 = n30320 | n30322 ;
  assign n30324 = n74029 & n30323 ;
  assign n75228 = ~n30093 ;
  assign n30097 = n75228 & n30096 ;
  assign n30325 = n29327 | n30096 ;
  assign n75229 = ~n30325 ;
  assign n30326 = n30277 & n75229 ;
  assign n30327 = n30097 | n30326 ;
  assign n30328 = n132 & n30327 ;
  assign n30329 = n29317 & n75213 ;
  assign n30330 = n30296 & n30329 ;
  assign n30331 = n30328 | n30330 ;
  assign n30332 = n74021 & n30331 ;
  assign n75230 = ~n30330 ;
  assign n31050 = x120 & n75230 ;
  assign n75231 = ~n30328 ;
  assign n31051 = n75231 & n31050 ;
  assign n31052 = n30332 | n31051 ;
  assign n75232 = ~n30276 ;
  assign n30278 = n30091 & n75232 ;
  assign n30333 = n29335 | n30091 ;
  assign n75233 = ~n30333 ;
  assign n30334 = n30087 & n75233 ;
  assign n30335 = n30278 | n30334 ;
  assign n30336 = n132 & n30335 ;
  assign n30337 = n29326 & n75213 ;
  assign n30338 = n30296 & n30337 ;
  assign n30339 = n30336 | n30338 ;
  assign n30340 = n73617 & n30339 ;
  assign n75234 = ~n30082 ;
  assign n30086 = n75234 & n30085 ;
  assign n30341 = n29344 | n30085 ;
  assign n75235 = ~n30341 ;
  assign n30342 = n30272 & n75235 ;
  assign n30343 = n30086 | n30342 ;
  assign n30344 = n132 & n30343 ;
  assign n30345 = n29334 & n75213 ;
  assign n30346 = n30296 & n30345 ;
  assign n30347 = n30344 | n30346 ;
  assign n30348 = n73188 & n30347 ;
  assign n75236 = ~n30346 ;
  assign n31040 = x118 & n75236 ;
  assign n75237 = ~n30344 ;
  assign n31041 = n75237 & n31040 ;
  assign n31042 = n30348 | n31041 ;
  assign n75238 = ~n30271 ;
  assign n30273 = n30080 & n75238 ;
  assign n30349 = n29353 | n30080 ;
  assign n75239 = ~n30349 ;
  assign n30350 = n30076 & n75239 ;
  assign n30351 = n30273 | n30350 ;
  assign n30352 = n132 & n30351 ;
  assign n30353 = n29343 & n75213 ;
  assign n30354 = n30296 & n30353 ;
  assign n30355 = n30352 | n30354 ;
  assign n30356 = n73177 & n30355 ;
  assign n75240 = ~n30071 ;
  assign n30075 = n75240 & n30074 ;
  assign n30357 = n29362 | n30074 ;
  assign n75241 = ~n30357 ;
  assign n30358 = n30267 & n75241 ;
  assign n30359 = n30075 | n30358 ;
  assign n30360 = n132 & n30359 ;
  assign n30361 = n29352 & n75213 ;
  assign n30362 = n30296 & n30361 ;
  assign n30363 = n30360 | n30362 ;
  assign n30364 = n72752 & n30363 ;
  assign n75242 = ~n30362 ;
  assign n31030 = x116 & n75242 ;
  assign n75243 = ~n30360 ;
  assign n31031 = n75243 & n31030 ;
  assign n31032 = n30364 | n31031 ;
  assign n75244 = ~n30266 ;
  assign n30268 = n30069 & n75244 ;
  assign n30365 = n29371 | n30069 ;
  assign n75245 = ~n30365 ;
  assign n30366 = n30065 & n75245 ;
  assign n30367 = n30268 | n30366 ;
  assign n30368 = n132 & n30367 ;
  assign n30369 = n29361 & n75213 ;
  assign n30370 = n30296 & n30369 ;
  assign n30371 = n30368 | n30370 ;
  assign n30372 = n72393 & n30371 ;
  assign n75246 = ~n30060 ;
  assign n30064 = n75246 & n30063 ;
  assign n30373 = n29380 | n30063 ;
  assign n75247 = ~n30373 ;
  assign n30374 = n30262 & n75247 ;
  assign n30375 = n30064 | n30374 ;
  assign n30376 = n132 & n30375 ;
  assign n30377 = n29370 & n75213 ;
  assign n30378 = n30296 & n30377 ;
  assign n30379 = n30376 | n30378 ;
  assign n30380 = n72385 & n30379 ;
  assign n75248 = ~n30378 ;
  assign n31020 = x114 & n75248 ;
  assign n75249 = ~n30376 ;
  assign n31021 = n75249 & n31020 ;
  assign n31022 = n30380 | n31021 ;
  assign n75250 = ~n30261 ;
  assign n30263 = n30058 & n75250 ;
  assign n30381 = n29389 | n30058 ;
  assign n75251 = ~n30381 ;
  assign n30382 = n30054 & n75251 ;
  assign n30383 = n30263 | n30382 ;
  assign n30384 = n132 & n30383 ;
  assign n30385 = n29379 & n75213 ;
  assign n30386 = n30296 & n30385 ;
  assign n30387 = n30384 | n30386 ;
  assign n30388 = n72025 & n30387 ;
  assign n75252 = ~n30049 ;
  assign n30053 = n75252 & n30052 ;
  assign n30389 = n29398 | n30052 ;
  assign n75253 = ~n30389 ;
  assign n30390 = n30257 & n75253 ;
  assign n30391 = n30053 | n30390 ;
  assign n30392 = n132 & n30391 ;
  assign n30393 = n29388 & n75213 ;
  assign n30394 = n30296 & n30393 ;
  assign n30395 = n30392 | n30394 ;
  assign n30396 = n71645 & n30395 ;
  assign n75254 = ~n30394 ;
  assign n31009 = x112 & n75254 ;
  assign n75255 = ~n30392 ;
  assign n31010 = n75255 & n31009 ;
  assign n31011 = n30396 | n31010 ;
  assign n75256 = ~n30256 ;
  assign n30258 = n30047 & n75256 ;
  assign n30397 = n29406 | n30047 ;
  assign n75257 = ~n30397 ;
  assign n30398 = n30043 & n75257 ;
  assign n30399 = n30258 | n30398 ;
  assign n30400 = n132 & n30399 ;
  assign n30401 = n29397 & n75213 ;
  assign n30402 = n30296 & n30401 ;
  assign n30403 = n30400 | n30402 ;
  assign n30404 = n71633 & n30403 ;
  assign n75258 = ~n30038 ;
  assign n30042 = n75258 & n30041 ;
  assign n30405 = n29414 | n30041 ;
  assign n75259 = ~n30405 ;
  assign n30406 = n30252 & n75259 ;
  assign n30407 = n30042 | n30406 ;
  assign n30408 = n132 & n30407 ;
  assign n30409 = n29405 & n75213 ;
  assign n30410 = n30296 & n30409 ;
  assign n30411 = n30408 | n30410 ;
  assign n30412 = n71253 & n30411 ;
  assign n75260 = ~n30410 ;
  assign n30998 = x110 & n75260 ;
  assign n75261 = ~n30408 ;
  assign n30999 = n75261 & n30998 ;
  assign n31000 = n30412 | n30999 ;
  assign n75262 = ~n30251 ;
  assign n30253 = n30036 & n75262 ;
  assign n30413 = n29423 | n30036 ;
  assign n75263 = ~n30413 ;
  assign n30414 = n30032 & n75263 ;
  assign n30415 = n30253 | n30414 ;
  assign n30416 = n132 & n30415 ;
  assign n30417 = n29413 & n75213 ;
  assign n30418 = n30296 & n30417 ;
  assign n30419 = n30416 | n30418 ;
  assign n30420 = n70935 & n30419 ;
  assign n75264 = ~n30027 ;
  assign n30031 = n75264 & n30030 ;
  assign n30421 = n29431 | n30030 ;
  assign n75265 = ~n30421 ;
  assign n30422 = n30247 & n75265 ;
  assign n30423 = n30031 | n30422 ;
  assign n30424 = n132 & n30423 ;
  assign n30425 = n29422 & n75213 ;
  assign n30426 = n30296 & n30425 ;
  assign n30427 = n30424 | n30426 ;
  assign n30428 = n70927 & n30427 ;
  assign n75266 = ~n30426 ;
  assign n30988 = x108 & n75266 ;
  assign n75267 = ~n30424 ;
  assign n30989 = n75267 & n30988 ;
  assign n30990 = n30428 | n30989 ;
  assign n75268 = ~n30246 ;
  assign n30248 = n30025 & n75268 ;
  assign n30429 = n29440 | n30025 ;
  assign n75269 = ~n30429 ;
  assign n30430 = n30021 & n75269 ;
  assign n30431 = n30248 | n30430 ;
  assign n30432 = n132 & n30431 ;
  assign n30433 = n29430 & n75213 ;
  assign n30434 = n30296 & n30433 ;
  assign n30435 = n30432 | n30434 ;
  assign n30436 = n70609 & n30435 ;
  assign n75270 = ~n30016 ;
  assign n30020 = n75270 & n30019 ;
  assign n30437 = n29448 | n30019 ;
  assign n75271 = ~n30437 ;
  assign n30438 = n30242 & n75271 ;
  assign n30439 = n30020 | n30438 ;
  assign n30440 = n132 & n30439 ;
  assign n30441 = n29439 & n75213 ;
  assign n30442 = n30296 & n30441 ;
  assign n30443 = n30440 | n30442 ;
  assign n30444 = n70276 & n30443 ;
  assign n75272 = ~n30442 ;
  assign n30978 = x106 & n75272 ;
  assign n75273 = ~n30440 ;
  assign n30979 = n75273 & n30978 ;
  assign n30980 = n30444 | n30979 ;
  assign n75274 = ~n30241 ;
  assign n30243 = n30014 & n75274 ;
  assign n30445 = n29457 | n30014 ;
  assign n75275 = ~n30445 ;
  assign n30446 = n30010 & n75275 ;
  assign n30447 = n30243 | n30446 ;
  assign n30448 = n132 & n30447 ;
  assign n30449 = n29447 & n75213 ;
  assign n30450 = n30296 & n30449 ;
  assign n30451 = n30448 | n30450 ;
  assign n30452 = n70176 & n30451 ;
  assign n75276 = ~n30005 ;
  assign n30009 = n75276 & n30008 ;
  assign n30453 = n29466 | n30008 ;
  assign n75277 = ~n30453 ;
  assign n30454 = n30237 & n75277 ;
  assign n30455 = n30009 | n30454 ;
  assign n30456 = n132 & n30455 ;
  assign n30457 = n29456 & n75213 ;
  assign n30458 = n30296 & n30457 ;
  assign n30459 = n30456 | n30458 ;
  assign n30460 = n69857 & n30459 ;
  assign n75278 = ~n30458 ;
  assign n30968 = x104 & n75278 ;
  assign n75279 = ~n30456 ;
  assign n30969 = n75279 & n30968 ;
  assign n30970 = n30460 | n30969 ;
  assign n75280 = ~n30236 ;
  assign n30238 = n30003 & n75280 ;
  assign n30461 = n29475 | n30003 ;
  assign n75281 = ~n30461 ;
  assign n30462 = n29999 & n75281 ;
  assign n30463 = n30238 | n30462 ;
  assign n30464 = n132 & n30463 ;
  assign n30465 = n29465 & n75213 ;
  assign n30466 = n30296 & n30465 ;
  assign n30467 = n30464 | n30466 ;
  assign n30468 = n69656 & n30467 ;
  assign n75282 = ~n29994 ;
  assign n29998 = n75282 & n29997 ;
  assign n30469 = n29484 | n29997 ;
  assign n75283 = ~n30469 ;
  assign n30470 = n30232 & n75283 ;
  assign n30471 = n29998 | n30470 ;
  assign n30472 = n132 & n30471 ;
  assign n30473 = n29474 & n75213 ;
  assign n30474 = n30296 & n30473 ;
  assign n30475 = n30472 | n30474 ;
  assign n30476 = n69528 & n30475 ;
  assign n75284 = ~n30474 ;
  assign n30958 = x102 & n75284 ;
  assign n75285 = ~n30472 ;
  assign n30959 = n75285 & n30958 ;
  assign n30960 = n30476 | n30959 ;
  assign n75286 = ~n30231 ;
  assign n30233 = n29992 & n75286 ;
  assign n30477 = n29493 | n29992 ;
  assign n75287 = ~n30477 ;
  assign n30478 = n29988 & n75287 ;
  assign n30479 = n30233 | n30478 ;
  assign n30480 = n132 & n30479 ;
  assign n30481 = n29483 & n75213 ;
  assign n30482 = n30296 & n30481 ;
  assign n30483 = n30480 | n30482 ;
  assign n30484 = n69261 & n30483 ;
  assign n75288 = ~n29983 ;
  assign n29987 = n75288 & n29986 ;
  assign n30485 = n29502 | n29986 ;
  assign n75289 = ~n30485 ;
  assign n30486 = n30227 & n75289 ;
  assign n30487 = n29987 | n30486 ;
  assign n30488 = n132 & n30487 ;
  assign n30489 = n29492 & n75213 ;
  assign n30490 = n30296 & n30489 ;
  assign n30491 = n30488 | n30490 ;
  assign n30492 = n69075 & n30491 ;
  assign n75290 = ~n30490 ;
  assign n30948 = x100 & n75290 ;
  assign n75291 = ~n30488 ;
  assign n30949 = n75291 & n30948 ;
  assign n30950 = n30492 | n30949 ;
  assign n75292 = ~n30226 ;
  assign n30228 = n29981 & n75292 ;
  assign n30493 = n29511 | n29981 ;
  assign n75293 = ~n30493 ;
  assign n30494 = n29977 & n75293 ;
  assign n30495 = n30228 | n30494 ;
  assign n30496 = n132 & n30495 ;
  assign n30497 = n29501 & n75213 ;
  assign n30498 = n30296 & n30497 ;
  assign n30499 = n30496 | n30498 ;
  assign n30500 = n68993 & n30499 ;
  assign n75294 = ~n29972 ;
  assign n29976 = n75294 & n29975 ;
  assign n30501 = n29519 | n29975 ;
  assign n75295 = ~n30501 ;
  assign n30502 = n30222 & n75295 ;
  assign n30503 = n29976 | n30502 ;
  assign n30504 = n132 & n30503 ;
  assign n30505 = n29510 & n75213 ;
  assign n30506 = n30296 & n30505 ;
  assign n30507 = n30504 | n30506 ;
  assign n30508 = n68716 & n30507 ;
  assign n75296 = ~n30506 ;
  assign n30938 = x98 & n75296 ;
  assign n75297 = ~n30504 ;
  assign n30939 = n75297 & n30938 ;
  assign n30940 = n30508 | n30939 ;
  assign n75298 = ~n30221 ;
  assign n30223 = n29970 & n75298 ;
  assign n30509 = n29528 | n29970 ;
  assign n75299 = ~n30509 ;
  assign n30510 = n29966 & n75299 ;
  assign n30511 = n30223 | n30510 ;
  assign n30512 = n132 & n30511 ;
  assign n30513 = n29518 & n75213 ;
  assign n30514 = n30296 & n30513 ;
  assign n30515 = n30512 | n30514 ;
  assign n30516 = n68545 & n30515 ;
  assign n75300 = ~n29961 ;
  assign n29965 = n75300 & n29964 ;
  assign n30517 = n29537 | n29964 ;
  assign n75301 = ~n30517 ;
  assign n30518 = n30217 & n75301 ;
  assign n30519 = n29965 | n30518 ;
  assign n30520 = n132 & n30519 ;
  assign n30521 = n29527 & n75213 ;
  assign n30522 = n30296 & n30521 ;
  assign n30523 = n30520 | n30522 ;
  assign n30524 = n68438 & n30523 ;
  assign n75302 = ~n30522 ;
  assign n30928 = x96 & n75302 ;
  assign n75303 = ~n30520 ;
  assign n30929 = n75303 & n30928 ;
  assign n30930 = n30524 | n30929 ;
  assign n75304 = ~n30216 ;
  assign n30218 = n29959 & n75304 ;
  assign n30525 = n29546 | n29959 ;
  assign n75305 = ~n30525 ;
  assign n30526 = n29955 & n75305 ;
  assign n30527 = n30218 | n30526 ;
  assign n30528 = n132 & n30527 ;
  assign n30529 = n29536 & n75213 ;
  assign n30530 = n30296 & n30529 ;
  assign n30531 = n30528 | n30530 ;
  assign n30532 = n68214 & n30531 ;
  assign n75306 = ~n29950 ;
  assign n29954 = n75306 & n29953 ;
  assign n30533 = n29555 | n29953 ;
  assign n75307 = ~n30533 ;
  assign n30534 = n30212 & n75307 ;
  assign n30535 = n29954 | n30534 ;
  assign n30536 = n132 & n30535 ;
  assign n30537 = n29545 & n75213 ;
  assign n30538 = n30296 & n30537 ;
  assign n30539 = n30536 | n30538 ;
  assign n30540 = n68058 & n30539 ;
  assign n75308 = ~n30538 ;
  assign n30918 = x94 & n75308 ;
  assign n75309 = ~n30536 ;
  assign n30919 = n75309 & n30918 ;
  assign n30920 = n30540 | n30919 ;
  assign n75310 = ~n30211 ;
  assign n30213 = n29948 & n75310 ;
  assign n30541 = n29564 | n29948 ;
  assign n75311 = ~n30541 ;
  assign n30542 = n29944 & n75311 ;
  assign n30543 = n30213 | n30542 ;
  assign n30544 = n132 & n30543 ;
  assign n30545 = n29554 & n75213 ;
  assign n30546 = n30296 & n30545 ;
  assign n30547 = n30544 | n30546 ;
  assign n30548 = n67986 & n30547 ;
  assign n75312 = ~n29939 ;
  assign n29943 = n75312 & n29942 ;
  assign n30549 = n29573 | n29942 ;
  assign n75313 = ~n30549 ;
  assign n30550 = n30207 & n75313 ;
  assign n30551 = n29943 | n30550 ;
  assign n30552 = n132 & n30551 ;
  assign n30553 = n29563 & n75213 ;
  assign n30554 = n30296 & n30553 ;
  assign n30555 = n30552 | n30554 ;
  assign n30556 = n67763 & n30555 ;
  assign n75314 = ~n30554 ;
  assign n30908 = x92 & n75314 ;
  assign n75315 = ~n30552 ;
  assign n30909 = n75315 & n30908 ;
  assign n30910 = n30556 | n30909 ;
  assign n75316 = ~n30206 ;
  assign n30208 = n29937 & n75316 ;
  assign n30557 = n29582 | n29937 ;
  assign n75317 = ~n30557 ;
  assign n30558 = n29933 & n75317 ;
  assign n30559 = n30208 | n30558 ;
  assign n30560 = n132 & n30559 ;
  assign n30561 = n29572 & n75213 ;
  assign n30562 = n30296 & n30561 ;
  assign n30563 = n30560 | n30562 ;
  assign n30564 = n67622 & n30563 ;
  assign n75318 = ~n29928 ;
  assign n29932 = n75318 & n29931 ;
  assign n30565 = n29591 | n29931 ;
  assign n75319 = ~n30565 ;
  assign n30566 = n30202 & n75319 ;
  assign n30567 = n29932 | n30566 ;
  assign n30568 = n132 & n30567 ;
  assign n30569 = n29581 & n75213 ;
  assign n30570 = n30296 & n30569 ;
  assign n30571 = n30568 | n30570 ;
  assign n30572 = n67531 & n30571 ;
  assign n75320 = ~n30570 ;
  assign n30898 = x90 & n75320 ;
  assign n75321 = ~n30568 ;
  assign n30899 = n75321 & n30898 ;
  assign n30900 = n30572 | n30899 ;
  assign n75322 = ~n30201 ;
  assign n30203 = n29926 & n75322 ;
  assign n30573 = n29600 | n29926 ;
  assign n75323 = ~n30573 ;
  assign n30574 = n29922 & n75323 ;
  assign n30575 = n30203 | n30574 ;
  assign n30576 = n132 & n30575 ;
  assign n30577 = n29590 & n75213 ;
  assign n30578 = n30296 & n30577 ;
  assign n30579 = n30576 | n30578 ;
  assign n30580 = n67348 & n30579 ;
  assign n75324 = ~n29917 ;
  assign n29921 = n75324 & n29920 ;
  assign n30581 = n29609 | n29920 ;
  assign n75325 = ~n30581 ;
  assign n30582 = n30197 & n75325 ;
  assign n30583 = n29921 | n30582 ;
  assign n30584 = n132 & n30583 ;
  assign n30585 = n29599 & n75213 ;
  assign n30586 = n30296 & n30585 ;
  assign n30587 = n30584 | n30586 ;
  assign n30588 = n67222 & n30587 ;
  assign n75326 = ~n30586 ;
  assign n30888 = x88 & n75326 ;
  assign n75327 = ~n30584 ;
  assign n30889 = n75327 & n30888 ;
  assign n30890 = n30588 | n30889 ;
  assign n75328 = ~n30196 ;
  assign n30198 = n29915 & n75328 ;
  assign n30589 = n29618 | n29915 ;
  assign n75329 = ~n30589 ;
  assign n30590 = n29911 & n75329 ;
  assign n30591 = n30198 | n30590 ;
  assign n30592 = n132 & n30591 ;
  assign n30593 = n29608 & n75213 ;
  assign n30594 = n30296 & n30593 ;
  assign n30595 = n30592 | n30594 ;
  assign n30596 = n67164 & n30595 ;
  assign n75330 = ~n29906 ;
  assign n29910 = n75330 & n29909 ;
  assign n30597 = n29627 | n29909 ;
  assign n75331 = ~n30597 ;
  assign n30598 = n30192 & n75331 ;
  assign n30599 = n29910 | n30598 ;
  assign n30600 = n132 & n30599 ;
  assign n30601 = n29617 & n75213 ;
  assign n30602 = n30296 & n30601 ;
  assign n30603 = n30600 | n30602 ;
  assign n30604 = n66979 & n30603 ;
  assign n75332 = ~n30602 ;
  assign n30878 = x86 & n75332 ;
  assign n75333 = ~n30600 ;
  assign n30879 = n75333 & n30878 ;
  assign n30880 = n30604 | n30879 ;
  assign n75334 = ~n30191 ;
  assign n30193 = n29904 & n75334 ;
  assign n30605 = n29636 | n29904 ;
  assign n75335 = ~n30605 ;
  assign n30606 = n29900 & n75335 ;
  assign n30607 = n30193 | n30606 ;
  assign n30608 = n132 & n30607 ;
  assign n30609 = n29626 & n75213 ;
  assign n30610 = n30296 & n30609 ;
  assign n30611 = n30608 | n30610 ;
  assign n30612 = n66868 & n30611 ;
  assign n75336 = ~n29895 ;
  assign n29899 = n75336 & n29898 ;
  assign n30613 = n29645 | n29898 ;
  assign n75337 = ~n30613 ;
  assign n30614 = n30187 & n75337 ;
  assign n30615 = n29899 | n30614 ;
  assign n30616 = n132 & n30615 ;
  assign n30617 = n29635 & n75213 ;
  assign n30618 = n30296 & n30617 ;
  assign n30619 = n30616 | n30618 ;
  assign n30620 = n66797 & n30619 ;
  assign n75338 = ~n30618 ;
  assign n30868 = x84 & n75338 ;
  assign n75339 = ~n30616 ;
  assign n30869 = n75339 & n30868 ;
  assign n30870 = n30620 | n30869 ;
  assign n75340 = ~n30186 ;
  assign n30188 = n29893 & n75340 ;
  assign n30621 = n29654 | n29893 ;
  assign n75341 = ~n30621 ;
  assign n30622 = n29889 & n75341 ;
  assign n30623 = n30188 | n30622 ;
  assign n30624 = n132 & n30623 ;
  assign n30625 = n29644 & n75213 ;
  assign n30626 = n30296 & n30625 ;
  assign n30627 = n30624 | n30626 ;
  assign n30628 = n66654 & n30627 ;
  assign n75342 = ~n29884 ;
  assign n29888 = n75342 & n29887 ;
  assign n30629 = n29663 | n29887 ;
  assign n75343 = ~n30629 ;
  assign n30630 = n30182 & n75343 ;
  assign n30631 = n29888 | n30630 ;
  assign n30632 = n132 & n30631 ;
  assign n30633 = n29653 & n75213 ;
  assign n30634 = n30296 & n30633 ;
  assign n30635 = n30632 | n30634 ;
  assign n30636 = n66560 & n30635 ;
  assign n75344 = ~n30634 ;
  assign n30858 = x82 & n75344 ;
  assign n75345 = ~n30632 ;
  assign n30859 = n75345 & n30858 ;
  assign n30860 = n30636 | n30859 ;
  assign n75346 = ~n30181 ;
  assign n30183 = n29882 & n75346 ;
  assign n30637 = n29672 | n29882 ;
  assign n75347 = ~n30637 ;
  assign n30638 = n29878 & n75347 ;
  assign n30639 = n30183 | n30638 ;
  assign n30640 = n132 & n30639 ;
  assign n30641 = n29662 & n75213 ;
  assign n30642 = n30296 & n30641 ;
  assign n30643 = n30640 | n30642 ;
  assign n30644 = n66505 & n30643 ;
  assign n75348 = ~n29873 ;
  assign n29877 = n75348 & n29876 ;
  assign n30645 = n29681 | n29876 ;
  assign n75349 = ~n30645 ;
  assign n30646 = n30177 & n75349 ;
  assign n30647 = n29877 | n30646 ;
  assign n30648 = n132 & n30647 ;
  assign n30649 = n29671 & n75213 ;
  assign n30650 = n30296 & n30649 ;
  assign n30651 = n30648 | n30650 ;
  assign n30652 = n66379 & n30651 ;
  assign n75350 = ~n30650 ;
  assign n30848 = x80 & n75350 ;
  assign n75351 = ~n30648 ;
  assign n30849 = n75351 & n30848 ;
  assign n30850 = n30652 | n30849 ;
  assign n75352 = ~n30176 ;
  assign n30178 = n29871 & n75352 ;
  assign n30653 = n29690 | n29871 ;
  assign n75353 = ~n30653 ;
  assign n30654 = n29867 & n75353 ;
  assign n30655 = n30178 | n30654 ;
  assign n30656 = n132 & n30655 ;
  assign n30657 = n29680 & n75213 ;
  assign n30658 = n30296 & n30657 ;
  assign n30659 = n30656 | n30658 ;
  assign n30660 = n66299 & n30659 ;
  assign n75354 = ~n29862 ;
  assign n29866 = n75354 & n29865 ;
  assign n30661 = n29699 | n29865 ;
  assign n75355 = ~n30661 ;
  assign n30662 = n30172 & n75355 ;
  assign n30663 = n29866 | n30662 ;
  assign n30664 = n132 & n30663 ;
  assign n30665 = n29689 & n75213 ;
  assign n30666 = n30296 & n30665 ;
  assign n30667 = n30664 | n30666 ;
  assign n30668 = n66244 & n30667 ;
  assign n75356 = ~n30666 ;
  assign n30837 = x78 & n75356 ;
  assign n75357 = ~n30664 ;
  assign n30838 = n75357 & n30837 ;
  assign n30839 = n30668 | n30838 ;
  assign n75358 = ~n30171 ;
  assign n30173 = n29860 & n75358 ;
  assign n30669 = n29708 | n29860 ;
  assign n75359 = ~n30669 ;
  assign n30670 = n29856 & n75359 ;
  assign n30671 = n30173 | n30670 ;
  assign n30672 = n132 & n30671 ;
  assign n30673 = n29698 & n75213 ;
  assign n30674 = n30296 & n30673 ;
  assign n30675 = n30672 | n30674 ;
  assign n30676 = n66145 & n30675 ;
  assign n75360 = ~n29851 ;
  assign n29855 = n75360 & n29854 ;
  assign n30677 = n29717 | n29854 ;
  assign n75361 = ~n30677 ;
  assign n30678 = n30167 & n75361 ;
  assign n30679 = n29855 | n30678 ;
  assign n30680 = n132 & n30679 ;
  assign n30681 = n29707 & n75213 ;
  assign n30682 = n30296 & n30681 ;
  assign n30683 = n30680 | n30682 ;
  assign n30684 = n66081 & n30683 ;
  assign n75362 = ~n30682 ;
  assign n30827 = x76 & n75362 ;
  assign n75363 = ~n30680 ;
  assign n30828 = n75363 & n30827 ;
  assign n30829 = n30684 | n30828 ;
  assign n75364 = ~n30166 ;
  assign n30168 = n29849 & n75364 ;
  assign n30685 = n29726 | n29849 ;
  assign n75365 = ~n30685 ;
  assign n30686 = n29845 & n75365 ;
  assign n30687 = n30168 | n30686 ;
  assign n30688 = n132 & n30687 ;
  assign n30689 = n29716 & n75213 ;
  assign n30690 = n30296 & n30689 ;
  assign n30691 = n30688 | n30690 ;
  assign n30692 = n66043 & n30691 ;
  assign n75366 = ~n29840 ;
  assign n29844 = n75366 & n29843 ;
  assign n30693 = n29735 | n29843 ;
  assign n75367 = ~n30693 ;
  assign n30694 = n30162 & n75367 ;
  assign n30695 = n29844 | n30694 ;
  assign n30696 = n132 & n30695 ;
  assign n30697 = n29725 & n75213 ;
  assign n30698 = n30296 & n30697 ;
  assign n30699 = n30696 | n30698 ;
  assign n30700 = n65960 & n30699 ;
  assign n75368 = ~n30698 ;
  assign n30817 = x74 & n75368 ;
  assign n75369 = ~n30696 ;
  assign n30818 = n75369 & n30817 ;
  assign n30819 = n30700 | n30818 ;
  assign n75370 = ~n30161 ;
  assign n30163 = n29838 & n75370 ;
  assign n30701 = n29744 | n29838 ;
  assign n75371 = ~n30701 ;
  assign n30702 = n29834 & n75371 ;
  assign n30703 = n30163 | n30702 ;
  assign n30704 = n132 & n30703 ;
  assign n30705 = n29734 & n75213 ;
  assign n30706 = n30296 & n30705 ;
  assign n30707 = n30704 | n30706 ;
  assign n30708 = n65909 & n30707 ;
  assign n75372 = ~n29829 ;
  assign n29833 = n75372 & n29832 ;
  assign n30709 = n29752 | n29832 ;
  assign n75373 = ~n30709 ;
  assign n30710 = n30157 & n75373 ;
  assign n30711 = n29833 | n30710 ;
  assign n30712 = n132 & n30711 ;
  assign n30713 = n29743 & n75213 ;
  assign n30714 = n30296 & n30713 ;
  assign n30715 = n30712 | n30714 ;
  assign n30716 = n65877 & n30715 ;
  assign n75374 = ~n30714 ;
  assign n30807 = x72 & n75374 ;
  assign n75375 = ~n30712 ;
  assign n30808 = n75375 & n30807 ;
  assign n30809 = n30716 | n30808 ;
  assign n75376 = ~n30156 ;
  assign n30158 = n29827 & n75376 ;
  assign n30717 = n29761 | n29827 ;
  assign n75377 = ~n30717 ;
  assign n30718 = n29823 & n75377 ;
  assign n30719 = n30158 | n30718 ;
  assign n30720 = n132 & n30719 ;
  assign n30721 = n29751 & n75213 ;
  assign n30722 = n30296 & n30721 ;
  assign n30723 = n30720 | n30722 ;
  assign n30724 = n65820 & n30723 ;
  assign n75378 = ~n29818 ;
  assign n29822 = n75378 & n29821 ;
  assign n30725 = n29770 | n29821 ;
  assign n75379 = ~n30725 ;
  assign n30726 = n30153 & n75379 ;
  assign n30727 = n29822 | n30726 ;
  assign n30728 = n132 & n30727 ;
  assign n30729 = n29760 & n75213 ;
  assign n30730 = n30296 & n30729 ;
  assign n30731 = n30728 | n30730 ;
  assign n30732 = n65791 & n30731 ;
  assign n75380 = ~n30730 ;
  assign n30797 = x70 & n75380 ;
  assign n75381 = ~n30728 ;
  assign n30798 = n75381 & n30797 ;
  assign n30799 = n30732 | n30798 ;
  assign n75382 = ~n30151 ;
  assign n30152 = n29816 & n75382 ;
  assign n30733 = n29778 | n29816 ;
  assign n75383 = ~n30733 ;
  assign n30734 = n29812 & n75383 ;
  assign n30735 = n30152 | n30734 ;
  assign n30736 = n132 & n30735 ;
  assign n30737 = n29769 & n75213 ;
  assign n30738 = n30296 & n30737 ;
  assign n30739 = n30736 | n30738 ;
  assign n30740 = n65772 & n30739 ;
  assign n75384 = ~n29808 ;
  assign n30149 = n75384 & n29811 ;
  assign n30741 = n29786 | n29811 ;
  assign n75385 = ~n30741 ;
  assign n30742 = n29807 & n75385 ;
  assign n30743 = n30149 | n30742 ;
  assign n30744 = n132 & n30743 ;
  assign n30745 = n29777 & n75213 ;
  assign n30746 = n30296 & n30745 ;
  assign n30747 = n30744 | n30746 ;
  assign n30748 = n65746 & n30747 ;
  assign n75386 = ~n30746 ;
  assign n30787 = x68 & n75386 ;
  assign n75387 = ~n30744 ;
  assign n30788 = n75387 & n30787 ;
  assign n30789 = n30748 | n30788 ;
  assign n75388 = ~n29803 ;
  assign n30750 = n75388 & n29806 ;
  assign n30749 = n29802 | n29806 ;
  assign n75389 = ~n30749 ;
  assign n30751 = n29801 & n75389 ;
  assign n30752 = n30750 | n30751 ;
  assign n30753 = n132 & n30752 ;
  assign n30754 = n29785 & n75213 ;
  assign n30755 = n30296 & n30754 ;
  assign n30756 = n30753 | n30755 ;
  assign n30757 = n65721 & n30756 ;
  assign n30758 = n29798 & n29800 ;
  assign n30759 = n75033 & n30758 ;
  assign n75390 = ~n30759 ;
  assign n30760 = n30145 & n75390 ;
  assign n30761 = n132 & n30760 ;
  assign n30762 = n29795 & n75213 ;
  assign n30763 = n30296 & n30762 ;
  assign n30764 = n30761 | n30763 ;
  assign n30765 = n65686 & n30764 ;
  assign n75391 = ~n30763 ;
  assign n30777 = x66 & n75391 ;
  assign n75392 = ~n30761 ;
  assign n30778 = n75392 & n30777 ;
  assign n30779 = n30765 | n30778 ;
  assign n30141 = n29800 & n132 ;
  assign n30140 = x64 & n132 ;
  assign n75393 = ~n30140 ;
  assign n30766 = x3 & n75393 ;
  assign n30767 = n30141 | n30766 ;
  assign n30768 = x65 & n30767 ;
  assign n30769 = n75213 & n30296 ;
  assign n75394 = ~n30769 ;
  assign n30770 = n29800 & n75394 ;
  assign n30771 = x65 | n30770 ;
  assign n30772 = n30766 | n30771 ;
  assign n75395 = ~n30768 ;
  assign n30773 = n75395 & n30772 ;
  assign n75396 = ~x2 ;
  assign n30774 = n75396 & x64 ;
  assign n30775 = n30773 | n30774 ;
  assign n30776 = n65670 & n30767 ;
  assign n75397 = ~n30776 ;
  assign n30780 = n30775 & n75397 ;
  assign n30781 = n30779 | n30780 ;
  assign n75398 = ~n30765 ;
  assign n30782 = n75398 & n30781 ;
  assign n75399 = ~n30755 ;
  assign n30783 = x67 & n75399 ;
  assign n75400 = ~n30753 ;
  assign n30784 = n75400 & n30783 ;
  assign n30785 = n30757 | n30784 ;
  assign n30786 = n30782 | n30785 ;
  assign n75401 = ~n30757 ;
  assign n30790 = n75401 & n30786 ;
  assign n30791 = n30789 | n30790 ;
  assign n75402 = ~n30748 ;
  assign n30792 = n75402 & n30791 ;
  assign n75403 = ~n30738 ;
  assign n30793 = x69 & n75403 ;
  assign n75404 = ~n30736 ;
  assign n30794 = n75404 & n30793 ;
  assign n30795 = n30740 | n30794 ;
  assign n30796 = n30792 | n30795 ;
  assign n75405 = ~n30740 ;
  assign n30800 = n75405 & n30796 ;
  assign n30801 = n30799 | n30800 ;
  assign n75406 = ~n30732 ;
  assign n30802 = n75406 & n30801 ;
  assign n75407 = ~n30722 ;
  assign n30803 = x71 & n75407 ;
  assign n75408 = ~n30720 ;
  assign n30804 = n75408 & n30803 ;
  assign n30805 = n30724 | n30804 ;
  assign n30806 = n30802 | n30805 ;
  assign n75409 = ~n30724 ;
  assign n30810 = n75409 & n30806 ;
  assign n30811 = n30809 | n30810 ;
  assign n75410 = ~n30716 ;
  assign n30812 = n75410 & n30811 ;
  assign n75411 = ~n30706 ;
  assign n30813 = x73 & n75411 ;
  assign n75412 = ~n30704 ;
  assign n30814 = n75412 & n30813 ;
  assign n30815 = n30708 | n30814 ;
  assign n30816 = n30812 | n30815 ;
  assign n75413 = ~n30708 ;
  assign n30820 = n75413 & n30816 ;
  assign n30821 = n30819 | n30820 ;
  assign n75414 = ~n30700 ;
  assign n30822 = n75414 & n30821 ;
  assign n75415 = ~n30690 ;
  assign n30823 = x75 & n75415 ;
  assign n75416 = ~n30688 ;
  assign n30824 = n75416 & n30823 ;
  assign n30825 = n30692 | n30824 ;
  assign n30826 = n30822 | n30825 ;
  assign n75417 = ~n30692 ;
  assign n30830 = n75417 & n30826 ;
  assign n30831 = n30829 | n30830 ;
  assign n75418 = ~n30684 ;
  assign n30832 = n75418 & n30831 ;
  assign n75419 = ~n30674 ;
  assign n30833 = x77 & n75419 ;
  assign n75420 = ~n30672 ;
  assign n30834 = n75420 & n30833 ;
  assign n30835 = n30676 | n30834 ;
  assign n30836 = n30832 | n30835 ;
  assign n75421 = ~n30676 ;
  assign n30841 = n75421 & n30836 ;
  assign n30842 = n30839 | n30841 ;
  assign n75422 = ~n30668 ;
  assign n30843 = n75422 & n30842 ;
  assign n75423 = ~n30658 ;
  assign n30844 = x79 & n75423 ;
  assign n75424 = ~n30656 ;
  assign n30845 = n75424 & n30844 ;
  assign n30846 = n30660 | n30845 ;
  assign n30847 = n30843 | n30846 ;
  assign n75425 = ~n30660 ;
  assign n30851 = n75425 & n30847 ;
  assign n30852 = n30850 | n30851 ;
  assign n75426 = ~n30652 ;
  assign n30853 = n75426 & n30852 ;
  assign n75427 = ~n30642 ;
  assign n30854 = x81 & n75427 ;
  assign n75428 = ~n30640 ;
  assign n30855 = n75428 & n30854 ;
  assign n30856 = n30644 | n30855 ;
  assign n30857 = n30853 | n30856 ;
  assign n75429 = ~n30644 ;
  assign n30861 = n75429 & n30857 ;
  assign n30862 = n30860 | n30861 ;
  assign n75430 = ~n30636 ;
  assign n30863 = n75430 & n30862 ;
  assign n75431 = ~n30626 ;
  assign n30864 = x83 & n75431 ;
  assign n75432 = ~n30624 ;
  assign n30865 = n75432 & n30864 ;
  assign n30866 = n30628 | n30865 ;
  assign n30867 = n30863 | n30866 ;
  assign n75433 = ~n30628 ;
  assign n30871 = n75433 & n30867 ;
  assign n30872 = n30870 | n30871 ;
  assign n75434 = ~n30620 ;
  assign n30873 = n75434 & n30872 ;
  assign n75435 = ~n30610 ;
  assign n30874 = x85 & n75435 ;
  assign n75436 = ~n30608 ;
  assign n30875 = n75436 & n30874 ;
  assign n30876 = n30612 | n30875 ;
  assign n30877 = n30873 | n30876 ;
  assign n75437 = ~n30612 ;
  assign n30881 = n75437 & n30877 ;
  assign n30882 = n30880 | n30881 ;
  assign n75438 = ~n30604 ;
  assign n30883 = n75438 & n30882 ;
  assign n75439 = ~n30594 ;
  assign n30884 = x87 & n75439 ;
  assign n75440 = ~n30592 ;
  assign n30885 = n75440 & n30884 ;
  assign n30886 = n30596 | n30885 ;
  assign n30887 = n30883 | n30886 ;
  assign n75441 = ~n30596 ;
  assign n30891 = n75441 & n30887 ;
  assign n30892 = n30890 | n30891 ;
  assign n75442 = ~n30588 ;
  assign n30893 = n75442 & n30892 ;
  assign n75443 = ~n30578 ;
  assign n30894 = x89 & n75443 ;
  assign n75444 = ~n30576 ;
  assign n30895 = n75444 & n30894 ;
  assign n30896 = n30580 | n30895 ;
  assign n30897 = n30893 | n30896 ;
  assign n75445 = ~n30580 ;
  assign n30901 = n75445 & n30897 ;
  assign n30902 = n30900 | n30901 ;
  assign n75446 = ~n30572 ;
  assign n30903 = n75446 & n30902 ;
  assign n75447 = ~n30562 ;
  assign n30904 = x91 & n75447 ;
  assign n75448 = ~n30560 ;
  assign n30905 = n75448 & n30904 ;
  assign n30906 = n30564 | n30905 ;
  assign n30907 = n30903 | n30906 ;
  assign n75449 = ~n30564 ;
  assign n30911 = n75449 & n30907 ;
  assign n30912 = n30910 | n30911 ;
  assign n75450 = ~n30556 ;
  assign n30913 = n75450 & n30912 ;
  assign n75451 = ~n30546 ;
  assign n30914 = x93 & n75451 ;
  assign n75452 = ~n30544 ;
  assign n30915 = n75452 & n30914 ;
  assign n30916 = n30548 | n30915 ;
  assign n30917 = n30913 | n30916 ;
  assign n75453 = ~n30548 ;
  assign n30921 = n75453 & n30917 ;
  assign n30922 = n30920 | n30921 ;
  assign n75454 = ~n30540 ;
  assign n30923 = n75454 & n30922 ;
  assign n75455 = ~n30530 ;
  assign n30924 = x95 & n75455 ;
  assign n75456 = ~n30528 ;
  assign n30925 = n75456 & n30924 ;
  assign n30926 = n30532 | n30925 ;
  assign n30927 = n30923 | n30926 ;
  assign n75457 = ~n30532 ;
  assign n30931 = n75457 & n30927 ;
  assign n30932 = n30930 | n30931 ;
  assign n75458 = ~n30524 ;
  assign n30933 = n75458 & n30932 ;
  assign n75459 = ~n30514 ;
  assign n30934 = x97 & n75459 ;
  assign n75460 = ~n30512 ;
  assign n30935 = n75460 & n30934 ;
  assign n30936 = n30516 | n30935 ;
  assign n30937 = n30933 | n30936 ;
  assign n75461 = ~n30516 ;
  assign n30941 = n75461 & n30937 ;
  assign n30942 = n30940 | n30941 ;
  assign n75462 = ~n30508 ;
  assign n30943 = n75462 & n30942 ;
  assign n75463 = ~n30498 ;
  assign n30944 = x99 & n75463 ;
  assign n75464 = ~n30496 ;
  assign n30945 = n75464 & n30944 ;
  assign n30946 = n30500 | n30945 ;
  assign n30947 = n30943 | n30946 ;
  assign n75465 = ~n30500 ;
  assign n30951 = n75465 & n30947 ;
  assign n30952 = n30950 | n30951 ;
  assign n75466 = ~n30492 ;
  assign n30953 = n75466 & n30952 ;
  assign n75467 = ~n30482 ;
  assign n30954 = x101 & n75467 ;
  assign n75468 = ~n30480 ;
  assign n30955 = n75468 & n30954 ;
  assign n30956 = n30484 | n30955 ;
  assign n30957 = n30953 | n30956 ;
  assign n75469 = ~n30484 ;
  assign n30961 = n75469 & n30957 ;
  assign n30962 = n30960 | n30961 ;
  assign n75470 = ~n30476 ;
  assign n30963 = n75470 & n30962 ;
  assign n75471 = ~n30466 ;
  assign n30964 = x103 & n75471 ;
  assign n75472 = ~n30464 ;
  assign n30965 = n75472 & n30964 ;
  assign n30966 = n30468 | n30965 ;
  assign n30967 = n30963 | n30966 ;
  assign n75473 = ~n30468 ;
  assign n30971 = n75473 & n30967 ;
  assign n30972 = n30970 | n30971 ;
  assign n75474 = ~n30460 ;
  assign n30973 = n75474 & n30972 ;
  assign n75475 = ~n30450 ;
  assign n30974 = x105 & n75475 ;
  assign n75476 = ~n30448 ;
  assign n30975 = n75476 & n30974 ;
  assign n30976 = n30452 | n30975 ;
  assign n30977 = n30973 | n30976 ;
  assign n75477 = ~n30452 ;
  assign n30981 = n75477 & n30977 ;
  assign n30982 = n30980 | n30981 ;
  assign n75478 = ~n30444 ;
  assign n30983 = n75478 & n30982 ;
  assign n75479 = ~n30434 ;
  assign n30984 = x107 & n75479 ;
  assign n75480 = ~n30432 ;
  assign n30985 = n75480 & n30984 ;
  assign n30986 = n30436 | n30985 ;
  assign n30987 = n30983 | n30986 ;
  assign n75481 = ~n30436 ;
  assign n30991 = n75481 & n30987 ;
  assign n30992 = n30990 | n30991 ;
  assign n75482 = ~n30428 ;
  assign n30993 = n75482 & n30992 ;
  assign n75483 = ~n30418 ;
  assign n30994 = x109 & n75483 ;
  assign n75484 = ~n30416 ;
  assign n30995 = n75484 & n30994 ;
  assign n30996 = n30420 | n30995 ;
  assign n30997 = n30993 | n30996 ;
  assign n75485 = ~n30420 ;
  assign n31001 = n75485 & n30997 ;
  assign n31002 = n31000 | n31001 ;
  assign n75486 = ~n30412 ;
  assign n31003 = n75486 & n31002 ;
  assign n75487 = ~n30402 ;
  assign n31004 = x111 & n75487 ;
  assign n75488 = ~n30400 ;
  assign n31005 = n75488 & n31004 ;
  assign n31006 = n30404 | n31005 ;
  assign n31008 = n31003 | n31006 ;
  assign n75489 = ~n30404 ;
  assign n31012 = n75489 & n31008 ;
  assign n31013 = n31011 | n31012 ;
  assign n75490 = ~n30396 ;
  assign n31014 = n75490 & n31013 ;
  assign n75491 = ~n30386 ;
  assign n31015 = x113 & n75491 ;
  assign n75492 = ~n30384 ;
  assign n31016 = n75492 & n31015 ;
  assign n31017 = n30388 | n31016 ;
  assign n31019 = n31014 | n31017 ;
  assign n75493 = ~n30388 ;
  assign n31023 = n75493 & n31019 ;
  assign n31024 = n31022 | n31023 ;
  assign n75494 = ~n30380 ;
  assign n31025 = n75494 & n31024 ;
  assign n75495 = ~n30370 ;
  assign n31026 = x115 & n75495 ;
  assign n75496 = ~n30368 ;
  assign n31027 = n75496 & n31026 ;
  assign n31028 = n30372 | n31027 ;
  assign n31029 = n31025 | n31028 ;
  assign n75497 = ~n30372 ;
  assign n31033 = n75497 & n31029 ;
  assign n31034 = n31032 | n31033 ;
  assign n75498 = ~n30364 ;
  assign n31035 = n75498 & n31034 ;
  assign n75499 = ~n30354 ;
  assign n31036 = x117 & n75499 ;
  assign n75500 = ~n30352 ;
  assign n31037 = n75500 & n31036 ;
  assign n31038 = n30356 | n31037 ;
  assign n31039 = n31035 | n31038 ;
  assign n75501 = ~n30356 ;
  assign n31043 = n75501 & n31039 ;
  assign n31044 = n31042 | n31043 ;
  assign n75502 = ~n30348 ;
  assign n31045 = n75502 & n31044 ;
  assign n75503 = ~n30338 ;
  assign n31046 = x119 & n75503 ;
  assign n75504 = ~n30336 ;
  assign n31047 = n75504 & n31046 ;
  assign n31048 = n30340 | n31047 ;
  assign n31049 = n31045 | n31048 ;
  assign n75505 = ~n30340 ;
  assign n31053 = n75505 & n31049 ;
  assign n31054 = n31052 | n31053 ;
  assign n75506 = ~n30332 ;
  assign n31055 = n75506 & n31054 ;
  assign n75507 = ~n30322 ;
  assign n31056 = x121 & n75507 ;
  assign n75508 = ~n30320 ;
  assign n31057 = n75508 & n31056 ;
  assign n31058 = n30324 | n31057 ;
  assign n31060 = n31055 | n31058 ;
  assign n75509 = ~n30324 ;
  assign n31064 = n75509 & n31060 ;
  assign n31065 = n31063 | n31064 ;
  assign n75510 = ~n30316 ;
  assign n31066 = n75510 & n31065 ;
  assign n75511 = ~n30306 ;
  assign n31067 = x123 & n75511 ;
  assign n75512 = ~n30304 ;
  assign n31068 = n75512 & n31067 ;
  assign n31069 = n30308 | n31068 ;
  assign n31070 = n31066 | n31069 ;
  assign n75513 = ~n30308 ;
  assign n31074 = n75513 & n31070 ;
  assign n31075 = n31073 | n31074 ;
  assign n75514 = ~n30300 ;
  assign n31076 = n75514 & n31075 ;
  assign n31077 = n29282 | n30134 ;
  assign n31078 = n30132 | n31077 ;
  assign n75515 = ~n31078 ;
  assign n31079 = n30120 & n75515 ;
  assign n31080 = n30132 | n30134 ;
  assign n75516 = ~n30295 ;
  assign n31081 = n75516 & n31080 ;
  assign n31082 = n31079 | n31081 ;
  assign n31083 = n132 & n31082 ;
  assign n31084 = n65369 & n30131 ;
  assign n31085 = n30296 & n31084 ;
  assign n31086 = n31083 | n31085 ;
  assign n75517 = ~x125 ;
  assign n31087 = n75517 & n31086 ;
  assign n75518 = ~n31085 ;
  assign n31088 = x125 & n75518 ;
  assign n75519 = ~n31083 ;
  assign n31089 = n75519 & n31088 ;
  assign n31090 = n65362 | n31089 ;
  assign n31091 = n31087 | n31090 ;
  assign n31092 = n31076 | n31091 ;
  assign n31093 = n73624 & n31086 ;
  assign n75520 = ~n31093 ;
  assign n31094 = n31092 & n75520 ;
  assign n32103 = n30300 | n31089 ;
  assign n32104 = n31087 | n32103 ;
  assign n75521 = ~n32104 ;
  assign n32105 = n31075 & n75521 ;
  assign n31096 = x64 & n75394 ;
  assign n75522 = ~n31096 ;
  assign n31097 = x3 & n75522 ;
  assign n31098 = n30141 | n31097 ;
  assign n31099 = x65 & n31098 ;
  assign n75523 = ~n31099 ;
  assign n31100 = n30772 & n75523 ;
  assign n31101 = n30774 | n31100 ;
  assign n31102 = n75397 & n31101 ;
  assign n31104 = n30779 | n31102 ;
  assign n31105 = n75398 & n31104 ;
  assign n31106 = n30785 | n31105 ;
  assign n31107 = n75401 & n31106 ;
  assign n31108 = n30789 | n31107 ;
  assign n31109 = n75402 & n31108 ;
  assign n31110 = n30795 | n31109 ;
  assign n31111 = n75405 & n31110 ;
  assign n31112 = n30799 | n31111 ;
  assign n31113 = n75406 & n31112 ;
  assign n31114 = n30805 | n31113 ;
  assign n31115 = n75409 & n31114 ;
  assign n31116 = n30809 | n31115 ;
  assign n31117 = n75410 & n31116 ;
  assign n31118 = n30815 | n31117 ;
  assign n31119 = n75413 & n31118 ;
  assign n31120 = n30819 | n31119 ;
  assign n31121 = n75414 & n31120 ;
  assign n31122 = n30825 | n31121 ;
  assign n31123 = n75417 & n31122 ;
  assign n31124 = n30829 | n31123 ;
  assign n31125 = n75418 & n31124 ;
  assign n31126 = n30835 | n31125 ;
  assign n31127 = n75421 & n31126 ;
  assign n31128 = n30839 | n31127 ;
  assign n31129 = n75422 & n31128 ;
  assign n31130 = n30846 | n31129 ;
  assign n31131 = n75425 & n31130 ;
  assign n31132 = n30850 | n31131 ;
  assign n31133 = n75426 & n31132 ;
  assign n31134 = n30856 | n31133 ;
  assign n31135 = n75429 & n31134 ;
  assign n31136 = n30860 | n31135 ;
  assign n31137 = n75430 & n31136 ;
  assign n31138 = n30866 | n31137 ;
  assign n31139 = n75433 & n31138 ;
  assign n31140 = n30870 | n31139 ;
  assign n31141 = n75434 & n31140 ;
  assign n31142 = n30876 | n31141 ;
  assign n31143 = n75437 & n31142 ;
  assign n31144 = n30880 | n31143 ;
  assign n31145 = n75438 & n31144 ;
  assign n31146 = n30886 | n31145 ;
  assign n31147 = n75441 & n31146 ;
  assign n31148 = n30890 | n31147 ;
  assign n31149 = n75442 & n31148 ;
  assign n31150 = n30896 | n31149 ;
  assign n31151 = n75445 & n31150 ;
  assign n31152 = n30900 | n31151 ;
  assign n31153 = n75446 & n31152 ;
  assign n31154 = n30906 | n31153 ;
  assign n31155 = n75449 & n31154 ;
  assign n31156 = n30910 | n31155 ;
  assign n31157 = n75450 & n31156 ;
  assign n31158 = n30916 | n31157 ;
  assign n31159 = n75453 & n31158 ;
  assign n31160 = n30920 | n31159 ;
  assign n31161 = n75454 & n31160 ;
  assign n31162 = n30926 | n31161 ;
  assign n31163 = n75457 & n31162 ;
  assign n31164 = n30930 | n31163 ;
  assign n31165 = n75458 & n31164 ;
  assign n31166 = n30936 | n31165 ;
  assign n31167 = n75461 & n31166 ;
  assign n31168 = n30940 | n31167 ;
  assign n31169 = n75462 & n31168 ;
  assign n31170 = n30946 | n31169 ;
  assign n31171 = n75465 & n31170 ;
  assign n31172 = n30950 | n31171 ;
  assign n31173 = n75466 & n31172 ;
  assign n31174 = n30956 | n31173 ;
  assign n31175 = n75469 & n31174 ;
  assign n31176 = n30960 | n31175 ;
  assign n31177 = n75470 & n31176 ;
  assign n31178 = n30966 | n31177 ;
  assign n31179 = n75473 & n31178 ;
  assign n31180 = n30970 | n31179 ;
  assign n31181 = n75474 & n31180 ;
  assign n31182 = n30976 | n31181 ;
  assign n31183 = n75477 & n31182 ;
  assign n31184 = n30980 | n31183 ;
  assign n31185 = n75478 & n31184 ;
  assign n31186 = n30986 | n31185 ;
  assign n31187 = n75481 & n31186 ;
  assign n31188 = n30990 | n31187 ;
  assign n31189 = n75482 & n31188 ;
  assign n31190 = n30996 | n31189 ;
  assign n31191 = n75485 & n31190 ;
  assign n31192 = n31000 | n31191 ;
  assign n31193 = n75486 & n31192 ;
  assign n31194 = n31006 | n31193 ;
  assign n31195 = n75489 & n31194 ;
  assign n31196 = n31011 | n31195 ;
  assign n31197 = n75490 & n31196 ;
  assign n31198 = n31017 | n31197 ;
  assign n31199 = n75493 & n31198 ;
  assign n31200 = n31022 | n31199 ;
  assign n31201 = n75494 & n31200 ;
  assign n31202 = n31028 | n31201 ;
  assign n31203 = n75497 & n31202 ;
  assign n31204 = n31032 | n31203 ;
  assign n31205 = n75498 & n31204 ;
  assign n31206 = n31038 | n31205 ;
  assign n31207 = n75501 & n31206 ;
  assign n31208 = n31042 | n31207 ;
  assign n31209 = n75502 & n31208 ;
  assign n31210 = n31048 | n31209 ;
  assign n31211 = n75505 & n31210 ;
  assign n31212 = n31052 | n31211 ;
  assign n31213 = n75506 & n31212 ;
  assign n31214 = n31058 | n31213 ;
  assign n31215 = n75509 & n31214 ;
  assign n31216 = n31063 | n31215 ;
  assign n31217 = n75510 & n31216 ;
  assign n31218 = n31069 | n31217 ;
  assign n31219 = n75513 & n31218 ;
  assign n31754 = n31073 | n31219 ;
  assign n31755 = n75514 & n31754 ;
  assign n32106 = n31087 | n31089 ;
  assign n75524 = ~n31755 ;
  assign n32107 = n75524 & n32106 ;
  assign n32108 = n32105 | n32107 ;
  assign n131 = ~n31094 ;
  assign n32109 = n131 & n32108 ;
  assign n32110 = n274 & n31086 ;
  assign n32111 = n31092 & n32110 ;
  assign n32112 = n32109 | n32111 ;
  assign n75526 = ~n65362 ;
  assign n32118 = n75526 & n32112 ;
  assign n75527 = ~n31074 ;
  assign n31220 = n31073 & n75527 ;
  assign n31221 = n30308 | n31073 ;
  assign n75528 = ~n31221 ;
  assign n31222 = n31218 & n75528 ;
  assign n31223 = n31220 | n31222 ;
  assign n31224 = n131 & n31223 ;
  assign n31225 = n30299 & n75520 ;
  assign n31226 = n31092 & n31225 ;
  assign n31227 = n31224 | n31226 ;
  assign n31228 = n75517 & n31227 ;
  assign n75529 = ~n31217 ;
  assign n31229 = n31069 & n75529 ;
  assign n31230 = n30316 | n31069 ;
  assign n75530 = ~n31230 ;
  assign n31231 = n31065 & n75530 ;
  assign n31232 = n31229 | n31231 ;
  assign n31233 = n131 & n31232 ;
  assign n31234 = n30307 & n75520 ;
  assign n31235 = n31092 & n31234 ;
  assign n31236 = n31233 | n31235 ;
  assign n31237 = n75210 & n31236 ;
  assign n75531 = ~n31064 ;
  assign n31238 = n31063 & n75531 ;
  assign n31239 = n30324 | n31063 ;
  assign n75532 = ~n31239 ;
  assign n31240 = n31214 & n75532 ;
  assign n31241 = n31238 | n31240 ;
  assign n31242 = n131 & n31241 ;
  assign n31243 = n30315 & n75520 ;
  assign n31244 = n31092 & n31243 ;
  assign n31245 = n31242 | n31244 ;
  assign n31246 = n74905 & n31245 ;
  assign n75533 = ~n31213 ;
  assign n31247 = n31058 & n75533 ;
  assign n31059 = n30332 | n31058 ;
  assign n75534 = ~n31059 ;
  assign n31248 = n75534 & n31212 ;
  assign n31249 = n31247 | n31248 ;
  assign n31250 = n131 & n31249 ;
  assign n31251 = n30323 & n75520 ;
  assign n31252 = n31092 & n31251 ;
  assign n31253 = n31250 | n31252 ;
  assign n31254 = n74431 & n31253 ;
  assign n75535 = ~n31053 ;
  assign n31255 = n31052 & n75535 ;
  assign n31256 = n30340 | n31052 ;
  assign n75536 = ~n31256 ;
  assign n31257 = n31210 & n75536 ;
  assign n31258 = n31255 | n31257 ;
  assign n31259 = n131 & n31258 ;
  assign n31260 = n30331 & n75520 ;
  assign n31261 = n31092 & n31260 ;
  assign n31262 = n31259 | n31261 ;
  assign n31263 = n74029 & n31262 ;
  assign n75537 = ~n31209 ;
  assign n31264 = n31048 & n75537 ;
  assign n31265 = n30348 | n31048 ;
  assign n75538 = ~n31265 ;
  assign n31266 = n31044 & n75538 ;
  assign n31267 = n31264 | n31266 ;
  assign n31268 = n131 & n31267 ;
  assign n31269 = n30339 & n75520 ;
  assign n31270 = n31092 & n31269 ;
  assign n31271 = n31268 | n31270 ;
  assign n31272 = n74021 & n31271 ;
  assign n75539 = ~n31043 ;
  assign n31273 = n31042 & n75539 ;
  assign n31274 = n30356 | n31042 ;
  assign n75540 = ~n31274 ;
  assign n31275 = n31206 & n75540 ;
  assign n31276 = n31273 | n31275 ;
  assign n31277 = n131 & n31276 ;
  assign n31278 = n30347 & n75520 ;
  assign n31279 = n31092 & n31278 ;
  assign n31280 = n31277 | n31279 ;
  assign n31281 = n73617 & n31280 ;
  assign n75541 = ~n31205 ;
  assign n31282 = n31038 & n75541 ;
  assign n31283 = n30364 | n31038 ;
  assign n75542 = ~n31283 ;
  assign n31284 = n31034 & n75542 ;
  assign n31285 = n31282 | n31284 ;
  assign n31286 = n131 & n31285 ;
  assign n31287 = n30355 & n75520 ;
  assign n31288 = n31092 & n31287 ;
  assign n31289 = n31286 | n31288 ;
  assign n31290 = n73188 & n31289 ;
  assign n75543 = ~n31033 ;
  assign n31291 = n31032 & n75543 ;
  assign n31292 = n30372 | n31032 ;
  assign n75544 = ~n31292 ;
  assign n31293 = n31202 & n75544 ;
  assign n31294 = n31291 | n31293 ;
  assign n31295 = n131 & n31294 ;
  assign n31296 = n30363 & n75520 ;
  assign n31297 = n31092 & n31296 ;
  assign n31298 = n31295 | n31297 ;
  assign n31299 = n73177 & n31298 ;
  assign n75545 = ~n31201 ;
  assign n31300 = n31028 & n75545 ;
  assign n31301 = n30380 | n31028 ;
  assign n75546 = ~n31301 ;
  assign n31302 = n31024 & n75546 ;
  assign n31303 = n31300 | n31302 ;
  assign n31304 = n131 & n31303 ;
  assign n31305 = n30371 & n75520 ;
  assign n31306 = n31092 & n31305 ;
  assign n31307 = n31304 | n31306 ;
  assign n31308 = n72752 & n31307 ;
  assign n75547 = ~n31023 ;
  assign n31309 = n31022 & n75547 ;
  assign n31310 = n30388 | n31022 ;
  assign n75548 = ~n31310 ;
  assign n31311 = n31198 & n75548 ;
  assign n31312 = n31309 | n31311 ;
  assign n31313 = n131 & n31312 ;
  assign n31314 = n30379 & n75520 ;
  assign n31315 = n31092 & n31314 ;
  assign n31316 = n31313 | n31315 ;
  assign n31317 = n72393 & n31316 ;
  assign n75549 = ~n31197 ;
  assign n31318 = n31017 & n75549 ;
  assign n31018 = n30396 | n31017 ;
  assign n75550 = ~n31018 ;
  assign n31319 = n75550 & n31196 ;
  assign n31320 = n31318 | n31319 ;
  assign n31321 = n131 & n31320 ;
  assign n31322 = n30387 & n75520 ;
  assign n31323 = n31092 & n31322 ;
  assign n31324 = n31321 | n31323 ;
  assign n31325 = n72385 & n31324 ;
  assign n75551 = ~n31012 ;
  assign n31326 = n31011 & n75551 ;
  assign n31327 = n30404 | n31011 ;
  assign n75552 = ~n31327 ;
  assign n31328 = n31194 & n75552 ;
  assign n31329 = n31326 | n31328 ;
  assign n31330 = n131 & n31329 ;
  assign n31331 = n30395 & n75520 ;
  assign n31332 = n31092 & n31331 ;
  assign n31333 = n31330 | n31332 ;
  assign n31334 = n72025 & n31333 ;
  assign n75553 = ~n31193 ;
  assign n31335 = n31006 & n75553 ;
  assign n31007 = n30412 | n31006 ;
  assign n75554 = ~n31007 ;
  assign n31336 = n75554 & n31192 ;
  assign n31337 = n31335 | n31336 ;
  assign n31338 = n131 & n31337 ;
  assign n31339 = n30403 & n75520 ;
  assign n31340 = n31092 & n31339 ;
  assign n31341 = n31338 | n31340 ;
  assign n31342 = n71645 & n31341 ;
  assign n75555 = ~n31001 ;
  assign n31343 = n31000 & n75555 ;
  assign n31344 = n30420 | n31000 ;
  assign n75556 = ~n31344 ;
  assign n31345 = n31190 & n75556 ;
  assign n31346 = n31343 | n31345 ;
  assign n31347 = n131 & n31346 ;
  assign n31348 = n30411 & n75520 ;
  assign n31349 = n31092 & n31348 ;
  assign n31350 = n31347 | n31349 ;
  assign n31351 = n71633 & n31350 ;
  assign n75557 = ~n31189 ;
  assign n31352 = n30996 & n75557 ;
  assign n31353 = n30428 | n30996 ;
  assign n75558 = ~n31353 ;
  assign n31354 = n30992 & n75558 ;
  assign n31355 = n31352 | n31354 ;
  assign n31356 = n131 & n31355 ;
  assign n31357 = n30419 & n75520 ;
  assign n31358 = n31092 & n31357 ;
  assign n31359 = n31356 | n31358 ;
  assign n31360 = n71253 & n31359 ;
  assign n75559 = ~n30991 ;
  assign n31361 = n30990 & n75559 ;
  assign n31362 = n30436 | n30990 ;
  assign n75560 = ~n31362 ;
  assign n31363 = n31186 & n75560 ;
  assign n31364 = n31361 | n31363 ;
  assign n31365 = n131 & n31364 ;
  assign n31366 = n30427 & n75520 ;
  assign n31367 = n31092 & n31366 ;
  assign n31368 = n31365 | n31367 ;
  assign n31369 = n70935 & n31368 ;
  assign n75561 = ~n31185 ;
  assign n31370 = n30986 & n75561 ;
  assign n31371 = n30444 | n30986 ;
  assign n75562 = ~n31371 ;
  assign n31372 = n30982 & n75562 ;
  assign n31373 = n31370 | n31372 ;
  assign n31374 = n131 & n31373 ;
  assign n31375 = n30435 & n75520 ;
  assign n31376 = n31092 & n31375 ;
  assign n31377 = n31374 | n31376 ;
  assign n31378 = n70927 & n31377 ;
  assign n75563 = ~n30981 ;
  assign n31379 = n30980 & n75563 ;
  assign n31380 = n30452 | n30980 ;
  assign n75564 = ~n31380 ;
  assign n31381 = n31182 & n75564 ;
  assign n31382 = n31379 | n31381 ;
  assign n31383 = n131 & n31382 ;
  assign n31384 = n30443 & n75520 ;
  assign n31385 = n31092 & n31384 ;
  assign n31386 = n31383 | n31385 ;
  assign n31387 = n70609 & n31386 ;
  assign n75565 = ~n31181 ;
  assign n31388 = n30976 & n75565 ;
  assign n31389 = n30460 | n30976 ;
  assign n75566 = ~n31389 ;
  assign n31390 = n30972 & n75566 ;
  assign n31391 = n31388 | n31390 ;
  assign n31392 = n131 & n31391 ;
  assign n31393 = n30451 & n75520 ;
  assign n31394 = n31092 & n31393 ;
  assign n31395 = n31392 | n31394 ;
  assign n31396 = n70276 & n31395 ;
  assign n75567 = ~n30971 ;
  assign n31397 = n30970 & n75567 ;
  assign n31398 = n30468 | n30970 ;
  assign n75568 = ~n31398 ;
  assign n31399 = n31178 & n75568 ;
  assign n31400 = n31397 | n31399 ;
  assign n31401 = n131 & n31400 ;
  assign n31402 = n30459 & n75520 ;
  assign n31403 = n31092 & n31402 ;
  assign n31404 = n31401 | n31403 ;
  assign n31405 = n70176 & n31404 ;
  assign n75569 = ~n31177 ;
  assign n31406 = n30966 & n75569 ;
  assign n31407 = n30476 | n30966 ;
  assign n75570 = ~n31407 ;
  assign n31408 = n30962 & n75570 ;
  assign n31409 = n31406 | n31408 ;
  assign n31410 = n131 & n31409 ;
  assign n31411 = n30467 & n75520 ;
  assign n31412 = n31092 & n31411 ;
  assign n31413 = n31410 | n31412 ;
  assign n31414 = n69857 & n31413 ;
  assign n75571 = ~n30961 ;
  assign n31415 = n30960 & n75571 ;
  assign n31416 = n30484 | n30960 ;
  assign n75572 = ~n31416 ;
  assign n31417 = n31174 & n75572 ;
  assign n31418 = n31415 | n31417 ;
  assign n31419 = n131 & n31418 ;
  assign n31420 = n30475 & n75520 ;
  assign n31421 = n31092 & n31420 ;
  assign n31422 = n31419 | n31421 ;
  assign n31423 = n69656 & n31422 ;
  assign n75573 = ~n31173 ;
  assign n31424 = n30956 & n75573 ;
  assign n31425 = n30492 | n30956 ;
  assign n75574 = ~n31425 ;
  assign n31426 = n30952 & n75574 ;
  assign n31427 = n31424 | n31426 ;
  assign n31428 = n131 & n31427 ;
  assign n31429 = n30483 & n75520 ;
  assign n31430 = n31092 & n31429 ;
  assign n31431 = n31428 | n31430 ;
  assign n31432 = n69528 & n31431 ;
  assign n75575 = ~n30951 ;
  assign n31433 = n30950 & n75575 ;
  assign n31434 = n30500 | n30950 ;
  assign n75576 = ~n31434 ;
  assign n31435 = n31170 & n75576 ;
  assign n31436 = n31433 | n31435 ;
  assign n31437 = n131 & n31436 ;
  assign n31438 = n30491 & n75520 ;
  assign n31439 = n31092 & n31438 ;
  assign n31440 = n31437 | n31439 ;
  assign n31441 = n69261 & n31440 ;
  assign n75577 = ~n31169 ;
  assign n31442 = n30946 & n75577 ;
  assign n31443 = n30508 | n30946 ;
  assign n75578 = ~n31443 ;
  assign n31444 = n30942 & n75578 ;
  assign n31445 = n31442 | n31444 ;
  assign n31446 = n131 & n31445 ;
  assign n31447 = n30499 & n75520 ;
  assign n31448 = n31092 & n31447 ;
  assign n31449 = n31446 | n31448 ;
  assign n31450 = n69075 & n31449 ;
  assign n75579 = ~n30941 ;
  assign n31451 = n30940 & n75579 ;
  assign n31452 = n30516 | n30940 ;
  assign n75580 = ~n31452 ;
  assign n31453 = n31166 & n75580 ;
  assign n31454 = n31451 | n31453 ;
  assign n31455 = n131 & n31454 ;
  assign n31456 = n30507 & n75520 ;
  assign n31457 = n31092 & n31456 ;
  assign n31458 = n31455 | n31457 ;
  assign n31459 = n68993 & n31458 ;
  assign n75581 = ~n31165 ;
  assign n31460 = n30936 & n75581 ;
  assign n31461 = n30524 | n30936 ;
  assign n75582 = ~n31461 ;
  assign n31462 = n30932 & n75582 ;
  assign n31463 = n31460 | n31462 ;
  assign n31464 = n131 & n31463 ;
  assign n31465 = n30515 & n75520 ;
  assign n31466 = n31092 & n31465 ;
  assign n31467 = n31464 | n31466 ;
  assign n31468 = n68716 & n31467 ;
  assign n75583 = ~n30931 ;
  assign n31469 = n30930 & n75583 ;
  assign n31470 = n30532 | n30930 ;
  assign n75584 = ~n31470 ;
  assign n31471 = n31162 & n75584 ;
  assign n31472 = n31469 | n31471 ;
  assign n31473 = n131 & n31472 ;
  assign n31474 = n30523 & n75520 ;
  assign n31475 = n31092 & n31474 ;
  assign n31476 = n31473 | n31475 ;
  assign n31477 = n68545 & n31476 ;
  assign n75585 = ~n31161 ;
  assign n31478 = n30926 & n75585 ;
  assign n31479 = n30540 | n30926 ;
  assign n75586 = ~n31479 ;
  assign n31480 = n30922 & n75586 ;
  assign n31481 = n31478 | n31480 ;
  assign n31482 = n131 & n31481 ;
  assign n31483 = n30531 & n75520 ;
  assign n31484 = n31092 & n31483 ;
  assign n31485 = n31482 | n31484 ;
  assign n31486 = n68438 & n31485 ;
  assign n75587 = ~n30921 ;
  assign n31487 = n30920 & n75587 ;
  assign n31488 = n30548 | n30920 ;
  assign n75588 = ~n31488 ;
  assign n31489 = n31158 & n75588 ;
  assign n31490 = n31487 | n31489 ;
  assign n31491 = n131 & n31490 ;
  assign n31492 = n30539 & n75520 ;
  assign n31493 = n31092 & n31492 ;
  assign n31494 = n31491 | n31493 ;
  assign n31495 = n68214 & n31494 ;
  assign n75589 = ~n31157 ;
  assign n31496 = n30916 & n75589 ;
  assign n31497 = n30556 | n30916 ;
  assign n75590 = ~n31497 ;
  assign n31498 = n30912 & n75590 ;
  assign n31499 = n31496 | n31498 ;
  assign n31500 = n131 & n31499 ;
  assign n31501 = n30547 & n75520 ;
  assign n31502 = n31092 & n31501 ;
  assign n31503 = n31500 | n31502 ;
  assign n31504 = n68058 & n31503 ;
  assign n75591 = ~n30911 ;
  assign n31505 = n30910 & n75591 ;
  assign n31506 = n30564 | n30910 ;
  assign n75592 = ~n31506 ;
  assign n31507 = n31154 & n75592 ;
  assign n31508 = n31505 | n31507 ;
  assign n31509 = n131 & n31508 ;
  assign n31510 = n30555 & n75520 ;
  assign n31511 = n31092 & n31510 ;
  assign n31512 = n31509 | n31511 ;
  assign n31513 = n67986 & n31512 ;
  assign n75593 = ~n31153 ;
  assign n31514 = n30906 & n75593 ;
  assign n31515 = n30572 | n30906 ;
  assign n75594 = ~n31515 ;
  assign n31516 = n30902 & n75594 ;
  assign n31517 = n31514 | n31516 ;
  assign n31518 = n131 & n31517 ;
  assign n31519 = n30563 & n75520 ;
  assign n31520 = n31092 & n31519 ;
  assign n31521 = n31518 | n31520 ;
  assign n31522 = n67763 & n31521 ;
  assign n75595 = ~n30901 ;
  assign n31523 = n30900 & n75595 ;
  assign n31524 = n30580 | n30900 ;
  assign n75596 = ~n31524 ;
  assign n31525 = n31150 & n75596 ;
  assign n31526 = n31523 | n31525 ;
  assign n31527 = n131 & n31526 ;
  assign n31528 = n30571 & n75520 ;
  assign n31529 = n31092 & n31528 ;
  assign n31530 = n31527 | n31529 ;
  assign n31531 = n67622 & n31530 ;
  assign n75597 = ~n31149 ;
  assign n31532 = n30896 & n75597 ;
  assign n31533 = n30588 | n30896 ;
  assign n75598 = ~n31533 ;
  assign n31534 = n30892 & n75598 ;
  assign n31535 = n31532 | n31534 ;
  assign n31536 = n131 & n31535 ;
  assign n31537 = n30579 & n75520 ;
  assign n31538 = n31092 & n31537 ;
  assign n31539 = n31536 | n31538 ;
  assign n31540 = n67531 & n31539 ;
  assign n75599 = ~n30891 ;
  assign n31541 = n30890 & n75599 ;
  assign n31542 = n30596 | n30890 ;
  assign n75600 = ~n31542 ;
  assign n31543 = n31146 & n75600 ;
  assign n31544 = n31541 | n31543 ;
  assign n31545 = n131 & n31544 ;
  assign n31546 = n30587 & n75520 ;
  assign n31547 = n31092 & n31546 ;
  assign n31548 = n31545 | n31547 ;
  assign n31549 = n67348 & n31548 ;
  assign n75601 = ~n31145 ;
  assign n31550 = n30886 & n75601 ;
  assign n31551 = n30604 | n30886 ;
  assign n75602 = ~n31551 ;
  assign n31552 = n30882 & n75602 ;
  assign n31553 = n31550 | n31552 ;
  assign n31554 = n131 & n31553 ;
  assign n31555 = n30595 & n75520 ;
  assign n31556 = n31092 & n31555 ;
  assign n31557 = n31554 | n31556 ;
  assign n31558 = n67222 & n31557 ;
  assign n75603 = ~n30881 ;
  assign n31559 = n30880 & n75603 ;
  assign n31560 = n30612 | n30880 ;
  assign n75604 = ~n31560 ;
  assign n31561 = n31142 & n75604 ;
  assign n31562 = n31559 | n31561 ;
  assign n31563 = n131 & n31562 ;
  assign n31564 = n30603 & n75520 ;
  assign n31565 = n31092 & n31564 ;
  assign n31566 = n31563 | n31565 ;
  assign n31567 = n67164 & n31566 ;
  assign n75605 = ~n31141 ;
  assign n31568 = n30876 & n75605 ;
  assign n31569 = n30620 | n30876 ;
  assign n75606 = ~n31569 ;
  assign n31570 = n30872 & n75606 ;
  assign n31571 = n31568 | n31570 ;
  assign n31572 = n131 & n31571 ;
  assign n31573 = n30611 & n75520 ;
  assign n31574 = n31092 & n31573 ;
  assign n31575 = n31572 | n31574 ;
  assign n31576 = n66979 & n31575 ;
  assign n75607 = ~n30871 ;
  assign n31577 = n30870 & n75607 ;
  assign n31578 = n30628 | n30870 ;
  assign n75608 = ~n31578 ;
  assign n31579 = n31138 & n75608 ;
  assign n31580 = n31577 | n31579 ;
  assign n31581 = n131 & n31580 ;
  assign n31582 = n30619 & n75520 ;
  assign n31583 = n31092 & n31582 ;
  assign n31584 = n31581 | n31583 ;
  assign n31585 = n66868 & n31584 ;
  assign n75609 = ~n31137 ;
  assign n31586 = n30866 & n75609 ;
  assign n31587 = n30636 | n30866 ;
  assign n75610 = ~n31587 ;
  assign n31588 = n30862 & n75610 ;
  assign n31589 = n31586 | n31588 ;
  assign n31590 = n131 & n31589 ;
  assign n31591 = n30627 & n75520 ;
  assign n31592 = n31092 & n31591 ;
  assign n31593 = n31590 | n31592 ;
  assign n31594 = n66797 & n31593 ;
  assign n75611 = ~n30861 ;
  assign n31595 = n30860 & n75611 ;
  assign n31596 = n30644 | n30860 ;
  assign n75612 = ~n31596 ;
  assign n31597 = n31134 & n75612 ;
  assign n31598 = n31595 | n31597 ;
  assign n31599 = n131 & n31598 ;
  assign n31600 = n30635 & n75520 ;
  assign n31601 = n31092 & n31600 ;
  assign n31602 = n31599 | n31601 ;
  assign n31603 = n66654 & n31602 ;
  assign n75613 = ~n31133 ;
  assign n31604 = n30856 & n75613 ;
  assign n31605 = n30652 | n30856 ;
  assign n75614 = ~n31605 ;
  assign n31606 = n30852 & n75614 ;
  assign n31607 = n31604 | n31606 ;
  assign n31608 = n131 & n31607 ;
  assign n31609 = n30643 & n75520 ;
  assign n31610 = n31092 & n31609 ;
  assign n31611 = n31608 | n31610 ;
  assign n31612 = n66560 & n31611 ;
  assign n75615 = ~n30851 ;
  assign n31613 = n30850 & n75615 ;
  assign n31614 = n30660 | n30850 ;
  assign n75616 = ~n31614 ;
  assign n31615 = n31130 & n75616 ;
  assign n31616 = n31613 | n31615 ;
  assign n31617 = n131 & n31616 ;
  assign n31618 = n30651 & n75520 ;
  assign n31619 = n31092 & n31618 ;
  assign n31620 = n31617 | n31619 ;
  assign n31621 = n66505 & n31620 ;
  assign n75617 = ~n31129 ;
  assign n31622 = n30846 & n75617 ;
  assign n31623 = n30668 | n30846 ;
  assign n75618 = ~n31623 ;
  assign n31624 = n30842 & n75618 ;
  assign n31625 = n31622 | n31624 ;
  assign n31626 = n131 & n31625 ;
  assign n31627 = n30659 & n75520 ;
  assign n31628 = n31092 & n31627 ;
  assign n31629 = n31626 | n31628 ;
  assign n31630 = n66379 & n31629 ;
  assign n75619 = ~n30841 ;
  assign n31631 = n30839 & n75619 ;
  assign n30840 = n30676 | n30839 ;
  assign n75620 = ~n30840 ;
  assign n31632 = n30836 & n75620 ;
  assign n31633 = n31631 | n31632 ;
  assign n31634 = n131 & n31633 ;
  assign n31635 = n30667 & n75520 ;
  assign n31636 = n31092 & n31635 ;
  assign n31637 = n31634 | n31636 ;
  assign n31638 = n66299 & n31637 ;
  assign n75621 = ~n31125 ;
  assign n31639 = n30835 & n75621 ;
  assign n31640 = n30684 | n30835 ;
  assign n75622 = ~n31640 ;
  assign n31641 = n30831 & n75622 ;
  assign n31642 = n31639 | n31641 ;
  assign n31643 = n131 & n31642 ;
  assign n31644 = n30675 & n75520 ;
  assign n31645 = n31092 & n31644 ;
  assign n31646 = n31643 | n31645 ;
  assign n31647 = n66244 & n31646 ;
  assign n75623 = ~n30830 ;
  assign n31648 = n30829 & n75623 ;
  assign n31649 = n30692 | n30829 ;
  assign n75624 = ~n31649 ;
  assign n31650 = n31122 & n75624 ;
  assign n31651 = n31648 | n31650 ;
  assign n31652 = n131 & n31651 ;
  assign n31653 = n30683 & n75520 ;
  assign n31654 = n31092 & n31653 ;
  assign n31655 = n31652 | n31654 ;
  assign n31656 = n66145 & n31655 ;
  assign n75625 = ~n31121 ;
  assign n31657 = n30825 & n75625 ;
  assign n31658 = n30700 | n30825 ;
  assign n75626 = ~n31658 ;
  assign n31659 = n30821 & n75626 ;
  assign n31660 = n31657 | n31659 ;
  assign n31661 = n131 & n31660 ;
  assign n31662 = n30691 & n75520 ;
  assign n31663 = n31092 & n31662 ;
  assign n31664 = n31661 | n31663 ;
  assign n31665 = n66081 & n31664 ;
  assign n75627 = ~n30820 ;
  assign n31666 = n30819 & n75627 ;
  assign n31667 = n30708 | n30819 ;
  assign n75628 = ~n31667 ;
  assign n31668 = n31118 & n75628 ;
  assign n31669 = n31666 | n31668 ;
  assign n31670 = n131 & n31669 ;
  assign n31671 = n30699 & n75520 ;
  assign n31672 = n31092 & n31671 ;
  assign n31673 = n31670 | n31672 ;
  assign n31674 = n66043 & n31673 ;
  assign n75629 = ~n31117 ;
  assign n31675 = n30815 & n75629 ;
  assign n31676 = n30716 | n30815 ;
  assign n75630 = ~n31676 ;
  assign n31677 = n30811 & n75630 ;
  assign n31678 = n31675 | n31677 ;
  assign n31679 = n131 & n31678 ;
  assign n31680 = n30707 & n75520 ;
  assign n31681 = n31092 & n31680 ;
  assign n31682 = n31679 | n31681 ;
  assign n31683 = n65960 & n31682 ;
  assign n75631 = ~n30810 ;
  assign n31684 = n30809 & n75631 ;
  assign n31685 = n30724 | n30809 ;
  assign n75632 = ~n31685 ;
  assign n31686 = n31114 & n75632 ;
  assign n31687 = n31684 | n31686 ;
  assign n31688 = n131 & n31687 ;
  assign n31689 = n30715 & n75520 ;
  assign n31690 = n31092 & n31689 ;
  assign n31691 = n31688 | n31690 ;
  assign n31692 = n65909 & n31691 ;
  assign n75633 = ~n31113 ;
  assign n31693 = n30805 & n75633 ;
  assign n31694 = n30732 | n30805 ;
  assign n75634 = ~n31694 ;
  assign n31695 = n30801 & n75634 ;
  assign n31696 = n31693 | n31695 ;
  assign n31697 = n131 & n31696 ;
  assign n31698 = n30723 & n75520 ;
  assign n31699 = n31092 & n31698 ;
  assign n31700 = n31697 | n31699 ;
  assign n31701 = n65877 & n31700 ;
  assign n75635 = ~n30800 ;
  assign n31702 = n30799 & n75635 ;
  assign n31703 = n30740 | n30799 ;
  assign n75636 = ~n31703 ;
  assign n31704 = n31110 & n75636 ;
  assign n31705 = n31702 | n31704 ;
  assign n31706 = n131 & n31705 ;
  assign n31707 = n30731 & n75520 ;
  assign n31708 = n31092 & n31707 ;
  assign n31709 = n31706 | n31708 ;
  assign n31710 = n65820 & n31709 ;
  assign n75637 = ~n31109 ;
  assign n31711 = n30795 & n75637 ;
  assign n31712 = n30748 | n30795 ;
  assign n75638 = ~n31712 ;
  assign n31713 = n30791 & n75638 ;
  assign n31714 = n31711 | n31713 ;
  assign n31715 = n131 & n31714 ;
  assign n31716 = n30739 & n75520 ;
  assign n31717 = n31092 & n31716 ;
  assign n31718 = n31715 | n31717 ;
  assign n31719 = n65791 & n31718 ;
  assign n75639 = ~n30790 ;
  assign n31721 = n30789 & n75639 ;
  assign n31720 = n30757 | n30789 ;
  assign n75640 = ~n31720 ;
  assign n31722 = n30786 & n75640 ;
  assign n31723 = n31721 | n31722 ;
  assign n31724 = n131 & n31723 ;
  assign n31725 = n30747 & n75520 ;
  assign n31726 = n31092 & n31725 ;
  assign n31727 = n31724 | n31726 ;
  assign n31728 = n65772 & n31727 ;
  assign n75641 = ~n31105 ;
  assign n31730 = n30785 & n75641 ;
  assign n31729 = n30765 | n30785 ;
  assign n75642 = ~n31729 ;
  assign n31731 = n31104 & n75642 ;
  assign n31732 = n31730 | n31731 ;
  assign n31733 = n131 & n31732 ;
  assign n31734 = n30756 & n75520 ;
  assign n31735 = n31092 & n31734 ;
  assign n31736 = n31733 | n31735 ;
  assign n31737 = n65746 & n31736 ;
  assign n75643 = ~n30780 ;
  assign n31738 = n30779 & n75643 ;
  assign n31103 = n30776 | n30779 ;
  assign n75644 = ~n31103 ;
  assign n31739 = n30775 & n75644 ;
  assign n31740 = n31738 | n31739 ;
  assign n31741 = n131 & n31740 ;
  assign n31742 = n30764 & n75520 ;
  assign n31743 = n31092 & n31742 ;
  assign n31744 = n31741 | n31743 ;
  assign n31745 = n65721 & n31744 ;
  assign n31746 = n30772 & n30774 ;
  assign n31747 = n75395 & n31746 ;
  assign n75645 = ~n31747 ;
  assign n31748 = n30775 & n75645 ;
  assign n31749 = n131 & n31748 ;
  assign n31750 = n30767 & n75520 ;
  assign n31751 = n31092 & n31750 ;
  assign n31752 = n31749 | n31751 ;
  assign n31753 = n65686 & n31752 ;
  assign n31095 = n30774 & n131 ;
  assign n31756 = n31091 | n31755 ;
  assign n31757 = n75520 & n31756 ;
  assign n75646 = ~n31757 ;
  assign n31758 = x64 & n75646 ;
  assign n75647 = ~n31758 ;
  assign n31759 = x2 & n75647 ;
  assign n31760 = n31095 | n31759 ;
  assign n31761 = n65670 & n31760 ;
  assign n31763 = x64 & n131 ;
  assign n75648 = ~n31763 ;
  assign n31764 = x2 & n75648 ;
  assign n31765 = n31095 | n31764 ;
  assign n31767 = x65 & n31765 ;
  assign n31766 = x65 | n31095 ;
  assign n31768 = n31759 | n31766 ;
  assign n75649 = ~n31767 ;
  assign n31769 = n75649 & n31768 ;
  assign n75650 = ~x1 ;
  assign n31770 = n75650 & x64 ;
  assign n31771 = n31769 | n31770 ;
  assign n75651 = ~n31761 ;
  assign n31772 = n75651 & n31771 ;
  assign n75652 = ~n31751 ;
  assign n31773 = x66 & n75652 ;
  assign n75653 = ~n31749 ;
  assign n31774 = n75653 & n31773 ;
  assign n31775 = n31753 | n31774 ;
  assign n31776 = n31772 | n31775 ;
  assign n75654 = ~n31753 ;
  assign n31777 = n75654 & n31776 ;
  assign n75655 = ~n31743 ;
  assign n31778 = x67 & n75655 ;
  assign n75656 = ~n31741 ;
  assign n31779 = n75656 & n31778 ;
  assign n31780 = n31745 | n31779 ;
  assign n31781 = n31777 | n31780 ;
  assign n75657 = ~n31745 ;
  assign n31782 = n75657 & n31781 ;
  assign n75658 = ~n31735 ;
  assign n31783 = x68 & n75658 ;
  assign n75659 = ~n31733 ;
  assign n31784 = n75659 & n31783 ;
  assign n31785 = n31737 | n31784 ;
  assign n31786 = n31782 | n31785 ;
  assign n75660 = ~n31737 ;
  assign n31787 = n75660 & n31786 ;
  assign n75661 = ~n31726 ;
  assign n31788 = x69 & n75661 ;
  assign n75662 = ~n31724 ;
  assign n31789 = n75662 & n31788 ;
  assign n31790 = n31728 | n31789 ;
  assign n31792 = n31787 | n31790 ;
  assign n75663 = ~n31728 ;
  assign n31793 = n75663 & n31792 ;
  assign n75664 = ~n31717 ;
  assign n31794 = x70 & n75664 ;
  assign n75665 = ~n31715 ;
  assign n31795 = n75665 & n31794 ;
  assign n31796 = n31719 | n31795 ;
  assign n31797 = n31793 | n31796 ;
  assign n75666 = ~n31719 ;
  assign n31798 = n75666 & n31797 ;
  assign n75667 = ~n31708 ;
  assign n31799 = x71 & n75667 ;
  assign n75668 = ~n31706 ;
  assign n31800 = n75668 & n31799 ;
  assign n31801 = n31710 | n31800 ;
  assign n31803 = n31798 | n31801 ;
  assign n75669 = ~n31710 ;
  assign n31804 = n75669 & n31803 ;
  assign n75670 = ~n31699 ;
  assign n31805 = x72 & n75670 ;
  assign n75671 = ~n31697 ;
  assign n31806 = n75671 & n31805 ;
  assign n31807 = n31701 | n31806 ;
  assign n31808 = n31804 | n31807 ;
  assign n75672 = ~n31701 ;
  assign n31809 = n75672 & n31808 ;
  assign n75673 = ~n31690 ;
  assign n31810 = x73 & n75673 ;
  assign n75674 = ~n31688 ;
  assign n31811 = n75674 & n31810 ;
  assign n31812 = n31692 | n31811 ;
  assign n31814 = n31809 | n31812 ;
  assign n75675 = ~n31692 ;
  assign n31815 = n75675 & n31814 ;
  assign n75676 = ~n31681 ;
  assign n31816 = x74 & n75676 ;
  assign n75677 = ~n31679 ;
  assign n31817 = n75677 & n31816 ;
  assign n31818 = n31683 | n31817 ;
  assign n31819 = n31815 | n31818 ;
  assign n75678 = ~n31683 ;
  assign n31820 = n75678 & n31819 ;
  assign n75679 = ~n31672 ;
  assign n31821 = x75 & n75679 ;
  assign n75680 = ~n31670 ;
  assign n31822 = n75680 & n31821 ;
  assign n31823 = n31674 | n31822 ;
  assign n31825 = n31820 | n31823 ;
  assign n75681 = ~n31674 ;
  assign n31826 = n75681 & n31825 ;
  assign n75682 = ~n31663 ;
  assign n31827 = x76 & n75682 ;
  assign n75683 = ~n31661 ;
  assign n31828 = n75683 & n31827 ;
  assign n31829 = n31665 | n31828 ;
  assign n31830 = n31826 | n31829 ;
  assign n75684 = ~n31665 ;
  assign n31831 = n75684 & n31830 ;
  assign n75685 = ~n31654 ;
  assign n31832 = x77 & n75685 ;
  assign n75686 = ~n31652 ;
  assign n31833 = n75686 & n31832 ;
  assign n31834 = n31656 | n31833 ;
  assign n31836 = n31831 | n31834 ;
  assign n75687 = ~n31656 ;
  assign n31837 = n75687 & n31836 ;
  assign n75688 = ~n31645 ;
  assign n31838 = x78 & n75688 ;
  assign n75689 = ~n31643 ;
  assign n31839 = n75689 & n31838 ;
  assign n31840 = n31647 | n31839 ;
  assign n31841 = n31837 | n31840 ;
  assign n75690 = ~n31647 ;
  assign n31842 = n75690 & n31841 ;
  assign n75691 = ~n31636 ;
  assign n31843 = x79 & n75691 ;
  assign n75692 = ~n31634 ;
  assign n31844 = n75692 & n31843 ;
  assign n31845 = n31638 | n31844 ;
  assign n31847 = n31842 | n31845 ;
  assign n75693 = ~n31638 ;
  assign n31848 = n75693 & n31847 ;
  assign n75694 = ~n31628 ;
  assign n31849 = x80 & n75694 ;
  assign n75695 = ~n31626 ;
  assign n31850 = n75695 & n31849 ;
  assign n31851 = n31630 | n31850 ;
  assign n31852 = n31848 | n31851 ;
  assign n75696 = ~n31630 ;
  assign n31853 = n75696 & n31852 ;
  assign n75697 = ~n31619 ;
  assign n31854 = x81 & n75697 ;
  assign n75698 = ~n31617 ;
  assign n31855 = n75698 & n31854 ;
  assign n31856 = n31621 | n31855 ;
  assign n31858 = n31853 | n31856 ;
  assign n75699 = ~n31621 ;
  assign n31859 = n75699 & n31858 ;
  assign n75700 = ~n31610 ;
  assign n31860 = x82 & n75700 ;
  assign n75701 = ~n31608 ;
  assign n31861 = n75701 & n31860 ;
  assign n31862 = n31612 | n31861 ;
  assign n31863 = n31859 | n31862 ;
  assign n75702 = ~n31612 ;
  assign n31864 = n75702 & n31863 ;
  assign n75703 = ~n31601 ;
  assign n31865 = x83 & n75703 ;
  assign n75704 = ~n31599 ;
  assign n31866 = n75704 & n31865 ;
  assign n31867 = n31603 | n31866 ;
  assign n31869 = n31864 | n31867 ;
  assign n75705 = ~n31603 ;
  assign n31870 = n75705 & n31869 ;
  assign n75706 = ~n31592 ;
  assign n31871 = x84 & n75706 ;
  assign n75707 = ~n31590 ;
  assign n31872 = n75707 & n31871 ;
  assign n31873 = n31594 | n31872 ;
  assign n31874 = n31870 | n31873 ;
  assign n75708 = ~n31594 ;
  assign n31875 = n75708 & n31874 ;
  assign n75709 = ~n31583 ;
  assign n31876 = x85 & n75709 ;
  assign n75710 = ~n31581 ;
  assign n31877 = n75710 & n31876 ;
  assign n31878 = n31585 | n31877 ;
  assign n31880 = n31875 | n31878 ;
  assign n75711 = ~n31585 ;
  assign n31881 = n75711 & n31880 ;
  assign n75712 = ~n31574 ;
  assign n31882 = x86 & n75712 ;
  assign n75713 = ~n31572 ;
  assign n31883 = n75713 & n31882 ;
  assign n31884 = n31576 | n31883 ;
  assign n31885 = n31881 | n31884 ;
  assign n75714 = ~n31576 ;
  assign n31886 = n75714 & n31885 ;
  assign n75715 = ~n31565 ;
  assign n31887 = x87 & n75715 ;
  assign n75716 = ~n31563 ;
  assign n31888 = n75716 & n31887 ;
  assign n31889 = n31567 | n31888 ;
  assign n31891 = n31886 | n31889 ;
  assign n75717 = ~n31567 ;
  assign n31892 = n75717 & n31891 ;
  assign n75718 = ~n31556 ;
  assign n31893 = x88 & n75718 ;
  assign n75719 = ~n31554 ;
  assign n31894 = n75719 & n31893 ;
  assign n31895 = n31558 | n31894 ;
  assign n31896 = n31892 | n31895 ;
  assign n75720 = ~n31558 ;
  assign n31897 = n75720 & n31896 ;
  assign n75721 = ~n31547 ;
  assign n31898 = x89 & n75721 ;
  assign n75722 = ~n31545 ;
  assign n31899 = n75722 & n31898 ;
  assign n31900 = n31549 | n31899 ;
  assign n31902 = n31897 | n31900 ;
  assign n75723 = ~n31549 ;
  assign n31903 = n75723 & n31902 ;
  assign n75724 = ~n31538 ;
  assign n31904 = x90 & n75724 ;
  assign n75725 = ~n31536 ;
  assign n31905 = n75725 & n31904 ;
  assign n31906 = n31540 | n31905 ;
  assign n31907 = n31903 | n31906 ;
  assign n75726 = ~n31540 ;
  assign n31908 = n75726 & n31907 ;
  assign n75727 = ~n31529 ;
  assign n31909 = x91 & n75727 ;
  assign n75728 = ~n31527 ;
  assign n31910 = n75728 & n31909 ;
  assign n31911 = n31531 | n31910 ;
  assign n31913 = n31908 | n31911 ;
  assign n75729 = ~n31531 ;
  assign n31914 = n75729 & n31913 ;
  assign n75730 = ~n31520 ;
  assign n31915 = x92 & n75730 ;
  assign n75731 = ~n31518 ;
  assign n31916 = n75731 & n31915 ;
  assign n31917 = n31522 | n31916 ;
  assign n31918 = n31914 | n31917 ;
  assign n75732 = ~n31522 ;
  assign n31919 = n75732 & n31918 ;
  assign n75733 = ~n31511 ;
  assign n31920 = x93 & n75733 ;
  assign n75734 = ~n31509 ;
  assign n31921 = n75734 & n31920 ;
  assign n31922 = n31513 | n31921 ;
  assign n31924 = n31919 | n31922 ;
  assign n75735 = ~n31513 ;
  assign n31925 = n75735 & n31924 ;
  assign n75736 = ~n31502 ;
  assign n31926 = x94 & n75736 ;
  assign n75737 = ~n31500 ;
  assign n31927 = n75737 & n31926 ;
  assign n31928 = n31504 | n31927 ;
  assign n31929 = n31925 | n31928 ;
  assign n75738 = ~n31504 ;
  assign n31930 = n75738 & n31929 ;
  assign n75739 = ~n31493 ;
  assign n31931 = x95 & n75739 ;
  assign n75740 = ~n31491 ;
  assign n31932 = n75740 & n31931 ;
  assign n31933 = n31495 | n31932 ;
  assign n31935 = n31930 | n31933 ;
  assign n75741 = ~n31495 ;
  assign n31936 = n75741 & n31935 ;
  assign n75742 = ~n31484 ;
  assign n31937 = x96 & n75742 ;
  assign n75743 = ~n31482 ;
  assign n31938 = n75743 & n31937 ;
  assign n31939 = n31486 | n31938 ;
  assign n31940 = n31936 | n31939 ;
  assign n75744 = ~n31486 ;
  assign n31941 = n75744 & n31940 ;
  assign n75745 = ~n31475 ;
  assign n31942 = x97 & n75745 ;
  assign n75746 = ~n31473 ;
  assign n31943 = n75746 & n31942 ;
  assign n31944 = n31477 | n31943 ;
  assign n31946 = n31941 | n31944 ;
  assign n75747 = ~n31477 ;
  assign n31947 = n75747 & n31946 ;
  assign n75748 = ~n31466 ;
  assign n31948 = x98 & n75748 ;
  assign n75749 = ~n31464 ;
  assign n31949 = n75749 & n31948 ;
  assign n31950 = n31468 | n31949 ;
  assign n31951 = n31947 | n31950 ;
  assign n75750 = ~n31468 ;
  assign n31952 = n75750 & n31951 ;
  assign n75751 = ~n31457 ;
  assign n31953 = x99 & n75751 ;
  assign n75752 = ~n31455 ;
  assign n31954 = n75752 & n31953 ;
  assign n31955 = n31459 | n31954 ;
  assign n31957 = n31952 | n31955 ;
  assign n75753 = ~n31459 ;
  assign n31958 = n75753 & n31957 ;
  assign n75754 = ~n31448 ;
  assign n31959 = x100 & n75754 ;
  assign n75755 = ~n31446 ;
  assign n31960 = n75755 & n31959 ;
  assign n31961 = n31450 | n31960 ;
  assign n31962 = n31958 | n31961 ;
  assign n75756 = ~n31450 ;
  assign n31963 = n75756 & n31962 ;
  assign n75757 = ~n31439 ;
  assign n31964 = x101 & n75757 ;
  assign n75758 = ~n31437 ;
  assign n31965 = n75758 & n31964 ;
  assign n31966 = n31441 | n31965 ;
  assign n31968 = n31963 | n31966 ;
  assign n75759 = ~n31441 ;
  assign n31969 = n75759 & n31968 ;
  assign n75760 = ~n31430 ;
  assign n31970 = x102 & n75760 ;
  assign n75761 = ~n31428 ;
  assign n31971 = n75761 & n31970 ;
  assign n31972 = n31432 | n31971 ;
  assign n31973 = n31969 | n31972 ;
  assign n75762 = ~n31432 ;
  assign n31974 = n75762 & n31973 ;
  assign n75763 = ~n31421 ;
  assign n31975 = x103 & n75763 ;
  assign n75764 = ~n31419 ;
  assign n31976 = n75764 & n31975 ;
  assign n31977 = n31423 | n31976 ;
  assign n31979 = n31974 | n31977 ;
  assign n75765 = ~n31423 ;
  assign n31980 = n75765 & n31979 ;
  assign n75766 = ~n31412 ;
  assign n31981 = x104 & n75766 ;
  assign n75767 = ~n31410 ;
  assign n31982 = n75767 & n31981 ;
  assign n31983 = n31414 | n31982 ;
  assign n31984 = n31980 | n31983 ;
  assign n75768 = ~n31414 ;
  assign n31985 = n75768 & n31984 ;
  assign n75769 = ~n31403 ;
  assign n31986 = x105 & n75769 ;
  assign n75770 = ~n31401 ;
  assign n31987 = n75770 & n31986 ;
  assign n31988 = n31405 | n31987 ;
  assign n31990 = n31985 | n31988 ;
  assign n75771 = ~n31405 ;
  assign n31991 = n75771 & n31990 ;
  assign n75772 = ~n31394 ;
  assign n31992 = x106 & n75772 ;
  assign n75773 = ~n31392 ;
  assign n31993 = n75773 & n31992 ;
  assign n31994 = n31396 | n31993 ;
  assign n31995 = n31991 | n31994 ;
  assign n75774 = ~n31396 ;
  assign n31996 = n75774 & n31995 ;
  assign n75775 = ~n31385 ;
  assign n31997 = x107 & n75775 ;
  assign n75776 = ~n31383 ;
  assign n31998 = n75776 & n31997 ;
  assign n31999 = n31387 | n31998 ;
  assign n32001 = n31996 | n31999 ;
  assign n75777 = ~n31387 ;
  assign n32002 = n75777 & n32001 ;
  assign n75778 = ~n31376 ;
  assign n32003 = x108 & n75778 ;
  assign n75779 = ~n31374 ;
  assign n32004 = n75779 & n32003 ;
  assign n32005 = n31378 | n32004 ;
  assign n32006 = n32002 | n32005 ;
  assign n75780 = ~n31378 ;
  assign n32007 = n75780 & n32006 ;
  assign n75781 = ~n31367 ;
  assign n32008 = x109 & n75781 ;
  assign n75782 = ~n31365 ;
  assign n32009 = n75782 & n32008 ;
  assign n32010 = n31369 | n32009 ;
  assign n32012 = n32007 | n32010 ;
  assign n75783 = ~n31369 ;
  assign n32013 = n75783 & n32012 ;
  assign n75784 = ~n31358 ;
  assign n32014 = x110 & n75784 ;
  assign n75785 = ~n31356 ;
  assign n32015 = n75785 & n32014 ;
  assign n32016 = n31360 | n32015 ;
  assign n32017 = n32013 | n32016 ;
  assign n75786 = ~n31360 ;
  assign n32018 = n75786 & n32017 ;
  assign n75787 = ~n31349 ;
  assign n32019 = x111 & n75787 ;
  assign n75788 = ~n31347 ;
  assign n32020 = n75788 & n32019 ;
  assign n32021 = n31351 | n32020 ;
  assign n32023 = n32018 | n32021 ;
  assign n75789 = ~n31351 ;
  assign n32024 = n75789 & n32023 ;
  assign n75790 = ~n31340 ;
  assign n32025 = x112 & n75790 ;
  assign n75791 = ~n31338 ;
  assign n32026 = n75791 & n32025 ;
  assign n32027 = n31342 | n32026 ;
  assign n32028 = n32024 | n32027 ;
  assign n75792 = ~n31342 ;
  assign n32029 = n75792 & n32028 ;
  assign n75793 = ~n31332 ;
  assign n32030 = x113 & n75793 ;
  assign n75794 = ~n31330 ;
  assign n32031 = n75794 & n32030 ;
  assign n32032 = n31334 | n32031 ;
  assign n32034 = n32029 | n32032 ;
  assign n75795 = ~n31334 ;
  assign n32035 = n75795 & n32034 ;
  assign n75796 = ~n31323 ;
  assign n32036 = x114 & n75796 ;
  assign n75797 = ~n31321 ;
  assign n32037 = n75797 & n32036 ;
  assign n32038 = n31325 | n32037 ;
  assign n32039 = n32035 | n32038 ;
  assign n75798 = ~n31325 ;
  assign n32040 = n75798 & n32039 ;
  assign n75799 = ~n31315 ;
  assign n32041 = x115 & n75799 ;
  assign n75800 = ~n31313 ;
  assign n32042 = n75800 & n32041 ;
  assign n32043 = n31317 | n32042 ;
  assign n32045 = n32040 | n32043 ;
  assign n75801 = ~n31317 ;
  assign n32046 = n75801 & n32045 ;
  assign n75802 = ~n31306 ;
  assign n32047 = x116 & n75802 ;
  assign n75803 = ~n31304 ;
  assign n32048 = n75803 & n32047 ;
  assign n32049 = n31308 | n32048 ;
  assign n32050 = n32046 | n32049 ;
  assign n75804 = ~n31308 ;
  assign n32051 = n75804 & n32050 ;
  assign n75805 = ~n31297 ;
  assign n32052 = x117 & n75805 ;
  assign n75806 = ~n31295 ;
  assign n32053 = n75806 & n32052 ;
  assign n32054 = n31299 | n32053 ;
  assign n32056 = n32051 | n32054 ;
  assign n75807 = ~n31299 ;
  assign n32057 = n75807 & n32056 ;
  assign n75808 = ~n31288 ;
  assign n32058 = x118 & n75808 ;
  assign n75809 = ~n31286 ;
  assign n32059 = n75809 & n32058 ;
  assign n32060 = n31290 | n32059 ;
  assign n32061 = n32057 | n32060 ;
  assign n75810 = ~n31290 ;
  assign n32062 = n75810 & n32061 ;
  assign n75811 = ~n31279 ;
  assign n32063 = x119 & n75811 ;
  assign n75812 = ~n31277 ;
  assign n32064 = n75812 & n32063 ;
  assign n32065 = n31281 | n32064 ;
  assign n32067 = n32062 | n32065 ;
  assign n75813 = ~n31281 ;
  assign n32068 = n75813 & n32067 ;
  assign n75814 = ~n31270 ;
  assign n32069 = x120 & n75814 ;
  assign n75815 = ~n31268 ;
  assign n32070 = n75815 & n32069 ;
  assign n32071 = n31272 | n32070 ;
  assign n32072 = n32068 | n32071 ;
  assign n75816 = ~n31272 ;
  assign n32073 = n75816 & n32072 ;
  assign n75817 = ~n31261 ;
  assign n32074 = x121 & n75817 ;
  assign n75818 = ~n31259 ;
  assign n32075 = n75818 & n32074 ;
  assign n32076 = n31263 | n32075 ;
  assign n32078 = n32073 | n32076 ;
  assign n75819 = ~n31263 ;
  assign n32079 = n75819 & n32078 ;
  assign n75820 = ~n31252 ;
  assign n32080 = x122 & n75820 ;
  assign n75821 = ~n31250 ;
  assign n32081 = n75821 & n32080 ;
  assign n32082 = n31254 | n32081 ;
  assign n32083 = n32079 | n32082 ;
  assign n75822 = ~n31254 ;
  assign n32084 = n75822 & n32083 ;
  assign n75823 = ~n31244 ;
  assign n32085 = x123 & n75823 ;
  assign n75824 = ~n31242 ;
  assign n32086 = n75824 & n32085 ;
  assign n32087 = n31246 | n32086 ;
  assign n32089 = n32084 | n32087 ;
  assign n75825 = ~n31246 ;
  assign n32090 = n75825 & n32089 ;
  assign n75826 = ~n31235 ;
  assign n32091 = x124 & n75826 ;
  assign n75827 = ~n31233 ;
  assign n32092 = n75827 & n32091 ;
  assign n32093 = n31237 | n32092 ;
  assign n32095 = n32090 | n32093 ;
  assign n75828 = ~n31237 ;
  assign n32096 = n75828 & n32095 ;
  assign n75829 = ~n31226 ;
  assign n32097 = x125 & n75829 ;
  assign n75830 = ~n31224 ;
  assign n32098 = n75830 & n32097 ;
  assign n32099 = n31228 | n32098 ;
  assign n32101 = n32096 | n32099 ;
  assign n75831 = ~n31228 ;
  assign n32102 = n75831 & n32101 ;
  assign n75832 = ~x126 ;
  assign n32113 = n75832 & n32112 ;
  assign n75833 = ~n32111 ;
  assign n32114 = x126 & n75833 ;
  assign n75834 = ~n32109 ;
  assign n32115 = n75834 & n32114 ;
  assign n32116 = x127 | n32115 ;
  assign n32117 = n32113 | n32116 ;
  assign n32119 = n32102 | n32117 ;
  assign n75835 = ~n32118 ;
  assign n32120 = n75835 & n32119 ;
  assign n75836 = ~n32090 ;
  assign n32123 = n75836 & n32093 ;
  assign n32094 = n31246 | n32093 ;
  assign n75837 = ~n32094 ;
  assign n32124 = n32089 & n75837 ;
  assign n32125 = n32123 | n32124 ;
  assign n130 = ~n32120 ;
  assign n32126 = n130 & n32125 ;
  assign n32127 = n31236 & n75835 ;
  assign n32128 = n32119 & n32127 ;
  assign n32129 = n32126 | n32128 ;
  assign n32131 = n65670 & n31765 ;
  assign n31762 = x65 & n31760 ;
  assign n75839 = ~n31762 ;
  assign n32130 = n75839 & n31768 ;
  assign n32132 = n31770 | n32130 ;
  assign n75840 = ~n32131 ;
  assign n32133 = n75840 & n32132 ;
  assign n32135 = n31775 | n32133 ;
  assign n32136 = n75654 & n32135 ;
  assign n32138 = n31780 | n32136 ;
  assign n32139 = n75657 & n32138 ;
  assign n32141 = n31785 | n32139 ;
  assign n32142 = n75660 & n32141 ;
  assign n32143 = n31790 | n32142 ;
  assign n32144 = n75663 & n32143 ;
  assign n32145 = n31796 | n32144 ;
  assign n32147 = n75666 & n32145 ;
  assign n32148 = n31801 | n32147 ;
  assign n32149 = n75669 & n32148 ;
  assign n32150 = n31807 | n32149 ;
  assign n32152 = n75672 & n32150 ;
  assign n32153 = n31812 | n32152 ;
  assign n32154 = n75675 & n32153 ;
  assign n32155 = n31818 | n32154 ;
  assign n32157 = n75678 & n32155 ;
  assign n32158 = n31823 | n32157 ;
  assign n32159 = n75681 & n32158 ;
  assign n32160 = n31829 | n32159 ;
  assign n32162 = n75684 & n32160 ;
  assign n32163 = n31834 | n32162 ;
  assign n32164 = n75687 & n32163 ;
  assign n32165 = n31840 | n32164 ;
  assign n32167 = n75690 & n32165 ;
  assign n32168 = n31845 | n32167 ;
  assign n32169 = n75693 & n32168 ;
  assign n32170 = n31851 | n32169 ;
  assign n32172 = n75696 & n32170 ;
  assign n32173 = n31856 | n32172 ;
  assign n32174 = n75699 & n32173 ;
  assign n32175 = n31862 | n32174 ;
  assign n32177 = n75702 & n32175 ;
  assign n32178 = n31867 | n32177 ;
  assign n32179 = n75705 & n32178 ;
  assign n32180 = n31873 | n32179 ;
  assign n32182 = n75708 & n32180 ;
  assign n32183 = n31878 | n32182 ;
  assign n32184 = n75711 & n32183 ;
  assign n32185 = n31884 | n32184 ;
  assign n32187 = n75714 & n32185 ;
  assign n32188 = n31889 | n32187 ;
  assign n32189 = n75717 & n32188 ;
  assign n32190 = n31895 | n32189 ;
  assign n32192 = n75720 & n32190 ;
  assign n32193 = n31900 | n32192 ;
  assign n32194 = n75723 & n32193 ;
  assign n32195 = n31906 | n32194 ;
  assign n32197 = n75726 & n32195 ;
  assign n32198 = n31911 | n32197 ;
  assign n32199 = n75729 & n32198 ;
  assign n32200 = n31917 | n32199 ;
  assign n32202 = n75732 & n32200 ;
  assign n32203 = n31922 | n32202 ;
  assign n32204 = n75735 & n32203 ;
  assign n32205 = n31928 | n32204 ;
  assign n32207 = n75738 & n32205 ;
  assign n32208 = n31933 | n32207 ;
  assign n32209 = n75741 & n32208 ;
  assign n32210 = n31939 | n32209 ;
  assign n32212 = n75744 & n32210 ;
  assign n32213 = n31944 | n32212 ;
  assign n32214 = n75747 & n32213 ;
  assign n32215 = n31950 | n32214 ;
  assign n32217 = n75750 & n32215 ;
  assign n32218 = n31955 | n32217 ;
  assign n32219 = n75753 & n32218 ;
  assign n32220 = n31961 | n32219 ;
  assign n32222 = n75756 & n32220 ;
  assign n32223 = n31966 | n32222 ;
  assign n32224 = n75759 & n32223 ;
  assign n32225 = n31972 | n32224 ;
  assign n32227 = n75762 & n32225 ;
  assign n32228 = n31977 | n32227 ;
  assign n32229 = n75765 & n32228 ;
  assign n32230 = n31983 | n32229 ;
  assign n32232 = n75768 & n32230 ;
  assign n32233 = n31988 | n32232 ;
  assign n32234 = n75771 & n32233 ;
  assign n32235 = n31994 | n32234 ;
  assign n32237 = n75774 & n32235 ;
  assign n32238 = n31999 | n32237 ;
  assign n32239 = n75777 & n32238 ;
  assign n32240 = n32005 | n32239 ;
  assign n32242 = n75780 & n32240 ;
  assign n32243 = n32010 | n32242 ;
  assign n32244 = n75783 & n32243 ;
  assign n32245 = n32016 | n32244 ;
  assign n32247 = n75786 & n32245 ;
  assign n32248 = n32021 | n32247 ;
  assign n32249 = n75789 & n32248 ;
  assign n32250 = n32027 | n32249 ;
  assign n32252 = n75792 & n32250 ;
  assign n32253 = n32032 | n32252 ;
  assign n32254 = n75795 & n32253 ;
  assign n32255 = n32038 | n32254 ;
  assign n32257 = n75798 & n32255 ;
  assign n32258 = n32043 | n32257 ;
  assign n32259 = n75801 & n32258 ;
  assign n32260 = n32049 | n32259 ;
  assign n32262 = n75804 & n32260 ;
  assign n32263 = n32054 | n32262 ;
  assign n32264 = n75807 & n32263 ;
  assign n32265 = n32060 | n32264 ;
  assign n32267 = n75810 & n32265 ;
  assign n32268 = n32065 | n32267 ;
  assign n32269 = n75813 & n32268 ;
  assign n32270 = n32071 | n32269 ;
  assign n32272 = n75816 & n32270 ;
  assign n32273 = n32076 | n32272 ;
  assign n32274 = n75819 & n32273 ;
  assign n75841 = ~n32274 ;
  assign n32275 = n32082 & n75841 ;
  assign n32277 = n31263 | n32082 ;
  assign n75842 = ~n32277 ;
  assign n32278 = n32078 & n75842 ;
  assign n32279 = n32275 | n32278 ;
  assign n32280 = n130 & n32279 ;
  assign n32281 = n31253 & n75835 ;
  assign n32282 = n32119 & n32281 ;
  assign n32283 = n32280 | n32282 ;
  assign n75843 = ~n32269 ;
  assign n32271 = n32071 & n75843 ;
  assign n32284 = n31281 | n32071 ;
  assign n75844 = ~n32284 ;
  assign n32285 = n32067 & n75844 ;
  assign n32286 = n32271 | n32285 ;
  assign n32287 = n130 & n32286 ;
  assign n32288 = n31271 & n75835 ;
  assign n32289 = n32119 & n32288 ;
  assign n32290 = n32287 | n32289 ;
  assign n75845 = ~n32264 ;
  assign n32266 = n32060 & n75845 ;
  assign n32291 = n31299 | n32060 ;
  assign n75846 = ~n32291 ;
  assign n32292 = n32056 & n75846 ;
  assign n32293 = n32266 | n32292 ;
  assign n32294 = n130 & n32293 ;
  assign n32295 = n31289 & n75835 ;
  assign n32296 = n32119 & n32295 ;
  assign n32297 = n32294 | n32296 ;
  assign n75847 = ~n32259 ;
  assign n32261 = n32049 & n75847 ;
  assign n32298 = n31317 | n32049 ;
  assign n75848 = ~n32298 ;
  assign n32299 = n32045 & n75848 ;
  assign n32300 = n32261 | n32299 ;
  assign n32301 = n130 & n32300 ;
  assign n32302 = n31307 & n75835 ;
  assign n32303 = n32119 & n32302 ;
  assign n32304 = n32301 | n32303 ;
  assign n75849 = ~n32254 ;
  assign n32256 = n32038 & n75849 ;
  assign n32305 = n31334 | n32038 ;
  assign n75850 = ~n32305 ;
  assign n32306 = n32034 & n75850 ;
  assign n32307 = n32256 | n32306 ;
  assign n32308 = n130 & n32307 ;
  assign n32309 = n31324 & n75835 ;
  assign n32310 = n32119 & n32309 ;
  assign n32311 = n32308 | n32310 ;
  assign n75851 = ~n32249 ;
  assign n32251 = n32027 & n75851 ;
  assign n32312 = n31351 | n32027 ;
  assign n75852 = ~n32312 ;
  assign n32313 = n32023 & n75852 ;
  assign n32314 = n32251 | n32313 ;
  assign n32315 = n130 & n32314 ;
  assign n32316 = n31341 & n75835 ;
  assign n32317 = n32119 & n32316 ;
  assign n32318 = n32315 | n32317 ;
  assign n75853 = ~n32244 ;
  assign n32246 = n32016 & n75853 ;
  assign n32319 = n31369 | n32016 ;
  assign n75854 = ~n32319 ;
  assign n32320 = n32012 & n75854 ;
  assign n32321 = n32246 | n32320 ;
  assign n32322 = n130 & n32321 ;
  assign n32323 = n31359 & n75835 ;
  assign n32324 = n32119 & n32323 ;
  assign n32325 = n32322 | n32324 ;
  assign n75855 = ~n32239 ;
  assign n32241 = n32005 & n75855 ;
  assign n32326 = n31387 | n32005 ;
  assign n75856 = ~n32326 ;
  assign n32327 = n32001 & n75856 ;
  assign n32328 = n32241 | n32327 ;
  assign n32329 = n130 & n32328 ;
  assign n32330 = n31377 & n75835 ;
  assign n32331 = n32119 & n32330 ;
  assign n32332 = n32329 | n32331 ;
  assign n75857 = ~n32234 ;
  assign n32236 = n31994 & n75857 ;
  assign n32333 = n31405 | n31994 ;
  assign n75858 = ~n32333 ;
  assign n32334 = n31990 & n75858 ;
  assign n32335 = n32236 | n32334 ;
  assign n32336 = n130 & n32335 ;
  assign n32337 = n31395 & n75835 ;
  assign n32338 = n32119 & n32337 ;
  assign n32339 = n32336 | n32338 ;
  assign n75859 = ~n32229 ;
  assign n32231 = n31983 & n75859 ;
  assign n32340 = n31423 | n31983 ;
  assign n75860 = ~n32340 ;
  assign n32341 = n31979 & n75860 ;
  assign n32342 = n32231 | n32341 ;
  assign n32343 = n130 & n32342 ;
  assign n32344 = n31413 & n75835 ;
  assign n32345 = n32119 & n32344 ;
  assign n32346 = n32343 | n32345 ;
  assign n75861 = ~n32224 ;
  assign n32226 = n31972 & n75861 ;
  assign n32347 = n31441 | n31972 ;
  assign n75862 = ~n32347 ;
  assign n32348 = n31968 & n75862 ;
  assign n32349 = n32226 | n32348 ;
  assign n32350 = n130 & n32349 ;
  assign n32351 = n31431 & n75835 ;
  assign n32352 = n32119 & n32351 ;
  assign n32353 = n32350 | n32352 ;
  assign n75863 = ~n32219 ;
  assign n32221 = n31961 & n75863 ;
  assign n32354 = n31459 | n31961 ;
  assign n75864 = ~n32354 ;
  assign n32355 = n31957 & n75864 ;
  assign n32356 = n32221 | n32355 ;
  assign n32357 = n130 & n32356 ;
  assign n32358 = n31449 & n75835 ;
  assign n32359 = n32119 & n32358 ;
  assign n32360 = n32357 | n32359 ;
  assign n75865 = ~n32214 ;
  assign n32216 = n31950 & n75865 ;
  assign n32361 = n31477 | n31950 ;
  assign n75866 = ~n32361 ;
  assign n32362 = n31946 & n75866 ;
  assign n32363 = n32216 | n32362 ;
  assign n32364 = n130 & n32363 ;
  assign n32365 = n31467 & n75835 ;
  assign n32366 = n32119 & n32365 ;
  assign n32367 = n32364 | n32366 ;
  assign n75867 = ~n32209 ;
  assign n32211 = n31939 & n75867 ;
  assign n32368 = n31495 | n31939 ;
  assign n75868 = ~n32368 ;
  assign n32369 = n31935 & n75868 ;
  assign n32370 = n32211 | n32369 ;
  assign n32371 = n130 & n32370 ;
  assign n32372 = n31485 & n75835 ;
  assign n32373 = n32119 & n32372 ;
  assign n32374 = n32371 | n32373 ;
  assign n75869 = ~n32204 ;
  assign n32206 = n31928 & n75869 ;
  assign n32375 = n31513 | n31928 ;
  assign n75870 = ~n32375 ;
  assign n32376 = n31924 & n75870 ;
  assign n32377 = n32206 | n32376 ;
  assign n32378 = n130 & n32377 ;
  assign n32379 = n31503 & n75835 ;
  assign n32380 = n32119 & n32379 ;
  assign n32381 = n32378 | n32380 ;
  assign n75871 = ~n32199 ;
  assign n32201 = n31917 & n75871 ;
  assign n32382 = n31531 | n31917 ;
  assign n75872 = ~n32382 ;
  assign n32383 = n31913 & n75872 ;
  assign n32384 = n32201 | n32383 ;
  assign n32385 = n130 & n32384 ;
  assign n32386 = n31521 & n75835 ;
  assign n32387 = n32119 & n32386 ;
  assign n32388 = n32385 | n32387 ;
  assign n75873 = ~n32194 ;
  assign n32196 = n31906 & n75873 ;
  assign n32389 = n31549 | n31906 ;
  assign n75874 = ~n32389 ;
  assign n32390 = n31902 & n75874 ;
  assign n32391 = n32196 | n32390 ;
  assign n32392 = n130 & n32391 ;
  assign n32393 = n31539 & n75835 ;
  assign n32394 = n32119 & n32393 ;
  assign n32395 = n32392 | n32394 ;
  assign n75875 = ~n32189 ;
  assign n32191 = n31895 & n75875 ;
  assign n32396 = n31567 | n31895 ;
  assign n75876 = ~n32396 ;
  assign n32397 = n31891 & n75876 ;
  assign n32398 = n32191 | n32397 ;
  assign n32399 = n130 & n32398 ;
  assign n32400 = n31557 & n75835 ;
  assign n32401 = n32119 & n32400 ;
  assign n32402 = n32399 | n32401 ;
  assign n75877 = ~n32184 ;
  assign n32186 = n31884 & n75877 ;
  assign n32403 = n31585 | n31884 ;
  assign n75878 = ~n32403 ;
  assign n32404 = n31880 & n75878 ;
  assign n32405 = n32186 | n32404 ;
  assign n32406 = n130 & n32405 ;
  assign n32407 = n31575 & n75835 ;
  assign n32408 = n32119 & n32407 ;
  assign n32409 = n32406 | n32408 ;
  assign n75879 = ~n32179 ;
  assign n32181 = n31873 & n75879 ;
  assign n32410 = n31603 | n31873 ;
  assign n75880 = ~n32410 ;
  assign n32411 = n31869 & n75880 ;
  assign n32412 = n32181 | n32411 ;
  assign n32413 = n130 & n32412 ;
  assign n32414 = n31593 & n75835 ;
  assign n32415 = n32119 & n32414 ;
  assign n32416 = n32413 | n32415 ;
  assign n75881 = ~n32174 ;
  assign n32176 = n31862 & n75881 ;
  assign n32417 = n31621 | n31862 ;
  assign n75882 = ~n32417 ;
  assign n32418 = n31858 & n75882 ;
  assign n32419 = n32176 | n32418 ;
  assign n32420 = n130 & n32419 ;
  assign n32421 = n31611 & n75835 ;
  assign n32422 = n32119 & n32421 ;
  assign n32423 = n32420 | n32422 ;
  assign n75883 = ~n32169 ;
  assign n32171 = n31851 & n75883 ;
  assign n32424 = n31638 | n31851 ;
  assign n75884 = ~n32424 ;
  assign n32425 = n31847 & n75884 ;
  assign n32426 = n32171 | n32425 ;
  assign n32427 = n130 & n32426 ;
  assign n32428 = n31629 & n75835 ;
  assign n32429 = n32119 & n32428 ;
  assign n32430 = n32427 | n32429 ;
  assign n75885 = ~n32164 ;
  assign n32166 = n31840 & n75885 ;
  assign n32431 = n31656 | n31840 ;
  assign n75886 = ~n32431 ;
  assign n32432 = n31836 & n75886 ;
  assign n32433 = n32166 | n32432 ;
  assign n32434 = n130 & n32433 ;
  assign n32435 = n31646 & n75835 ;
  assign n32436 = n32119 & n32435 ;
  assign n32437 = n32434 | n32436 ;
  assign n75887 = ~n32159 ;
  assign n32161 = n31829 & n75887 ;
  assign n32438 = n31674 | n31829 ;
  assign n75888 = ~n32438 ;
  assign n32439 = n31825 & n75888 ;
  assign n32440 = n32161 | n32439 ;
  assign n32441 = n130 & n32440 ;
  assign n32442 = n31664 & n75835 ;
  assign n32443 = n32119 & n32442 ;
  assign n32444 = n32441 | n32443 ;
  assign n75889 = ~n32154 ;
  assign n32156 = n31818 & n75889 ;
  assign n32445 = n31692 | n31818 ;
  assign n75890 = ~n32445 ;
  assign n32446 = n31814 & n75890 ;
  assign n32447 = n32156 | n32446 ;
  assign n32448 = n130 & n32447 ;
  assign n32449 = n31682 & n75835 ;
  assign n32450 = n32119 & n32449 ;
  assign n32451 = n32448 | n32450 ;
  assign n75891 = ~n32149 ;
  assign n32151 = n31807 & n75891 ;
  assign n32452 = n31710 | n31807 ;
  assign n75892 = ~n32452 ;
  assign n32453 = n31803 & n75892 ;
  assign n32454 = n32151 | n32453 ;
  assign n32455 = n130 & n32454 ;
  assign n32456 = n31700 & n75835 ;
  assign n32457 = n32119 & n32456 ;
  assign n32458 = n32455 | n32457 ;
  assign n75893 = ~n32144 ;
  assign n32146 = n31796 & n75893 ;
  assign n32459 = n31728 | n31796 ;
  assign n75894 = ~n32459 ;
  assign n32460 = n31792 & n75894 ;
  assign n32461 = n32146 | n32460 ;
  assign n32462 = n130 & n32461 ;
  assign n32463 = n31718 & n75835 ;
  assign n32464 = n32119 & n32463 ;
  assign n32465 = n32462 | n32464 ;
  assign n75895 = ~n32139 ;
  assign n32140 = n31785 & n75895 ;
  assign n32466 = n31745 | n31785 ;
  assign n75896 = ~n32466 ;
  assign n32467 = n32138 & n75896 ;
  assign n32468 = n32140 | n32467 ;
  assign n32469 = n130 & n32468 ;
  assign n32470 = n31736 & n75835 ;
  assign n32471 = n32119 & n32470 ;
  assign n32472 = n32469 | n32471 ;
  assign n75897 = ~n32133 ;
  assign n32134 = n31775 & n75897 ;
  assign n32473 = n31775 | n32131 ;
  assign n75898 = ~n32473 ;
  assign n32474 = n31771 & n75898 ;
  assign n32475 = n32134 | n32474 ;
  assign n32476 = n130 & n32475 ;
  assign n32477 = n31752 & n75835 ;
  assign n32478 = n32119 & n32477 ;
  assign n32479 = n32476 | n32478 ;
  assign n75899 = ~x0 ;
  assign n32480 = n75899 & x64 ;
  assign n32121 = n31770 & n130 ;
  assign n32122 = x64 & n130 ;
  assign n75900 = ~n32122 ;
  assign n32481 = x1 & n75900 ;
  assign n32482 = n32121 | n32481 ;
  assign n75901 = ~n32480 ;
  assign n32483 = n75901 & n32482 ;
  assign n32276 = n32082 | n32274 ;
  assign n32484 = n75822 & n32276 ;
  assign n32485 = n32087 | n32484 ;
  assign n32486 = n75825 & n32485 ;
  assign n32487 = n32093 | n32486 ;
  assign n32488 = n75828 & n32487 ;
  assign n32489 = n32099 | n32488 ;
  assign n32490 = n75831 & n32489 ;
  assign n32491 = n32117 | n32490 ;
  assign n32492 = n75835 & n32491 ;
  assign n75902 = ~n32492 ;
  assign n32493 = n31770 & n75902 ;
  assign n75903 = ~n32493 ;
  assign n32494 = n32480 & n75903 ;
  assign n75904 = ~n32481 ;
  assign n32495 = n75904 & n32494 ;
  assign n32496 = x65 | n32495 ;
  assign n32498 = n31768 & n31770 ;
  assign n32499 = n75649 & n32498 ;
  assign n75905 = ~n32499 ;
  assign n32500 = n31771 & n75905 ;
  assign n32501 = n130 & n32500 ;
  assign n32502 = n31765 & n75835 ;
  assign n32503 = n32119 & n32502 ;
  assign n32504 = n32501 | n32503 ;
  assign n75906 = ~n32504 ;
  assign n32505 = n32496 & n75906 ;
  assign n75907 = ~n32483 ;
  assign n32506 = n75907 & n32505 ;
  assign n32507 = x66 | n32506 ;
  assign n32497 = n75907 & n32496 ;
  assign n75908 = ~n32497 ;
  assign n32508 = n75908 & n32504 ;
  assign n75909 = ~n32508 ;
  assign n32509 = n32507 & n75909 ;
  assign n75910 = ~n32509 ;
  assign n32510 = n32479 & n75910 ;
  assign n32511 = n32479 | n32508 ;
  assign n75911 = ~n32511 ;
  assign n32512 = n32507 & n75911 ;
  assign n32513 = x67 | n32512 ;
  assign n75912 = ~n31777 ;
  assign n32137 = n75912 & n31780 ;
  assign n32515 = n31753 | n31780 ;
  assign n75913 = ~n32515 ;
  assign n32516 = n32135 & n75913 ;
  assign n32517 = n32137 | n32516 ;
  assign n32518 = n130 & n32517 ;
  assign n32519 = n31744 & n75835 ;
  assign n32520 = n32119 & n32519 ;
  assign n32521 = n32518 | n32520 ;
  assign n75914 = ~n32521 ;
  assign n32522 = n32513 & n75914 ;
  assign n75915 = ~n32510 ;
  assign n32523 = n75915 & n32522 ;
  assign n32524 = x68 | n32523 ;
  assign n32514 = n75915 & n32513 ;
  assign n75916 = ~n32514 ;
  assign n32525 = n75916 & n32521 ;
  assign n75917 = ~n32525 ;
  assign n32526 = n32524 & n75917 ;
  assign n75918 = ~n32526 ;
  assign n32527 = n32472 & n75918 ;
  assign n32528 = n32472 | n32525 ;
  assign n75919 = ~n32528 ;
  assign n32529 = n32524 & n75919 ;
  assign n32530 = x69 | n32529 ;
  assign n75920 = ~n31787 ;
  assign n31791 = n75920 & n31790 ;
  assign n32532 = n31737 | n31790 ;
  assign n75921 = ~n32532 ;
  assign n32533 = n32141 & n75921 ;
  assign n32534 = n31791 | n32533 ;
  assign n32535 = n130 & n32534 ;
  assign n32536 = n31727 & n75835 ;
  assign n32537 = n32119 & n32536 ;
  assign n32538 = n32535 | n32537 ;
  assign n75922 = ~n32538 ;
  assign n32539 = n32530 & n75922 ;
  assign n75923 = ~n32527 ;
  assign n32540 = n75923 & n32539 ;
  assign n32541 = x70 | n32540 ;
  assign n32531 = n75923 & n32530 ;
  assign n75924 = ~n32531 ;
  assign n32542 = n75924 & n32538 ;
  assign n75925 = ~n32542 ;
  assign n32543 = n32541 & n75925 ;
  assign n75926 = ~n32543 ;
  assign n32544 = n32465 & n75926 ;
  assign n32545 = n32465 | n32542 ;
  assign n75927 = ~n32545 ;
  assign n32546 = n32541 & n75927 ;
  assign n32547 = x71 | n32546 ;
  assign n75928 = ~n31798 ;
  assign n31802 = n75928 & n31801 ;
  assign n32549 = n31719 | n31801 ;
  assign n75929 = ~n32549 ;
  assign n32550 = n32145 & n75929 ;
  assign n32551 = n31802 | n32550 ;
  assign n32552 = n130 & n32551 ;
  assign n32553 = n31709 & n75835 ;
  assign n32554 = n32119 & n32553 ;
  assign n32555 = n32552 | n32554 ;
  assign n75930 = ~n32555 ;
  assign n32556 = n32547 & n75930 ;
  assign n75931 = ~n32544 ;
  assign n32557 = n75931 & n32556 ;
  assign n32558 = x72 | n32557 ;
  assign n32548 = n75931 & n32547 ;
  assign n75932 = ~n32548 ;
  assign n32559 = n75932 & n32555 ;
  assign n75933 = ~n32559 ;
  assign n32560 = n32558 & n75933 ;
  assign n75934 = ~n32560 ;
  assign n32561 = n32458 & n75934 ;
  assign n32562 = n32458 | n32559 ;
  assign n75935 = ~n32562 ;
  assign n32563 = n32558 & n75935 ;
  assign n32564 = x73 | n32563 ;
  assign n75936 = ~n31809 ;
  assign n31813 = n75936 & n31812 ;
  assign n32566 = n31701 | n31812 ;
  assign n75937 = ~n32566 ;
  assign n32567 = n32150 & n75937 ;
  assign n32568 = n31813 | n32567 ;
  assign n32569 = n130 & n32568 ;
  assign n32570 = n31691 & n75835 ;
  assign n32571 = n32119 & n32570 ;
  assign n32572 = n32569 | n32571 ;
  assign n75938 = ~n32572 ;
  assign n32573 = n32564 & n75938 ;
  assign n75939 = ~n32561 ;
  assign n32574 = n75939 & n32573 ;
  assign n32575 = x74 | n32574 ;
  assign n32565 = n75939 & n32564 ;
  assign n75940 = ~n32565 ;
  assign n32576 = n75940 & n32572 ;
  assign n75941 = ~n32576 ;
  assign n32577 = n32575 & n75941 ;
  assign n75942 = ~n32577 ;
  assign n32578 = n32451 & n75942 ;
  assign n32579 = n32451 | n32576 ;
  assign n75943 = ~n32579 ;
  assign n32580 = n32575 & n75943 ;
  assign n32581 = x75 | n32580 ;
  assign n75944 = ~n31820 ;
  assign n31824 = n75944 & n31823 ;
  assign n32583 = n31683 | n31823 ;
  assign n75945 = ~n32583 ;
  assign n32584 = n32155 & n75945 ;
  assign n32585 = n31824 | n32584 ;
  assign n32586 = n130 & n32585 ;
  assign n32587 = n31673 & n75835 ;
  assign n32588 = n32119 & n32587 ;
  assign n32589 = n32586 | n32588 ;
  assign n75946 = ~n32589 ;
  assign n32590 = n32581 & n75946 ;
  assign n75947 = ~n32578 ;
  assign n32591 = n75947 & n32590 ;
  assign n32592 = x76 | n32591 ;
  assign n32582 = n75947 & n32581 ;
  assign n75948 = ~n32582 ;
  assign n32593 = n75948 & n32589 ;
  assign n75949 = ~n32593 ;
  assign n32594 = n32592 & n75949 ;
  assign n75950 = ~n32594 ;
  assign n32595 = n32444 & n75950 ;
  assign n32596 = n32444 | n32593 ;
  assign n75951 = ~n32596 ;
  assign n32597 = n32592 & n75951 ;
  assign n32598 = x77 | n32597 ;
  assign n75952 = ~n31831 ;
  assign n31835 = n75952 & n31834 ;
  assign n32600 = n31665 | n31834 ;
  assign n75953 = ~n32600 ;
  assign n32601 = n32160 & n75953 ;
  assign n32602 = n31835 | n32601 ;
  assign n32603 = n130 & n32602 ;
  assign n32604 = n31655 & n75835 ;
  assign n32605 = n32119 & n32604 ;
  assign n32606 = n32603 | n32605 ;
  assign n75954 = ~n32606 ;
  assign n32607 = n32598 & n75954 ;
  assign n75955 = ~n32595 ;
  assign n32608 = n75955 & n32607 ;
  assign n32609 = x78 | n32608 ;
  assign n32599 = n75955 & n32598 ;
  assign n75956 = ~n32599 ;
  assign n32610 = n75956 & n32606 ;
  assign n75957 = ~n32610 ;
  assign n32611 = n32609 & n75957 ;
  assign n75958 = ~n32611 ;
  assign n32612 = n32437 & n75958 ;
  assign n32613 = n32437 | n32610 ;
  assign n75959 = ~n32613 ;
  assign n32614 = n32609 & n75959 ;
  assign n32615 = x79 | n32614 ;
  assign n75960 = ~n31842 ;
  assign n31846 = n75960 & n31845 ;
  assign n32617 = n31647 | n31845 ;
  assign n75961 = ~n32617 ;
  assign n32618 = n32165 & n75961 ;
  assign n32619 = n31846 | n32618 ;
  assign n32620 = n130 & n32619 ;
  assign n32621 = n31637 & n75835 ;
  assign n32622 = n32119 & n32621 ;
  assign n32623 = n32620 | n32622 ;
  assign n75962 = ~n32623 ;
  assign n32624 = n32615 & n75962 ;
  assign n75963 = ~n32612 ;
  assign n32625 = n75963 & n32624 ;
  assign n32626 = x80 | n32625 ;
  assign n32616 = n75963 & n32615 ;
  assign n75964 = ~n32616 ;
  assign n32627 = n75964 & n32623 ;
  assign n75965 = ~n32627 ;
  assign n32628 = n32626 & n75965 ;
  assign n75966 = ~n32628 ;
  assign n32629 = n32430 & n75966 ;
  assign n32630 = n32430 | n32627 ;
  assign n75967 = ~n32630 ;
  assign n32631 = n32626 & n75967 ;
  assign n32632 = x81 | n32631 ;
  assign n75968 = ~n31853 ;
  assign n31857 = n75968 & n31856 ;
  assign n32634 = n31630 | n31856 ;
  assign n75969 = ~n32634 ;
  assign n32635 = n32170 & n75969 ;
  assign n32636 = n31857 | n32635 ;
  assign n32637 = n130 & n32636 ;
  assign n32638 = n31620 & n75835 ;
  assign n32639 = n32119 & n32638 ;
  assign n32640 = n32637 | n32639 ;
  assign n75970 = ~n32640 ;
  assign n32641 = n32632 & n75970 ;
  assign n75971 = ~n32629 ;
  assign n32642 = n75971 & n32641 ;
  assign n32643 = x82 | n32642 ;
  assign n32633 = n75971 & n32632 ;
  assign n75972 = ~n32633 ;
  assign n32644 = n75972 & n32640 ;
  assign n75973 = ~n32644 ;
  assign n32645 = n32643 & n75973 ;
  assign n75974 = ~n32645 ;
  assign n32646 = n32423 & n75974 ;
  assign n32647 = n32423 | n32644 ;
  assign n75975 = ~n32647 ;
  assign n32648 = n32643 & n75975 ;
  assign n32649 = x83 | n32648 ;
  assign n75976 = ~n31864 ;
  assign n31868 = n75976 & n31867 ;
  assign n32651 = n31612 | n31867 ;
  assign n75977 = ~n32651 ;
  assign n32652 = n32175 & n75977 ;
  assign n32653 = n31868 | n32652 ;
  assign n32654 = n130 & n32653 ;
  assign n32655 = n31602 & n75835 ;
  assign n32656 = n32119 & n32655 ;
  assign n32657 = n32654 | n32656 ;
  assign n75978 = ~n32657 ;
  assign n32658 = n32649 & n75978 ;
  assign n75979 = ~n32646 ;
  assign n32659 = n75979 & n32658 ;
  assign n32660 = x84 | n32659 ;
  assign n32650 = n75979 & n32649 ;
  assign n75980 = ~n32650 ;
  assign n32661 = n75980 & n32657 ;
  assign n75981 = ~n32661 ;
  assign n32662 = n32660 & n75981 ;
  assign n75982 = ~n32662 ;
  assign n32663 = n32416 & n75982 ;
  assign n32664 = n32416 | n32661 ;
  assign n75983 = ~n32664 ;
  assign n32665 = n32660 & n75983 ;
  assign n32666 = x85 | n32665 ;
  assign n75984 = ~n31875 ;
  assign n31879 = n75984 & n31878 ;
  assign n32668 = n31594 | n31878 ;
  assign n75985 = ~n32668 ;
  assign n32669 = n32180 & n75985 ;
  assign n32670 = n31879 | n32669 ;
  assign n32671 = n130 & n32670 ;
  assign n32672 = n31584 & n75835 ;
  assign n32673 = n32119 & n32672 ;
  assign n32674 = n32671 | n32673 ;
  assign n75986 = ~n32674 ;
  assign n32675 = n32666 & n75986 ;
  assign n75987 = ~n32663 ;
  assign n32676 = n75987 & n32675 ;
  assign n32677 = x86 | n32676 ;
  assign n32667 = n75987 & n32666 ;
  assign n75988 = ~n32667 ;
  assign n32678 = n75988 & n32674 ;
  assign n75989 = ~n32678 ;
  assign n32679 = n32677 & n75989 ;
  assign n75990 = ~n32679 ;
  assign n32680 = n32409 & n75990 ;
  assign n32681 = n32409 | n32678 ;
  assign n75991 = ~n32681 ;
  assign n32682 = n32677 & n75991 ;
  assign n32683 = x87 | n32682 ;
  assign n75992 = ~n31886 ;
  assign n31890 = n75992 & n31889 ;
  assign n32685 = n31576 | n31889 ;
  assign n75993 = ~n32685 ;
  assign n32686 = n32185 & n75993 ;
  assign n32687 = n31890 | n32686 ;
  assign n32688 = n130 & n32687 ;
  assign n32689 = n31566 & n75835 ;
  assign n32690 = n32119 & n32689 ;
  assign n32691 = n32688 | n32690 ;
  assign n75994 = ~n32691 ;
  assign n32692 = n32683 & n75994 ;
  assign n75995 = ~n32680 ;
  assign n32693 = n75995 & n32692 ;
  assign n32694 = x88 | n32693 ;
  assign n32684 = n75995 & n32683 ;
  assign n75996 = ~n32684 ;
  assign n32695 = n75996 & n32691 ;
  assign n75997 = ~n32695 ;
  assign n32696 = n32694 & n75997 ;
  assign n75998 = ~n32696 ;
  assign n32697 = n32402 & n75998 ;
  assign n32698 = n32402 | n32695 ;
  assign n75999 = ~n32698 ;
  assign n32699 = n32694 & n75999 ;
  assign n32700 = x89 | n32699 ;
  assign n76000 = ~n31897 ;
  assign n31901 = n76000 & n31900 ;
  assign n32702 = n31558 | n31900 ;
  assign n76001 = ~n32702 ;
  assign n32703 = n32190 & n76001 ;
  assign n32704 = n31901 | n32703 ;
  assign n32705 = n130 & n32704 ;
  assign n32706 = n31548 & n75835 ;
  assign n32707 = n32119 & n32706 ;
  assign n32708 = n32705 | n32707 ;
  assign n76002 = ~n32708 ;
  assign n32709 = n32700 & n76002 ;
  assign n76003 = ~n32697 ;
  assign n32710 = n76003 & n32709 ;
  assign n32711 = x90 | n32710 ;
  assign n32701 = n76003 & n32700 ;
  assign n76004 = ~n32701 ;
  assign n32712 = n76004 & n32708 ;
  assign n76005 = ~n32712 ;
  assign n32713 = n32711 & n76005 ;
  assign n76006 = ~n32713 ;
  assign n32714 = n32395 & n76006 ;
  assign n32715 = n32395 | n32712 ;
  assign n76007 = ~n32715 ;
  assign n32716 = n32711 & n76007 ;
  assign n32717 = x91 | n32716 ;
  assign n76008 = ~n31908 ;
  assign n31912 = n76008 & n31911 ;
  assign n32719 = n31540 | n31911 ;
  assign n76009 = ~n32719 ;
  assign n32720 = n32195 & n76009 ;
  assign n32721 = n31912 | n32720 ;
  assign n32722 = n130 & n32721 ;
  assign n32723 = n31530 & n75835 ;
  assign n32724 = n32119 & n32723 ;
  assign n32725 = n32722 | n32724 ;
  assign n76010 = ~n32725 ;
  assign n32726 = n32717 & n76010 ;
  assign n76011 = ~n32714 ;
  assign n32727 = n76011 & n32726 ;
  assign n32728 = x92 | n32727 ;
  assign n32718 = n76011 & n32717 ;
  assign n76012 = ~n32718 ;
  assign n32729 = n76012 & n32725 ;
  assign n76013 = ~n32729 ;
  assign n32730 = n32728 & n76013 ;
  assign n76014 = ~n32730 ;
  assign n32731 = n32388 & n76014 ;
  assign n32732 = n32388 | n32729 ;
  assign n76015 = ~n32732 ;
  assign n32733 = n32728 & n76015 ;
  assign n32734 = x93 | n32733 ;
  assign n76016 = ~n31919 ;
  assign n31923 = n76016 & n31922 ;
  assign n32736 = n31522 | n31922 ;
  assign n76017 = ~n32736 ;
  assign n32737 = n32200 & n76017 ;
  assign n32738 = n31923 | n32737 ;
  assign n32739 = n130 & n32738 ;
  assign n32740 = n31512 & n75835 ;
  assign n32741 = n32119 & n32740 ;
  assign n32742 = n32739 | n32741 ;
  assign n76018 = ~n32742 ;
  assign n32743 = n32734 & n76018 ;
  assign n76019 = ~n32731 ;
  assign n32744 = n76019 & n32743 ;
  assign n32745 = x94 | n32744 ;
  assign n32735 = n76019 & n32734 ;
  assign n76020 = ~n32735 ;
  assign n32746 = n76020 & n32742 ;
  assign n76021 = ~n32746 ;
  assign n32747 = n32745 & n76021 ;
  assign n76022 = ~n32747 ;
  assign n32748 = n32381 & n76022 ;
  assign n32749 = n32381 | n32746 ;
  assign n76023 = ~n32749 ;
  assign n32750 = n32745 & n76023 ;
  assign n32751 = x95 | n32750 ;
  assign n76024 = ~n31930 ;
  assign n31934 = n76024 & n31933 ;
  assign n32753 = n31504 | n31933 ;
  assign n76025 = ~n32753 ;
  assign n32754 = n32205 & n76025 ;
  assign n32755 = n31934 | n32754 ;
  assign n32756 = n130 & n32755 ;
  assign n32757 = n31494 & n75835 ;
  assign n32758 = n32119 & n32757 ;
  assign n32759 = n32756 | n32758 ;
  assign n76026 = ~n32759 ;
  assign n32760 = n32751 & n76026 ;
  assign n76027 = ~n32748 ;
  assign n32761 = n76027 & n32760 ;
  assign n32762 = x96 | n32761 ;
  assign n32752 = n76027 & n32751 ;
  assign n76028 = ~n32752 ;
  assign n32763 = n76028 & n32759 ;
  assign n76029 = ~n32763 ;
  assign n32764 = n32762 & n76029 ;
  assign n76030 = ~n32764 ;
  assign n32765 = n32374 & n76030 ;
  assign n32766 = n32374 | n32763 ;
  assign n76031 = ~n32766 ;
  assign n32767 = n32762 & n76031 ;
  assign n32768 = x97 | n32767 ;
  assign n76032 = ~n31941 ;
  assign n31945 = n76032 & n31944 ;
  assign n32770 = n31486 | n31944 ;
  assign n76033 = ~n32770 ;
  assign n32771 = n32210 & n76033 ;
  assign n32772 = n31945 | n32771 ;
  assign n32773 = n130 & n32772 ;
  assign n32774 = n31476 & n75835 ;
  assign n32775 = n32119 & n32774 ;
  assign n32776 = n32773 | n32775 ;
  assign n76034 = ~n32776 ;
  assign n32777 = n32768 & n76034 ;
  assign n76035 = ~n32765 ;
  assign n32778 = n76035 & n32777 ;
  assign n32779 = x98 | n32778 ;
  assign n32769 = n76035 & n32768 ;
  assign n76036 = ~n32769 ;
  assign n32780 = n76036 & n32776 ;
  assign n76037 = ~n32780 ;
  assign n32781 = n32779 & n76037 ;
  assign n76038 = ~n32781 ;
  assign n32782 = n32367 & n76038 ;
  assign n32783 = n32367 | n32780 ;
  assign n76039 = ~n32783 ;
  assign n32784 = n32779 & n76039 ;
  assign n32785 = x99 | n32784 ;
  assign n76040 = ~n31952 ;
  assign n31956 = n76040 & n31955 ;
  assign n32787 = n31468 | n31955 ;
  assign n76041 = ~n32787 ;
  assign n32788 = n32215 & n76041 ;
  assign n32789 = n31956 | n32788 ;
  assign n32790 = n130 & n32789 ;
  assign n32791 = n31458 & n75835 ;
  assign n32792 = n32119 & n32791 ;
  assign n32793 = n32790 | n32792 ;
  assign n76042 = ~n32793 ;
  assign n32794 = n32785 & n76042 ;
  assign n76043 = ~n32782 ;
  assign n32795 = n76043 & n32794 ;
  assign n32796 = x100 | n32795 ;
  assign n32786 = n76043 & n32785 ;
  assign n76044 = ~n32786 ;
  assign n32797 = n76044 & n32793 ;
  assign n76045 = ~n32797 ;
  assign n32798 = n32796 & n76045 ;
  assign n76046 = ~n32798 ;
  assign n32799 = n32360 & n76046 ;
  assign n32800 = n32360 | n32797 ;
  assign n76047 = ~n32800 ;
  assign n32801 = n32796 & n76047 ;
  assign n32802 = x101 | n32801 ;
  assign n76048 = ~n31963 ;
  assign n31967 = n76048 & n31966 ;
  assign n32804 = n31450 | n31966 ;
  assign n76049 = ~n32804 ;
  assign n32805 = n32220 & n76049 ;
  assign n32806 = n31967 | n32805 ;
  assign n32807 = n130 & n32806 ;
  assign n32808 = n31440 & n75835 ;
  assign n32809 = n32119 & n32808 ;
  assign n32810 = n32807 | n32809 ;
  assign n76050 = ~n32810 ;
  assign n32811 = n32802 & n76050 ;
  assign n76051 = ~n32799 ;
  assign n32812 = n76051 & n32811 ;
  assign n32813 = x102 | n32812 ;
  assign n32803 = n76051 & n32802 ;
  assign n76052 = ~n32803 ;
  assign n32814 = n76052 & n32810 ;
  assign n76053 = ~n32814 ;
  assign n32815 = n32813 & n76053 ;
  assign n76054 = ~n32815 ;
  assign n32816 = n32353 & n76054 ;
  assign n32817 = n32353 | n32814 ;
  assign n76055 = ~n32817 ;
  assign n32818 = n32813 & n76055 ;
  assign n32819 = x103 | n32818 ;
  assign n76056 = ~n31974 ;
  assign n31978 = n76056 & n31977 ;
  assign n32821 = n31432 | n31977 ;
  assign n76057 = ~n32821 ;
  assign n32822 = n32225 & n76057 ;
  assign n32823 = n31978 | n32822 ;
  assign n32824 = n130 & n32823 ;
  assign n32825 = n31422 & n75835 ;
  assign n32826 = n32119 & n32825 ;
  assign n32827 = n32824 | n32826 ;
  assign n76058 = ~n32827 ;
  assign n32828 = n32819 & n76058 ;
  assign n76059 = ~n32816 ;
  assign n32829 = n76059 & n32828 ;
  assign n32830 = x104 | n32829 ;
  assign n32820 = n76059 & n32819 ;
  assign n76060 = ~n32820 ;
  assign n32831 = n76060 & n32827 ;
  assign n76061 = ~n32831 ;
  assign n32832 = n32830 & n76061 ;
  assign n76062 = ~n32832 ;
  assign n32833 = n32346 & n76062 ;
  assign n32834 = n32346 | n32831 ;
  assign n76063 = ~n32834 ;
  assign n32835 = n32830 & n76063 ;
  assign n32836 = x105 | n32835 ;
  assign n76064 = ~n31985 ;
  assign n31989 = n76064 & n31988 ;
  assign n32838 = n31414 | n31988 ;
  assign n76065 = ~n32838 ;
  assign n32839 = n32230 & n76065 ;
  assign n32840 = n31989 | n32839 ;
  assign n32841 = n130 & n32840 ;
  assign n32842 = n31404 & n75835 ;
  assign n32843 = n32119 & n32842 ;
  assign n32844 = n32841 | n32843 ;
  assign n76066 = ~n32844 ;
  assign n32845 = n32836 & n76066 ;
  assign n76067 = ~n32833 ;
  assign n32846 = n76067 & n32845 ;
  assign n32847 = x106 | n32846 ;
  assign n32837 = n76067 & n32836 ;
  assign n76068 = ~n32837 ;
  assign n32848 = n76068 & n32844 ;
  assign n76069 = ~n32848 ;
  assign n32849 = n32847 & n76069 ;
  assign n76070 = ~n32849 ;
  assign n32850 = n32339 & n76070 ;
  assign n32851 = n32339 | n32848 ;
  assign n76071 = ~n32851 ;
  assign n32852 = n32847 & n76071 ;
  assign n32853 = x107 | n32852 ;
  assign n76072 = ~n31996 ;
  assign n32000 = n76072 & n31999 ;
  assign n32855 = n31396 | n31999 ;
  assign n76073 = ~n32855 ;
  assign n32856 = n32235 & n76073 ;
  assign n32857 = n32000 | n32856 ;
  assign n32858 = n130 & n32857 ;
  assign n32859 = n31386 & n75835 ;
  assign n32860 = n32119 & n32859 ;
  assign n32861 = n32858 | n32860 ;
  assign n76074 = ~n32861 ;
  assign n32862 = n32853 & n76074 ;
  assign n76075 = ~n32850 ;
  assign n32863 = n76075 & n32862 ;
  assign n32864 = x108 | n32863 ;
  assign n32854 = n76075 & n32853 ;
  assign n76076 = ~n32854 ;
  assign n32865 = n76076 & n32861 ;
  assign n76077 = ~n32865 ;
  assign n32866 = n32864 & n76077 ;
  assign n76078 = ~n32866 ;
  assign n32867 = n32332 & n76078 ;
  assign n32868 = n32332 | n32865 ;
  assign n76079 = ~n32868 ;
  assign n32869 = n32864 & n76079 ;
  assign n32870 = x109 | n32869 ;
  assign n76080 = ~n32007 ;
  assign n32011 = n76080 & n32010 ;
  assign n32872 = n31378 | n32010 ;
  assign n76081 = ~n32872 ;
  assign n32873 = n32240 & n76081 ;
  assign n32874 = n32011 | n32873 ;
  assign n32875 = n130 & n32874 ;
  assign n32876 = n31368 & n75835 ;
  assign n32877 = n32119 & n32876 ;
  assign n32878 = n32875 | n32877 ;
  assign n76082 = ~n32878 ;
  assign n32879 = n32870 & n76082 ;
  assign n76083 = ~n32867 ;
  assign n32880 = n76083 & n32879 ;
  assign n32881 = x110 | n32880 ;
  assign n32871 = n76083 & n32870 ;
  assign n76084 = ~n32871 ;
  assign n32882 = n76084 & n32878 ;
  assign n76085 = ~n32882 ;
  assign n32883 = n32881 & n76085 ;
  assign n76086 = ~n32883 ;
  assign n32884 = n32325 & n76086 ;
  assign n32885 = n32325 | n32882 ;
  assign n76087 = ~n32885 ;
  assign n32886 = n32881 & n76087 ;
  assign n32887 = x111 | n32886 ;
  assign n76088 = ~n32018 ;
  assign n32022 = n76088 & n32021 ;
  assign n32889 = n31360 | n32021 ;
  assign n76089 = ~n32889 ;
  assign n32890 = n32245 & n76089 ;
  assign n32891 = n32022 | n32890 ;
  assign n32892 = n130 & n32891 ;
  assign n32893 = n31350 & n75835 ;
  assign n32894 = n32119 & n32893 ;
  assign n32895 = n32892 | n32894 ;
  assign n76090 = ~n32895 ;
  assign n32896 = n32887 & n76090 ;
  assign n76091 = ~n32884 ;
  assign n32897 = n76091 & n32896 ;
  assign n32898 = x112 | n32897 ;
  assign n32888 = n76091 & n32887 ;
  assign n76092 = ~n32888 ;
  assign n32899 = n76092 & n32895 ;
  assign n76093 = ~n32899 ;
  assign n32900 = n32898 & n76093 ;
  assign n76094 = ~n32900 ;
  assign n32901 = n32318 & n76094 ;
  assign n32902 = n32318 | n32899 ;
  assign n76095 = ~n32902 ;
  assign n32903 = n32898 & n76095 ;
  assign n32904 = x113 | n32903 ;
  assign n76096 = ~n32029 ;
  assign n32033 = n76096 & n32032 ;
  assign n32906 = n31342 | n32032 ;
  assign n76097 = ~n32906 ;
  assign n32907 = n32250 & n76097 ;
  assign n32908 = n32033 | n32907 ;
  assign n32909 = n130 & n32908 ;
  assign n32910 = n31333 & n75835 ;
  assign n32911 = n32119 & n32910 ;
  assign n32912 = n32909 | n32911 ;
  assign n76098 = ~n32912 ;
  assign n32913 = n32904 & n76098 ;
  assign n76099 = ~n32901 ;
  assign n32914 = n76099 & n32913 ;
  assign n32915 = x114 | n32914 ;
  assign n32905 = n76099 & n32904 ;
  assign n76100 = ~n32905 ;
  assign n32916 = n76100 & n32912 ;
  assign n76101 = ~n32916 ;
  assign n32917 = n32915 & n76101 ;
  assign n76102 = ~n32917 ;
  assign n32918 = n32311 & n76102 ;
  assign n32919 = n32311 | n32916 ;
  assign n76103 = ~n32919 ;
  assign n32920 = n32915 & n76103 ;
  assign n32921 = x115 | n32920 ;
  assign n76104 = ~n32040 ;
  assign n32044 = n76104 & n32043 ;
  assign n32923 = n31325 | n32043 ;
  assign n76105 = ~n32923 ;
  assign n32924 = n32255 & n76105 ;
  assign n32925 = n32044 | n32924 ;
  assign n32926 = n130 & n32925 ;
  assign n32927 = n31316 & n75835 ;
  assign n32928 = n32119 & n32927 ;
  assign n32929 = n32926 | n32928 ;
  assign n76106 = ~n32929 ;
  assign n32930 = n32921 & n76106 ;
  assign n76107 = ~n32918 ;
  assign n32931 = n76107 & n32930 ;
  assign n32932 = x116 | n32931 ;
  assign n32922 = n76107 & n32921 ;
  assign n76108 = ~n32922 ;
  assign n32933 = n76108 & n32929 ;
  assign n76109 = ~n32933 ;
  assign n32934 = n32932 & n76109 ;
  assign n76110 = ~n32934 ;
  assign n32935 = n32304 & n76110 ;
  assign n32936 = n32304 | n32933 ;
  assign n76111 = ~n32936 ;
  assign n32937 = n32932 & n76111 ;
  assign n32938 = x117 | n32937 ;
  assign n76112 = ~n32051 ;
  assign n32055 = n76112 & n32054 ;
  assign n32940 = n31308 | n32054 ;
  assign n76113 = ~n32940 ;
  assign n32941 = n32260 & n76113 ;
  assign n32942 = n32055 | n32941 ;
  assign n32943 = n130 & n32942 ;
  assign n32944 = n31298 & n75835 ;
  assign n32945 = n32119 & n32944 ;
  assign n32946 = n32943 | n32945 ;
  assign n76114 = ~n32946 ;
  assign n32947 = n32938 & n76114 ;
  assign n76115 = ~n32935 ;
  assign n32948 = n76115 & n32947 ;
  assign n32949 = x118 | n32948 ;
  assign n32939 = n76115 & n32938 ;
  assign n76116 = ~n32939 ;
  assign n32950 = n76116 & n32946 ;
  assign n76117 = ~n32950 ;
  assign n32951 = n32949 & n76117 ;
  assign n76118 = ~n32951 ;
  assign n32952 = n32297 & n76118 ;
  assign n32953 = n32297 | n32950 ;
  assign n76119 = ~n32953 ;
  assign n32954 = n32949 & n76119 ;
  assign n32955 = x119 | n32954 ;
  assign n76120 = ~n32062 ;
  assign n32066 = n76120 & n32065 ;
  assign n32957 = n31290 | n32065 ;
  assign n76121 = ~n32957 ;
  assign n32958 = n32265 & n76121 ;
  assign n32959 = n32066 | n32958 ;
  assign n32960 = n130 & n32959 ;
  assign n32961 = n31280 & n75835 ;
  assign n32962 = n32119 & n32961 ;
  assign n32963 = n32960 | n32962 ;
  assign n76122 = ~n32963 ;
  assign n32964 = n32955 & n76122 ;
  assign n76123 = ~n32952 ;
  assign n32965 = n76123 & n32964 ;
  assign n32966 = x120 | n32965 ;
  assign n32956 = n76123 & n32955 ;
  assign n76124 = ~n32956 ;
  assign n32967 = n76124 & n32963 ;
  assign n76125 = ~n32967 ;
  assign n32968 = n32966 & n76125 ;
  assign n76126 = ~n32968 ;
  assign n32969 = n32290 & n76126 ;
  assign n32970 = n32290 | n32967 ;
  assign n76127 = ~n32970 ;
  assign n32971 = n32966 & n76127 ;
  assign n32972 = x121 | n32971 ;
  assign n76128 = ~n32073 ;
  assign n32077 = n76128 & n32076 ;
  assign n32974 = n31272 | n32076 ;
  assign n76129 = ~n32974 ;
  assign n32975 = n32270 & n76129 ;
  assign n32976 = n32077 | n32975 ;
  assign n32977 = n130 & n32976 ;
  assign n32978 = n31262 & n75835 ;
  assign n32979 = n32119 & n32978 ;
  assign n32980 = n32977 | n32979 ;
  assign n76130 = ~n32980 ;
  assign n32981 = n32972 & n76130 ;
  assign n76131 = ~n32969 ;
  assign n32982 = n76131 & n32981 ;
  assign n32983 = x122 | n32982 ;
  assign n32973 = n76131 & n32972 ;
  assign n76132 = ~n32973 ;
  assign n32984 = n76132 & n32980 ;
  assign n76133 = ~n32984 ;
  assign n32985 = n32983 & n76133 ;
  assign n76134 = ~n32985 ;
  assign n32986 = n32283 & n76134 ;
  assign n32987 = n32283 | n32984 ;
  assign n76135 = ~n32987 ;
  assign n32988 = n32983 & n76135 ;
  assign n32989 = x123 | n32988 ;
  assign n76136 = ~n32084 ;
  assign n32088 = n76136 & n32087 ;
  assign n32990 = n31254 | n32087 ;
  assign n76137 = ~n32990 ;
  assign n32991 = n32276 & n76137 ;
  assign n32992 = n32088 | n32991 ;
  assign n32993 = n130 & n32992 ;
  assign n32994 = n31245 & n75835 ;
  assign n32995 = n32119 & n32994 ;
  assign n32996 = n32993 | n32995 ;
  assign n76138 = ~n32996 ;
  assign n32997 = n32989 & n76138 ;
  assign n76139 = ~n32986 ;
  assign n32998 = n76139 & n32997 ;
  assign n32999 = x124 | n32998 ;
  assign n33000 = n76139 & n32989 ;
  assign n76140 = ~n33000 ;
  assign n33001 = n32996 & n76140 ;
  assign n76141 = ~n33001 ;
  assign n33002 = n32999 & n76141 ;
  assign n76142 = ~n33002 ;
  assign n33003 = n32129 & n76142 ;
  assign n33004 = n32129 | n33001 ;
  assign n76143 = ~n33004 ;
  assign n33005 = n32999 & n76143 ;
  assign n33006 = x125 | n33005 ;
  assign n76144 = ~n32096 ;
  assign n32100 = n76144 & n32099 ;
  assign n33007 = n31237 | n32099 ;
  assign n76145 = ~n33007 ;
  assign n33008 = n32095 & n76145 ;
  assign n33009 = n32100 | n33008 ;
  assign n33011 = n75902 & n33009 ;
  assign n33010 = n31227 & n75835 ;
  assign n33012 = n32119 & n33010 ;
  assign n33013 = n33011 | n33012 ;
  assign n76146 = ~n33013 ;
  assign n33014 = n33006 & n76146 ;
  assign n76147 = ~n33003 ;
  assign n33015 = n76147 & n33014 ;
  assign n33016 = x126 | n33015 ;
  assign n33017 = n76147 & n33006 ;
  assign n76148 = ~n33017 ;
  assign n33018 = n33013 & n76148 ;
  assign n33020 = n31228 | n32115 ;
  assign n33021 = n32113 | n33020 ;
  assign n76149 = ~n33021 ;
  assign n33023 = n32101 & n76149 ;
  assign n33022 = n32113 | n32115 ;
  assign n76150 = ~n32102 ;
  assign n33024 = n76150 & n33022 ;
  assign n33025 = n33023 | n33024 ;
  assign n33026 = n130 & n33025 ;
  assign n33027 = n65362 & n32112 ;
  assign n33028 = n32119 & n33027 ;
  assign n33029 = n33026 | n33028 ;
  assign n33030 = n33018 | n33029 ;
  assign n76151 = ~n33030 ;
  assign n33031 = n33016 & n76151 ;
  assign n33032 = x127 | n33031 ;
  assign n76152 = ~n33018 ;
  assign n33019 = n33016 & n76152 ;
  assign n76153 = ~n33019 ;
  assign n33033 = n76153 & n33029 ;
  assign n76154 = ~n33033 ;
  assign n33034 = n33032 & n76154 ;
  assign n471 = n453 | n470 ;
  assign n33035 = n66453 | n67612 ;
  assign n33036 = n303 | n33035 ;
  assign n33037 = n66070 | n33036 ;
  assign n33038 = x65 | x66 ;
  assign n33039 = n86486 | n33038 ;
  assign n33040 = n65199 | n33039 ;
  assign n33041 = n462 | n33040 ;
  assign n33042 = n513 | n33041 ;
  assign n33043 = n65221 & n65693 ;
  assign n33044 = n65694 & n33043 ;
  assign n33045 = n65695 & n33044 ;
  assign n33046 = n65696 & n33045 ;
  assign n76155 = ~n33046 ;
  assign n33047 = n65821 & n76155 ;
  assign n76156 = ~n33047 ;
  assign n33048 = n66008 & n76156 ;
  assign n33052 = x63 & n76155 ;
  assign n76157 = ~n33052 ;
  assign n33053 = n68051 & n76157 ;
  assign n76158 = ~n33048 ;
  assign n33054 = n76158 & n33053 ;
  assign n33049 = n69653 & n76158 ;
  assign n76159 = ~n33049 ;
  assign n33055 = n76159 & n33052 ;
  assign n33056 = n33054 | n33055 ;
  assign n33051 = n304 & n76158 ;
  assign n33050 = n296 & n76158 ;
  assign n76160 = ~n33050 ;
  assign n33057 = x62 & n76160 ;
  assign n33059 = n33051 | n33057 ;
  assign n33060 = n65697 & n33059 ;
  assign n76161 = ~n33060 ;
  assign n33061 = n307 & n76161 ;
  assign n76162 = ~n33054 ;
  assign n33062 = x66 & n76162 ;
  assign n76163 = ~n33055 ;
  assign n33063 = n76163 & n33062 ;
  assign n33064 = n65686 & n33056 ;
  assign n33065 = n33063 | n33064 ;
  assign n33066 = n33061 & n33065 ;
  assign n33067 = x66 | n33066 ;
  assign n33068 = n33061 | n33063 ;
  assign n76164 = ~n33064 ;
  assign n33069 = n76164 & n33068 ;
  assign n33071 = n320 | n33069 ;
  assign n76165 = ~n33071 ;
  assign n33072 = n33067 & n76165 ;
  assign n76166 = ~n33072 ;
  assign n33073 = n33056 & n76166 ;
  assign n33074 = n65704 & n33068 ;
  assign n76167 = ~n33066 ;
  assign n33075 = n76167 & n33074 ;
  assign n76168 = ~n33069 ;
  assign n33076 = n76168 & n33075 ;
  assign n76169 = ~n33076 ;
  assign n33077 = x67 & n76169 ;
  assign n76170 = ~n33073 ;
  assign n33078 = n76170 & n33077 ;
  assign n33079 = n337 & n76168 ;
  assign n76171 = ~n33079 ;
  assign n33080 = n33059 & n76171 ;
  assign n76172 = ~n33051 ;
  assign n33058 = n345 & n76172 ;
  assign n76173 = ~n33057 ;
  assign n33081 = n76173 & n33058 ;
  assign n33082 = n76168 & n33081 ;
  assign n33083 = n33080 | n33082 ;
  assign n33084 = n65686 & n33083 ;
  assign n76174 = ~n33082 ;
  assign n33085 = x66 & n76174 ;
  assign n76175 = ~n33080 ;
  assign n33086 = n76175 & n33085 ;
  assign n33070 = n357 & n76168 ;
  assign n76176 = ~n33070 ;
  assign n33087 = x61 & n76176 ;
  assign n33088 = n364 & n76168 ;
  assign n33090 = n33087 | n33088 ;
  assign n33091 = n65723 & n33090 ;
  assign n76177 = ~n33091 ;
  assign n33092 = n371 & n76177 ;
  assign n33093 = n33086 | n33092 ;
  assign n76178 = ~n33084 ;
  assign n33094 = n76178 & n33093 ;
  assign n33095 = n33078 | n33094 ;
  assign n33096 = n33073 | n33076 ;
  assign n33097 = n65721 & n33096 ;
  assign n76179 = ~n33097 ;
  assign n33098 = n33095 & n76179 ;
  assign n33100 = n33084 | n33086 ;
  assign n33101 = n33092 & n33100 ;
  assign n33103 = n65727 & n33093 ;
  assign n76180 = ~n33101 ;
  assign n33104 = n76180 & n33103 ;
  assign n76181 = ~n33098 ;
  assign n33105 = n76181 & n33104 ;
  assign n33102 = x66 | n33101 ;
  assign n33106 = n65727 & n33102 ;
  assign n33107 = n76181 & n33106 ;
  assign n76182 = ~n33107 ;
  assign n33108 = n33083 & n76182 ;
  assign n33109 = n33105 | n33108 ;
  assign n33110 = n33078 | n33097 ;
  assign n33111 = n33094 & n33110 ;
  assign n33112 = n381 | n33111 ;
  assign n33113 = n33094 | n33110 ;
  assign n76183 = ~n33112 ;
  assign n33114 = n76183 & n33113 ;
  assign n33115 = n76181 & n33114 ;
  assign n33099 = n381 | n33098 ;
  assign n33116 = n33096 & n33099 ;
  assign n76184 = ~n33116 ;
  assign n33117 = x68 & n76184 ;
  assign n76185 = ~n33115 ;
  assign n33118 = n76185 & n33117 ;
  assign n33119 = n65721 & n33109 ;
  assign n76186 = ~n33105 ;
  assign n33120 = x67 & n76186 ;
  assign n76187 = ~n33108 ;
  assign n33121 = n76187 & n33120 ;
  assign n33123 = n413 & n76181 ;
  assign n76188 = ~n33123 ;
  assign n33124 = n33090 & n76188 ;
  assign n76189 = ~n33088 ;
  assign n33089 = n419 & n76189 ;
  assign n76190 = ~n33087 ;
  assign n33125 = n76190 & n33089 ;
  assign n33126 = n76181 & n33125 ;
  assign n33127 = n33124 | n33126 ;
  assign n33128 = n65686 & n33127 ;
  assign n76191 = ~n33126 ;
  assign n33129 = x66 & n76191 ;
  assign n76192 = ~n33124 ;
  assign n33130 = n76192 & n33129 ;
  assign n33131 = n434 & n76181 ;
  assign n76193 = ~n33131 ;
  assign n33132 = x60 & n76193 ;
  assign n33133 = n439 & n76181 ;
  assign n33134 = n33132 | n33133 ;
  assign n33135 = n65748 & n33134 ;
  assign n76194 = ~n33135 ;
  assign n33136 = n444 & n76194 ;
  assign n33137 = n33130 | n33136 ;
  assign n76195 = ~n33128 ;
  assign n33138 = n76195 & n33137 ;
  assign n33139 = n33121 | n33138 ;
  assign n76196 = ~n33119 ;
  assign n33140 = n76196 & n33139 ;
  assign n33141 = n33118 | n33140 ;
  assign n33142 = n33115 | n33116 ;
  assign n33143 = n65746 & n33142 ;
  assign n76197 = ~n33143 ;
  assign n33144 = n33141 & n76197 ;
  assign n33122 = n33119 | n33121 ;
  assign n33145 = n33122 & n76195 ;
  assign n33146 = n33137 & n33145 ;
  assign n33147 = x67 | n33146 ;
  assign n33148 = n65753 & n33147 ;
  assign n76198 = ~n33144 ;
  assign n33149 = n76198 & n33148 ;
  assign n76199 = ~n33149 ;
  assign n33150 = n33109 & n76199 ;
  assign n33152 = n470 | n33146 ;
  assign n76200 = ~n33152 ;
  assign n33153 = n33139 & n76200 ;
  assign n33154 = n76198 & n33153 ;
  assign n33155 = n33150 | n33154 ;
  assign n33157 = x68 & n33155 ;
  assign n33156 = x68 | n33154 ;
  assign n33158 = n33150 | n33156 ;
  assign n76201 = ~n33157 ;
  assign n33159 = n76201 & n33158 ;
  assign n33160 = n33128 | n33130 ;
  assign n33161 = n33136 & n33160 ;
  assign n33162 = x66 | n33161 ;
  assign n33163 = n65753 & n33162 ;
  assign n33164 = n76198 & n33163 ;
  assign n76202 = ~n33164 ;
  assign n33165 = n33127 & n76202 ;
  assign n33166 = n65753 & n33137 ;
  assign n76203 = ~n33161 ;
  assign n33167 = n76203 & n33166 ;
  assign n33168 = n76198 & n33167 ;
  assign n33169 = n33165 | n33168 ;
  assign n33171 = x67 & n33169 ;
  assign n33170 = x67 | n33168 ;
  assign n33172 = n33165 | n33170 ;
  assign n76204 = ~n33171 ;
  assign n33173 = n76204 & n33172 ;
  assign n33151 = n506 & n76198 ;
  assign n76205 = ~n33151 ;
  assign n33174 = n33134 & n76205 ;
  assign n76206 = ~n33133 ;
  assign n33175 = n514 & n76206 ;
  assign n76207 = ~n33132 ;
  assign n33176 = n76207 & n33175 ;
  assign n33177 = n76198 & n33176 ;
  assign n33178 = n33174 | n33177 ;
  assign n33179 = n65686 & n33178 ;
  assign n33180 = n525 & n76198 ;
  assign n76208 = ~n33180 ;
  assign n33181 = x59 & n76208 ;
  assign n33182 = n531 & n76198 ;
  assign n33183 = n33181 | n33182 ;
  assign n33184 = x65 & n33183 ;
  assign n33185 = x65 | n33182 ;
  assign n33186 = n33181 | n33185 ;
  assign n76209 = ~n33184 ;
  assign n33187 = n76209 & n33186 ;
  assign n33188 = n538 | n33187 ;
  assign n33189 = n65670 & n33183 ;
  assign n76210 = ~n33189 ;
  assign n33190 = n33188 & n76210 ;
  assign n76211 = ~n33177 ;
  assign n33191 = x66 & n76211 ;
  assign n76212 = ~n33174 ;
  assign n33192 = n76212 & n33191 ;
  assign n33193 = n33179 | n33192 ;
  assign n33195 = n33190 | n33193 ;
  assign n76213 = ~n33179 ;
  assign n33196 = n76213 & n33195 ;
  assign n33197 = n33173 | n33196 ;
  assign n33198 = n65721 & n33169 ;
  assign n76214 = ~n33198 ;
  assign n33199 = n33197 & n76214 ;
  assign n33200 = n33159 | n33199 ;
  assign n33201 = n65746 & n33155 ;
  assign n76215 = ~n33201 ;
  assign n33202 = n33200 & n76215 ;
  assign n33203 = n33118 | n33143 ;
  assign n33204 = n76196 & n33203 ;
  assign n33205 = n33139 & n33204 ;
  assign n33206 = x68 | n33205 ;
  assign n33208 = n65753 & n33206 ;
  assign n33209 = n76198 & n33208 ;
  assign n76216 = ~n33209 ;
  assign n33210 = n33142 & n76216 ;
  assign n33207 = n470 | n33205 ;
  assign n76217 = ~n33207 ;
  assign n33211 = n33141 & n76217 ;
  assign n33212 = n76198 & n33211 ;
  assign n33213 = n33210 | n33212 ;
  assign n33215 = x69 & n33213 ;
  assign n33214 = x69 | n33212 ;
  assign n33216 = n33210 | n33214 ;
  assign n76218 = ~n33215 ;
  assign n33217 = n76218 & n33216 ;
  assign n33218 = n570 | n33217 ;
  assign n33219 = n33202 | n33218 ;
  assign n33220 = n65753 & n33213 ;
  assign n76219 = ~n33220 ;
  assign n33221 = n33219 & n76219 ;
  assign n33222 = n33159 & n76214 ;
  assign n33223 = n33197 & n33222 ;
  assign n76220 = ~n33223 ;
  assign n33224 = n33200 & n76220 ;
  assign n76221 = ~n33221 ;
  assign n33225 = n76221 & n33224 ;
  assign n33226 = n33155 & n76219 ;
  assign n33227 = n33219 & n33226 ;
  assign n33228 = n33225 | n33227 ;
  assign n33229 = n76215 & n33217 ;
  assign n33230 = n33200 & n33229 ;
  assign n33231 = n33202 | n33217 ;
  assign n76222 = ~n33230 ;
  assign n33232 = n76222 & n33231 ;
  assign n33233 = n76221 & n33232 ;
  assign n33234 = n470 & n33213 ;
  assign n33235 = n33219 & n33234 ;
  assign n33236 = n33233 | n33235 ;
  assign n33237 = n65791 & n33236 ;
  assign n33238 = n65772 & n33228 ;
  assign n33239 = n33173 & n76213 ;
  assign n33240 = n33195 & n33239 ;
  assign n76223 = ~n33240 ;
  assign n33241 = n33197 & n76223 ;
  assign n33242 = n76221 & n33241 ;
  assign n33243 = n33169 & n76219 ;
  assign n33244 = n33219 & n33243 ;
  assign n33245 = n33242 | n33244 ;
  assign n33246 = n65746 & n33245 ;
  assign n76224 = ~n33190 ;
  assign n33194 = n76224 & n33193 ;
  assign n33247 = n33189 | n33193 ;
  assign n76225 = ~n33247 ;
  assign n33248 = n33188 & n76225 ;
  assign n33249 = n33194 | n33248 ;
  assign n33250 = n76221 & n33249 ;
  assign n33251 = n33178 & n76219 ;
  assign n33252 = n33219 & n33251 ;
  assign n33253 = n33250 | n33252 ;
  assign n33254 = n65721 & n33253 ;
  assign n33255 = n538 & n33186 ;
  assign n33256 = n76209 & n33255 ;
  assign n76226 = ~n33256 ;
  assign n33257 = n33188 & n76226 ;
  assign n33258 = n76221 & n33257 ;
  assign n33259 = n33183 & n76219 ;
  assign n33260 = n33219 & n33259 ;
  assign n33261 = n33258 | n33260 ;
  assign n33262 = n65686 & n33261 ;
  assign n33263 = x64 & n76221 ;
  assign n76227 = ~n33263 ;
  assign n33264 = x58 & n76227 ;
  assign n33265 = n538 & n76221 ;
  assign n33266 = n33264 | n33265 ;
  assign n33267 = x65 & n33266 ;
  assign n33268 = x65 | n33265 ;
  assign n33269 = n33264 | n33268 ;
  assign n76228 = ~n33267 ;
  assign n33270 = n76228 & n33269 ;
  assign n33271 = n626 | n33270 ;
  assign n33272 = n65670 & n33266 ;
  assign n76229 = ~n33272 ;
  assign n33273 = n33271 & n76229 ;
  assign n76230 = ~n33260 ;
  assign n33274 = x66 & n76230 ;
  assign n76231 = ~n33258 ;
  assign n33275 = n76231 & n33274 ;
  assign n33276 = n33262 | n33275 ;
  assign n33277 = n33273 | n33276 ;
  assign n76232 = ~n33262 ;
  assign n33278 = n76232 & n33277 ;
  assign n76233 = ~n33252 ;
  assign n33279 = x67 & n76233 ;
  assign n76234 = ~n33250 ;
  assign n33280 = n76234 & n33279 ;
  assign n33281 = n33254 | n33280 ;
  assign n33283 = n33278 | n33281 ;
  assign n76235 = ~n33254 ;
  assign n33284 = n76235 & n33283 ;
  assign n76236 = ~n33244 ;
  assign n33285 = x68 & n76236 ;
  assign n76237 = ~n33242 ;
  assign n33286 = n76237 & n33285 ;
  assign n33287 = n33246 | n33286 ;
  assign n33289 = n33284 | n33287 ;
  assign n76238 = ~n33246 ;
  assign n33290 = n76238 & n33289 ;
  assign n76239 = ~n33227 ;
  assign n33291 = x69 & n76239 ;
  assign n76240 = ~n33225 ;
  assign n33292 = n76240 & n33291 ;
  assign n33293 = n33238 | n33292 ;
  assign n33295 = n33290 | n33293 ;
  assign n76241 = ~n33238 ;
  assign n33296 = n76241 & n33295 ;
  assign n76242 = ~n33235 ;
  assign n33297 = x70 & n76242 ;
  assign n76243 = ~n33233 ;
  assign n33298 = n76243 & n33297 ;
  assign n33299 = n33237 | n33298 ;
  assign n33301 = n33296 | n33299 ;
  assign n76244 = ~n33237 ;
  assign n33302 = n76244 & n33301 ;
  assign n33303 = n659 | n33302 ;
  assign n33306 = n33228 & n33303 ;
  assign n76245 = ~n33290 ;
  assign n33294 = n76245 & n33293 ;
  assign n33307 = n33246 | n33293 ;
  assign n76246 = ~n33307 ;
  assign n33308 = n33289 & n76246 ;
  assign n33309 = n33294 | n33308 ;
  assign n33310 = n65826 & n33309 ;
  assign n76247 = ~n33302 ;
  assign n33311 = n76247 & n33310 ;
  assign n33312 = n33306 | n33311 ;
  assign n76248 = ~n33236 ;
  assign n33305 = n76248 & n33303 ;
  assign n76249 = ~n33296 ;
  assign n33300 = n76249 & n33299 ;
  assign n33313 = n33238 | n33299 ;
  assign n76250 = ~n33313 ;
  assign n33314 = n33295 & n76250 ;
  assign n33315 = n33300 | n33314 ;
  assign n33316 = n33303 | n33315 ;
  assign n76251 = ~n33305 ;
  assign n33317 = n76251 & n33316 ;
  assign n33318 = n65820 & n33317 ;
  assign n33319 = n65791 & n33312 ;
  assign n33320 = n33245 & n33303 ;
  assign n76252 = ~n33284 ;
  assign n33288 = n76252 & n33287 ;
  assign n33321 = n33254 | n33287 ;
  assign n76253 = ~n33321 ;
  assign n33322 = n33283 & n76253 ;
  assign n33323 = n33288 | n33322 ;
  assign n33324 = n65826 & n33323 ;
  assign n33325 = n76247 & n33324 ;
  assign n33326 = n33320 | n33325 ;
  assign n33327 = n65772 & n33326 ;
  assign n33328 = n33253 & n33303 ;
  assign n76254 = ~n33278 ;
  assign n33282 = n76254 & n33281 ;
  assign n33329 = n33262 | n33281 ;
  assign n76255 = ~n33329 ;
  assign n33330 = n33277 & n76255 ;
  assign n33331 = n33282 | n33330 ;
  assign n33332 = n65826 & n33331 ;
  assign n33333 = n76247 & n33332 ;
  assign n33334 = n33328 | n33333 ;
  assign n33335 = n65746 & n33334 ;
  assign n33336 = n33261 & n33303 ;
  assign n33337 = n33272 | n33276 ;
  assign n76256 = ~n33337 ;
  assign n33338 = n33271 & n76256 ;
  assign n76257 = ~n33273 ;
  assign n33339 = n76257 & n33276 ;
  assign n33340 = n33338 | n33339 ;
  assign n33341 = n65826 & n33340 ;
  assign n33342 = n76247 & n33341 ;
  assign n33343 = n33336 | n33342 ;
  assign n33344 = n65721 & n33343 ;
  assign n33345 = n33266 & n33303 ;
  assign n33346 = n626 & n33269 ;
  assign n33347 = n76228 & n33346 ;
  assign n33348 = n659 | n33347 ;
  assign n76258 = ~n33348 ;
  assign n33349 = n33271 & n76258 ;
  assign n33350 = n76247 & n33349 ;
  assign n33351 = n33345 | n33350 ;
  assign n33352 = n65686 & n33351 ;
  assign n33304 = n716 & n76247 ;
  assign n76259 = ~n33304 ;
  assign n33353 = x57 & n76259 ;
  assign n33354 = n723 & n76247 ;
  assign n33355 = n33353 | n33354 ;
  assign n33356 = x65 & n33355 ;
  assign n33357 = x65 | n33354 ;
  assign n33358 = n33353 | n33357 ;
  assign n76260 = ~n33356 ;
  assign n33359 = n76260 & n33358 ;
  assign n33361 = n729 | n33359 ;
  assign n33362 = n65670 & n33355 ;
  assign n76261 = ~n33362 ;
  assign n33363 = n33361 & n76261 ;
  assign n76262 = ~n33350 ;
  assign n33364 = x66 & n76262 ;
  assign n76263 = ~n33345 ;
  assign n33365 = n76263 & n33364 ;
  assign n33366 = n33352 | n33365 ;
  assign n33367 = n33363 | n33366 ;
  assign n76264 = ~n33352 ;
  assign n33368 = n76264 & n33367 ;
  assign n76265 = ~n33342 ;
  assign n33369 = x67 & n76265 ;
  assign n76266 = ~n33336 ;
  assign n33370 = n76266 & n33369 ;
  assign n33371 = n33344 | n33370 ;
  assign n33372 = n33368 | n33371 ;
  assign n76267 = ~n33344 ;
  assign n33373 = n76267 & n33372 ;
  assign n76268 = ~n33333 ;
  assign n33374 = x68 & n76268 ;
  assign n76269 = ~n33328 ;
  assign n33375 = n76269 & n33374 ;
  assign n33376 = n33335 | n33375 ;
  assign n33377 = n33373 | n33376 ;
  assign n76270 = ~n33335 ;
  assign n33378 = n76270 & n33377 ;
  assign n76271 = ~n33325 ;
  assign n33379 = x69 & n76271 ;
  assign n76272 = ~n33320 ;
  assign n33380 = n76272 & n33379 ;
  assign n33381 = n33327 | n33380 ;
  assign n33382 = n33378 | n33381 ;
  assign n76273 = ~n33327 ;
  assign n33383 = n76273 & n33382 ;
  assign n76274 = ~n33311 ;
  assign n33384 = x70 & n76274 ;
  assign n76275 = ~n33306 ;
  assign n33385 = n76275 & n33384 ;
  assign n33386 = n33319 | n33385 ;
  assign n33388 = n33383 | n33386 ;
  assign n76276 = ~n33319 ;
  assign n33389 = n76276 & n33388 ;
  assign n76277 = ~n33303 ;
  assign n33390 = n76277 & n33315 ;
  assign n33391 = n33236 & n33303 ;
  assign n76278 = ~n33391 ;
  assign n33392 = x71 & n76278 ;
  assign n76279 = ~n33390 ;
  assign n33393 = n76279 & n33392 ;
  assign n33394 = n33318 | n33393 ;
  assign n33396 = n33389 | n33394 ;
  assign n76280 = ~n33318 ;
  assign n33397 = n76280 & n33396 ;
  assign n33398 = n768 | n33397 ;
  assign n33399 = n33312 & n33398 ;
  assign n76281 = ~n33383 ;
  assign n33387 = n76281 & n33386 ;
  assign n33400 = n33327 | n33386 ;
  assign n76282 = ~n33400 ;
  assign n33401 = n33382 & n76282 ;
  assign n33402 = n33387 | n33401 ;
  assign n33403 = n65864 & n33402 ;
  assign n76283 = ~n33397 ;
  assign n33404 = n76283 & n33403 ;
  assign n33405 = n33399 | n33404 ;
  assign n33406 = n65820 & n33405 ;
  assign n76284 = ~n33404 ;
  assign n33489 = x71 & n76284 ;
  assign n76285 = ~n33399 ;
  assign n33490 = n76285 & n33489 ;
  assign n33491 = n33406 | n33490 ;
  assign n33407 = n33326 & n33398 ;
  assign n33408 = n33335 | n33381 ;
  assign n76286 = ~n33408 ;
  assign n33409 = n33377 & n76286 ;
  assign n76287 = ~n33378 ;
  assign n33410 = n76287 & n33381 ;
  assign n33411 = n33409 | n33410 ;
  assign n33412 = n65864 & n33411 ;
  assign n33413 = n76283 & n33412 ;
  assign n33414 = n33407 | n33413 ;
  assign n33415 = n65791 & n33414 ;
  assign n33416 = n33334 & n33398 ;
  assign n33417 = n33344 | n33376 ;
  assign n76288 = ~n33417 ;
  assign n33418 = n33372 & n76288 ;
  assign n76289 = ~n33373 ;
  assign n33419 = n76289 & n33376 ;
  assign n33420 = n33418 | n33419 ;
  assign n33421 = n65864 & n33420 ;
  assign n33422 = n76283 & n33421 ;
  assign n33423 = n33416 | n33422 ;
  assign n33424 = n65772 & n33423 ;
  assign n76290 = ~n33422 ;
  assign n33478 = x69 & n76290 ;
  assign n76291 = ~n33416 ;
  assign n33479 = n76291 & n33478 ;
  assign n33480 = n33424 | n33479 ;
  assign n33425 = n33343 & n33398 ;
  assign n33426 = n33352 | n33371 ;
  assign n76292 = ~n33426 ;
  assign n33427 = n33367 & n76292 ;
  assign n76293 = ~n33368 ;
  assign n33428 = n76293 & n33371 ;
  assign n33429 = n33427 | n33428 ;
  assign n33430 = n65864 & n33429 ;
  assign n33431 = n76283 & n33430 ;
  assign n33432 = n33425 | n33431 ;
  assign n33433 = n65746 & n33432 ;
  assign n33434 = n33351 & n33398 ;
  assign n33435 = n33362 | n33366 ;
  assign n76294 = ~n33435 ;
  assign n33436 = n33361 & n76294 ;
  assign n76295 = ~n33363 ;
  assign n33437 = n76295 & n33366 ;
  assign n33438 = n33436 | n33437 ;
  assign n33439 = n65864 & n33438 ;
  assign n33440 = n76283 & n33439 ;
  assign n33441 = n33434 | n33440 ;
  assign n33442 = n65721 & n33441 ;
  assign n33443 = n33355 & n33398 ;
  assign n33360 = n729 & n33358 ;
  assign n33444 = n76260 & n33360 ;
  assign n33445 = n768 | n33444 ;
  assign n76296 = ~n33445 ;
  assign n33446 = n33361 & n76296 ;
  assign n33447 = n76283 & n33446 ;
  assign n33448 = n33443 | n33447 ;
  assign n33449 = n65686 & n33448 ;
  assign n33450 = n827 & n76283 ;
  assign n76297 = ~n33450 ;
  assign n33451 = x56 & n76297 ;
  assign n33452 = n833 & n76283 ;
  assign n33453 = n33451 | n33452 ;
  assign n33454 = x65 & n33453 ;
  assign n33455 = x65 | n33452 ;
  assign n33456 = n33451 | n33455 ;
  assign n76298 = ~n33454 ;
  assign n33457 = n76298 & n33456 ;
  assign n33458 = n840 | n33457 ;
  assign n33459 = n65670 & n33453 ;
  assign n76299 = ~n33459 ;
  assign n33460 = n33458 & n76299 ;
  assign n76300 = ~n33447 ;
  assign n33461 = x66 & n76300 ;
  assign n76301 = ~n33443 ;
  assign n33462 = n76301 & n33461 ;
  assign n33463 = n33449 | n33462 ;
  assign n33465 = n33460 | n33463 ;
  assign n76302 = ~n33449 ;
  assign n33466 = n76302 & n33465 ;
  assign n76303 = ~n33440 ;
  assign n33467 = x67 & n76303 ;
  assign n76304 = ~n33434 ;
  assign n33468 = n76304 & n33467 ;
  assign n33469 = n33442 | n33468 ;
  assign n33471 = n33466 | n33469 ;
  assign n76305 = ~n33442 ;
  assign n33472 = n76305 & n33471 ;
  assign n76306 = ~n33431 ;
  assign n33473 = x68 & n76306 ;
  assign n76307 = ~n33425 ;
  assign n33474 = n76307 & n33473 ;
  assign n33475 = n33433 | n33474 ;
  assign n33477 = n33472 | n33475 ;
  assign n76308 = ~n33433 ;
  assign n33481 = n76308 & n33477 ;
  assign n33482 = n33480 | n33481 ;
  assign n76309 = ~n33424 ;
  assign n33483 = n76309 & n33482 ;
  assign n76310 = ~n33413 ;
  assign n33484 = x70 & n76310 ;
  assign n76311 = ~n33407 ;
  assign n33485 = n76311 & n33484 ;
  assign n33486 = n33415 | n33485 ;
  assign n33488 = n33483 | n33486 ;
  assign n76312 = ~n33415 ;
  assign n33493 = n76312 & n33488 ;
  assign n33494 = n33491 | n33493 ;
  assign n76313 = ~n33406 ;
  assign n33495 = n76313 & n33494 ;
  assign n76314 = ~n33389 ;
  assign n33395 = n76314 & n33394 ;
  assign n33496 = n33319 | n33394 ;
  assign n76315 = ~n33496 ;
  assign n33497 = n33388 & n76315 ;
  assign n33498 = n33395 | n33497 ;
  assign n33499 = n33398 | n33498 ;
  assign n76316 = ~n33317 ;
  assign n33500 = n76316 & n33398 ;
  assign n76317 = ~n33500 ;
  assign n33501 = n33499 & n76317 ;
  assign n33502 = n65877 & n33501 ;
  assign n76318 = ~n33398 ;
  assign n33503 = n76318 & n33498 ;
  assign n33504 = n33317 & n33398 ;
  assign n76319 = ~n33504 ;
  assign n33505 = x72 & n76319 ;
  assign n76320 = ~n33503 ;
  assign n33506 = n76320 & n33505 ;
  assign n33507 = n886 | n33506 ;
  assign n33508 = n33502 | n33507 ;
  assign n33509 = n33495 | n33508 ;
  assign n33510 = n65864 & n33501 ;
  assign n76321 = ~n33510 ;
  assign n33511 = n33509 & n76321 ;
  assign n33520 = n33406 | n33506 ;
  assign n33521 = n33502 | n33520 ;
  assign n76322 = ~n33521 ;
  assign n33522 = n33494 & n76322 ;
  assign n33523 = n33502 | n33506 ;
  assign n76323 = ~n33495 ;
  assign n33524 = n76323 & n33523 ;
  assign n33525 = n33522 | n33524 ;
  assign n76324 = ~n33511 ;
  assign n33526 = n76324 & n33525 ;
  assign n33527 = n768 & n33317 ;
  assign n33528 = n33509 & n33527 ;
  assign n33529 = n33526 | n33528 ;
  assign n33530 = n65909 & n33529 ;
  assign n76325 = ~n33493 ;
  assign n33513 = n33491 & n76325 ;
  assign n33492 = n33415 | n33491 ;
  assign n76326 = ~n33492 ;
  assign n33514 = n33488 & n76326 ;
  assign n33515 = n33513 | n33514 ;
  assign n33516 = n76324 & n33515 ;
  assign n33517 = n33405 & n76321 ;
  assign n33518 = n33509 & n33517 ;
  assign n33519 = n33516 | n33518 ;
  assign n33531 = n65877 & n33519 ;
  assign n76327 = ~n33483 ;
  assign n33532 = n76327 & n33486 ;
  assign n33487 = n33424 | n33486 ;
  assign n76328 = ~n33487 ;
  assign n33533 = n33482 & n76328 ;
  assign n33534 = n33532 | n33533 ;
  assign n33535 = n76324 & n33534 ;
  assign n33536 = n33414 & n76321 ;
  assign n33537 = n33509 & n33536 ;
  assign n33538 = n33535 | n33537 ;
  assign n33539 = n65820 & n33538 ;
  assign n76329 = ~n33481 ;
  assign n33540 = n33480 & n76329 ;
  assign n33541 = n33433 | n33480 ;
  assign n76330 = ~n33541 ;
  assign n33542 = n33477 & n76330 ;
  assign n33543 = n33540 | n33542 ;
  assign n33544 = n76324 & n33543 ;
  assign n33545 = n33423 & n76321 ;
  assign n33546 = n33509 & n33545 ;
  assign n33547 = n33544 | n33546 ;
  assign n33548 = n65791 & n33547 ;
  assign n76331 = ~n33472 ;
  assign n33476 = n76331 & n33475 ;
  assign n33549 = n33442 | n33475 ;
  assign n76332 = ~n33549 ;
  assign n33550 = n33471 & n76332 ;
  assign n33551 = n33476 | n33550 ;
  assign n33552 = n76324 & n33551 ;
  assign n33553 = n33432 & n76321 ;
  assign n33554 = n33509 & n33553 ;
  assign n33555 = n33552 | n33554 ;
  assign n33556 = n65772 & n33555 ;
  assign n76333 = ~n33466 ;
  assign n33470 = n76333 & n33469 ;
  assign n33557 = n33449 | n33469 ;
  assign n76334 = ~n33557 ;
  assign n33558 = n33465 & n76334 ;
  assign n33559 = n33470 | n33558 ;
  assign n33560 = n76324 & n33559 ;
  assign n33561 = n33441 & n76321 ;
  assign n33562 = n33509 & n33561 ;
  assign n33563 = n33560 | n33562 ;
  assign n33564 = n65746 & n33563 ;
  assign n76335 = ~n33460 ;
  assign n33464 = n76335 & n33463 ;
  assign n33565 = n33459 | n33463 ;
  assign n76336 = ~n33565 ;
  assign n33566 = n33458 & n76336 ;
  assign n33567 = n33464 | n33566 ;
  assign n33568 = n76324 & n33567 ;
  assign n33569 = n33448 & n76321 ;
  assign n33570 = n33509 & n33569 ;
  assign n33571 = n33568 | n33570 ;
  assign n33572 = n65721 & n33571 ;
  assign n33573 = n840 & n33456 ;
  assign n33574 = n76298 & n33573 ;
  assign n76337 = ~n33574 ;
  assign n33575 = n33458 & n76337 ;
  assign n33576 = n76324 & n33575 ;
  assign n33577 = n33453 & n76321 ;
  assign n33578 = n33509 & n33577 ;
  assign n33579 = n33576 | n33578 ;
  assign n33580 = n65686 & n33579 ;
  assign n33512 = n840 & n76324 ;
  assign n33581 = x64 & n76324 ;
  assign n76338 = ~n33581 ;
  assign n33582 = x55 & n76338 ;
  assign n33583 = n33512 | n33582 ;
  assign n33585 = x65 & n33583 ;
  assign n33584 = x65 | n33512 ;
  assign n33586 = n33582 | n33584 ;
  assign n76339 = ~n33585 ;
  assign n33587 = n76339 & n33586 ;
  assign n33588 = n990 | n33587 ;
  assign n33589 = n65670 & n33583 ;
  assign n76340 = ~n33589 ;
  assign n33590 = n33588 & n76340 ;
  assign n76341 = ~n33578 ;
  assign n33591 = x66 & n76341 ;
  assign n76342 = ~n33576 ;
  assign n33592 = n76342 & n33591 ;
  assign n33593 = n33580 | n33592 ;
  assign n33594 = n33590 | n33593 ;
  assign n76343 = ~n33580 ;
  assign n33595 = n76343 & n33594 ;
  assign n76344 = ~n33570 ;
  assign n33596 = x67 & n76344 ;
  assign n76345 = ~n33568 ;
  assign n33597 = n76345 & n33596 ;
  assign n33598 = n33572 | n33597 ;
  assign n33599 = n33595 | n33598 ;
  assign n76346 = ~n33572 ;
  assign n33600 = n76346 & n33599 ;
  assign n76347 = ~n33562 ;
  assign n33601 = x68 & n76347 ;
  assign n76348 = ~n33560 ;
  assign n33602 = n76348 & n33601 ;
  assign n33603 = n33564 | n33602 ;
  assign n33604 = n33600 | n33603 ;
  assign n76349 = ~n33564 ;
  assign n33605 = n76349 & n33604 ;
  assign n76350 = ~n33554 ;
  assign n33606 = x69 & n76350 ;
  assign n76351 = ~n33552 ;
  assign n33607 = n76351 & n33606 ;
  assign n33608 = n33556 | n33607 ;
  assign n33610 = n33605 | n33608 ;
  assign n76352 = ~n33556 ;
  assign n33611 = n76352 & n33610 ;
  assign n76353 = ~n33546 ;
  assign n33612 = x70 & n76353 ;
  assign n76354 = ~n33544 ;
  assign n33613 = n76354 & n33612 ;
  assign n33614 = n33548 | n33613 ;
  assign n33615 = n33611 | n33614 ;
  assign n76355 = ~n33548 ;
  assign n33616 = n76355 & n33615 ;
  assign n76356 = ~n33537 ;
  assign n33617 = x71 & n76356 ;
  assign n76357 = ~n33535 ;
  assign n33618 = n76357 & n33617 ;
  assign n33619 = n33539 | n33618 ;
  assign n33621 = n33616 | n33619 ;
  assign n76358 = ~n33539 ;
  assign n33622 = n76358 & n33621 ;
  assign n76359 = ~n33518 ;
  assign n33623 = x72 & n76359 ;
  assign n76360 = ~n33516 ;
  assign n33624 = n76360 & n33623 ;
  assign n33625 = n33531 | n33624 ;
  assign n33626 = n33622 | n33625 ;
  assign n76361 = ~n33531 ;
  assign n33627 = n76361 & n33626 ;
  assign n76362 = ~n33528 ;
  assign n33628 = x73 & n76362 ;
  assign n76363 = ~n33526 ;
  assign n33629 = n76363 & n33628 ;
  assign n33630 = n33530 | n33629 ;
  assign n33632 = n33627 | n33630 ;
  assign n76364 = ~n33530 ;
  assign n33633 = n76364 & n33632 ;
  assign n33634 = n1041 | n33633 ;
  assign n76365 = ~n33529 ;
  assign n33635 = n76365 & n33634 ;
  assign n76366 = ~n33627 ;
  assign n33631 = n76366 & n33630 ;
  assign n33648 = n33531 | n33630 ;
  assign n76367 = ~n33648 ;
  assign n33649 = n33626 & n76367 ;
  assign n33650 = n33631 | n33649 ;
  assign n33651 = n33634 | n33650 ;
  assign n76368 = ~n33635 ;
  assign n33652 = n76368 & n33651 ;
  assign n33653 = n65960 & n33652 ;
  assign n76369 = ~n33634 ;
  assign n33765 = n76369 & n33650 ;
  assign n33766 = n33529 & n33634 ;
  assign n76370 = ~n33766 ;
  assign n33767 = x74 & n76370 ;
  assign n76371 = ~n33765 ;
  assign n33768 = n76371 & n33767 ;
  assign n33769 = n33653 | n33768 ;
  assign n33636 = n33519 & n33634 ;
  assign n76372 = ~n33622 ;
  assign n33641 = n76372 & n33625 ;
  assign n33642 = n33539 | n33625 ;
  assign n76373 = ~n33642 ;
  assign n33643 = n33621 & n76373 ;
  assign n33644 = n33641 | n33643 ;
  assign n33645 = n65954 & n33644 ;
  assign n76374 = ~n33633 ;
  assign n33646 = n76374 & n33645 ;
  assign n33647 = n33636 | n33646 ;
  assign n33654 = n65909 & n33647 ;
  assign n33655 = n33538 & n33634 ;
  assign n76375 = ~n33616 ;
  assign n33620 = n76375 & n33619 ;
  assign n33656 = n33548 | n33619 ;
  assign n76376 = ~n33656 ;
  assign n33657 = n33615 & n76376 ;
  assign n33658 = n33620 | n33657 ;
  assign n33659 = n65954 & n33658 ;
  assign n33660 = n76374 & n33659 ;
  assign n33661 = n33655 | n33660 ;
  assign n33662 = n65877 & n33661 ;
  assign n76377 = ~n33660 ;
  assign n33753 = x72 & n76377 ;
  assign n76378 = ~n33655 ;
  assign n33754 = n76378 & n33753 ;
  assign n33755 = n33662 | n33754 ;
  assign n33663 = n33547 & n33634 ;
  assign n76379 = ~n33611 ;
  assign n33640 = n76379 & n33614 ;
  assign n33664 = n33556 | n33614 ;
  assign n76380 = ~n33664 ;
  assign n33665 = n33610 & n76380 ;
  assign n33666 = n33640 | n33665 ;
  assign n33667 = n65954 & n33666 ;
  assign n33668 = n76374 & n33667 ;
  assign n33669 = n33663 | n33668 ;
  assign n33670 = n65820 & n33669 ;
  assign n33671 = n33555 & n33634 ;
  assign n76381 = ~n33605 ;
  assign n33609 = n76381 & n33608 ;
  assign n33672 = n33564 | n33608 ;
  assign n76382 = ~n33672 ;
  assign n33673 = n33604 & n76382 ;
  assign n33674 = n33609 | n33673 ;
  assign n33675 = n65954 & n33674 ;
  assign n33676 = n76374 & n33675 ;
  assign n33677 = n33671 | n33676 ;
  assign n33678 = n65791 & n33677 ;
  assign n76383 = ~n33676 ;
  assign n33742 = x70 & n76383 ;
  assign n76384 = ~n33671 ;
  assign n33743 = n76384 & n33742 ;
  assign n33744 = n33678 | n33743 ;
  assign n33679 = n33563 & n33634 ;
  assign n76385 = ~n33600 ;
  assign n33639 = n76385 & n33603 ;
  assign n33680 = n33572 | n33603 ;
  assign n76386 = ~n33680 ;
  assign n33681 = n33599 & n76386 ;
  assign n33682 = n33639 | n33681 ;
  assign n33683 = n65954 & n33682 ;
  assign n33684 = n76374 & n33683 ;
  assign n33685 = n33679 | n33684 ;
  assign n33686 = n65772 & n33685 ;
  assign n33687 = n33571 & n33634 ;
  assign n76387 = ~n33595 ;
  assign n33638 = n76387 & n33598 ;
  assign n33688 = n33580 | n33598 ;
  assign n76388 = ~n33688 ;
  assign n33689 = n33594 & n76388 ;
  assign n33690 = n33638 | n33689 ;
  assign n33691 = n65954 & n33690 ;
  assign n33692 = n76374 & n33691 ;
  assign n33693 = n33687 | n33692 ;
  assign n33694 = n65746 & n33693 ;
  assign n76389 = ~n33692 ;
  assign n33732 = x68 & n76389 ;
  assign n76390 = ~n33687 ;
  assign n33733 = n76390 & n33732 ;
  assign n33734 = n33694 | n33733 ;
  assign n33637 = n33579 & n33634 ;
  assign n33695 = n33589 | n33593 ;
  assign n76391 = ~n33695 ;
  assign n33696 = n33588 & n76391 ;
  assign n76392 = ~n33590 ;
  assign n33697 = n76392 & n33593 ;
  assign n33698 = n33696 | n33697 ;
  assign n33699 = n65954 & n33698 ;
  assign n33700 = n76374 & n33699 ;
  assign n33701 = n33637 | n33700 ;
  assign n33702 = n65721 & n33701 ;
  assign n33703 = n33583 & n33634 ;
  assign n33704 = n990 & n33586 ;
  assign n33705 = n76339 & n33704 ;
  assign n33706 = n1041 | n33705 ;
  assign n76393 = ~n33706 ;
  assign n33707 = n33588 & n76393 ;
  assign n33708 = n76374 & n33707 ;
  assign n33709 = n33703 | n33708 ;
  assign n33710 = n65686 & n33709 ;
  assign n76394 = ~n33708 ;
  assign n33722 = x66 & n76394 ;
  assign n76395 = ~n33703 ;
  assign n33723 = n76395 & n33722 ;
  assign n33724 = n33710 | n33723 ;
  assign n33711 = n1141 & n76374 ;
  assign n76396 = ~n33711 ;
  assign n33712 = x54 & n76396 ;
  assign n33713 = n1146 & n76374 ;
  assign n33714 = n33712 | n33713 ;
  assign n33715 = x65 & n33714 ;
  assign n33716 = x65 | n33713 ;
  assign n33717 = n33712 | n33716 ;
  assign n76397 = ~n33715 ;
  assign n33718 = n76397 & n33717 ;
  assign n33720 = n1161 | n33718 ;
  assign n33721 = n65670 & n33714 ;
  assign n76398 = ~n33721 ;
  assign n33725 = n33720 & n76398 ;
  assign n33726 = n33724 | n33725 ;
  assign n76399 = ~n33710 ;
  assign n33727 = n76399 & n33726 ;
  assign n76400 = ~n33700 ;
  assign n33728 = x67 & n76400 ;
  assign n76401 = ~n33637 ;
  assign n33729 = n76401 & n33728 ;
  assign n33730 = n33702 | n33729 ;
  assign n33731 = n33727 | n33730 ;
  assign n76402 = ~n33702 ;
  assign n33735 = n76402 & n33731 ;
  assign n33736 = n33734 | n33735 ;
  assign n76403 = ~n33694 ;
  assign n33737 = n76403 & n33736 ;
  assign n76404 = ~n33684 ;
  assign n33738 = x69 & n76404 ;
  assign n76405 = ~n33679 ;
  assign n33739 = n76405 & n33738 ;
  assign n33740 = n33686 | n33739 ;
  assign n33741 = n33737 | n33740 ;
  assign n76406 = ~n33686 ;
  assign n33745 = n76406 & n33741 ;
  assign n33746 = n33744 | n33745 ;
  assign n76407 = ~n33678 ;
  assign n33747 = n76407 & n33746 ;
  assign n76408 = ~n33668 ;
  assign n33748 = x71 & n76408 ;
  assign n76409 = ~n33663 ;
  assign n33749 = n76409 & n33748 ;
  assign n33750 = n33670 | n33749 ;
  assign n33752 = n33747 | n33750 ;
  assign n76410 = ~n33670 ;
  assign n33757 = n76410 & n33752 ;
  assign n33758 = n33755 | n33757 ;
  assign n76411 = ~n33662 ;
  assign n33759 = n76411 & n33758 ;
  assign n76412 = ~n33646 ;
  assign n33760 = x73 & n76412 ;
  assign n76413 = ~n33636 ;
  assign n33761 = n76413 & n33760 ;
  assign n33762 = n33654 | n33761 ;
  assign n33764 = n33759 | n33762 ;
  assign n76414 = ~n33654 ;
  assign n33770 = n76414 & n33764 ;
  assign n33771 = n33769 | n33770 ;
  assign n76415 = ~n33653 ;
  assign n33772 = n76415 & n33771 ;
  assign n33773 = n1214 | n33772 ;
  assign n76416 = ~n33652 ;
  assign n33775 = n76416 & n33773 ;
  assign n76417 = ~n33770 ;
  assign n33909 = n33769 & n76417 ;
  assign n33910 = n33654 | n33769 ;
  assign n76418 = ~n33910 ;
  assign n33911 = n33764 & n76418 ;
  assign n33912 = n33909 | n33911 ;
  assign n33913 = n33773 | n33912 ;
  assign n76419 = ~n33775 ;
  assign n33914 = n76419 & n33913 ;
  assign n33922 = n66016 & n33914 ;
  assign n33776 = n33647 & n33773 ;
  assign n33763 = n33662 | n33762 ;
  assign n76420 = ~n33763 ;
  assign n33778 = n33758 & n76420 ;
  assign n76421 = ~n33759 ;
  assign n33779 = n76421 & n33762 ;
  assign n33780 = n33778 | n33779 ;
  assign n33781 = n66016 & n33780 ;
  assign n76422 = ~n33772 ;
  assign n33782 = n76422 & n33781 ;
  assign n33783 = n33776 | n33782 ;
  assign n33784 = n65960 & n33783 ;
  assign n33785 = n33661 & n33773 ;
  assign n33756 = n33670 | n33755 ;
  assign n76423 = ~n33756 ;
  assign n33786 = n33752 & n76423 ;
  assign n76424 = ~n33757 ;
  assign n33787 = n33755 & n76424 ;
  assign n33788 = n33786 | n33787 ;
  assign n33789 = n66016 & n33788 ;
  assign n33790 = n76422 & n33789 ;
  assign n33791 = n33785 | n33790 ;
  assign n33792 = n65909 & n33791 ;
  assign n33793 = n33669 & n33773 ;
  assign n33751 = n33678 | n33750 ;
  assign n76425 = ~n33751 ;
  assign n33794 = n33746 & n76425 ;
  assign n76426 = ~n33747 ;
  assign n33795 = n76426 & n33750 ;
  assign n33796 = n33794 | n33795 ;
  assign n33797 = n66016 & n33796 ;
  assign n33798 = n76422 & n33797 ;
  assign n33799 = n33793 | n33798 ;
  assign n33800 = n65877 & n33799 ;
  assign n33801 = n33677 & n33773 ;
  assign n33777 = n33686 | n33744 ;
  assign n76427 = ~n33777 ;
  assign n33802 = n33741 & n76427 ;
  assign n76428 = ~n33745 ;
  assign n33803 = n33744 & n76428 ;
  assign n33804 = n33802 | n33803 ;
  assign n33805 = n66016 & n33804 ;
  assign n33806 = n76422 & n33805 ;
  assign n33807 = n33801 | n33806 ;
  assign n33808 = n65820 & n33807 ;
  assign n33809 = n33685 & n33773 ;
  assign n33810 = n33694 | n33740 ;
  assign n76429 = ~n33810 ;
  assign n33811 = n33736 & n76429 ;
  assign n76430 = ~n33737 ;
  assign n33812 = n76430 & n33740 ;
  assign n33813 = n33811 | n33812 ;
  assign n33814 = n66016 & n33813 ;
  assign n33815 = n76422 & n33814 ;
  assign n33816 = n33809 | n33815 ;
  assign n33817 = n65791 & n33816 ;
  assign n33818 = n33693 & n33773 ;
  assign n33819 = n33702 | n33734 ;
  assign n76431 = ~n33819 ;
  assign n33820 = n33731 & n76431 ;
  assign n76432 = ~n33735 ;
  assign n33821 = n33734 & n76432 ;
  assign n33822 = n33820 | n33821 ;
  assign n33823 = n66016 & n33822 ;
  assign n33824 = n76422 & n33823 ;
  assign n33825 = n33818 | n33824 ;
  assign n33826 = n65772 & n33825 ;
  assign n33827 = n33701 & n33773 ;
  assign n33828 = n33710 | n33730 ;
  assign n76433 = ~n33828 ;
  assign n33829 = n33726 & n76433 ;
  assign n76434 = ~n33727 ;
  assign n33830 = n76434 & n33730 ;
  assign n33831 = n33829 | n33830 ;
  assign n33832 = n66016 & n33831 ;
  assign n33833 = n76422 & n33832 ;
  assign n33834 = n33827 | n33833 ;
  assign n33835 = n65746 & n33834 ;
  assign n33836 = n33709 & n33773 ;
  assign n76435 = ~n33725 ;
  assign n33837 = n33724 & n76435 ;
  assign n33838 = n33721 | n33724 ;
  assign n76436 = ~n33838 ;
  assign n33839 = n33720 & n76436 ;
  assign n33840 = n33837 | n33839 ;
  assign n33841 = n66016 & n33840 ;
  assign n33842 = n76422 & n33841 ;
  assign n33843 = n33836 | n33842 ;
  assign n33844 = n65721 & n33843 ;
  assign n33774 = n33714 & n33773 ;
  assign n33719 = n1161 & n33717 ;
  assign n33845 = n76397 & n33719 ;
  assign n33846 = n1214 | n33845 ;
  assign n76437 = ~n33846 ;
  assign n33847 = n33720 & n76437 ;
  assign n33848 = n76422 & n33847 ;
  assign n33849 = n33774 | n33848 ;
  assign n33850 = n65686 & n33849 ;
  assign n33851 = n1323 & n76422 ;
  assign n33852 = n1317 & n76422 ;
  assign n76438 = ~n33852 ;
  assign n33853 = x53 & n76438 ;
  assign n33854 = n33851 | n33853 ;
  assign n33859 = n65670 & n33854 ;
  assign n33855 = x65 & n33854 ;
  assign n33856 = x65 | n33851 ;
  assign n33857 = n33853 | n33856 ;
  assign n76439 = ~n33855 ;
  assign n33858 = n76439 & n33857 ;
  assign n33860 = n1337 | n33858 ;
  assign n76440 = ~n33859 ;
  assign n33861 = n76440 & n33860 ;
  assign n76441 = ~n33848 ;
  assign n33862 = x66 & n76441 ;
  assign n76442 = ~n33774 ;
  assign n33863 = n76442 & n33862 ;
  assign n33864 = n33861 | n33863 ;
  assign n76443 = ~n33850 ;
  assign n33865 = n76443 & n33864 ;
  assign n76444 = ~n33842 ;
  assign n33866 = x67 & n76444 ;
  assign n76445 = ~n33836 ;
  assign n33867 = n76445 & n33866 ;
  assign n33868 = n33844 | n33867 ;
  assign n33869 = n33865 | n33868 ;
  assign n76446 = ~n33844 ;
  assign n33870 = n76446 & n33869 ;
  assign n76447 = ~n33833 ;
  assign n33871 = x68 & n76447 ;
  assign n76448 = ~n33827 ;
  assign n33872 = n76448 & n33871 ;
  assign n33873 = n33835 | n33872 ;
  assign n33874 = n33870 | n33873 ;
  assign n76449 = ~n33835 ;
  assign n33875 = n76449 & n33874 ;
  assign n76450 = ~n33824 ;
  assign n33876 = x69 & n76450 ;
  assign n76451 = ~n33818 ;
  assign n33877 = n76451 & n33876 ;
  assign n33878 = n33826 | n33877 ;
  assign n33879 = n33875 | n33878 ;
  assign n76452 = ~n33826 ;
  assign n33880 = n76452 & n33879 ;
  assign n76453 = ~n33815 ;
  assign n33881 = x70 & n76453 ;
  assign n76454 = ~n33809 ;
  assign n33882 = n76454 & n33881 ;
  assign n33883 = n33817 | n33882 ;
  assign n33885 = n33880 | n33883 ;
  assign n76455 = ~n33817 ;
  assign n33886 = n76455 & n33885 ;
  assign n76456 = ~n33806 ;
  assign n33887 = x71 & n76456 ;
  assign n76457 = ~n33801 ;
  assign n33888 = n76457 & n33887 ;
  assign n33889 = n33808 | n33888 ;
  assign n33890 = n33886 | n33889 ;
  assign n76458 = ~n33808 ;
  assign n33891 = n76458 & n33890 ;
  assign n76459 = ~n33798 ;
  assign n33892 = x72 & n76459 ;
  assign n76460 = ~n33793 ;
  assign n33893 = n76460 & n33892 ;
  assign n33894 = n33800 | n33893 ;
  assign n33896 = n33891 | n33894 ;
  assign n76461 = ~n33800 ;
  assign n33897 = n76461 & n33896 ;
  assign n76462 = ~n33790 ;
  assign n33898 = x73 & n76462 ;
  assign n76463 = ~n33785 ;
  assign n33899 = n76463 & n33898 ;
  assign n33900 = n33792 | n33899 ;
  assign n33901 = n33897 | n33900 ;
  assign n76464 = ~n33792 ;
  assign n33902 = n76464 & n33901 ;
  assign n76465 = ~n33782 ;
  assign n33903 = x74 & n76465 ;
  assign n76466 = ~n33776 ;
  assign n33904 = n76466 & n33903 ;
  assign n33905 = n33784 | n33904 ;
  assign n33907 = n33902 | n33905 ;
  assign n76467 = ~n33784 ;
  assign n33908 = n76467 & n33907 ;
  assign n33915 = n66043 & n33914 ;
  assign n76468 = ~n33773 ;
  assign n33916 = n76468 & n33912 ;
  assign n33917 = n33652 & n33773 ;
  assign n76469 = ~n33917 ;
  assign n33918 = x75 & n76469 ;
  assign n76470 = ~n33916 ;
  assign n33919 = n76470 & n33918 ;
  assign n33920 = n1405 | n33919 ;
  assign n33921 = n33915 | n33920 ;
  assign n33923 = n33908 | n33921 ;
  assign n76471 = ~n33922 ;
  assign n33924 = n76471 & n33923 ;
  assign n76472 = ~n33902 ;
  assign n33906 = n76472 & n33905 ;
  assign n33927 = n33850 | n33863 ;
  assign n33929 = n33861 | n33927 ;
  assign n33930 = n76443 & n33929 ;
  assign n33931 = n33867 | n33930 ;
  assign n33933 = n76446 & n33931 ;
  assign n33935 = n33873 | n33933 ;
  assign n33936 = n76449 & n33935 ;
  assign n33938 = n33878 | n33936 ;
  assign n33939 = n76452 & n33938 ;
  assign n33940 = n33883 | n33939 ;
  assign n33941 = n76455 & n33940 ;
  assign n33942 = n33889 | n33941 ;
  assign n33944 = n76458 & n33942 ;
  assign n33945 = n33894 | n33944 ;
  assign n33946 = n76461 & n33945 ;
  assign n33947 = n33900 | n33946 ;
  assign n33949 = n33792 | n33905 ;
  assign n76473 = ~n33949 ;
  assign n33950 = n33947 & n76473 ;
  assign n33951 = n33906 | n33950 ;
  assign n76474 = ~n33924 ;
  assign n33952 = n76474 & n33951 ;
  assign n33953 = n76464 & n33947 ;
  assign n33954 = n33905 | n33953 ;
  assign n33955 = n76467 & n33954 ;
  assign n33956 = n33921 | n33955 ;
  assign n33957 = n33783 & n76471 ;
  assign n33958 = n33956 & n33957 ;
  assign n33959 = n33952 | n33958 ;
  assign n33960 = n33784 | n33919 ;
  assign n33961 = n33915 | n33960 ;
  assign n76475 = ~n33961 ;
  assign n33962 = n33907 & n76475 ;
  assign n33963 = n33915 | n33919 ;
  assign n76476 = ~n33955 ;
  assign n33964 = n76476 & n33963 ;
  assign n33965 = n33962 | n33964 ;
  assign n33966 = n76474 & n33965 ;
  assign n33967 = n1214 & n33652 ;
  assign n33968 = n33956 & n33967 ;
  assign n33969 = n33966 | n33968 ;
  assign n33970 = n66081 & n33969 ;
  assign n76477 = ~n33968 ;
  assign n34113 = x76 & n76477 ;
  assign n76478 = ~n33966 ;
  assign n34114 = n76478 & n34113 ;
  assign n34115 = n33970 | n34114 ;
  assign n33971 = n66043 & n33959 ;
  assign n76479 = ~n33946 ;
  assign n33948 = n33900 & n76479 ;
  assign n33972 = n33800 | n33900 ;
  assign n76480 = ~n33972 ;
  assign n33973 = n33896 & n76480 ;
  assign n33974 = n33948 | n33973 ;
  assign n33975 = n76474 & n33974 ;
  assign n33976 = n33791 & n76471 ;
  assign n33977 = n33956 & n33976 ;
  assign n33978 = n33975 | n33977 ;
  assign n33979 = n65960 & n33978 ;
  assign n76481 = ~n33977 ;
  assign n34101 = x74 & n76481 ;
  assign n76482 = ~n33975 ;
  assign n34102 = n76482 & n34101 ;
  assign n34103 = n33979 | n34102 ;
  assign n76483 = ~n33891 ;
  assign n33895 = n76483 & n33894 ;
  assign n33980 = n33808 | n33894 ;
  assign n76484 = ~n33980 ;
  assign n33981 = n33942 & n76484 ;
  assign n33982 = n33895 | n33981 ;
  assign n33983 = n76474 & n33982 ;
  assign n33984 = n33799 & n76471 ;
  assign n33985 = n33956 & n33984 ;
  assign n33986 = n33983 | n33985 ;
  assign n33987 = n65909 & n33986 ;
  assign n76485 = ~n33941 ;
  assign n33943 = n33889 & n76485 ;
  assign n33988 = n33817 | n33889 ;
  assign n76486 = ~n33988 ;
  assign n33989 = n33885 & n76486 ;
  assign n33990 = n33943 | n33989 ;
  assign n33991 = n76474 & n33990 ;
  assign n33992 = n33807 & n76471 ;
  assign n33993 = n33956 & n33992 ;
  assign n33994 = n33991 | n33993 ;
  assign n33995 = n65877 & n33994 ;
  assign n76487 = ~n33993 ;
  assign n34089 = x72 & n76487 ;
  assign n76488 = ~n33991 ;
  assign n34090 = n76488 & n34089 ;
  assign n34091 = n33995 | n34090 ;
  assign n76489 = ~n33880 ;
  assign n33884 = n76489 & n33883 ;
  assign n33996 = n33826 | n33883 ;
  assign n76490 = ~n33996 ;
  assign n33997 = n33938 & n76490 ;
  assign n33998 = n33884 | n33997 ;
  assign n33999 = n76474 & n33998 ;
  assign n34000 = n33816 & n76471 ;
  assign n34001 = n33956 & n34000 ;
  assign n34002 = n33999 | n34001 ;
  assign n34003 = n65820 & n34002 ;
  assign n76491 = ~n33936 ;
  assign n33937 = n33878 & n76491 ;
  assign n34004 = n33835 | n33878 ;
  assign n76492 = ~n34004 ;
  assign n34005 = n33874 & n76492 ;
  assign n34006 = n33937 | n34005 ;
  assign n34007 = n76474 & n34006 ;
  assign n34008 = n33825 & n76471 ;
  assign n34009 = n33956 & n34008 ;
  assign n34010 = n34007 | n34009 ;
  assign n34011 = n65791 & n34010 ;
  assign n76493 = ~n34009 ;
  assign n34077 = x70 & n76493 ;
  assign n76494 = ~n34007 ;
  assign n34078 = n76494 & n34077 ;
  assign n34079 = n34011 | n34078 ;
  assign n76495 = ~n33870 ;
  assign n33934 = n76495 & n33873 ;
  assign n34012 = n33868 | n33930 ;
  assign n34013 = n33844 | n33873 ;
  assign n76496 = ~n34013 ;
  assign n34014 = n34012 & n76496 ;
  assign n34015 = n33934 | n34014 ;
  assign n34016 = n76474 & n34015 ;
  assign n34017 = n33834 & n76471 ;
  assign n34018 = n33956 & n34017 ;
  assign n34019 = n34016 | n34018 ;
  assign n34020 = n65772 & n34019 ;
  assign n76497 = ~n33930 ;
  assign n33932 = n33868 & n76497 ;
  assign n34021 = n33850 | n33868 ;
  assign n76498 = ~n34021 ;
  assign n34022 = n33929 & n76498 ;
  assign n34023 = n33932 | n34022 ;
  assign n34024 = n76474 & n34023 ;
  assign n34025 = n33843 & n76471 ;
  assign n34026 = n33956 & n34025 ;
  assign n34027 = n34024 | n34026 ;
  assign n34028 = n65746 & n34027 ;
  assign n76499 = ~n34026 ;
  assign n34066 = x68 & n76499 ;
  assign n76500 = ~n34024 ;
  assign n34067 = n76500 & n34066 ;
  assign n34068 = n34028 | n34067 ;
  assign n76501 = ~n33861 ;
  assign n33928 = n76501 & n33927 ;
  assign n34029 = n33859 | n33927 ;
  assign n76502 = ~n34029 ;
  assign n34030 = n33860 & n76502 ;
  assign n34031 = n33928 | n34030 ;
  assign n34032 = n76474 & n34031 ;
  assign n34033 = n33849 & n76471 ;
  assign n34034 = n33956 & n34033 ;
  assign n34035 = n34032 | n34034 ;
  assign n34036 = n65721 & n34035 ;
  assign n34037 = n1337 & n33857 ;
  assign n34038 = n76439 & n34037 ;
  assign n76503 = ~n34038 ;
  assign n34039 = n33860 & n76503 ;
  assign n34040 = n76474 & n34039 ;
  assign n34041 = n33854 & n76471 ;
  assign n34042 = n33956 & n34041 ;
  assign n34043 = n34040 | n34042 ;
  assign n34044 = n65686 & n34043 ;
  assign n76504 = ~n34042 ;
  assign n34056 = x66 & n76504 ;
  assign n76505 = ~n34040 ;
  assign n34057 = n76505 & n34056 ;
  assign n34058 = n34044 | n34057 ;
  assign n33926 = n1337 & n76474 ;
  assign n33925 = x64 & n76474 ;
  assign n76506 = ~n33925 ;
  assign n34045 = x52 & n76506 ;
  assign n34046 = n33926 | n34045 ;
  assign n34047 = x65 & n34046 ;
  assign n34048 = n76471 & n33956 ;
  assign n76507 = ~n34048 ;
  assign n34049 = n1337 & n76507 ;
  assign n34050 = x65 | n34049 ;
  assign n34051 = n34045 | n34050 ;
  assign n76508 = ~n34047 ;
  assign n34052 = n76508 & n34051 ;
  assign n34054 = n1547 | n34052 ;
  assign n34055 = n65670 & n34046 ;
  assign n76509 = ~n34055 ;
  assign n34059 = n34054 & n76509 ;
  assign n34060 = n34058 | n34059 ;
  assign n76510 = ~n34044 ;
  assign n34061 = n76510 & n34060 ;
  assign n76511 = ~n34034 ;
  assign n34062 = x67 & n76511 ;
  assign n76512 = ~n34032 ;
  assign n34063 = n76512 & n34062 ;
  assign n34064 = n34036 | n34063 ;
  assign n34065 = n34061 | n34064 ;
  assign n76513 = ~n34036 ;
  assign n34069 = n76513 & n34065 ;
  assign n34070 = n34068 | n34069 ;
  assign n76514 = ~n34028 ;
  assign n34071 = n76514 & n34070 ;
  assign n76515 = ~n34018 ;
  assign n34072 = x69 & n76515 ;
  assign n76516 = ~n34016 ;
  assign n34073 = n76516 & n34072 ;
  assign n34074 = n34020 | n34073 ;
  assign n34076 = n34071 | n34074 ;
  assign n76517 = ~n34020 ;
  assign n34081 = n76517 & n34076 ;
  assign n34082 = n34079 | n34081 ;
  assign n76518 = ~n34011 ;
  assign n34083 = n76518 & n34082 ;
  assign n76519 = ~n34001 ;
  assign n34084 = x71 & n76519 ;
  assign n76520 = ~n33999 ;
  assign n34085 = n76520 & n34084 ;
  assign n34086 = n34003 | n34085 ;
  assign n34088 = n34083 | n34086 ;
  assign n76521 = ~n34003 ;
  assign n34093 = n76521 & n34088 ;
  assign n34094 = n34091 | n34093 ;
  assign n76522 = ~n33995 ;
  assign n34095 = n76522 & n34094 ;
  assign n76523 = ~n33985 ;
  assign n34096 = x73 & n76523 ;
  assign n76524 = ~n33983 ;
  assign n34097 = n76524 & n34096 ;
  assign n34098 = n33987 | n34097 ;
  assign n34100 = n34095 | n34098 ;
  assign n76525 = ~n33987 ;
  assign n34105 = n76525 & n34100 ;
  assign n34106 = n34103 | n34105 ;
  assign n76526 = ~n33979 ;
  assign n34107 = n76526 & n34106 ;
  assign n76527 = ~n33958 ;
  assign n34108 = x75 & n76527 ;
  assign n76528 = ~n33952 ;
  assign n34109 = n76528 & n34108 ;
  assign n34110 = n33971 | n34109 ;
  assign n34112 = n34107 | n34110 ;
  assign n76529 = ~n33971 ;
  assign n34116 = n76529 & n34112 ;
  assign n34117 = n34115 | n34116 ;
  assign n76530 = ~n33970 ;
  assign n34118 = n76530 & n34117 ;
  assign n34119 = n1611 | n34118 ;
  assign n34122 = n33959 & n34119 ;
  assign n34111 = n33979 | n34110 ;
  assign n34124 = x64 & n76507 ;
  assign n76531 = ~n34124 ;
  assign n34125 = x52 & n76531 ;
  assign n34126 = n33926 | n34125 ;
  assign n34127 = x65 & n34126 ;
  assign n76532 = ~n34127 ;
  assign n34128 = n34051 & n76532 ;
  assign n34129 = n1547 | n34128 ;
  assign n34130 = n76509 & n34129 ;
  assign n34132 = n34058 | n34130 ;
  assign n34133 = n76510 & n34132 ;
  assign n34134 = n34064 | n34133 ;
  assign n34135 = n76513 & n34134 ;
  assign n34136 = n34068 | n34135 ;
  assign n34137 = n76514 & n34136 ;
  assign n34138 = n34074 | n34137 ;
  assign n34139 = n76517 & n34138 ;
  assign n34140 = n34079 | n34139 ;
  assign n34141 = n76518 & n34140 ;
  assign n34142 = n34086 | n34141 ;
  assign n34143 = n76521 & n34142 ;
  assign n34144 = n34091 | n34143 ;
  assign n34145 = n76522 & n34144 ;
  assign n34146 = n34098 | n34145 ;
  assign n34147 = n76525 & n34146 ;
  assign n34148 = n34103 | n34147 ;
  assign n76533 = ~n34111 ;
  assign n34149 = n76533 & n34148 ;
  assign n76534 = ~n34107 ;
  assign n34150 = n76534 & n34110 ;
  assign n34151 = n34149 | n34150 ;
  assign n34152 = n66151 & n34151 ;
  assign n76535 = ~n34118 ;
  assign n34153 = n76535 & n34152 ;
  assign n34154 = n34122 | n34153 ;
  assign n76536 = ~n33969 ;
  assign n34121 = n76536 & n34119 ;
  assign n76537 = ~n34116 ;
  assign n34158 = n34115 & n76537 ;
  assign n34155 = n76526 & n34148 ;
  assign n34156 = n34110 | n34155 ;
  assign n34159 = n33971 | n34115 ;
  assign n76538 = ~n34159 ;
  assign n34160 = n34156 & n76538 ;
  assign n34161 = n34158 | n34160 ;
  assign n34162 = n34119 | n34161 ;
  assign n76539 = ~n34121 ;
  assign n34163 = n76539 & n34162 ;
  assign n34164 = n66145 & n34163 ;
  assign n34165 = n66081 & n34154 ;
  assign n34166 = n33978 & n34119 ;
  assign n34104 = n33987 | n34103 ;
  assign n76540 = ~n34104 ;
  assign n34167 = n34100 & n76540 ;
  assign n76541 = ~n34147 ;
  assign n34168 = n34103 & n76541 ;
  assign n34169 = n34167 | n34168 ;
  assign n34170 = n66151 & n34169 ;
  assign n34171 = n76535 & n34170 ;
  assign n34172 = n34166 | n34171 ;
  assign n34173 = n66043 & n34172 ;
  assign n34174 = n33986 & n34119 ;
  assign n34099 = n33995 | n34098 ;
  assign n76542 = ~n34099 ;
  assign n34175 = n76542 & n34144 ;
  assign n76543 = ~n34095 ;
  assign n34176 = n76543 & n34098 ;
  assign n34177 = n34175 | n34176 ;
  assign n34178 = n66151 & n34177 ;
  assign n34179 = n76535 & n34178 ;
  assign n34180 = n34174 | n34179 ;
  assign n34181 = n65960 & n34180 ;
  assign n34182 = n33994 & n34119 ;
  assign n34092 = n34003 | n34091 ;
  assign n76544 = ~n34092 ;
  assign n34183 = n34088 & n76544 ;
  assign n76545 = ~n34143 ;
  assign n34184 = n34091 & n76545 ;
  assign n34185 = n34183 | n34184 ;
  assign n34186 = n66151 & n34185 ;
  assign n34187 = n76535 & n34186 ;
  assign n34188 = n34182 | n34187 ;
  assign n34189 = n65909 & n34188 ;
  assign n34190 = n34002 & n34119 ;
  assign n34087 = n34011 | n34086 ;
  assign n76546 = ~n34087 ;
  assign n34191 = n76546 & n34140 ;
  assign n76547 = ~n34083 ;
  assign n34192 = n76547 & n34086 ;
  assign n34193 = n34191 | n34192 ;
  assign n34194 = n66151 & n34193 ;
  assign n34195 = n76535 & n34194 ;
  assign n34196 = n34190 | n34195 ;
  assign n34197 = n65877 & n34196 ;
  assign n34198 = n34010 & n34119 ;
  assign n34080 = n34020 | n34079 ;
  assign n76548 = ~n34080 ;
  assign n34199 = n34076 & n76548 ;
  assign n76549 = ~n34139 ;
  assign n34200 = n34079 & n76549 ;
  assign n34201 = n34199 | n34200 ;
  assign n34202 = n66151 & n34201 ;
  assign n34203 = n76535 & n34202 ;
  assign n34204 = n34198 | n34203 ;
  assign n34205 = n65820 & n34204 ;
  assign n34206 = n34019 & n34119 ;
  assign n34075 = n34028 | n34074 ;
  assign n76550 = ~n34075 ;
  assign n34207 = n76550 & n34136 ;
  assign n76551 = ~n34071 ;
  assign n34208 = n76551 & n34074 ;
  assign n34209 = n34207 | n34208 ;
  assign n34210 = n66151 & n34209 ;
  assign n34211 = n76535 & n34210 ;
  assign n34212 = n34206 | n34211 ;
  assign n34213 = n65791 & n34212 ;
  assign n34214 = n34027 & n34119 ;
  assign n34215 = n34036 | n34068 ;
  assign n76552 = ~n34215 ;
  assign n34216 = n34065 & n76552 ;
  assign n76553 = ~n34135 ;
  assign n34217 = n34068 & n76553 ;
  assign n34218 = n34216 | n34217 ;
  assign n34219 = n66151 & n34218 ;
  assign n34220 = n76535 & n34219 ;
  assign n34221 = n34214 | n34220 ;
  assign n34222 = n65772 & n34221 ;
  assign n34223 = n34035 & n34119 ;
  assign n34224 = n34044 | n34064 ;
  assign n76554 = ~n34224 ;
  assign n34225 = n34060 & n76554 ;
  assign n76555 = ~n34061 ;
  assign n34226 = n76555 & n34064 ;
  assign n34227 = n34225 | n34226 ;
  assign n34228 = n66151 & n34227 ;
  assign n34229 = n76535 & n34228 ;
  assign n34230 = n34223 | n34229 ;
  assign n34231 = n65746 & n34230 ;
  assign n34232 = n34043 & n34119 ;
  assign n34131 = n34055 | n34058 ;
  assign n76556 = ~n34131 ;
  assign n34233 = n34129 & n76556 ;
  assign n76557 = ~n34130 ;
  assign n34234 = n34058 & n76557 ;
  assign n34235 = n34233 | n34234 ;
  assign n34236 = n66151 & n34235 ;
  assign n34237 = n76535 & n34236 ;
  assign n34238 = n34232 | n34237 ;
  assign n34239 = n65721 & n34238 ;
  assign n34120 = n34046 & n34119 ;
  assign n34053 = n1547 & n34051 ;
  assign n34240 = n34053 & n76532 ;
  assign n34241 = n1611 | n34240 ;
  assign n76558 = ~n34241 ;
  assign n34242 = n34129 & n76558 ;
  assign n34243 = n76535 & n34242 ;
  assign n34244 = n34120 | n34243 ;
  assign n34245 = n65686 & n34244 ;
  assign n34123 = n1753 & n76535 ;
  assign n34246 = n1747 & n76535 ;
  assign n76559 = ~n34246 ;
  assign n34247 = x51 & n76559 ;
  assign n34248 = n34123 | n34247 ;
  assign n34249 = n65670 & n34248 ;
  assign n34157 = n76529 & n34156 ;
  assign n34251 = n34115 | n34157 ;
  assign n34252 = n76530 & n34251 ;
  assign n76560 = ~n34252 ;
  assign n34253 = n1747 & n76560 ;
  assign n76561 = ~n34253 ;
  assign n34254 = x51 & n76561 ;
  assign n34255 = n34123 | n34254 ;
  assign n34257 = x65 & n34255 ;
  assign n34256 = x65 | n34123 ;
  assign n34258 = n34247 | n34256 ;
  assign n76562 = ~n34257 ;
  assign n34259 = n76562 & n34258 ;
  assign n34260 = n1761 | n34259 ;
  assign n76563 = ~n34249 ;
  assign n34261 = n76563 & n34260 ;
  assign n76564 = ~n34243 ;
  assign n34262 = x66 & n76564 ;
  assign n76565 = ~n34120 ;
  assign n34263 = n76565 & n34262 ;
  assign n34264 = n34245 | n34263 ;
  assign n34265 = n34261 | n34264 ;
  assign n76566 = ~n34245 ;
  assign n34266 = n76566 & n34265 ;
  assign n76567 = ~n34237 ;
  assign n34267 = x67 & n76567 ;
  assign n76568 = ~n34232 ;
  assign n34268 = n76568 & n34267 ;
  assign n34269 = n34266 | n34268 ;
  assign n76569 = ~n34239 ;
  assign n34270 = n76569 & n34269 ;
  assign n76570 = ~n34229 ;
  assign n34271 = x68 & n76570 ;
  assign n76571 = ~n34223 ;
  assign n34272 = n76571 & n34271 ;
  assign n34273 = n34231 | n34272 ;
  assign n34274 = n34270 | n34273 ;
  assign n76572 = ~n34231 ;
  assign n34275 = n76572 & n34274 ;
  assign n76573 = ~n34220 ;
  assign n34276 = x69 & n76573 ;
  assign n76574 = ~n34214 ;
  assign n34277 = n76574 & n34276 ;
  assign n34278 = n34222 | n34277 ;
  assign n34279 = n34275 | n34278 ;
  assign n76575 = ~n34222 ;
  assign n34280 = n76575 & n34279 ;
  assign n76576 = ~n34211 ;
  assign n34281 = x70 & n76576 ;
  assign n76577 = ~n34206 ;
  assign n34282 = n76577 & n34281 ;
  assign n34283 = n34213 | n34282 ;
  assign n34284 = n34280 | n34283 ;
  assign n76578 = ~n34213 ;
  assign n34285 = n76578 & n34284 ;
  assign n76579 = ~n34203 ;
  assign n34286 = x71 & n76579 ;
  assign n76580 = ~n34198 ;
  assign n34287 = n76580 & n34286 ;
  assign n34288 = n34205 | n34287 ;
  assign n34290 = n34285 | n34288 ;
  assign n76581 = ~n34205 ;
  assign n34291 = n76581 & n34290 ;
  assign n76582 = ~n34195 ;
  assign n34292 = x72 & n76582 ;
  assign n76583 = ~n34190 ;
  assign n34293 = n76583 & n34292 ;
  assign n34294 = n34197 | n34293 ;
  assign n34295 = n34291 | n34294 ;
  assign n76584 = ~n34197 ;
  assign n34296 = n76584 & n34295 ;
  assign n76585 = ~n34187 ;
  assign n34297 = x73 & n76585 ;
  assign n76586 = ~n34182 ;
  assign n34298 = n76586 & n34297 ;
  assign n34299 = n34189 | n34298 ;
  assign n34301 = n34296 | n34299 ;
  assign n76587 = ~n34189 ;
  assign n34302 = n76587 & n34301 ;
  assign n76588 = ~n34179 ;
  assign n34303 = x74 & n76588 ;
  assign n76589 = ~n34174 ;
  assign n34304 = n76589 & n34303 ;
  assign n34305 = n34181 | n34304 ;
  assign n34306 = n34302 | n34305 ;
  assign n76590 = ~n34181 ;
  assign n34307 = n76590 & n34306 ;
  assign n76591 = ~n34171 ;
  assign n34308 = x75 & n76591 ;
  assign n76592 = ~n34166 ;
  assign n34309 = n76592 & n34308 ;
  assign n34310 = n34173 | n34309 ;
  assign n34312 = n34307 | n34310 ;
  assign n76593 = ~n34173 ;
  assign n34313 = n76593 & n34312 ;
  assign n76594 = ~n34153 ;
  assign n34314 = x76 & n76594 ;
  assign n76595 = ~n34122 ;
  assign n34315 = n76595 & n34314 ;
  assign n34316 = n34165 | n34315 ;
  assign n34317 = n34313 | n34316 ;
  assign n76596 = ~n34165 ;
  assign n34318 = n76596 & n34317 ;
  assign n76597 = ~n34119 ;
  assign n34319 = n76597 & n34161 ;
  assign n34320 = n33969 & n34119 ;
  assign n76598 = ~n34320 ;
  assign n34321 = x77 & n76598 ;
  assign n76599 = ~n34319 ;
  assign n34322 = n76599 & n34321 ;
  assign n34323 = n34164 | n34322 ;
  assign n34325 = n34318 | n34323 ;
  assign n76600 = ~n34164 ;
  assign n34326 = n76600 & n34325 ;
  assign n34327 = n1839 | n34326 ;
  assign n34329 = n34154 & n34327 ;
  assign n34331 = n65670 & n34255 ;
  assign n34250 = x65 & n34248 ;
  assign n76601 = ~n34250 ;
  assign n34330 = n76601 & n34258 ;
  assign n34332 = n1761 | n34330 ;
  assign n76602 = ~n34331 ;
  assign n34333 = n76602 & n34332 ;
  assign n34334 = n34264 | n34333 ;
  assign n34335 = n76566 & n34334 ;
  assign n34336 = n34239 | n34268 ;
  assign n34338 = n34335 | n34336 ;
  assign n34339 = n76569 & n34338 ;
  assign n34341 = n34273 | n34339 ;
  assign n34342 = n76572 & n34341 ;
  assign n34344 = n34278 | n34342 ;
  assign n34345 = n76575 & n34344 ;
  assign n34346 = n34283 | n34345 ;
  assign n34348 = n76578 & n34346 ;
  assign n34349 = n34288 | n34348 ;
  assign n34350 = n76581 & n34349 ;
  assign n34351 = n34294 | n34350 ;
  assign n34353 = n76584 & n34351 ;
  assign n34354 = n34299 | n34353 ;
  assign n34355 = n76587 & n34354 ;
  assign n34356 = n34305 | n34355 ;
  assign n34358 = n76590 & n34356 ;
  assign n34359 = n34310 | n34358 ;
  assign n34360 = n76593 & n34359 ;
  assign n76603 = ~n34360 ;
  assign n34361 = n34316 & n76603 ;
  assign n34363 = n34173 | n34316 ;
  assign n76604 = ~n34363 ;
  assign n34364 = n34312 & n76604 ;
  assign n34365 = n34361 | n34364 ;
  assign n34366 = n66219 & n34365 ;
  assign n76605 = ~n34326 ;
  assign n34367 = n76605 & n34366 ;
  assign n34368 = n34329 | n34367 ;
  assign n34369 = n66145 & n34368 ;
  assign n76606 = ~n34367 ;
  assign n34542 = x77 & n76606 ;
  assign n76607 = ~n34329 ;
  assign n34543 = n76607 & n34542 ;
  assign n34544 = n34369 | n34543 ;
  assign n34370 = n34172 & n34327 ;
  assign n76608 = ~n34307 ;
  assign n34311 = n76608 & n34310 ;
  assign n34371 = n34181 | n34310 ;
  assign n76609 = ~n34371 ;
  assign n34372 = n34356 & n76609 ;
  assign n34373 = n34311 | n34372 ;
  assign n34374 = n66219 & n34373 ;
  assign n34375 = n76605 & n34374 ;
  assign n34376 = n34370 | n34375 ;
  assign n34377 = n66081 & n34376 ;
  assign n34378 = n34180 & n34327 ;
  assign n76610 = ~n34355 ;
  assign n34357 = n34305 & n76610 ;
  assign n34379 = n34189 | n34305 ;
  assign n76611 = ~n34379 ;
  assign n34380 = n34301 & n76611 ;
  assign n34381 = n34357 | n34380 ;
  assign n34382 = n66219 & n34381 ;
  assign n34383 = n76605 & n34382 ;
  assign n34384 = n34378 | n34383 ;
  assign n34385 = n66043 & n34384 ;
  assign n76612 = ~n34383 ;
  assign n34530 = x75 & n76612 ;
  assign n76613 = ~n34378 ;
  assign n34531 = n76613 & n34530 ;
  assign n34532 = n34385 | n34531 ;
  assign n34386 = n34188 & n34327 ;
  assign n76614 = ~n34296 ;
  assign n34300 = n76614 & n34299 ;
  assign n34387 = n34197 | n34299 ;
  assign n76615 = ~n34387 ;
  assign n34388 = n34351 & n76615 ;
  assign n34389 = n34300 | n34388 ;
  assign n34390 = n66219 & n34389 ;
  assign n34391 = n76605 & n34390 ;
  assign n34392 = n34386 | n34391 ;
  assign n34393 = n65960 & n34392 ;
  assign n34394 = n34196 & n34327 ;
  assign n76616 = ~n34350 ;
  assign n34352 = n34294 & n76616 ;
  assign n34395 = n34205 | n34294 ;
  assign n76617 = ~n34395 ;
  assign n34396 = n34290 & n76617 ;
  assign n34397 = n34352 | n34396 ;
  assign n34398 = n66219 & n34397 ;
  assign n34399 = n76605 & n34398 ;
  assign n34400 = n34394 | n34399 ;
  assign n34401 = n65909 & n34400 ;
  assign n76618 = ~n34399 ;
  assign n34518 = x73 & n76618 ;
  assign n76619 = ~n34394 ;
  assign n34519 = n76619 & n34518 ;
  assign n34520 = n34401 | n34519 ;
  assign n34402 = n34204 & n34327 ;
  assign n76620 = ~n34285 ;
  assign n34289 = n76620 & n34288 ;
  assign n34403 = n34213 | n34288 ;
  assign n76621 = ~n34403 ;
  assign n34404 = n34346 & n76621 ;
  assign n34405 = n34289 | n34404 ;
  assign n34406 = n66219 & n34405 ;
  assign n34407 = n76605 & n34406 ;
  assign n34408 = n34402 | n34407 ;
  assign n34409 = n65877 & n34408 ;
  assign n34410 = n34212 & n34327 ;
  assign n76622 = ~n34345 ;
  assign n34347 = n34283 & n76622 ;
  assign n34411 = n34222 | n34283 ;
  assign n76623 = ~n34411 ;
  assign n34412 = n34279 & n76623 ;
  assign n34413 = n34347 | n34412 ;
  assign n34414 = n66219 & n34413 ;
  assign n34415 = n76605 & n34414 ;
  assign n34416 = n34410 | n34415 ;
  assign n34417 = n65820 & n34416 ;
  assign n76624 = ~n34415 ;
  assign n34506 = x71 & n76624 ;
  assign n76625 = ~n34410 ;
  assign n34507 = n76625 & n34506 ;
  assign n34508 = n34417 | n34507 ;
  assign n34418 = n34221 & n34327 ;
  assign n76626 = ~n34275 ;
  assign n34343 = n76626 & n34278 ;
  assign n34419 = n34231 | n34278 ;
  assign n76627 = ~n34419 ;
  assign n34420 = n34274 & n76627 ;
  assign n34421 = n34343 | n34420 ;
  assign n34422 = n66219 & n34421 ;
  assign n34423 = n76605 & n34422 ;
  assign n34424 = n34418 | n34423 ;
  assign n34425 = n65791 & n34424 ;
  assign n34426 = n34230 & n34327 ;
  assign n76628 = ~n34339 ;
  assign n34340 = n34273 & n76628 ;
  assign n34427 = n34266 | n34336 ;
  assign n34428 = n34239 | n34273 ;
  assign n76629 = ~n34428 ;
  assign n34429 = n34427 & n76629 ;
  assign n34430 = n34340 | n34429 ;
  assign n34431 = n66219 & n34430 ;
  assign n34432 = n76605 & n34431 ;
  assign n34433 = n34426 | n34432 ;
  assign n34434 = n65772 & n34433 ;
  assign n76630 = ~n34432 ;
  assign n34495 = x69 & n76630 ;
  assign n76631 = ~n34426 ;
  assign n34496 = n76631 & n34495 ;
  assign n34497 = n34434 | n34496 ;
  assign n34435 = n34238 & n34327 ;
  assign n76632 = ~n34266 ;
  assign n34337 = n76632 & n34336 ;
  assign n34436 = n34245 | n34336 ;
  assign n76633 = ~n34436 ;
  assign n34437 = n34265 & n76633 ;
  assign n34438 = n34337 | n34437 ;
  assign n34439 = n66219 & n34438 ;
  assign n34440 = n76605 & n34439 ;
  assign n34441 = n34435 | n34440 ;
  assign n34442 = n65746 & n34441 ;
  assign n34443 = n34244 & n34327 ;
  assign n34444 = n34264 | n34331 ;
  assign n76634 = ~n34444 ;
  assign n34445 = n34332 & n76634 ;
  assign n76635 = ~n34333 ;
  assign n34446 = n34264 & n76635 ;
  assign n34447 = n34445 | n34446 ;
  assign n34448 = n66219 & n34447 ;
  assign n34449 = n76605 & n34448 ;
  assign n34450 = n34443 | n34449 ;
  assign n34451 = n65721 & n34450 ;
  assign n76636 = ~n34449 ;
  assign n34485 = x67 & n76636 ;
  assign n76637 = ~n34443 ;
  assign n34486 = n76637 & n34485 ;
  assign n34487 = n34451 | n34486 ;
  assign n34452 = n34248 & n34327 ;
  assign n34453 = n1761 & n34258 ;
  assign n34454 = n76562 & n34453 ;
  assign n34455 = n1839 | n34454 ;
  assign n76638 = ~n34455 ;
  assign n34456 = n34332 & n76638 ;
  assign n34457 = n76605 & n34456 ;
  assign n34458 = n34452 | n34457 ;
  assign n34459 = n65686 & n34458 ;
  assign n34460 = n1969 & n76605 ;
  assign n76639 = ~n34460 ;
  assign n34461 = x50 & n76639 ;
  assign n34462 = n1982 & n76605 ;
  assign n34463 = n34461 | n34462 ;
  assign n34464 = x65 & n34463 ;
  assign n34362 = n34316 | n34360 ;
  assign n34465 = n76596 & n34362 ;
  assign n34466 = n34323 | n34465 ;
  assign n34467 = n76600 & n34466 ;
  assign n76640 = ~n34467 ;
  assign n34468 = n1969 & n76640 ;
  assign n76641 = ~n34468 ;
  assign n34470 = x50 & n76641 ;
  assign n34471 = x65 | n34462 ;
  assign n34472 = n34470 | n34471 ;
  assign n76642 = ~n34464 ;
  assign n34473 = n76642 & n34472 ;
  assign n34474 = n1989 | n34473 ;
  assign n34475 = n34462 | n34470 ;
  assign n34476 = n65670 & n34475 ;
  assign n76643 = ~n34476 ;
  assign n34477 = n34474 & n76643 ;
  assign n34469 = n1839 | n34467 ;
  assign n34478 = n34255 & n34469 ;
  assign n34479 = n34457 | n34478 ;
  assign n34480 = n65686 & n34479 ;
  assign n76644 = ~n34457 ;
  assign n34481 = x66 & n76644 ;
  assign n76645 = ~n34478 ;
  assign n34482 = n76645 & n34481 ;
  assign n34483 = n34480 | n34482 ;
  assign n34484 = n34477 | n34483 ;
  assign n76646 = ~n34459 ;
  assign n34488 = n76646 & n34484 ;
  assign n34489 = n34487 | n34488 ;
  assign n76647 = ~n34451 ;
  assign n34490 = n76647 & n34489 ;
  assign n76648 = ~n34440 ;
  assign n34491 = x68 & n76648 ;
  assign n76649 = ~n34435 ;
  assign n34492 = n76649 & n34491 ;
  assign n34493 = n34442 | n34492 ;
  assign n34494 = n34490 | n34493 ;
  assign n76650 = ~n34442 ;
  assign n34498 = n76650 & n34494 ;
  assign n34499 = n34497 | n34498 ;
  assign n76651 = ~n34434 ;
  assign n34500 = n76651 & n34499 ;
  assign n76652 = ~n34423 ;
  assign n34501 = x70 & n76652 ;
  assign n76653 = ~n34418 ;
  assign n34502 = n76653 & n34501 ;
  assign n34503 = n34425 | n34502 ;
  assign n34505 = n34500 | n34503 ;
  assign n76654 = ~n34425 ;
  assign n34510 = n76654 & n34505 ;
  assign n34511 = n34508 | n34510 ;
  assign n76655 = ~n34417 ;
  assign n34512 = n76655 & n34511 ;
  assign n76656 = ~n34407 ;
  assign n34513 = x72 & n76656 ;
  assign n76657 = ~n34402 ;
  assign n34514 = n76657 & n34513 ;
  assign n34515 = n34409 | n34514 ;
  assign n34517 = n34512 | n34515 ;
  assign n76658 = ~n34409 ;
  assign n34522 = n76658 & n34517 ;
  assign n34523 = n34520 | n34522 ;
  assign n76659 = ~n34401 ;
  assign n34524 = n76659 & n34523 ;
  assign n76660 = ~n34391 ;
  assign n34525 = x74 & n76660 ;
  assign n76661 = ~n34386 ;
  assign n34526 = n76661 & n34525 ;
  assign n34527 = n34393 | n34526 ;
  assign n34529 = n34524 | n34527 ;
  assign n76662 = ~n34393 ;
  assign n34534 = n76662 & n34529 ;
  assign n34535 = n34532 | n34534 ;
  assign n76663 = ~n34385 ;
  assign n34536 = n76663 & n34535 ;
  assign n76664 = ~n34375 ;
  assign n34537 = x76 & n76664 ;
  assign n76665 = ~n34370 ;
  assign n34538 = n76665 & n34537 ;
  assign n34539 = n34377 | n34538 ;
  assign n34541 = n34536 | n34539 ;
  assign n76666 = ~n34377 ;
  assign n34546 = n76666 & n34541 ;
  assign n34547 = n34544 | n34546 ;
  assign n76667 = ~n34369 ;
  assign n34548 = n76667 & n34547 ;
  assign n76668 = ~n34163 ;
  assign n34328 = n76668 & n34327 ;
  assign n76669 = ~n34318 ;
  assign n34324 = n76669 & n34323 ;
  assign n34549 = n34165 | n34323 ;
  assign n76670 = ~n34549 ;
  assign n34550 = n34362 & n76670 ;
  assign n34551 = n34324 | n34550 ;
  assign n34552 = n34327 | n34551 ;
  assign n76671 = ~n34328 ;
  assign n34553 = n76671 & n34552 ;
  assign n34554 = n66244 & n34553 ;
  assign n76672 = ~n34327 ;
  assign n34555 = n76672 & n34551 ;
  assign n34556 = n34163 & n34327 ;
  assign n76673 = ~n34556 ;
  assign n34557 = x78 & n76673 ;
  assign n76674 = ~n34555 ;
  assign n34558 = n76674 & n34557 ;
  assign n34559 = n2069 | n34558 ;
  assign n34560 = n34554 | n34559 ;
  assign n34561 = n34548 | n34560 ;
  assign n34562 = n66219 & n34553 ;
  assign n76675 = ~n34562 ;
  assign n34563 = n34561 & n76675 ;
  assign n34572 = n34369 | n34558 ;
  assign n34573 = n34554 | n34572 ;
  assign n76676 = ~n34573 ;
  assign n34574 = n34547 & n76676 ;
  assign n76677 = ~n34452 ;
  assign n34578 = n76677 & n34481 ;
  assign n34579 = n34459 | n34578 ;
  assign n34575 = x65 & n34475 ;
  assign n76678 = ~n34575 ;
  assign n34576 = n34472 & n76678 ;
  assign n34577 = n1989 | n34576 ;
  assign n34580 = n76643 & n34577 ;
  assign n34581 = n34579 | n34580 ;
  assign n76679 = ~n34480 ;
  assign n34582 = n76679 & n34581 ;
  assign n34583 = n34487 | n34582 ;
  assign n34584 = n76647 & n34583 ;
  assign n34585 = n34493 | n34584 ;
  assign n34586 = n76650 & n34585 ;
  assign n34587 = n34497 | n34586 ;
  assign n34588 = n76651 & n34587 ;
  assign n34589 = n34503 | n34588 ;
  assign n34590 = n76654 & n34589 ;
  assign n34591 = n34508 | n34590 ;
  assign n34592 = n76655 & n34591 ;
  assign n34593 = n34515 | n34592 ;
  assign n34594 = n76658 & n34593 ;
  assign n34595 = n34520 | n34594 ;
  assign n34596 = n76659 & n34595 ;
  assign n34597 = n34527 | n34596 ;
  assign n34598 = n76662 & n34597 ;
  assign n34599 = n34532 | n34598 ;
  assign n34600 = n76663 & n34599 ;
  assign n34601 = n34539 | n34600 ;
  assign n34602 = n76666 & n34601 ;
  assign n34603 = n34544 | n34602 ;
  assign n34604 = n76667 & n34603 ;
  assign n34605 = n34554 | n34558 ;
  assign n76680 = ~n34604 ;
  assign n34606 = n76680 & n34605 ;
  assign n34607 = n34574 | n34606 ;
  assign n76681 = ~n34563 ;
  assign n34608 = n76681 & n34607 ;
  assign n34609 = n1839 & n34163 ;
  assign n34610 = n34561 & n34609 ;
  assign n34611 = n34608 | n34610 ;
  assign n34612 = n66299 & n34611 ;
  assign n76682 = ~n34546 ;
  assign n34565 = n34544 & n76682 ;
  assign n34545 = n34377 | n34544 ;
  assign n76683 = ~n34545 ;
  assign n34566 = n34541 & n76683 ;
  assign n34567 = n34565 | n34566 ;
  assign n34568 = n76681 & n34567 ;
  assign n34569 = n34368 & n76675 ;
  assign n34570 = n34561 & n34569 ;
  assign n34571 = n34568 | n34570 ;
  assign n34613 = n66244 & n34571 ;
  assign n76684 = ~n34600 ;
  assign n34614 = n34539 & n76684 ;
  assign n34540 = n34385 | n34539 ;
  assign n76685 = ~n34540 ;
  assign n34615 = n76685 & n34599 ;
  assign n34616 = n34614 | n34615 ;
  assign n34617 = n76681 & n34616 ;
  assign n34618 = n34376 & n76675 ;
  assign n34619 = n34561 & n34618 ;
  assign n34620 = n34617 | n34619 ;
  assign n34621 = n66145 & n34620 ;
  assign n76686 = ~n34534 ;
  assign n34622 = n34532 & n76686 ;
  assign n34533 = n34393 | n34532 ;
  assign n76687 = ~n34533 ;
  assign n34623 = n34529 & n76687 ;
  assign n34624 = n34622 | n34623 ;
  assign n34625 = n76681 & n34624 ;
  assign n34626 = n34384 & n76675 ;
  assign n34627 = n34561 & n34626 ;
  assign n34628 = n34625 | n34627 ;
  assign n34629 = n66081 & n34628 ;
  assign n76688 = ~n34596 ;
  assign n34630 = n34527 & n76688 ;
  assign n34528 = n34401 | n34527 ;
  assign n76689 = ~n34528 ;
  assign n34631 = n76689 & n34595 ;
  assign n34632 = n34630 | n34631 ;
  assign n34633 = n76681 & n34632 ;
  assign n34634 = n34392 & n76675 ;
  assign n34635 = n34561 & n34634 ;
  assign n34636 = n34633 | n34635 ;
  assign n34637 = n66043 & n34636 ;
  assign n76690 = ~n34522 ;
  assign n34638 = n34520 & n76690 ;
  assign n34521 = n34409 | n34520 ;
  assign n76691 = ~n34521 ;
  assign n34639 = n34517 & n76691 ;
  assign n34640 = n34638 | n34639 ;
  assign n34641 = n76681 & n34640 ;
  assign n34642 = n34400 & n76675 ;
  assign n34643 = n34561 & n34642 ;
  assign n34644 = n34641 | n34643 ;
  assign n34645 = n65960 & n34644 ;
  assign n76692 = ~n34592 ;
  assign n34646 = n34515 & n76692 ;
  assign n34516 = n34417 | n34515 ;
  assign n76693 = ~n34516 ;
  assign n34647 = n76693 & n34591 ;
  assign n34648 = n34646 | n34647 ;
  assign n34649 = n76681 & n34648 ;
  assign n34650 = n34408 & n76675 ;
  assign n34651 = n34561 & n34650 ;
  assign n34652 = n34649 | n34651 ;
  assign n34653 = n65909 & n34652 ;
  assign n76694 = ~n34510 ;
  assign n34654 = n34508 & n76694 ;
  assign n34509 = n34425 | n34508 ;
  assign n76695 = ~n34509 ;
  assign n34655 = n34505 & n76695 ;
  assign n34656 = n34654 | n34655 ;
  assign n34657 = n76681 & n34656 ;
  assign n34658 = n34416 & n76675 ;
  assign n34659 = n34561 & n34658 ;
  assign n34660 = n34657 | n34659 ;
  assign n34661 = n65877 & n34660 ;
  assign n76696 = ~n34588 ;
  assign n34662 = n34503 & n76696 ;
  assign n34504 = n34434 | n34503 ;
  assign n76697 = ~n34504 ;
  assign n34663 = n76697 & n34587 ;
  assign n34664 = n34662 | n34663 ;
  assign n34665 = n76681 & n34664 ;
  assign n34666 = n34424 & n76675 ;
  assign n34667 = n34561 & n34666 ;
  assign n34668 = n34665 | n34667 ;
  assign n34669 = n65820 & n34668 ;
  assign n76698 = ~n34498 ;
  assign n34671 = n34497 & n76698 ;
  assign n34670 = n34442 | n34497 ;
  assign n76699 = ~n34670 ;
  assign n34672 = n34494 & n76699 ;
  assign n34673 = n34671 | n34672 ;
  assign n34674 = n76681 & n34673 ;
  assign n34675 = n34433 & n76675 ;
  assign n34676 = n34561 & n34675 ;
  assign n34677 = n34674 | n34676 ;
  assign n34678 = n65791 & n34677 ;
  assign n76700 = ~n34584 ;
  assign n34680 = n34493 & n76700 ;
  assign n34679 = n34451 | n34493 ;
  assign n76701 = ~n34679 ;
  assign n34681 = n34583 & n76701 ;
  assign n34682 = n34680 | n34681 ;
  assign n34683 = n76681 & n34682 ;
  assign n34684 = n34441 & n76675 ;
  assign n34685 = n34561 & n34684 ;
  assign n34686 = n34683 | n34685 ;
  assign n34687 = n65772 & n34686 ;
  assign n34688 = n76679 & n34484 ;
  assign n76702 = ~n34688 ;
  assign n34690 = n34487 & n76702 ;
  assign n34689 = n34480 | n34487 ;
  assign n76703 = ~n34689 ;
  assign n34691 = n34484 & n76703 ;
  assign n34692 = n34690 | n34691 ;
  assign n34693 = n76681 & n34692 ;
  assign n34694 = n34450 & n76675 ;
  assign n34695 = n34561 & n34694 ;
  assign n34696 = n34693 | n34695 ;
  assign n34697 = n65746 & n34696 ;
  assign n76704 = ~n34580 ;
  assign n34699 = n34579 & n76704 ;
  assign n34698 = n34476 | n34483 ;
  assign n76705 = ~n34698 ;
  assign n34700 = n34577 & n76705 ;
  assign n34701 = n34699 | n34700 ;
  assign n34702 = n76681 & n34701 ;
  assign n34703 = n34479 & n76675 ;
  assign n34704 = n34561 & n34703 ;
  assign n34705 = n34702 | n34704 ;
  assign n34706 = n65721 & n34705 ;
  assign n34707 = n1989 & n34472 ;
  assign n34708 = n76678 & n34707 ;
  assign n76706 = ~n34708 ;
  assign n34709 = n34577 & n76706 ;
  assign n34710 = n76681 & n34709 ;
  assign n34711 = n34475 & n76675 ;
  assign n34712 = n34561 & n34711 ;
  assign n34713 = n34710 | n34712 ;
  assign n34714 = n65686 & n34713 ;
  assign n34564 = n1989 & n76681 ;
  assign n34719 = x64 & n76681 ;
  assign n76707 = ~n34719 ;
  assign n34720 = x49 & n76707 ;
  assign n34721 = n34564 | n34720 ;
  assign n34723 = x65 & n34721 ;
  assign n34715 = n34560 | n34604 ;
  assign n34716 = n76675 & n34715 ;
  assign n76708 = ~n34716 ;
  assign n34717 = x64 & n76708 ;
  assign n76709 = ~n34717 ;
  assign n34718 = x49 & n76709 ;
  assign n34722 = x65 | n34564 ;
  assign n34724 = n34718 | n34722 ;
  assign n76710 = ~n34723 ;
  assign n34725 = n76710 & n34724 ;
  assign n34726 = n2241 | n34725 ;
  assign n34727 = n65670 & n34721 ;
  assign n76711 = ~n34727 ;
  assign n34728 = n34726 & n76711 ;
  assign n76712 = ~n34712 ;
  assign n34729 = x66 & n76712 ;
  assign n76713 = ~n34710 ;
  assign n34730 = n76713 & n34729 ;
  assign n34731 = n34714 | n34730 ;
  assign n34732 = n34728 | n34731 ;
  assign n76714 = ~n34714 ;
  assign n34733 = n76714 & n34732 ;
  assign n76715 = ~n34704 ;
  assign n34734 = x67 & n76715 ;
  assign n76716 = ~n34702 ;
  assign n34735 = n76716 & n34734 ;
  assign n34736 = n34706 | n34735 ;
  assign n34737 = n34733 | n34736 ;
  assign n76717 = ~n34706 ;
  assign n34738 = n76717 & n34737 ;
  assign n76718 = ~n34695 ;
  assign n34739 = x68 & n76718 ;
  assign n76719 = ~n34693 ;
  assign n34740 = n76719 & n34739 ;
  assign n34741 = n34697 | n34740 ;
  assign n34742 = n34738 | n34741 ;
  assign n76720 = ~n34697 ;
  assign n34743 = n76720 & n34742 ;
  assign n76721 = ~n34685 ;
  assign n34744 = x69 & n76721 ;
  assign n76722 = ~n34683 ;
  assign n34745 = n76722 & n34744 ;
  assign n34746 = n34687 | n34745 ;
  assign n34748 = n34743 | n34746 ;
  assign n76723 = ~n34687 ;
  assign n34749 = n76723 & n34748 ;
  assign n76724 = ~n34676 ;
  assign n34750 = x70 & n76724 ;
  assign n76725 = ~n34674 ;
  assign n34751 = n76725 & n34750 ;
  assign n34752 = n34678 | n34751 ;
  assign n34753 = n34749 | n34752 ;
  assign n76726 = ~n34678 ;
  assign n34754 = n76726 & n34753 ;
  assign n76727 = ~n34667 ;
  assign n34755 = x71 & n76727 ;
  assign n76728 = ~n34665 ;
  assign n34756 = n76728 & n34755 ;
  assign n34757 = n34669 | n34756 ;
  assign n34759 = n34754 | n34757 ;
  assign n76729 = ~n34669 ;
  assign n34760 = n76729 & n34759 ;
  assign n76730 = ~n34659 ;
  assign n34761 = x72 & n76730 ;
  assign n76731 = ~n34657 ;
  assign n34762 = n76731 & n34761 ;
  assign n34763 = n34661 | n34762 ;
  assign n34764 = n34760 | n34763 ;
  assign n76732 = ~n34661 ;
  assign n34765 = n76732 & n34764 ;
  assign n76733 = ~n34651 ;
  assign n34766 = x73 & n76733 ;
  assign n76734 = ~n34649 ;
  assign n34767 = n76734 & n34766 ;
  assign n34768 = n34653 | n34767 ;
  assign n34770 = n34765 | n34768 ;
  assign n76735 = ~n34653 ;
  assign n34771 = n76735 & n34770 ;
  assign n76736 = ~n34643 ;
  assign n34772 = x74 & n76736 ;
  assign n76737 = ~n34641 ;
  assign n34773 = n76737 & n34772 ;
  assign n34774 = n34645 | n34773 ;
  assign n34775 = n34771 | n34774 ;
  assign n76738 = ~n34645 ;
  assign n34776 = n76738 & n34775 ;
  assign n76739 = ~n34635 ;
  assign n34777 = x75 & n76739 ;
  assign n76740 = ~n34633 ;
  assign n34778 = n76740 & n34777 ;
  assign n34779 = n34637 | n34778 ;
  assign n34781 = n34776 | n34779 ;
  assign n76741 = ~n34637 ;
  assign n34782 = n76741 & n34781 ;
  assign n76742 = ~n34627 ;
  assign n34783 = x76 & n76742 ;
  assign n76743 = ~n34625 ;
  assign n34784 = n76743 & n34783 ;
  assign n34785 = n34629 | n34784 ;
  assign n34786 = n34782 | n34785 ;
  assign n76744 = ~n34629 ;
  assign n34787 = n76744 & n34786 ;
  assign n76745 = ~n34619 ;
  assign n34788 = x77 & n76745 ;
  assign n76746 = ~n34617 ;
  assign n34789 = n76746 & n34788 ;
  assign n34790 = n34621 | n34789 ;
  assign n34792 = n34787 | n34790 ;
  assign n76747 = ~n34621 ;
  assign n34793 = n76747 & n34792 ;
  assign n76748 = ~n34570 ;
  assign n34794 = x78 & n76748 ;
  assign n76749 = ~n34568 ;
  assign n34795 = n76749 & n34794 ;
  assign n34796 = n34613 | n34795 ;
  assign n34797 = n34793 | n34796 ;
  assign n76750 = ~n34613 ;
  assign n34798 = n76750 & n34797 ;
  assign n76751 = ~n34610 ;
  assign n34799 = x79 & n76751 ;
  assign n76752 = ~n34608 ;
  assign n34800 = n76752 & n34799 ;
  assign n34801 = n34612 | n34800 ;
  assign n34803 = n34798 | n34801 ;
  assign n76753 = ~n34612 ;
  assign n34804 = n76753 & n34803 ;
  assign n34805 = n67897 | n34804 ;
  assign n76754 = ~n34611 ;
  assign n34806 = n76754 & n34805 ;
  assign n76755 = ~n34798 ;
  assign n34802 = n76755 & n34801 ;
  assign n34809 = n34564 | n34718 ;
  assign n34810 = x65 & n34809 ;
  assign n76756 = ~n34810 ;
  assign n34811 = n34724 & n76756 ;
  assign n34812 = n2241 | n34811 ;
  assign n34813 = n76711 & n34812 ;
  assign n34814 = n34731 | n34813 ;
  assign n34815 = n76714 & n34814 ;
  assign n34817 = n34736 | n34815 ;
  assign n34818 = n76717 & n34817 ;
  assign n34820 = n34741 | n34818 ;
  assign n34821 = n76720 & n34820 ;
  assign n34822 = n34746 | n34821 ;
  assign n34823 = n76723 & n34822 ;
  assign n34824 = n34752 | n34823 ;
  assign n34826 = n76726 & n34824 ;
  assign n34827 = n34757 | n34826 ;
  assign n34828 = n76729 & n34827 ;
  assign n34829 = n34763 | n34828 ;
  assign n34831 = n76732 & n34829 ;
  assign n34832 = n34768 | n34831 ;
  assign n34833 = n76735 & n34832 ;
  assign n34834 = n34774 | n34833 ;
  assign n34836 = n76738 & n34834 ;
  assign n34837 = n34779 | n34836 ;
  assign n34838 = n76741 & n34837 ;
  assign n34839 = n34785 | n34838 ;
  assign n34841 = n76744 & n34839 ;
  assign n34842 = n34790 | n34841 ;
  assign n34843 = n76747 & n34842 ;
  assign n34845 = n34796 | n34843 ;
  assign n34852 = n34613 | n34801 ;
  assign n76757 = ~n34852 ;
  assign n34853 = n34845 & n76757 ;
  assign n34854 = n34802 | n34853 ;
  assign n34855 = n34805 | n34854 ;
  assign n76758 = ~n34806 ;
  assign n34856 = n76758 & n34855 ;
  assign n34857 = n66379 & n34856 ;
  assign n76759 = ~n34805 ;
  assign n35056 = n76759 & n34854 ;
  assign n35057 = n34611 & n34805 ;
  assign n76760 = ~n35057 ;
  assign n35058 = x80 & n76760 ;
  assign n76761 = ~n35056 ;
  assign n35059 = n76761 & n35058 ;
  assign n35060 = n34857 | n35059 ;
  assign n34807 = n34571 & n34805 ;
  assign n76762 = ~n34843 ;
  assign n34844 = n34796 & n76762 ;
  assign n34846 = n34621 | n34796 ;
  assign n76763 = ~n34846 ;
  assign n34847 = n34792 & n76763 ;
  assign n34848 = n34844 | n34847 ;
  assign n34849 = n65678 & n34848 ;
  assign n76764 = ~n34804 ;
  assign n34850 = n76764 & n34849 ;
  assign n34851 = n34807 | n34850 ;
  assign n34858 = n66299 & n34851 ;
  assign n34859 = n34620 & n34805 ;
  assign n76765 = ~n34787 ;
  assign n34791 = n76765 & n34790 ;
  assign n34860 = n34629 | n34790 ;
  assign n76766 = ~n34860 ;
  assign n34861 = n34839 & n76766 ;
  assign n34862 = n34791 | n34861 ;
  assign n34863 = n65678 & n34862 ;
  assign n34864 = n76764 & n34863 ;
  assign n34865 = n34859 | n34864 ;
  assign n34866 = n66244 & n34865 ;
  assign n76767 = ~n34864 ;
  assign n35044 = x78 & n76767 ;
  assign n76768 = ~n34859 ;
  assign n35045 = n76768 & n35044 ;
  assign n35046 = n34866 | n35045 ;
  assign n34867 = n34628 & n34805 ;
  assign n76769 = ~n34838 ;
  assign n34840 = n34785 & n76769 ;
  assign n34868 = n34637 | n34785 ;
  assign n76770 = ~n34868 ;
  assign n34869 = n34781 & n76770 ;
  assign n34870 = n34840 | n34869 ;
  assign n34871 = n65678 & n34870 ;
  assign n34872 = n76764 & n34871 ;
  assign n34873 = n34867 | n34872 ;
  assign n34874 = n66145 & n34873 ;
  assign n34875 = n34636 & n34805 ;
  assign n76771 = ~n34776 ;
  assign n34780 = n76771 & n34779 ;
  assign n34876 = n34645 | n34779 ;
  assign n76772 = ~n34876 ;
  assign n34877 = n34834 & n76772 ;
  assign n34878 = n34780 | n34877 ;
  assign n34879 = n65678 & n34878 ;
  assign n34880 = n76764 & n34879 ;
  assign n34881 = n34875 | n34880 ;
  assign n34882 = n66081 & n34881 ;
  assign n76773 = ~n34880 ;
  assign n35032 = x76 & n76773 ;
  assign n76774 = ~n34875 ;
  assign n35033 = n76774 & n35032 ;
  assign n35034 = n34882 | n35033 ;
  assign n34883 = n34644 & n34805 ;
  assign n76775 = ~n34833 ;
  assign n34835 = n34774 & n76775 ;
  assign n34884 = n34653 | n34774 ;
  assign n76776 = ~n34884 ;
  assign n34885 = n34770 & n76776 ;
  assign n34886 = n34835 | n34885 ;
  assign n34887 = n65678 & n34886 ;
  assign n34888 = n76764 & n34887 ;
  assign n34889 = n34883 | n34888 ;
  assign n34890 = n66043 & n34889 ;
  assign n34891 = n34652 & n34805 ;
  assign n76777 = ~n34765 ;
  assign n34769 = n76777 & n34768 ;
  assign n34892 = n34661 | n34768 ;
  assign n76778 = ~n34892 ;
  assign n34893 = n34829 & n76778 ;
  assign n34894 = n34769 | n34893 ;
  assign n34895 = n65678 & n34894 ;
  assign n34896 = n76764 & n34895 ;
  assign n34897 = n34891 | n34896 ;
  assign n34898 = n65960 & n34897 ;
  assign n76779 = ~n34896 ;
  assign n35020 = x74 & n76779 ;
  assign n76780 = ~n34891 ;
  assign n35021 = n76780 & n35020 ;
  assign n35022 = n34898 | n35021 ;
  assign n34899 = n34660 & n34805 ;
  assign n76781 = ~n34828 ;
  assign n34830 = n34763 & n76781 ;
  assign n34900 = n34669 | n34763 ;
  assign n76782 = ~n34900 ;
  assign n34901 = n34759 & n76782 ;
  assign n34902 = n34830 | n34901 ;
  assign n34903 = n65678 & n34902 ;
  assign n34904 = n76764 & n34903 ;
  assign n34905 = n34899 | n34904 ;
  assign n34906 = n65909 & n34905 ;
  assign n34907 = n34668 & n34805 ;
  assign n76783 = ~n34754 ;
  assign n34758 = n76783 & n34757 ;
  assign n34908 = n34678 | n34757 ;
  assign n76784 = ~n34908 ;
  assign n34909 = n34824 & n76784 ;
  assign n34910 = n34758 | n34909 ;
  assign n34911 = n65678 & n34910 ;
  assign n34912 = n76764 & n34911 ;
  assign n34913 = n34907 | n34912 ;
  assign n34914 = n65877 & n34913 ;
  assign n76785 = ~n34912 ;
  assign n35008 = x72 & n76785 ;
  assign n76786 = ~n34907 ;
  assign n35009 = n76786 & n35008 ;
  assign n35010 = n34914 | n35009 ;
  assign n34915 = n34677 & n34805 ;
  assign n76787 = ~n34823 ;
  assign n34825 = n34752 & n76787 ;
  assign n34916 = n34687 | n34752 ;
  assign n76788 = ~n34916 ;
  assign n34917 = n34748 & n76788 ;
  assign n34918 = n34825 | n34917 ;
  assign n34919 = n65678 & n34918 ;
  assign n34920 = n76764 & n34919 ;
  assign n34921 = n34915 | n34920 ;
  assign n34922 = n65820 & n34921 ;
  assign n34923 = n34686 & n34805 ;
  assign n76789 = ~n34743 ;
  assign n34747 = n76789 & n34746 ;
  assign n34924 = n34697 | n34746 ;
  assign n76790 = ~n34924 ;
  assign n34925 = n34820 & n76790 ;
  assign n34926 = n34747 | n34925 ;
  assign n34927 = n65678 & n34926 ;
  assign n34928 = n76764 & n34927 ;
  assign n34929 = n34923 | n34928 ;
  assign n34930 = n65791 & n34929 ;
  assign n76791 = ~n34928 ;
  assign n34997 = x70 & n76791 ;
  assign n76792 = ~n34923 ;
  assign n34998 = n76792 & n34997 ;
  assign n34999 = n34930 | n34998 ;
  assign n34931 = n34696 & n34805 ;
  assign n76793 = ~n34818 ;
  assign n34819 = n34741 & n76793 ;
  assign n34932 = n34706 | n34741 ;
  assign n76794 = ~n34932 ;
  assign n34933 = n34737 & n76794 ;
  assign n34934 = n34819 | n34933 ;
  assign n34935 = n65678 & n34934 ;
  assign n34936 = n76764 & n34935 ;
  assign n34937 = n34931 | n34936 ;
  assign n34938 = n65772 & n34937 ;
  assign n34939 = n34705 & n34805 ;
  assign n76795 = ~n34733 ;
  assign n34816 = n76795 & n34736 ;
  assign n34940 = n34714 | n34736 ;
  assign n76796 = ~n34940 ;
  assign n34941 = n34732 & n76796 ;
  assign n34942 = n34816 | n34941 ;
  assign n34943 = n65678 & n34942 ;
  assign n34944 = n76764 & n34943 ;
  assign n34945 = n34939 | n34944 ;
  assign n34946 = n65746 & n34945 ;
  assign n76797 = ~n34944 ;
  assign n34987 = x68 & n76797 ;
  assign n76798 = ~n34939 ;
  assign n34988 = n76798 & n34987 ;
  assign n34989 = n34946 | n34988 ;
  assign n34808 = n34713 & n34805 ;
  assign n34947 = n34727 | n34731 ;
  assign n76799 = ~n34947 ;
  assign n34948 = n34812 & n76799 ;
  assign n76800 = ~n34813 ;
  assign n34949 = n34731 & n76800 ;
  assign n34950 = n34948 | n34949 ;
  assign n34951 = n65678 & n34950 ;
  assign n34952 = n76764 & n34951 ;
  assign n34953 = n34808 | n34952 ;
  assign n34954 = n65721 & n34953 ;
  assign n34955 = n34805 & n34809 ;
  assign n34956 = n2241 & n34724 ;
  assign n34957 = n76710 & n34956 ;
  assign n34958 = n67897 | n34957 ;
  assign n76801 = ~n34958 ;
  assign n34959 = n34812 & n76801 ;
  assign n34960 = n76764 & n34959 ;
  assign n34961 = n34955 | n34960 ;
  assign n34962 = n65686 & n34961 ;
  assign n76802 = ~n34960 ;
  assign n34977 = x66 & n76802 ;
  assign n76803 = ~n34955 ;
  assign n34978 = n76803 & n34977 ;
  assign n34979 = n34962 | n34978 ;
  assign n34963 = n76750 & n34845 ;
  assign n34964 = n34801 | n34963 ;
  assign n34965 = n76753 & n34964 ;
  assign n76804 = ~n34965 ;
  assign n34966 = n2484 & n76804 ;
  assign n76805 = ~n34966 ;
  assign n34967 = x48 & n76805 ;
  assign n34968 = n2489 & n76764 ;
  assign n34969 = n34967 | n34968 ;
  assign n34970 = x65 & n34969 ;
  assign n34971 = x65 | n34968 ;
  assign n34972 = n34967 | n34971 ;
  assign n76806 = ~n34970 ;
  assign n34973 = n76806 & n34972 ;
  assign n34975 = n2497 | n34973 ;
  assign n34976 = n65670 & n34969 ;
  assign n76807 = ~n34976 ;
  assign n34980 = n34975 & n76807 ;
  assign n34981 = n34979 | n34980 ;
  assign n76808 = ~n34962 ;
  assign n34982 = n76808 & n34981 ;
  assign n76809 = ~n34952 ;
  assign n34983 = x67 & n76809 ;
  assign n76810 = ~n34808 ;
  assign n34984 = n76810 & n34983 ;
  assign n34985 = n34954 | n34984 ;
  assign n34986 = n34982 | n34985 ;
  assign n76811 = ~n34954 ;
  assign n34990 = n76811 & n34986 ;
  assign n34991 = n34989 | n34990 ;
  assign n76812 = ~n34946 ;
  assign n34992 = n76812 & n34991 ;
  assign n76813 = ~n34936 ;
  assign n34993 = x69 & n76813 ;
  assign n76814 = ~n34931 ;
  assign n34994 = n76814 & n34993 ;
  assign n34995 = n34938 | n34994 ;
  assign n34996 = n34992 | n34995 ;
  assign n76815 = ~n34938 ;
  assign n35000 = n76815 & n34996 ;
  assign n35001 = n34999 | n35000 ;
  assign n76816 = ~n34930 ;
  assign n35002 = n76816 & n35001 ;
  assign n76817 = ~n34920 ;
  assign n35003 = x71 & n76817 ;
  assign n76818 = ~n34915 ;
  assign n35004 = n76818 & n35003 ;
  assign n35005 = n34922 | n35004 ;
  assign n35007 = n35002 | n35005 ;
  assign n76819 = ~n34922 ;
  assign n35012 = n76819 & n35007 ;
  assign n35013 = n35010 | n35012 ;
  assign n76820 = ~n34914 ;
  assign n35014 = n76820 & n35013 ;
  assign n76821 = ~n34904 ;
  assign n35015 = x73 & n76821 ;
  assign n76822 = ~n34899 ;
  assign n35016 = n76822 & n35015 ;
  assign n35017 = n34906 | n35016 ;
  assign n35019 = n35014 | n35017 ;
  assign n76823 = ~n34906 ;
  assign n35024 = n76823 & n35019 ;
  assign n35025 = n35022 | n35024 ;
  assign n76824 = ~n34898 ;
  assign n35026 = n76824 & n35025 ;
  assign n76825 = ~n34888 ;
  assign n35027 = x75 & n76825 ;
  assign n76826 = ~n34883 ;
  assign n35028 = n76826 & n35027 ;
  assign n35029 = n34890 | n35028 ;
  assign n35031 = n35026 | n35029 ;
  assign n76827 = ~n34890 ;
  assign n35036 = n76827 & n35031 ;
  assign n35037 = n35034 | n35036 ;
  assign n76828 = ~n34882 ;
  assign n35038 = n76828 & n35037 ;
  assign n76829 = ~n34872 ;
  assign n35039 = x77 & n76829 ;
  assign n76830 = ~n34867 ;
  assign n35040 = n76830 & n35039 ;
  assign n35041 = n34874 | n35040 ;
  assign n35043 = n35038 | n35041 ;
  assign n76831 = ~n34874 ;
  assign n35048 = n76831 & n35043 ;
  assign n35049 = n35046 | n35048 ;
  assign n76832 = ~n34866 ;
  assign n35050 = n76832 & n35049 ;
  assign n76833 = ~n34850 ;
  assign n35051 = x79 & n76833 ;
  assign n76834 = ~n34807 ;
  assign n35052 = n76834 & n35051 ;
  assign n35053 = n34858 | n35052 ;
  assign n35055 = n35050 | n35053 ;
  assign n76835 = ~n34858 ;
  assign n35061 = n76835 & n35055 ;
  assign n35062 = n35060 | n35061 ;
  assign n76836 = ~n34857 ;
  assign n35063 = n76836 & n35062 ;
  assign n35064 = n344 | n35063 ;
  assign n76837 = ~n34856 ;
  assign n35066 = n76837 & n35064 ;
  assign n76838 = ~n35061 ;
  assign n35321 = n35060 & n76838 ;
  assign n35069 = n2484 & n76764 ;
  assign n76839 = ~n35069 ;
  assign n35070 = x48 & n76839 ;
  assign n35071 = n34968 | n35070 ;
  assign n35072 = x65 & n35071 ;
  assign n76840 = ~n35072 ;
  assign n35073 = n34972 & n76840 ;
  assign n35074 = n2497 | n35073 ;
  assign n35075 = n76807 & n35074 ;
  assign n35076 = n34979 | n35075 ;
  assign n35077 = n76808 & n35076 ;
  assign n35078 = n34985 | n35077 ;
  assign n35079 = n76811 & n35078 ;
  assign n35080 = n34989 | n35079 ;
  assign n35081 = n76812 & n35080 ;
  assign n35082 = n34995 | n35081 ;
  assign n35083 = n76815 & n35082 ;
  assign n35084 = n34999 | n35083 ;
  assign n35085 = n76816 & n35084 ;
  assign n35086 = n35005 | n35085 ;
  assign n35087 = n76819 & n35086 ;
  assign n35088 = n35010 | n35087 ;
  assign n35089 = n76820 & n35088 ;
  assign n35090 = n35017 | n35089 ;
  assign n35091 = n76823 & n35090 ;
  assign n35092 = n35022 | n35091 ;
  assign n35093 = n76824 & n35092 ;
  assign n35094 = n35029 | n35093 ;
  assign n35095 = n76827 & n35094 ;
  assign n35096 = n35034 | n35095 ;
  assign n35097 = n76828 & n35096 ;
  assign n35098 = n35041 | n35097 ;
  assign n35099 = n76831 & n35098 ;
  assign n35100 = n35046 | n35099 ;
  assign n35102 = n76832 & n35100 ;
  assign n35224 = n35053 | n35102 ;
  assign n35322 = n34858 | n35060 ;
  assign n76841 = ~n35322 ;
  assign n35323 = n35224 & n76841 ;
  assign n35324 = n35321 | n35323 ;
  assign n35325 = n35064 | n35324 ;
  assign n76842 = ~n35066 ;
  assign n35326 = n76842 & n35325 ;
  assign n35334 = n65715 & n35326 ;
  assign n35067 = n34851 & n35064 ;
  assign n35054 = n34866 | n35053 ;
  assign n76843 = ~n35054 ;
  assign n35101 = n76843 & n35100 ;
  assign n76844 = ~n35102 ;
  assign n35103 = n35053 & n76844 ;
  assign n35104 = n35101 | n35103 ;
  assign n35105 = n65715 & n35104 ;
  assign n76845 = ~n35063 ;
  assign n35106 = n76845 & n35105 ;
  assign n35107 = n35067 | n35106 ;
  assign n35108 = n66379 & n35107 ;
  assign n35109 = n34865 & n35064 ;
  assign n35047 = n34874 | n35046 ;
  assign n76846 = ~n35047 ;
  assign n35110 = n35043 & n76846 ;
  assign n76847 = ~n35048 ;
  assign n35111 = n35046 & n76847 ;
  assign n35112 = n35110 | n35111 ;
  assign n35113 = n65715 & n35112 ;
  assign n35114 = n76845 & n35113 ;
  assign n35115 = n35109 | n35114 ;
  assign n35116 = n66299 & n35115 ;
  assign n35117 = n34873 & n35064 ;
  assign n35042 = n34882 | n35041 ;
  assign n76848 = ~n35042 ;
  assign n35118 = n76848 & n35096 ;
  assign n76849 = ~n35097 ;
  assign n35119 = n35041 & n76849 ;
  assign n35120 = n35118 | n35119 ;
  assign n35121 = n65715 & n35120 ;
  assign n35122 = n76845 & n35121 ;
  assign n35123 = n35117 | n35122 ;
  assign n35124 = n66244 & n35123 ;
  assign n35125 = n34881 & n35064 ;
  assign n35035 = n34890 | n35034 ;
  assign n76850 = ~n35035 ;
  assign n35126 = n35031 & n76850 ;
  assign n76851 = ~n35036 ;
  assign n35127 = n35034 & n76851 ;
  assign n35128 = n35126 | n35127 ;
  assign n35129 = n65715 & n35128 ;
  assign n35130 = n76845 & n35129 ;
  assign n35131 = n35125 | n35130 ;
  assign n35132 = n66145 & n35131 ;
  assign n35133 = n34889 & n35064 ;
  assign n35030 = n34898 | n35029 ;
  assign n76852 = ~n35030 ;
  assign n35134 = n76852 & n35092 ;
  assign n76853 = ~n35093 ;
  assign n35135 = n35029 & n76853 ;
  assign n35136 = n35134 | n35135 ;
  assign n35137 = n65715 & n35136 ;
  assign n35138 = n76845 & n35137 ;
  assign n35139 = n35133 | n35138 ;
  assign n35140 = n66081 & n35139 ;
  assign n35141 = n34897 & n35064 ;
  assign n35023 = n34906 | n35022 ;
  assign n76854 = ~n35023 ;
  assign n35142 = n35019 & n76854 ;
  assign n76855 = ~n35024 ;
  assign n35143 = n35022 & n76855 ;
  assign n35144 = n35142 | n35143 ;
  assign n35145 = n65715 & n35144 ;
  assign n35146 = n76845 & n35145 ;
  assign n35147 = n35141 | n35146 ;
  assign n35148 = n66043 & n35147 ;
  assign n35149 = n34905 & n35064 ;
  assign n35018 = n34914 | n35017 ;
  assign n76856 = ~n35018 ;
  assign n35150 = n76856 & n35088 ;
  assign n76857 = ~n35089 ;
  assign n35151 = n35017 & n76857 ;
  assign n35152 = n35150 | n35151 ;
  assign n35153 = n65715 & n35152 ;
  assign n35154 = n76845 & n35153 ;
  assign n35155 = n35149 | n35154 ;
  assign n35156 = n65960 & n35155 ;
  assign n35157 = n34913 & n35064 ;
  assign n35011 = n34922 | n35010 ;
  assign n76858 = ~n35011 ;
  assign n35158 = n35007 & n76858 ;
  assign n76859 = ~n35012 ;
  assign n35159 = n35010 & n76859 ;
  assign n35160 = n35158 | n35159 ;
  assign n35161 = n65715 & n35160 ;
  assign n35162 = n76845 & n35161 ;
  assign n35163 = n35157 | n35162 ;
  assign n35164 = n65909 & n35163 ;
  assign n35165 = n34921 & n35064 ;
  assign n35006 = n34930 | n35005 ;
  assign n76860 = ~n35006 ;
  assign n35166 = n76860 & n35084 ;
  assign n76861 = ~n35085 ;
  assign n35167 = n35005 & n76861 ;
  assign n35168 = n35166 | n35167 ;
  assign n35169 = n65715 & n35168 ;
  assign n35170 = n76845 & n35169 ;
  assign n35171 = n35165 | n35170 ;
  assign n35172 = n65877 & n35171 ;
  assign n35173 = n34929 & n35064 ;
  assign n35068 = n34938 | n34999 ;
  assign n76862 = ~n35068 ;
  assign n35174 = n34996 & n76862 ;
  assign n76863 = ~n35000 ;
  assign n35175 = n34999 & n76863 ;
  assign n35176 = n35174 | n35175 ;
  assign n35177 = n65715 & n35176 ;
  assign n35178 = n76845 & n35177 ;
  assign n35179 = n35173 | n35178 ;
  assign n35180 = n65820 & n35179 ;
  assign n35181 = n34937 & n35064 ;
  assign n35182 = n34946 | n34995 ;
  assign n76864 = ~n35182 ;
  assign n35183 = n35080 & n76864 ;
  assign n76865 = ~n35081 ;
  assign n35184 = n34995 & n76865 ;
  assign n35185 = n35183 | n35184 ;
  assign n35186 = n65715 & n35185 ;
  assign n35187 = n76845 & n35186 ;
  assign n35188 = n35181 | n35187 ;
  assign n35189 = n65791 & n35188 ;
  assign n35190 = n34945 & n35064 ;
  assign n35191 = n34954 | n34989 ;
  assign n76866 = ~n35191 ;
  assign n35192 = n35078 & n76866 ;
  assign n76867 = ~n34990 ;
  assign n35193 = n34989 & n76867 ;
  assign n35194 = n35192 | n35193 ;
  assign n35195 = n65715 & n35194 ;
  assign n35196 = n76845 & n35195 ;
  assign n35197 = n35190 | n35196 ;
  assign n35198 = n65772 & n35197 ;
  assign n35199 = n34953 & n35064 ;
  assign n35200 = n34962 | n34985 ;
  assign n76868 = ~n35200 ;
  assign n35201 = n35076 & n76868 ;
  assign n76869 = ~n35077 ;
  assign n35202 = n34985 & n76869 ;
  assign n35203 = n35201 | n35202 ;
  assign n35204 = n65715 & n35203 ;
  assign n35205 = n76845 & n35204 ;
  assign n35206 = n35199 | n35205 ;
  assign n35207 = n65746 & n35206 ;
  assign n35208 = n34961 & n35064 ;
  assign n76870 = ~n35075 ;
  assign n35209 = n34979 & n76870 ;
  assign n35210 = n34976 | n34979 ;
  assign n76871 = ~n35210 ;
  assign n35211 = n35074 & n76871 ;
  assign n35212 = n35209 | n35211 ;
  assign n35213 = n65715 & n35212 ;
  assign n35214 = n76845 & n35213 ;
  assign n35215 = n35208 | n35214 ;
  assign n35216 = n65721 & n35215 ;
  assign n35065 = n34969 & n35064 ;
  assign n34974 = n2497 & n34972 ;
  assign n35217 = n34974 & n76840 ;
  assign n35218 = n344 | n35217 ;
  assign n76872 = ~n35218 ;
  assign n35219 = n35074 & n76872 ;
  assign n35220 = n76845 & n35219 ;
  assign n35221 = n35065 | n35220 ;
  assign n35222 = n65686 & n35221 ;
  assign n35223 = n2766 & n76845 ;
  assign n35225 = n76835 & n35224 ;
  assign n35226 = n35060 | n35225 ;
  assign n35227 = n76836 & n35226 ;
  assign n76873 = ~n35227 ;
  assign n35228 = n2761 & n76873 ;
  assign n76874 = ~n35228 ;
  assign n35229 = x47 & n76874 ;
  assign n35230 = n35223 | n35229 ;
  assign n35238 = n65670 & n35230 ;
  assign n35231 = n2761 & n76845 ;
  assign n76875 = ~n35231 ;
  assign n35232 = x47 & n76875 ;
  assign n35233 = n35223 | n35232 ;
  assign n35234 = x65 & n35233 ;
  assign n35235 = x65 | n35223 ;
  assign n35236 = n35232 | n35235 ;
  assign n76876 = ~n35234 ;
  assign n35237 = n76876 & n35236 ;
  assign n35239 = n2773 | n35237 ;
  assign n76877 = ~n35238 ;
  assign n35240 = n76877 & n35239 ;
  assign n76878 = ~n35220 ;
  assign n35241 = x66 & n76878 ;
  assign n76879 = ~n35065 ;
  assign n35242 = n76879 & n35241 ;
  assign n35243 = n35240 | n35242 ;
  assign n76880 = ~n35222 ;
  assign n35244 = n76880 & n35243 ;
  assign n76881 = ~n35214 ;
  assign n35245 = x67 & n76881 ;
  assign n76882 = ~n35208 ;
  assign n35246 = n76882 & n35245 ;
  assign n35247 = n35216 | n35246 ;
  assign n35248 = n35244 | n35247 ;
  assign n76883 = ~n35216 ;
  assign n35249 = n76883 & n35248 ;
  assign n76884 = ~n35205 ;
  assign n35250 = x68 & n76884 ;
  assign n76885 = ~n35199 ;
  assign n35251 = n76885 & n35250 ;
  assign n35252 = n35207 | n35251 ;
  assign n35253 = n35249 | n35252 ;
  assign n76886 = ~n35207 ;
  assign n35254 = n76886 & n35253 ;
  assign n76887 = ~n35196 ;
  assign n35255 = x69 & n76887 ;
  assign n76888 = ~n35190 ;
  assign n35256 = n76888 & n35255 ;
  assign n35257 = n35198 | n35256 ;
  assign n35258 = n35254 | n35257 ;
  assign n76889 = ~n35198 ;
  assign n35259 = n76889 & n35258 ;
  assign n76890 = ~n35187 ;
  assign n35260 = x70 & n76890 ;
  assign n76891 = ~n35181 ;
  assign n35261 = n76891 & n35260 ;
  assign n35262 = n35189 | n35261 ;
  assign n35264 = n35259 | n35262 ;
  assign n76892 = ~n35189 ;
  assign n35265 = n76892 & n35264 ;
  assign n76893 = ~n35178 ;
  assign n35266 = x71 & n76893 ;
  assign n76894 = ~n35173 ;
  assign n35267 = n76894 & n35266 ;
  assign n35268 = n35180 | n35267 ;
  assign n35269 = n35265 | n35268 ;
  assign n76895 = ~n35180 ;
  assign n35270 = n76895 & n35269 ;
  assign n76896 = ~n35170 ;
  assign n35271 = x72 & n76896 ;
  assign n76897 = ~n35165 ;
  assign n35272 = n76897 & n35271 ;
  assign n35273 = n35172 | n35272 ;
  assign n35275 = n35270 | n35273 ;
  assign n76898 = ~n35172 ;
  assign n35276 = n76898 & n35275 ;
  assign n76899 = ~n35162 ;
  assign n35277 = x73 & n76899 ;
  assign n76900 = ~n35157 ;
  assign n35278 = n76900 & n35277 ;
  assign n35279 = n35164 | n35278 ;
  assign n35280 = n35276 | n35279 ;
  assign n76901 = ~n35164 ;
  assign n35281 = n76901 & n35280 ;
  assign n76902 = ~n35154 ;
  assign n35282 = x74 & n76902 ;
  assign n76903 = ~n35149 ;
  assign n35283 = n76903 & n35282 ;
  assign n35284 = n35156 | n35283 ;
  assign n35286 = n35281 | n35284 ;
  assign n76904 = ~n35156 ;
  assign n35287 = n76904 & n35286 ;
  assign n76905 = ~n35146 ;
  assign n35288 = x75 & n76905 ;
  assign n76906 = ~n35141 ;
  assign n35289 = n76906 & n35288 ;
  assign n35290 = n35148 | n35289 ;
  assign n35291 = n35287 | n35290 ;
  assign n76907 = ~n35148 ;
  assign n35292 = n76907 & n35291 ;
  assign n76908 = ~n35138 ;
  assign n35293 = x76 & n76908 ;
  assign n76909 = ~n35133 ;
  assign n35294 = n76909 & n35293 ;
  assign n35295 = n35140 | n35294 ;
  assign n35297 = n35292 | n35295 ;
  assign n76910 = ~n35140 ;
  assign n35298 = n76910 & n35297 ;
  assign n76911 = ~n35130 ;
  assign n35299 = x77 & n76911 ;
  assign n76912 = ~n35125 ;
  assign n35300 = n76912 & n35299 ;
  assign n35301 = n35132 | n35300 ;
  assign n35302 = n35298 | n35301 ;
  assign n76913 = ~n35132 ;
  assign n35303 = n76913 & n35302 ;
  assign n76914 = ~n35122 ;
  assign n35304 = x78 & n76914 ;
  assign n76915 = ~n35117 ;
  assign n35305 = n76915 & n35304 ;
  assign n35306 = n35124 | n35305 ;
  assign n35308 = n35303 | n35306 ;
  assign n76916 = ~n35124 ;
  assign n35309 = n76916 & n35308 ;
  assign n76917 = ~n35114 ;
  assign n35310 = x79 & n76917 ;
  assign n76918 = ~n35109 ;
  assign n35311 = n76918 & n35310 ;
  assign n35312 = n35116 | n35311 ;
  assign n35313 = n35309 | n35312 ;
  assign n76919 = ~n35116 ;
  assign n35314 = n76919 & n35313 ;
  assign n76920 = ~n35106 ;
  assign n35315 = x80 & n76920 ;
  assign n76921 = ~n35067 ;
  assign n35316 = n76921 & n35315 ;
  assign n35317 = n35108 | n35316 ;
  assign n35319 = n35314 | n35317 ;
  assign n76922 = ~n35108 ;
  assign n35320 = n76922 & n35319 ;
  assign n35327 = n66505 & n35326 ;
  assign n76923 = ~n35064 ;
  assign n35328 = n76923 & n35324 ;
  assign n35329 = n34856 & n35064 ;
  assign n76924 = ~n35329 ;
  assign n35330 = x81 & n76924 ;
  assign n76925 = ~n35328 ;
  assign n35331 = n76925 & n35330 ;
  assign n35332 = n2875 | n35331 ;
  assign n35333 = n35327 | n35332 ;
  assign n35335 = n35320 | n35333 ;
  assign n76926 = ~n35334 ;
  assign n35336 = n76926 & n35335 ;
  assign n76927 = ~n35314 ;
  assign n35318 = n76927 & n35317 ;
  assign n35339 = x65 & n35230 ;
  assign n76928 = ~n35339 ;
  assign n35340 = n35236 & n76928 ;
  assign n35341 = n2773 | n35340 ;
  assign n35342 = n76877 & n35341 ;
  assign n35343 = n35222 | n35242 ;
  assign n35345 = n35342 | n35343 ;
  assign n35346 = n76880 & n35345 ;
  assign n35347 = n35246 | n35346 ;
  assign n35349 = n76883 & n35347 ;
  assign n35351 = n35252 | n35349 ;
  assign n35352 = n76886 & n35351 ;
  assign n35354 = n35257 | n35352 ;
  assign n35355 = n76889 & n35354 ;
  assign n35356 = n35262 | n35355 ;
  assign n35357 = n76892 & n35356 ;
  assign n35358 = n35268 | n35357 ;
  assign n35360 = n76895 & n35358 ;
  assign n35361 = n35273 | n35360 ;
  assign n35362 = n76898 & n35361 ;
  assign n35363 = n35279 | n35362 ;
  assign n35365 = n76901 & n35363 ;
  assign n35366 = n35284 | n35365 ;
  assign n35367 = n76904 & n35366 ;
  assign n35368 = n35290 | n35367 ;
  assign n35370 = n76907 & n35368 ;
  assign n35371 = n35295 | n35370 ;
  assign n35372 = n76910 & n35371 ;
  assign n35373 = n35301 | n35372 ;
  assign n35375 = n76913 & n35373 ;
  assign n35376 = n35306 | n35375 ;
  assign n35377 = n76916 & n35376 ;
  assign n35378 = n35312 | n35377 ;
  assign n35380 = n35116 | n35317 ;
  assign n76929 = ~n35380 ;
  assign n35381 = n35378 & n76929 ;
  assign n35382 = n35318 | n35381 ;
  assign n76930 = ~n35336 ;
  assign n35383 = n76930 & n35382 ;
  assign n35384 = n76919 & n35378 ;
  assign n35385 = n35317 | n35384 ;
  assign n35386 = n76922 & n35385 ;
  assign n35387 = n35333 | n35386 ;
  assign n35388 = n35107 & n76926 ;
  assign n35389 = n35387 & n35388 ;
  assign n35390 = n35383 | n35389 ;
  assign n35391 = n35108 | n35331 ;
  assign n35392 = n35327 | n35391 ;
  assign n76931 = ~n35392 ;
  assign n35393 = n35319 & n76931 ;
  assign n35394 = n35327 | n35331 ;
  assign n76932 = ~n35386 ;
  assign n35395 = n76932 & n35394 ;
  assign n35396 = n35393 | n35395 ;
  assign n35397 = n76930 & n35396 ;
  assign n35398 = n344 & n34856 ;
  assign n35399 = n35387 & n35398 ;
  assign n35400 = n35397 | n35399 ;
  assign n35401 = n66560 & n35400 ;
  assign n76933 = ~n35399 ;
  assign n35628 = x82 & n76933 ;
  assign n76934 = ~n35397 ;
  assign n35629 = n76934 & n35628 ;
  assign n35630 = n35401 | n35629 ;
  assign n35402 = n66505 & n35390 ;
  assign n76935 = ~n35377 ;
  assign n35379 = n35312 & n76935 ;
  assign n35403 = n35124 | n35312 ;
  assign n76936 = ~n35403 ;
  assign n35404 = n35308 & n76936 ;
  assign n35405 = n35379 | n35404 ;
  assign n35406 = n76930 & n35405 ;
  assign n35407 = n35115 & n76926 ;
  assign n35408 = n35387 & n35407 ;
  assign n35409 = n35406 | n35408 ;
  assign n35410 = n66379 & n35409 ;
  assign n76937 = ~n35408 ;
  assign n35616 = x80 & n76937 ;
  assign n76938 = ~n35406 ;
  assign n35617 = n76938 & n35616 ;
  assign n35618 = n35410 | n35617 ;
  assign n76939 = ~n35303 ;
  assign n35307 = n76939 & n35306 ;
  assign n35411 = n35132 | n35306 ;
  assign n76940 = ~n35411 ;
  assign n35412 = n35373 & n76940 ;
  assign n35413 = n35307 | n35412 ;
  assign n35414 = n76930 & n35413 ;
  assign n35415 = n35123 & n76926 ;
  assign n35416 = n35387 & n35415 ;
  assign n35417 = n35414 | n35416 ;
  assign n35418 = n66299 & n35417 ;
  assign n76941 = ~n35372 ;
  assign n35374 = n35301 & n76941 ;
  assign n35419 = n35140 | n35301 ;
  assign n76942 = ~n35419 ;
  assign n35420 = n35297 & n76942 ;
  assign n35421 = n35374 | n35420 ;
  assign n35422 = n76930 & n35421 ;
  assign n35423 = n35131 & n76926 ;
  assign n35424 = n35387 & n35423 ;
  assign n35425 = n35422 | n35424 ;
  assign n35426 = n66244 & n35425 ;
  assign n76943 = ~n35424 ;
  assign n35604 = x78 & n76943 ;
  assign n76944 = ~n35422 ;
  assign n35605 = n76944 & n35604 ;
  assign n35606 = n35426 | n35605 ;
  assign n76945 = ~n35292 ;
  assign n35296 = n76945 & n35295 ;
  assign n35427 = n35148 | n35295 ;
  assign n76946 = ~n35427 ;
  assign n35428 = n35368 & n76946 ;
  assign n35429 = n35296 | n35428 ;
  assign n35430 = n76930 & n35429 ;
  assign n35431 = n35139 & n76926 ;
  assign n35432 = n35387 & n35431 ;
  assign n35433 = n35430 | n35432 ;
  assign n35434 = n66145 & n35433 ;
  assign n76947 = ~n35367 ;
  assign n35369 = n35290 & n76947 ;
  assign n35435 = n35156 | n35290 ;
  assign n76948 = ~n35435 ;
  assign n35436 = n35286 & n76948 ;
  assign n35437 = n35369 | n35436 ;
  assign n35438 = n76930 & n35437 ;
  assign n35439 = n35147 & n76926 ;
  assign n35440 = n35387 & n35439 ;
  assign n35441 = n35438 | n35440 ;
  assign n35442 = n66081 & n35441 ;
  assign n76949 = ~n35440 ;
  assign n35592 = x76 & n76949 ;
  assign n76950 = ~n35438 ;
  assign n35593 = n76950 & n35592 ;
  assign n35594 = n35442 | n35593 ;
  assign n76951 = ~n35281 ;
  assign n35285 = n76951 & n35284 ;
  assign n35443 = n35164 | n35284 ;
  assign n76952 = ~n35443 ;
  assign n35444 = n35363 & n76952 ;
  assign n35445 = n35285 | n35444 ;
  assign n35446 = n76930 & n35445 ;
  assign n35447 = n35155 & n76926 ;
  assign n35448 = n35387 & n35447 ;
  assign n35449 = n35446 | n35448 ;
  assign n35450 = n66043 & n35449 ;
  assign n76953 = ~n35362 ;
  assign n35364 = n35279 & n76953 ;
  assign n35451 = n35172 | n35279 ;
  assign n76954 = ~n35451 ;
  assign n35452 = n35275 & n76954 ;
  assign n35453 = n35364 | n35452 ;
  assign n35454 = n76930 & n35453 ;
  assign n35455 = n35163 & n76926 ;
  assign n35456 = n35387 & n35455 ;
  assign n35457 = n35454 | n35456 ;
  assign n35458 = n65960 & n35457 ;
  assign n76955 = ~n35456 ;
  assign n35580 = x74 & n76955 ;
  assign n76956 = ~n35454 ;
  assign n35581 = n76956 & n35580 ;
  assign n35582 = n35458 | n35581 ;
  assign n76957 = ~n35270 ;
  assign n35274 = n76957 & n35273 ;
  assign n35459 = n35180 | n35273 ;
  assign n76958 = ~n35459 ;
  assign n35460 = n35358 & n76958 ;
  assign n35461 = n35274 | n35460 ;
  assign n35462 = n76930 & n35461 ;
  assign n35463 = n35171 & n76926 ;
  assign n35464 = n35387 & n35463 ;
  assign n35465 = n35462 | n35464 ;
  assign n35466 = n65909 & n35465 ;
  assign n76959 = ~n35357 ;
  assign n35359 = n35268 & n76959 ;
  assign n35467 = n35189 | n35268 ;
  assign n76960 = ~n35467 ;
  assign n35468 = n35264 & n76960 ;
  assign n35469 = n35359 | n35468 ;
  assign n35470 = n76930 & n35469 ;
  assign n35471 = n35179 & n76926 ;
  assign n35472 = n35387 & n35471 ;
  assign n35473 = n35470 | n35472 ;
  assign n35474 = n65877 & n35473 ;
  assign n76961 = ~n35472 ;
  assign n35568 = x72 & n76961 ;
  assign n76962 = ~n35470 ;
  assign n35569 = n76962 & n35568 ;
  assign n35570 = n35474 | n35569 ;
  assign n76963 = ~n35259 ;
  assign n35263 = n76963 & n35262 ;
  assign n35475 = n35198 | n35262 ;
  assign n76964 = ~n35475 ;
  assign n35476 = n35354 & n76964 ;
  assign n35477 = n35263 | n35476 ;
  assign n35478 = n76930 & n35477 ;
  assign n35479 = n35188 & n76926 ;
  assign n35480 = n35387 & n35479 ;
  assign n35481 = n35478 | n35480 ;
  assign n35482 = n65820 & n35481 ;
  assign n76965 = ~n35352 ;
  assign n35353 = n35257 & n76965 ;
  assign n35483 = n35207 | n35257 ;
  assign n76966 = ~n35483 ;
  assign n35484 = n35253 & n76966 ;
  assign n35485 = n35353 | n35484 ;
  assign n35486 = n76930 & n35485 ;
  assign n35487 = n35197 & n76926 ;
  assign n35488 = n35387 & n35487 ;
  assign n35489 = n35486 | n35488 ;
  assign n35490 = n65791 & n35489 ;
  assign n76967 = ~n35488 ;
  assign n35556 = x70 & n76967 ;
  assign n76968 = ~n35486 ;
  assign n35557 = n76968 & n35556 ;
  assign n35558 = n35490 | n35557 ;
  assign n76969 = ~n35249 ;
  assign n35350 = n76969 & n35252 ;
  assign n35491 = n35247 | n35346 ;
  assign n35492 = n35216 | n35252 ;
  assign n76970 = ~n35492 ;
  assign n35493 = n35491 & n76970 ;
  assign n35494 = n35350 | n35493 ;
  assign n35495 = n76930 & n35494 ;
  assign n35496 = n35206 & n76926 ;
  assign n35497 = n35387 & n35496 ;
  assign n35498 = n35495 | n35497 ;
  assign n35499 = n65772 & n35498 ;
  assign n76971 = ~n35346 ;
  assign n35348 = n35247 & n76971 ;
  assign n35500 = n35222 | n35247 ;
  assign n76972 = ~n35500 ;
  assign n35501 = n35345 & n76972 ;
  assign n35502 = n35348 | n35501 ;
  assign n35503 = n76930 & n35502 ;
  assign n35504 = n35215 & n76926 ;
  assign n35505 = n35387 & n35504 ;
  assign n35506 = n35503 | n35505 ;
  assign n35507 = n65746 & n35506 ;
  assign n76973 = ~n35505 ;
  assign n35545 = x68 & n76973 ;
  assign n76974 = ~n35503 ;
  assign n35546 = n76974 & n35545 ;
  assign n35547 = n35507 | n35546 ;
  assign n76975 = ~n35240 ;
  assign n35344 = n76975 & n35343 ;
  assign n35508 = n35238 | n35343 ;
  assign n76976 = ~n35508 ;
  assign n35509 = n35239 & n76976 ;
  assign n35510 = n35344 | n35509 ;
  assign n35511 = n76930 & n35510 ;
  assign n35512 = n35221 & n76926 ;
  assign n35513 = n35387 & n35512 ;
  assign n35514 = n35511 | n35513 ;
  assign n35515 = n65721 & n35514 ;
  assign n35516 = n2773 & n35236 ;
  assign n35517 = n76928 & n35516 ;
  assign n76977 = ~n35517 ;
  assign n35518 = n35239 & n76977 ;
  assign n35519 = n76930 & n35518 ;
  assign n35520 = n35230 & n76926 ;
  assign n35521 = n35387 & n35520 ;
  assign n35522 = n35519 | n35521 ;
  assign n35523 = n65686 & n35522 ;
  assign n76978 = ~n35521 ;
  assign n35535 = x66 & n76978 ;
  assign n76979 = ~n35519 ;
  assign n35536 = n76979 & n35535 ;
  assign n35537 = n35523 | n35536 ;
  assign n35338 = n2773 & n76930 ;
  assign n35337 = x64 & n76930 ;
  assign n76980 = ~n35337 ;
  assign n35524 = x46 & n76980 ;
  assign n35525 = n35338 | n35524 ;
  assign n35526 = x65 & n35525 ;
  assign n35527 = n76926 & n35387 ;
  assign n76981 = ~n35527 ;
  assign n35528 = n2773 & n76981 ;
  assign n35529 = x65 | n35528 ;
  assign n35530 = n35524 | n35529 ;
  assign n76982 = ~n35526 ;
  assign n35531 = n76982 & n35530 ;
  assign n35533 = n3081 | n35531 ;
  assign n35534 = n65670 & n35525 ;
  assign n76983 = ~n35534 ;
  assign n35538 = n35533 & n76983 ;
  assign n35539 = n35537 | n35538 ;
  assign n76984 = ~n35523 ;
  assign n35540 = n76984 & n35539 ;
  assign n76985 = ~n35513 ;
  assign n35541 = x67 & n76985 ;
  assign n76986 = ~n35511 ;
  assign n35542 = n76986 & n35541 ;
  assign n35543 = n35515 | n35542 ;
  assign n35544 = n35540 | n35543 ;
  assign n76987 = ~n35515 ;
  assign n35548 = n76987 & n35544 ;
  assign n35549 = n35547 | n35548 ;
  assign n76988 = ~n35507 ;
  assign n35550 = n76988 & n35549 ;
  assign n76989 = ~n35497 ;
  assign n35551 = x69 & n76989 ;
  assign n76990 = ~n35495 ;
  assign n35552 = n76990 & n35551 ;
  assign n35553 = n35499 | n35552 ;
  assign n35555 = n35550 | n35553 ;
  assign n76991 = ~n35499 ;
  assign n35560 = n76991 & n35555 ;
  assign n35561 = n35558 | n35560 ;
  assign n76992 = ~n35490 ;
  assign n35562 = n76992 & n35561 ;
  assign n76993 = ~n35480 ;
  assign n35563 = x71 & n76993 ;
  assign n76994 = ~n35478 ;
  assign n35564 = n76994 & n35563 ;
  assign n35565 = n35482 | n35564 ;
  assign n35567 = n35562 | n35565 ;
  assign n76995 = ~n35482 ;
  assign n35572 = n76995 & n35567 ;
  assign n35573 = n35570 | n35572 ;
  assign n76996 = ~n35474 ;
  assign n35574 = n76996 & n35573 ;
  assign n76997 = ~n35464 ;
  assign n35575 = x73 & n76997 ;
  assign n76998 = ~n35462 ;
  assign n35576 = n76998 & n35575 ;
  assign n35577 = n35466 | n35576 ;
  assign n35579 = n35574 | n35577 ;
  assign n76999 = ~n35466 ;
  assign n35584 = n76999 & n35579 ;
  assign n35585 = n35582 | n35584 ;
  assign n77000 = ~n35458 ;
  assign n35586 = n77000 & n35585 ;
  assign n77001 = ~n35448 ;
  assign n35587 = x75 & n77001 ;
  assign n77002 = ~n35446 ;
  assign n35588 = n77002 & n35587 ;
  assign n35589 = n35450 | n35588 ;
  assign n35591 = n35586 | n35589 ;
  assign n77003 = ~n35450 ;
  assign n35596 = n77003 & n35591 ;
  assign n35597 = n35594 | n35596 ;
  assign n77004 = ~n35442 ;
  assign n35598 = n77004 & n35597 ;
  assign n77005 = ~n35432 ;
  assign n35599 = x77 & n77005 ;
  assign n77006 = ~n35430 ;
  assign n35600 = n77006 & n35599 ;
  assign n35601 = n35434 | n35600 ;
  assign n35603 = n35598 | n35601 ;
  assign n77007 = ~n35434 ;
  assign n35608 = n77007 & n35603 ;
  assign n35609 = n35606 | n35608 ;
  assign n77008 = ~n35426 ;
  assign n35610 = n77008 & n35609 ;
  assign n77009 = ~n35416 ;
  assign n35611 = x79 & n77009 ;
  assign n77010 = ~n35414 ;
  assign n35612 = n77010 & n35611 ;
  assign n35613 = n35418 | n35612 ;
  assign n35615 = n35610 | n35613 ;
  assign n77011 = ~n35418 ;
  assign n35620 = n77011 & n35615 ;
  assign n35621 = n35618 | n35620 ;
  assign n77012 = ~n35410 ;
  assign n35622 = n77012 & n35621 ;
  assign n77013 = ~n35389 ;
  assign n35623 = x81 & n77013 ;
  assign n77014 = ~n35383 ;
  assign n35624 = n77014 & n35623 ;
  assign n35625 = n35402 | n35624 ;
  assign n35627 = n35622 | n35625 ;
  assign n77015 = ~n35402 ;
  assign n35631 = n77015 & n35627 ;
  assign n35632 = n35630 | n35631 ;
  assign n77016 = ~n35401 ;
  assign n35633 = n77016 & n35632 ;
  assign n35634 = n3180 | n35633 ;
  assign n35637 = n35390 & n35634 ;
  assign n35626 = n35410 | n35625 ;
  assign n35638 = x64 & n76981 ;
  assign n77017 = ~n35638 ;
  assign n35639 = x46 & n77017 ;
  assign n35640 = n35338 | n35639 ;
  assign n35641 = x65 & n35640 ;
  assign n77018 = ~n35641 ;
  assign n35642 = n35530 & n77018 ;
  assign n35643 = n3081 | n35642 ;
  assign n35644 = n76983 & n35643 ;
  assign n35646 = n35537 | n35644 ;
  assign n35647 = n76984 & n35646 ;
  assign n35648 = n35543 | n35647 ;
  assign n35649 = n76987 & n35648 ;
  assign n35650 = n35547 | n35649 ;
  assign n35651 = n76988 & n35650 ;
  assign n35652 = n35553 | n35651 ;
  assign n35653 = n76991 & n35652 ;
  assign n35654 = n35558 | n35653 ;
  assign n35655 = n76992 & n35654 ;
  assign n35656 = n35565 | n35655 ;
  assign n35657 = n76995 & n35656 ;
  assign n35658 = n35570 | n35657 ;
  assign n35659 = n76996 & n35658 ;
  assign n35660 = n35577 | n35659 ;
  assign n35661 = n76999 & n35660 ;
  assign n35662 = n35582 | n35661 ;
  assign n35663 = n77000 & n35662 ;
  assign n35664 = n35589 | n35663 ;
  assign n35665 = n77003 & n35664 ;
  assign n35666 = n35594 | n35665 ;
  assign n35667 = n77004 & n35666 ;
  assign n35668 = n35601 | n35667 ;
  assign n35669 = n77007 & n35668 ;
  assign n35670 = n35606 | n35669 ;
  assign n35671 = n77008 & n35670 ;
  assign n35672 = n35613 | n35671 ;
  assign n35673 = n77011 & n35672 ;
  assign n35674 = n35618 | n35673 ;
  assign n77019 = ~n35626 ;
  assign n35675 = n77019 & n35674 ;
  assign n35676 = n77012 & n35674 ;
  assign n77020 = ~n35676 ;
  assign n35677 = n35625 & n77020 ;
  assign n35678 = n35675 | n35677 ;
  assign n35679 = n66660 & n35678 ;
  assign n77021 = ~n35633 ;
  assign n35680 = n77021 & n35679 ;
  assign n35681 = n35637 | n35680 ;
  assign n77022 = ~n35400 ;
  assign n35635 = n77022 & n35634 ;
  assign n77023 = ~n35631 ;
  assign n35684 = n35630 & n77023 ;
  assign n35682 = n35625 | n35676 ;
  assign n35685 = n35402 | n35630 ;
  assign n77024 = ~n35685 ;
  assign n35686 = n35682 & n77024 ;
  assign n35687 = n35684 | n35686 ;
  assign n35688 = n35634 | n35687 ;
  assign n77025 = ~n35635 ;
  assign n35689 = n77025 & n35688 ;
  assign n35690 = n66654 & n35689 ;
  assign n35691 = n66560 & n35681 ;
  assign n35692 = n35409 & n35634 ;
  assign n35619 = n35418 | n35618 ;
  assign n77026 = ~n35619 ;
  assign n35693 = n35615 & n77026 ;
  assign n77027 = ~n35620 ;
  assign n35694 = n35618 & n77027 ;
  assign n35695 = n35693 | n35694 ;
  assign n35696 = n66660 & n35695 ;
  assign n35697 = n77021 & n35696 ;
  assign n35698 = n35692 | n35697 ;
  assign n35699 = n66505 & n35698 ;
  assign n35700 = n35417 & n35634 ;
  assign n35614 = n35426 | n35613 ;
  assign n77028 = ~n35614 ;
  assign n35701 = n77028 & n35670 ;
  assign n77029 = ~n35671 ;
  assign n35702 = n35613 & n77029 ;
  assign n35703 = n35701 | n35702 ;
  assign n35704 = n66660 & n35703 ;
  assign n35705 = n77021 & n35704 ;
  assign n35706 = n35700 | n35705 ;
  assign n35707 = n66379 & n35706 ;
  assign n35708 = n35425 & n35634 ;
  assign n35607 = n35434 | n35606 ;
  assign n77030 = ~n35607 ;
  assign n35709 = n35603 & n77030 ;
  assign n77031 = ~n35608 ;
  assign n35710 = n35606 & n77031 ;
  assign n35711 = n35709 | n35710 ;
  assign n35712 = n66660 & n35711 ;
  assign n35713 = n77021 & n35712 ;
  assign n35714 = n35708 | n35713 ;
  assign n35715 = n66299 & n35714 ;
  assign n35716 = n35433 & n35634 ;
  assign n35602 = n35442 | n35601 ;
  assign n77032 = ~n35602 ;
  assign n35717 = n77032 & n35666 ;
  assign n77033 = ~n35667 ;
  assign n35718 = n35601 & n77033 ;
  assign n35719 = n35717 | n35718 ;
  assign n35720 = n66660 & n35719 ;
  assign n35721 = n77021 & n35720 ;
  assign n35722 = n35716 | n35721 ;
  assign n35723 = n66244 & n35722 ;
  assign n35724 = n35441 & n35634 ;
  assign n35595 = n35450 | n35594 ;
  assign n77034 = ~n35595 ;
  assign n35725 = n35591 & n77034 ;
  assign n77035 = ~n35596 ;
  assign n35726 = n35594 & n77035 ;
  assign n35727 = n35725 | n35726 ;
  assign n35728 = n66660 & n35727 ;
  assign n35729 = n77021 & n35728 ;
  assign n35730 = n35724 | n35729 ;
  assign n35731 = n66145 & n35730 ;
  assign n35732 = n35449 & n35634 ;
  assign n35590 = n35458 | n35589 ;
  assign n77036 = ~n35590 ;
  assign n35733 = n77036 & n35662 ;
  assign n77037 = ~n35663 ;
  assign n35734 = n35589 & n77037 ;
  assign n35735 = n35733 | n35734 ;
  assign n35736 = n66660 & n35735 ;
  assign n35737 = n77021 & n35736 ;
  assign n35738 = n35732 | n35737 ;
  assign n35739 = n66081 & n35738 ;
  assign n35740 = n35457 & n35634 ;
  assign n35583 = n35466 | n35582 ;
  assign n77038 = ~n35583 ;
  assign n35741 = n35579 & n77038 ;
  assign n77039 = ~n35584 ;
  assign n35742 = n35582 & n77039 ;
  assign n35743 = n35741 | n35742 ;
  assign n35744 = n66660 & n35743 ;
  assign n35745 = n77021 & n35744 ;
  assign n35746 = n35740 | n35745 ;
  assign n35747 = n66043 & n35746 ;
  assign n35748 = n35465 & n35634 ;
  assign n35578 = n35474 | n35577 ;
  assign n77040 = ~n35578 ;
  assign n35749 = n77040 & n35658 ;
  assign n77041 = ~n35659 ;
  assign n35750 = n35577 & n77041 ;
  assign n35751 = n35749 | n35750 ;
  assign n35752 = n66660 & n35751 ;
  assign n35753 = n77021 & n35752 ;
  assign n35754 = n35748 | n35753 ;
  assign n35755 = n65960 & n35754 ;
  assign n35756 = n35473 & n35634 ;
  assign n35571 = n35482 | n35570 ;
  assign n77042 = ~n35571 ;
  assign n35757 = n35567 & n77042 ;
  assign n77043 = ~n35572 ;
  assign n35758 = n35570 & n77043 ;
  assign n35759 = n35757 | n35758 ;
  assign n35760 = n66660 & n35759 ;
  assign n35761 = n77021 & n35760 ;
  assign n35762 = n35756 | n35761 ;
  assign n35763 = n65909 & n35762 ;
  assign n35764 = n35481 & n35634 ;
  assign n35566 = n35490 | n35565 ;
  assign n77044 = ~n35566 ;
  assign n35765 = n77044 & n35654 ;
  assign n77045 = ~n35655 ;
  assign n35766 = n35565 & n77045 ;
  assign n35767 = n35765 | n35766 ;
  assign n35768 = n66660 & n35767 ;
  assign n35769 = n77021 & n35768 ;
  assign n35770 = n35764 | n35769 ;
  assign n35771 = n65877 & n35770 ;
  assign n35772 = n35489 & n35634 ;
  assign n35559 = n35499 | n35558 ;
  assign n77046 = ~n35559 ;
  assign n35773 = n35555 & n77046 ;
  assign n77047 = ~n35560 ;
  assign n35774 = n35558 & n77047 ;
  assign n35775 = n35773 | n35774 ;
  assign n35776 = n66660 & n35775 ;
  assign n35777 = n77021 & n35776 ;
  assign n35778 = n35772 | n35777 ;
  assign n35779 = n65820 & n35778 ;
  assign n35780 = n35498 & n35634 ;
  assign n35554 = n35507 | n35553 ;
  assign n77048 = ~n35554 ;
  assign n35781 = n77048 & n35650 ;
  assign n77049 = ~n35651 ;
  assign n35782 = n35553 & n77049 ;
  assign n35783 = n35781 | n35782 ;
  assign n35784 = n66660 & n35783 ;
  assign n35785 = n77021 & n35784 ;
  assign n35786 = n35780 | n35785 ;
  assign n35787 = n65791 & n35786 ;
  assign n35788 = n35506 & n35634 ;
  assign n35789 = n35515 | n35547 ;
  assign n77050 = ~n35789 ;
  assign n35790 = n35544 & n77050 ;
  assign n77051 = ~n35548 ;
  assign n35791 = n35547 & n77051 ;
  assign n35792 = n35790 | n35791 ;
  assign n35793 = n66660 & n35792 ;
  assign n35794 = n77021 & n35793 ;
  assign n35795 = n35788 | n35794 ;
  assign n35796 = n65772 & n35795 ;
  assign n35797 = n35514 & n35634 ;
  assign n35798 = n35523 | n35543 ;
  assign n77052 = ~n35798 ;
  assign n35799 = n35539 & n77052 ;
  assign n77053 = ~n35647 ;
  assign n35800 = n35543 & n77053 ;
  assign n35801 = n35799 | n35800 ;
  assign n35802 = n66660 & n35801 ;
  assign n35803 = n77021 & n35802 ;
  assign n35804 = n35797 | n35803 ;
  assign n35805 = n65746 & n35804 ;
  assign n35806 = n35522 & n35634 ;
  assign n35645 = n35534 | n35537 ;
  assign n77054 = ~n35645 ;
  assign n35807 = n35643 & n77054 ;
  assign n77055 = ~n35538 ;
  assign n35808 = n35537 & n77055 ;
  assign n35809 = n35807 | n35808 ;
  assign n35810 = n66660 & n35809 ;
  assign n35811 = n77021 & n35810 ;
  assign n35812 = n35806 | n35811 ;
  assign n35813 = n65721 & n35812 ;
  assign n35636 = n35525 & n35634 ;
  assign n35532 = n3081 & n35530 ;
  assign n35815 = n35532 & n77018 ;
  assign n35816 = n3180 | n35815 ;
  assign n77056 = ~n35816 ;
  assign n35817 = n35643 & n77056 ;
  assign n35818 = n77021 & n35817 ;
  assign n35819 = n35636 | n35818 ;
  assign n35820 = n65686 & n35819 ;
  assign n35814 = n3382 & n77021 ;
  assign n35821 = n3375 & n77021 ;
  assign n77057 = ~n35821 ;
  assign n35822 = x45 & n77057 ;
  assign n35823 = n35814 | n35822 ;
  assign n35824 = n65670 & n35823 ;
  assign n35683 = n77015 & n35682 ;
  assign n35826 = n35630 | n35683 ;
  assign n35827 = n77016 & n35826 ;
  assign n77058 = ~n35827 ;
  assign n35828 = n3375 & n77058 ;
  assign n77059 = ~n35828 ;
  assign n35829 = x45 & n77059 ;
  assign n35830 = n35814 | n35829 ;
  assign n35832 = x65 & n35830 ;
  assign n35831 = x65 | n35814 ;
  assign n35833 = n35822 | n35831 ;
  assign n77060 = ~n35832 ;
  assign n35834 = n77060 & n35833 ;
  assign n35835 = n3393 | n35834 ;
  assign n77061 = ~n35824 ;
  assign n35836 = n77061 & n35835 ;
  assign n77062 = ~n35818 ;
  assign n35837 = x66 & n77062 ;
  assign n77063 = ~n35636 ;
  assign n35838 = n77063 & n35837 ;
  assign n35839 = n35820 | n35838 ;
  assign n35840 = n35836 | n35839 ;
  assign n77064 = ~n35820 ;
  assign n35841 = n77064 & n35840 ;
  assign n77065 = ~n35811 ;
  assign n35842 = x67 & n77065 ;
  assign n77066 = ~n35806 ;
  assign n35843 = n77066 & n35842 ;
  assign n35844 = n35841 | n35843 ;
  assign n77067 = ~n35813 ;
  assign n35845 = n77067 & n35844 ;
  assign n77068 = ~n35803 ;
  assign n35846 = x68 & n77068 ;
  assign n77069 = ~n35797 ;
  assign n35847 = n77069 & n35846 ;
  assign n35848 = n35805 | n35847 ;
  assign n35849 = n35845 | n35848 ;
  assign n77070 = ~n35805 ;
  assign n35850 = n77070 & n35849 ;
  assign n77071 = ~n35794 ;
  assign n35851 = x69 & n77071 ;
  assign n77072 = ~n35788 ;
  assign n35852 = n77072 & n35851 ;
  assign n35853 = n35796 | n35852 ;
  assign n35854 = n35850 | n35853 ;
  assign n77073 = ~n35796 ;
  assign n35855 = n77073 & n35854 ;
  assign n77074 = ~n35785 ;
  assign n35856 = x70 & n77074 ;
  assign n77075 = ~n35780 ;
  assign n35857 = n77075 & n35856 ;
  assign n35858 = n35787 | n35857 ;
  assign n35859 = n35855 | n35858 ;
  assign n77076 = ~n35787 ;
  assign n35860 = n77076 & n35859 ;
  assign n77077 = ~n35777 ;
  assign n35861 = x71 & n77077 ;
  assign n77078 = ~n35772 ;
  assign n35862 = n77078 & n35861 ;
  assign n35863 = n35779 | n35862 ;
  assign n35865 = n35860 | n35863 ;
  assign n77079 = ~n35779 ;
  assign n35866 = n77079 & n35865 ;
  assign n77080 = ~n35769 ;
  assign n35867 = x72 & n77080 ;
  assign n77081 = ~n35764 ;
  assign n35868 = n77081 & n35867 ;
  assign n35869 = n35771 | n35868 ;
  assign n35870 = n35866 | n35869 ;
  assign n77082 = ~n35771 ;
  assign n35871 = n77082 & n35870 ;
  assign n77083 = ~n35761 ;
  assign n35872 = x73 & n77083 ;
  assign n77084 = ~n35756 ;
  assign n35873 = n77084 & n35872 ;
  assign n35874 = n35763 | n35873 ;
  assign n35876 = n35871 | n35874 ;
  assign n77085 = ~n35763 ;
  assign n35877 = n77085 & n35876 ;
  assign n77086 = ~n35753 ;
  assign n35878 = x74 & n77086 ;
  assign n77087 = ~n35748 ;
  assign n35879 = n77087 & n35878 ;
  assign n35880 = n35755 | n35879 ;
  assign n35881 = n35877 | n35880 ;
  assign n77088 = ~n35755 ;
  assign n35882 = n77088 & n35881 ;
  assign n77089 = ~n35745 ;
  assign n35883 = x75 & n77089 ;
  assign n77090 = ~n35740 ;
  assign n35884 = n77090 & n35883 ;
  assign n35885 = n35747 | n35884 ;
  assign n35887 = n35882 | n35885 ;
  assign n77091 = ~n35747 ;
  assign n35888 = n77091 & n35887 ;
  assign n77092 = ~n35737 ;
  assign n35889 = x76 & n77092 ;
  assign n77093 = ~n35732 ;
  assign n35890 = n77093 & n35889 ;
  assign n35891 = n35739 | n35890 ;
  assign n35892 = n35888 | n35891 ;
  assign n77094 = ~n35739 ;
  assign n35893 = n77094 & n35892 ;
  assign n77095 = ~n35729 ;
  assign n35894 = x77 & n77095 ;
  assign n77096 = ~n35724 ;
  assign n35895 = n77096 & n35894 ;
  assign n35896 = n35731 | n35895 ;
  assign n35898 = n35893 | n35896 ;
  assign n77097 = ~n35731 ;
  assign n35899 = n77097 & n35898 ;
  assign n77098 = ~n35721 ;
  assign n35900 = x78 & n77098 ;
  assign n77099 = ~n35716 ;
  assign n35901 = n77099 & n35900 ;
  assign n35902 = n35723 | n35901 ;
  assign n35903 = n35899 | n35902 ;
  assign n77100 = ~n35723 ;
  assign n35904 = n77100 & n35903 ;
  assign n77101 = ~n35713 ;
  assign n35905 = x79 & n77101 ;
  assign n77102 = ~n35708 ;
  assign n35906 = n77102 & n35905 ;
  assign n35907 = n35715 | n35906 ;
  assign n35909 = n35904 | n35907 ;
  assign n77103 = ~n35715 ;
  assign n35910 = n77103 & n35909 ;
  assign n77104 = ~n35705 ;
  assign n35911 = x80 & n77104 ;
  assign n77105 = ~n35700 ;
  assign n35912 = n77105 & n35911 ;
  assign n35913 = n35707 | n35912 ;
  assign n35914 = n35910 | n35913 ;
  assign n77106 = ~n35707 ;
  assign n35915 = n77106 & n35914 ;
  assign n77107 = ~n35697 ;
  assign n35916 = x81 & n77107 ;
  assign n77108 = ~n35692 ;
  assign n35917 = n77108 & n35916 ;
  assign n35918 = n35699 | n35917 ;
  assign n35920 = n35915 | n35918 ;
  assign n77109 = ~n35699 ;
  assign n35921 = n77109 & n35920 ;
  assign n77110 = ~n35680 ;
  assign n35922 = x82 & n77110 ;
  assign n77111 = ~n35637 ;
  assign n35923 = n77111 & n35922 ;
  assign n35924 = n35691 | n35923 ;
  assign n35925 = n35921 | n35924 ;
  assign n77112 = ~n35691 ;
  assign n35926 = n77112 & n35925 ;
  assign n77113 = ~n35634 ;
  assign n35927 = n77113 & n35687 ;
  assign n35928 = n35400 & n35634 ;
  assign n77114 = ~n35928 ;
  assign n35929 = x83 & n77114 ;
  assign n77115 = ~n35927 ;
  assign n35930 = n77115 & n35929 ;
  assign n35931 = n35690 | n35930 ;
  assign n35933 = n35926 | n35931 ;
  assign n77116 = ~n35690 ;
  assign n35934 = n77116 & n35933 ;
  assign n35935 = n65666 | n35934 ;
  assign n35936 = n35681 & n35935 ;
  assign n35938 = n65670 & n35830 ;
  assign n35825 = x65 & n35823 ;
  assign n77117 = ~n35825 ;
  assign n35937 = n77117 & n35833 ;
  assign n35939 = n3393 | n35937 ;
  assign n77118 = ~n35938 ;
  assign n35940 = n77118 & n35939 ;
  assign n35941 = n35839 | n35940 ;
  assign n35942 = n77064 & n35941 ;
  assign n35943 = n35813 | n35843 ;
  assign n35945 = n35942 | n35943 ;
  assign n35946 = n77067 & n35945 ;
  assign n35948 = n35848 | n35946 ;
  assign n35949 = n77070 & n35948 ;
  assign n35951 = n35853 | n35949 ;
  assign n35952 = n77073 & n35951 ;
  assign n35953 = n35858 | n35952 ;
  assign n35955 = n77076 & n35953 ;
  assign n35956 = n35863 | n35955 ;
  assign n35957 = n77079 & n35956 ;
  assign n35958 = n35869 | n35957 ;
  assign n35960 = n77082 & n35958 ;
  assign n35961 = n35874 | n35960 ;
  assign n35962 = n77085 & n35961 ;
  assign n35963 = n35880 | n35962 ;
  assign n35965 = n77088 & n35963 ;
  assign n35966 = n35885 | n35965 ;
  assign n35967 = n77091 & n35966 ;
  assign n35968 = n35891 | n35967 ;
  assign n35970 = n77094 & n35968 ;
  assign n35971 = n35896 | n35970 ;
  assign n35972 = n77097 & n35971 ;
  assign n35973 = n35902 | n35972 ;
  assign n35975 = n77100 & n35973 ;
  assign n35976 = n35907 | n35975 ;
  assign n35977 = n77103 & n35976 ;
  assign n35978 = n35913 | n35977 ;
  assign n35980 = n77106 & n35978 ;
  assign n35981 = n35918 | n35980 ;
  assign n35982 = n77109 & n35981 ;
  assign n77119 = ~n35982 ;
  assign n35983 = n35924 & n77119 ;
  assign n35985 = n35699 | n35924 ;
  assign n77120 = ~n35985 ;
  assign n35986 = n35920 & n77120 ;
  assign n35987 = n35983 | n35986 ;
  assign n35988 = n65674 & n35987 ;
  assign n77121 = ~n35934 ;
  assign n35989 = n77121 & n35988 ;
  assign n35990 = n35936 | n35989 ;
  assign n35991 = n66654 & n35990 ;
  assign n77122 = ~n35989 ;
  assign n36238 = x83 & n77122 ;
  assign n77123 = ~n35936 ;
  assign n36239 = n77123 & n36238 ;
  assign n36240 = n35991 | n36239 ;
  assign n35992 = n35698 & n35935 ;
  assign n77124 = ~n35915 ;
  assign n35919 = n77124 & n35918 ;
  assign n35993 = n35707 | n35918 ;
  assign n77125 = ~n35993 ;
  assign n35994 = n35978 & n77125 ;
  assign n35995 = n35919 | n35994 ;
  assign n35996 = n65674 & n35995 ;
  assign n35997 = n77121 & n35996 ;
  assign n35998 = n35992 | n35997 ;
  assign n35999 = n66560 & n35998 ;
  assign n36000 = n35706 & n35935 ;
  assign n77126 = ~n35977 ;
  assign n35979 = n35913 & n77126 ;
  assign n36001 = n35715 | n35913 ;
  assign n77127 = ~n36001 ;
  assign n36002 = n35909 & n77127 ;
  assign n36003 = n35979 | n36002 ;
  assign n36004 = n65674 & n36003 ;
  assign n36005 = n77121 & n36004 ;
  assign n36006 = n36000 | n36005 ;
  assign n36007 = n66505 & n36006 ;
  assign n77128 = ~n36005 ;
  assign n36228 = x81 & n77128 ;
  assign n77129 = ~n36000 ;
  assign n36229 = n77129 & n36228 ;
  assign n36230 = n36007 | n36229 ;
  assign n36008 = n35714 & n35935 ;
  assign n77130 = ~n35904 ;
  assign n35908 = n77130 & n35907 ;
  assign n36009 = n35723 | n35907 ;
  assign n77131 = ~n36009 ;
  assign n36010 = n35973 & n77131 ;
  assign n36011 = n35908 | n36010 ;
  assign n36012 = n65674 & n36011 ;
  assign n36013 = n77121 & n36012 ;
  assign n36014 = n36008 | n36013 ;
  assign n36015 = n66379 & n36014 ;
  assign n36016 = n35722 & n35935 ;
  assign n77132 = ~n35972 ;
  assign n35974 = n35902 & n77132 ;
  assign n36017 = n35731 | n35902 ;
  assign n77133 = ~n36017 ;
  assign n36018 = n35898 & n77133 ;
  assign n36019 = n35974 | n36018 ;
  assign n36020 = n65674 & n36019 ;
  assign n36021 = n77121 & n36020 ;
  assign n36022 = n36016 | n36021 ;
  assign n36023 = n66299 & n36022 ;
  assign n77134 = ~n36021 ;
  assign n36218 = x79 & n77134 ;
  assign n77135 = ~n36016 ;
  assign n36219 = n77135 & n36218 ;
  assign n36220 = n36023 | n36219 ;
  assign n36024 = n35730 & n35935 ;
  assign n77136 = ~n35893 ;
  assign n35897 = n77136 & n35896 ;
  assign n36025 = n35739 | n35896 ;
  assign n77137 = ~n36025 ;
  assign n36026 = n35968 & n77137 ;
  assign n36027 = n35897 | n36026 ;
  assign n36028 = n65674 & n36027 ;
  assign n36029 = n77121 & n36028 ;
  assign n36030 = n36024 | n36029 ;
  assign n36031 = n66244 & n36030 ;
  assign n36032 = n35738 & n35935 ;
  assign n77138 = ~n35967 ;
  assign n35969 = n35891 & n77138 ;
  assign n36033 = n35747 | n35891 ;
  assign n77139 = ~n36033 ;
  assign n36034 = n35887 & n77139 ;
  assign n36035 = n35969 | n36034 ;
  assign n36036 = n65674 & n36035 ;
  assign n36037 = n77121 & n36036 ;
  assign n36038 = n36032 | n36037 ;
  assign n36039 = n66145 & n36038 ;
  assign n77140 = ~n36037 ;
  assign n36207 = x77 & n77140 ;
  assign n77141 = ~n36032 ;
  assign n36208 = n77141 & n36207 ;
  assign n36209 = n36039 | n36208 ;
  assign n36040 = n35746 & n35935 ;
  assign n77142 = ~n35882 ;
  assign n35886 = n77142 & n35885 ;
  assign n36041 = n35755 | n35885 ;
  assign n77143 = ~n36041 ;
  assign n36042 = n35963 & n77143 ;
  assign n36043 = n35886 | n36042 ;
  assign n36044 = n65674 & n36043 ;
  assign n36045 = n77121 & n36044 ;
  assign n36046 = n36040 | n36045 ;
  assign n36047 = n66081 & n36046 ;
  assign n36048 = n35754 & n35935 ;
  assign n77144 = ~n35962 ;
  assign n35964 = n35880 & n77144 ;
  assign n36049 = n35763 | n35880 ;
  assign n77145 = ~n36049 ;
  assign n36050 = n35876 & n77145 ;
  assign n36051 = n35964 | n36050 ;
  assign n36052 = n65674 & n36051 ;
  assign n36053 = n77121 & n36052 ;
  assign n36054 = n36048 | n36053 ;
  assign n36055 = n66043 & n36054 ;
  assign n77146 = ~n36053 ;
  assign n36196 = x75 & n77146 ;
  assign n77147 = ~n36048 ;
  assign n36197 = n77147 & n36196 ;
  assign n36198 = n36055 | n36197 ;
  assign n36056 = n35762 & n35935 ;
  assign n77148 = ~n35871 ;
  assign n35875 = n77148 & n35874 ;
  assign n36057 = n35771 | n35874 ;
  assign n77149 = ~n36057 ;
  assign n36058 = n35958 & n77149 ;
  assign n36059 = n35875 | n36058 ;
  assign n36060 = n65674 & n36059 ;
  assign n36061 = n77121 & n36060 ;
  assign n36062 = n36056 | n36061 ;
  assign n36063 = n65960 & n36062 ;
  assign n36064 = n35770 & n35935 ;
  assign n77150 = ~n35957 ;
  assign n35959 = n35869 & n77150 ;
  assign n36065 = n35779 | n35869 ;
  assign n77151 = ~n36065 ;
  assign n36066 = n35865 & n77151 ;
  assign n36067 = n35959 | n36066 ;
  assign n36068 = n65674 & n36067 ;
  assign n36069 = n77121 & n36068 ;
  assign n36070 = n36064 | n36069 ;
  assign n36071 = n65909 & n36070 ;
  assign n77152 = ~n36069 ;
  assign n36186 = x73 & n77152 ;
  assign n77153 = ~n36064 ;
  assign n36187 = n77153 & n36186 ;
  assign n36188 = n36071 | n36187 ;
  assign n36072 = n35778 & n35935 ;
  assign n77154 = ~n35860 ;
  assign n35864 = n77154 & n35863 ;
  assign n36073 = n35787 | n35863 ;
  assign n77155 = ~n36073 ;
  assign n36074 = n35953 & n77155 ;
  assign n36075 = n35864 | n36074 ;
  assign n36076 = n65674 & n36075 ;
  assign n36077 = n77121 & n36076 ;
  assign n36078 = n36072 | n36077 ;
  assign n36079 = n65877 & n36078 ;
  assign n36080 = n35786 & n35935 ;
  assign n77156 = ~n35952 ;
  assign n35954 = n35858 & n77156 ;
  assign n36081 = n35796 | n35858 ;
  assign n77157 = ~n36081 ;
  assign n36082 = n35854 & n77157 ;
  assign n36083 = n35954 | n36082 ;
  assign n36084 = n65674 & n36083 ;
  assign n36085 = n77121 & n36084 ;
  assign n36086 = n36080 | n36085 ;
  assign n36087 = n65820 & n36086 ;
  assign n77158 = ~n36085 ;
  assign n36176 = x71 & n77158 ;
  assign n77159 = ~n36080 ;
  assign n36177 = n77159 & n36176 ;
  assign n36178 = n36087 | n36177 ;
  assign n36088 = n35795 & n35935 ;
  assign n77160 = ~n35850 ;
  assign n35950 = n77160 & n35853 ;
  assign n36089 = n35805 | n35853 ;
  assign n77161 = ~n36089 ;
  assign n36090 = n35849 & n77161 ;
  assign n36091 = n35950 | n36090 ;
  assign n36092 = n65674 & n36091 ;
  assign n36093 = n77121 & n36092 ;
  assign n36094 = n36088 | n36093 ;
  assign n36095 = n65791 & n36094 ;
  assign n36096 = n35804 & n35935 ;
  assign n77162 = ~n35946 ;
  assign n35947 = n35848 & n77162 ;
  assign n36097 = n35841 | n35943 ;
  assign n36098 = n35813 | n35848 ;
  assign n77163 = ~n36098 ;
  assign n36099 = n36097 & n77163 ;
  assign n36100 = n35947 | n36099 ;
  assign n36101 = n65674 & n36100 ;
  assign n36102 = n77121 & n36101 ;
  assign n36103 = n36096 | n36102 ;
  assign n36104 = n65772 & n36103 ;
  assign n77164 = ~n36102 ;
  assign n36165 = x69 & n77164 ;
  assign n77165 = ~n36096 ;
  assign n36166 = n77165 & n36165 ;
  assign n36167 = n36104 | n36166 ;
  assign n36105 = n35812 & n35935 ;
  assign n77166 = ~n35841 ;
  assign n35944 = n77166 & n35943 ;
  assign n36106 = n35820 | n35943 ;
  assign n77167 = ~n36106 ;
  assign n36107 = n35840 & n77167 ;
  assign n36108 = n35944 | n36107 ;
  assign n36109 = n65674 & n36108 ;
  assign n36110 = n77121 & n36109 ;
  assign n36111 = n36105 | n36110 ;
  assign n36112 = n65746 & n36111 ;
  assign n36113 = n35819 & n35935 ;
  assign n36114 = n35839 | n35938 ;
  assign n77168 = ~n36114 ;
  assign n36115 = n35939 & n77168 ;
  assign n77169 = ~n35940 ;
  assign n36116 = n35839 & n77169 ;
  assign n36117 = n36115 | n36116 ;
  assign n36118 = n65674 & n36117 ;
  assign n36119 = n77121 & n36118 ;
  assign n36120 = n36113 | n36119 ;
  assign n36122 = n65721 & n36120 ;
  assign n77170 = ~n36119 ;
  assign n36121 = x67 & n77170 ;
  assign n77171 = ~n36113 ;
  assign n36156 = n77171 & n36121 ;
  assign n36157 = n36122 | n36156 ;
  assign n36123 = n35823 & n35935 ;
  assign n36124 = n3393 & n35833 ;
  assign n36125 = n77060 & n36124 ;
  assign n36126 = n65666 | n36125 ;
  assign n77172 = ~n36126 ;
  assign n36127 = n35939 & n77172 ;
  assign n36128 = n77121 & n36127 ;
  assign n36129 = n36123 | n36128 ;
  assign n36130 = n65686 & n36129 ;
  assign n36131 = n3694 & n77121 ;
  assign n77173 = ~n36131 ;
  assign n36132 = x44 & n77173 ;
  assign n36133 = n3706 & n77121 ;
  assign n36134 = n36132 | n36133 ;
  assign n36135 = x65 & n36134 ;
  assign n35984 = n35924 | n35982 ;
  assign n36136 = n77112 & n35984 ;
  assign n36137 = n35931 | n36136 ;
  assign n36138 = n77116 & n36137 ;
  assign n77174 = ~n36138 ;
  assign n36139 = n3694 & n77174 ;
  assign n77175 = ~n36139 ;
  assign n36141 = x44 & n77175 ;
  assign n36142 = x65 | n36133 ;
  assign n36143 = n36141 | n36142 ;
  assign n77176 = ~n36135 ;
  assign n36144 = n77176 & n36143 ;
  assign n36145 = n3713 | n36144 ;
  assign n36146 = n36133 | n36141 ;
  assign n36147 = n65670 & n36146 ;
  assign n77177 = ~n36147 ;
  assign n36148 = n36145 & n77177 ;
  assign n36140 = n65666 | n36138 ;
  assign n36149 = n35830 & n36140 ;
  assign n36150 = n36128 | n36149 ;
  assign n36151 = n65686 & n36150 ;
  assign n77178 = ~n36128 ;
  assign n36152 = x66 & n77178 ;
  assign n77179 = ~n36149 ;
  assign n36153 = n77179 & n36152 ;
  assign n36154 = n36151 | n36153 ;
  assign n36155 = n36148 | n36154 ;
  assign n77180 = ~n36130 ;
  assign n36158 = n77180 & n36155 ;
  assign n36159 = n36157 | n36158 ;
  assign n77181 = ~n36122 ;
  assign n36160 = n77181 & n36159 ;
  assign n77182 = ~n36110 ;
  assign n36161 = x68 & n77182 ;
  assign n77183 = ~n36105 ;
  assign n36162 = n77183 & n36161 ;
  assign n36163 = n36112 | n36162 ;
  assign n36164 = n36160 | n36163 ;
  assign n77184 = ~n36112 ;
  assign n36168 = n77184 & n36164 ;
  assign n36169 = n36167 | n36168 ;
  assign n77185 = ~n36104 ;
  assign n36170 = n77185 & n36169 ;
  assign n77186 = ~n36093 ;
  assign n36171 = x70 & n77186 ;
  assign n77187 = ~n36088 ;
  assign n36172 = n77187 & n36171 ;
  assign n36173 = n36095 | n36172 ;
  assign n36175 = n36170 | n36173 ;
  assign n77188 = ~n36095 ;
  assign n36179 = n77188 & n36175 ;
  assign n36180 = n36178 | n36179 ;
  assign n77189 = ~n36087 ;
  assign n36181 = n77189 & n36180 ;
  assign n77190 = ~n36077 ;
  assign n36182 = x72 & n77190 ;
  assign n77191 = ~n36072 ;
  assign n36183 = n77191 & n36182 ;
  assign n36184 = n36079 | n36183 ;
  assign n36185 = n36181 | n36184 ;
  assign n77192 = ~n36079 ;
  assign n36189 = n77192 & n36185 ;
  assign n36190 = n36188 | n36189 ;
  assign n77193 = ~n36071 ;
  assign n36191 = n77193 & n36190 ;
  assign n77194 = ~n36061 ;
  assign n36192 = x74 & n77194 ;
  assign n77195 = ~n36056 ;
  assign n36193 = n77195 & n36192 ;
  assign n36194 = n36063 | n36193 ;
  assign n36195 = n36191 | n36194 ;
  assign n77196 = ~n36063 ;
  assign n36199 = n77196 & n36195 ;
  assign n36200 = n36198 | n36199 ;
  assign n77197 = ~n36055 ;
  assign n36201 = n77197 & n36200 ;
  assign n77198 = ~n36045 ;
  assign n36202 = x76 & n77198 ;
  assign n77199 = ~n36040 ;
  assign n36203 = n77199 & n36202 ;
  assign n36204 = n36047 | n36203 ;
  assign n36206 = n36201 | n36204 ;
  assign n77200 = ~n36047 ;
  assign n36211 = n77200 & n36206 ;
  assign n36212 = n36209 | n36211 ;
  assign n77201 = ~n36039 ;
  assign n36213 = n77201 & n36212 ;
  assign n77202 = ~n36029 ;
  assign n36214 = x78 & n77202 ;
  assign n77203 = ~n36024 ;
  assign n36215 = n77203 & n36214 ;
  assign n36216 = n36031 | n36215 ;
  assign n36217 = n36213 | n36216 ;
  assign n77204 = ~n36031 ;
  assign n36221 = n77204 & n36217 ;
  assign n36222 = n36220 | n36221 ;
  assign n77205 = ~n36023 ;
  assign n36223 = n77205 & n36222 ;
  assign n77206 = ~n36013 ;
  assign n36224 = x80 & n77206 ;
  assign n77207 = ~n36008 ;
  assign n36225 = n77207 & n36224 ;
  assign n36226 = n36015 | n36225 ;
  assign n36227 = n36223 | n36226 ;
  assign n77208 = ~n36015 ;
  assign n36231 = n77208 & n36227 ;
  assign n36232 = n36230 | n36231 ;
  assign n77209 = ~n36007 ;
  assign n36233 = n77209 & n36232 ;
  assign n77210 = ~n35997 ;
  assign n36234 = x82 & n77210 ;
  assign n77211 = ~n35992 ;
  assign n36235 = n77211 & n36234 ;
  assign n36236 = n35999 | n36235 ;
  assign n36237 = n36233 | n36236 ;
  assign n77212 = ~n35999 ;
  assign n36241 = n77212 & n36237 ;
  assign n36242 = n36240 | n36241 ;
  assign n77213 = ~n35991 ;
  assign n36243 = n77213 & n36242 ;
  assign n77214 = ~n35926 ;
  assign n35932 = n77214 & n35931 ;
  assign n36244 = n35691 | n35931 ;
  assign n77215 = ~n36244 ;
  assign n36245 = n35984 & n77215 ;
  assign n36246 = n35932 | n36245 ;
  assign n36247 = n35935 | n36246 ;
  assign n77216 = ~n35689 ;
  assign n36248 = n77216 & n35935 ;
  assign n77217 = ~n36248 ;
  assign n36249 = n36247 & n77217 ;
  assign n36250 = n66797 & n36249 ;
  assign n77218 = ~n35935 ;
  assign n36251 = n77218 & n36246 ;
  assign n36252 = n35689 & n35935 ;
  assign n77219 = ~n36252 ;
  assign n36253 = x84 & n77219 ;
  assign n77220 = ~n36251 ;
  assign n36254 = n77220 & n36253 ;
  assign n36255 = n513 | n36254 ;
  assign n36256 = n36250 | n36255 ;
  assign n36257 = n36243 | n36256 ;
  assign n36258 = n65674 & n36249 ;
  assign n77221 = ~n36258 ;
  assign n36259 = n36257 & n77221 ;
  assign n36309 = n35991 | n36254 ;
  assign n36310 = n36250 | n36309 ;
  assign n77222 = ~n36310 ;
  assign n36311 = n36242 & n77222 ;
  assign n77223 = ~n36123 ;
  assign n36264 = n77223 & n36152 ;
  assign n36265 = n36130 | n36264 ;
  assign n36261 = x65 & n36146 ;
  assign n77224 = ~n36261 ;
  assign n36262 = n36143 & n77224 ;
  assign n36263 = n3713 | n36262 ;
  assign n36266 = n77177 & n36263 ;
  assign n36267 = n36265 | n36266 ;
  assign n77225 = ~n36151 ;
  assign n36268 = n77225 & n36267 ;
  assign n36269 = n36157 | n36268 ;
  assign n36270 = n77181 & n36269 ;
  assign n36271 = n36163 | n36270 ;
  assign n36272 = n77184 & n36271 ;
  assign n36273 = n36167 | n36272 ;
  assign n36274 = n77185 & n36273 ;
  assign n36275 = n36173 | n36274 ;
  assign n36276 = n77188 & n36275 ;
  assign n36277 = n36178 | n36276 ;
  assign n36278 = n77189 & n36277 ;
  assign n36279 = n36184 | n36278 ;
  assign n36280 = n77192 & n36279 ;
  assign n36281 = n36188 | n36280 ;
  assign n36282 = n77193 & n36281 ;
  assign n36283 = n36194 | n36282 ;
  assign n36284 = n77196 & n36283 ;
  assign n36285 = n36198 | n36284 ;
  assign n36286 = n77197 & n36285 ;
  assign n36287 = n36204 | n36286 ;
  assign n36288 = n77200 & n36287 ;
  assign n36289 = n36209 | n36288 ;
  assign n36290 = n77201 & n36289 ;
  assign n36291 = n36216 | n36290 ;
  assign n36292 = n77204 & n36291 ;
  assign n36293 = n36220 | n36292 ;
  assign n36294 = n77205 & n36293 ;
  assign n36295 = n36226 | n36294 ;
  assign n36296 = n77208 & n36295 ;
  assign n36297 = n36230 | n36296 ;
  assign n36298 = n77209 & n36297 ;
  assign n36299 = n36236 | n36298 ;
  assign n36300 = n77212 & n36299 ;
  assign n36312 = n36240 | n36300 ;
  assign n36313 = n77213 & n36312 ;
  assign n36314 = n36250 | n36254 ;
  assign n77226 = ~n36313 ;
  assign n36315 = n77226 & n36314 ;
  assign n36316 = n36311 | n36315 ;
  assign n77227 = ~n36259 ;
  assign n36317 = n77227 & n36316 ;
  assign n36318 = n65666 & n35689 ;
  assign n36319 = n36257 & n36318 ;
  assign n36320 = n36317 | n36319 ;
  assign n36321 = n66868 & n36320 ;
  assign n77228 = ~n36241 ;
  assign n36301 = n36240 & n77228 ;
  assign n36302 = n35999 | n36240 ;
  assign n77229 = ~n36302 ;
  assign n36303 = n36299 & n77229 ;
  assign n36304 = n36301 | n36303 ;
  assign n36305 = n77227 & n36304 ;
  assign n36306 = n35990 & n77221 ;
  assign n36307 = n36257 & n36306 ;
  assign n36308 = n36305 | n36307 ;
  assign n36322 = n66797 & n36308 ;
  assign n77230 = ~n36298 ;
  assign n36323 = n36236 & n77230 ;
  assign n36324 = n36007 | n36236 ;
  assign n77231 = ~n36324 ;
  assign n36325 = n36232 & n77231 ;
  assign n36326 = n36323 | n36325 ;
  assign n36327 = n77227 & n36326 ;
  assign n36328 = n35998 & n77221 ;
  assign n36329 = n36257 & n36328 ;
  assign n36330 = n36327 | n36329 ;
  assign n36331 = n66654 & n36330 ;
  assign n77232 = ~n36231 ;
  assign n36332 = n36230 & n77232 ;
  assign n36333 = n36015 | n36230 ;
  assign n77233 = ~n36333 ;
  assign n36334 = n36295 & n77233 ;
  assign n36335 = n36332 | n36334 ;
  assign n36336 = n77227 & n36335 ;
  assign n36337 = n36006 & n77221 ;
  assign n36338 = n36257 & n36337 ;
  assign n36339 = n36336 | n36338 ;
  assign n36340 = n66560 & n36339 ;
  assign n77234 = ~n36294 ;
  assign n36341 = n36226 & n77234 ;
  assign n36342 = n36023 | n36226 ;
  assign n77235 = ~n36342 ;
  assign n36343 = n36222 & n77235 ;
  assign n36344 = n36341 | n36343 ;
  assign n36345 = n77227 & n36344 ;
  assign n36346 = n36014 & n77221 ;
  assign n36347 = n36257 & n36346 ;
  assign n36348 = n36345 | n36347 ;
  assign n36349 = n66505 & n36348 ;
  assign n77236 = ~n36221 ;
  assign n36350 = n36220 & n77236 ;
  assign n36351 = n36031 | n36220 ;
  assign n77237 = ~n36351 ;
  assign n36352 = n36291 & n77237 ;
  assign n36353 = n36350 | n36352 ;
  assign n36354 = n77227 & n36353 ;
  assign n36355 = n36022 & n77221 ;
  assign n36356 = n36257 & n36355 ;
  assign n36357 = n36354 | n36356 ;
  assign n36358 = n66379 & n36357 ;
  assign n77238 = ~n36290 ;
  assign n36359 = n36216 & n77238 ;
  assign n36360 = n36039 | n36216 ;
  assign n77239 = ~n36360 ;
  assign n36361 = n36212 & n77239 ;
  assign n36362 = n36359 | n36361 ;
  assign n36363 = n77227 & n36362 ;
  assign n36364 = n36030 & n77221 ;
  assign n36365 = n36257 & n36364 ;
  assign n36366 = n36363 | n36365 ;
  assign n36367 = n66299 & n36366 ;
  assign n77240 = ~n36211 ;
  assign n36368 = n36209 & n77240 ;
  assign n36210 = n36047 | n36209 ;
  assign n77241 = ~n36210 ;
  assign n36369 = n36206 & n77241 ;
  assign n36370 = n36368 | n36369 ;
  assign n36371 = n77227 & n36370 ;
  assign n36372 = n36038 & n77221 ;
  assign n36373 = n36257 & n36372 ;
  assign n36374 = n36371 | n36373 ;
  assign n36375 = n66244 & n36374 ;
  assign n77242 = ~n36286 ;
  assign n36376 = n36204 & n77242 ;
  assign n36205 = n36055 | n36204 ;
  assign n77243 = ~n36205 ;
  assign n36377 = n77243 & n36285 ;
  assign n36378 = n36376 | n36377 ;
  assign n36379 = n77227 & n36378 ;
  assign n36380 = n36046 & n77221 ;
  assign n36381 = n36257 & n36380 ;
  assign n36382 = n36379 | n36381 ;
  assign n36383 = n66145 & n36382 ;
  assign n77244 = ~n36199 ;
  assign n36384 = n36198 & n77244 ;
  assign n36385 = n36063 | n36198 ;
  assign n77245 = ~n36385 ;
  assign n36386 = n36283 & n77245 ;
  assign n36387 = n36384 | n36386 ;
  assign n36388 = n77227 & n36387 ;
  assign n36389 = n36054 & n77221 ;
  assign n36390 = n36257 & n36389 ;
  assign n36391 = n36388 | n36390 ;
  assign n36392 = n66081 & n36391 ;
  assign n77246 = ~n36282 ;
  assign n36393 = n36194 & n77246 ;
  assign n36394 = n36071 | n36194 ;
  assign n77247 = ~n36394 ;
  assign n36395 = n36190 & n77247 ;
  assign n36396 = n36393 | n36395 ;
  assign n36397 = n77227 & n36396 ;
  assign n36398 = n36062 & n77221 ;
  assign n36399 = n36257 & n36398 ;
  assign n36400 = n36397 | n36399 ;
  assign n36401 = n66043 & n36400 ;
  assign n77248 = ~n36189 ;
  assign n36402 = n36188 & n77248 ;
  assign n36403 = n36079 | n36188 ;
  assign n77249 = ~n36403 ;
  assign n36404 = n36279 & n77249 ;
  assign n36405 = n36402 | n36404 ;
  assign n36406 = n77227 & n36405 ;
  assign n36407 = n36070 & n77221 ;
  assign n36408 = n36257 & n36407 ;
  assign n36409 = n36406 | n36408 ;
  assign n36410 = n65960 & n36409 ;
  assign n77250 = ~n36278 ;
  assign n36411 = n36184 & n77250 ;
  assign n36412 = n36087 | n36184 ;
  assign n77251 = ~n36412 ;
  assign n36413 = n36180 & n77251 ;
  assign n36414 = n36411 | n36413 ;
  assign n36415 = n77227 & n36414 ;
  assign n36416 = n36078 & n77221 ;
  assign n36417 = n36257 & n36416 ;
  assign n36418 = n36415 | n36417 ;
  assign n36419 = n65909 & n36418 ;
  assign n77252 = ~n36179 ;
  assign n36420 = n36178 & n77252 ;
  assign n36421 = n36095 | n36178 ;
  assign n77253 = ~n36421 ;
  assign n36422 = n36275 & n77253 ;
  assign n36423 = n36420 | n36422 ;
  assign n36424 = n77227 & n36423 ;
  assign n36425 = n36086 & n77221 ;
  assign n36426 = n36257 & n36425 ;
  assign n36427 = n36424 | n36426 ;
  assign n36428 = n65877 & n36427 ;
  assign n77254 = ~n36274 ;
  assign n36429 = n36173 & n77254 ;
  assign n36174 = n36104 | n36173 ;
  assign n77255 = ~n36174 ;
  assign n36430 = n77255 & n36273 ;
  assign n36431 = n36429 | n36430 ;
  assign n36432 = n77227 & n36431 ;
  assign n36433 = n36094 & n77221 ;
  assign n36434 = n36257 & n36433 ;
  assign n36435 = n36432 | n36434 ;
  assign n36436 = n65820 & n36435 ;
  assign n77256 = ~n36168 ;
  assign n36437 = n36167 & n77256 ;
  assign n36438 = n36112 | n36167 ;
  assign n77257 = ~n36438 ;
  assign n36439 = n36271 & n77257 ;
  assign n36440 = n36437 | n36439 ;
  assign n36441 = n77227 & n36440 ;
  assign n36442 = n36103 & n77221 ;
  assign n36443 = n36257 & n36442 ;
  assign n36444 = n36441 | n36443 ;
  assign n36445 = n65791 & n36444 ;
  assign n77258 = ~n36270 ;
  assign n36446 = n36163 & n77258 ;
  assign n36447 = n36122 | n36163 ;
  assign n77259 = ~n36447 ;
  assign n36448 = n36159 & n77259 ;
  assign n36449 = n36446 | n36448 ;
  assign n36450 = n77227 & n36449 ;
  assign n36451 = n36111 & n77221 ;
  assign n36452 = n36257 & n36451 ;
  assign n36453 = n36450 | n36452 ;
  assign n36454 = n65772 & n36453 ;
  assign n36455 = n77225 & n36155 ;
  assign n77260 = ~n36455 ;
  assign n36457 = n36157 & n77260 ;
  assign n36456 = n36151 | n36157 ;
  assign n77261 = ~n36456 ;
  assign n36458 = n36155 & n77261 ;
  assign n36459 = n36457 | n36458 ;
  assign n36460 = n77227 & n36459 ;
  assign n36461 = n36120 & n77221 ;
  assign n36462 = n36257 & n36461 ;
  assign n36463 = n36460 | n36462 ;
  assign n36464 = n65746 & n36463 ;
  assign n77262 = ~n36266 ;
  assign n36466 = n36265 & n77262 ;
  assign n36465 = n36147 | n36154 ;
  assign n77263 = ~n36465 ;
  assign n36467 = n36263 & n77263 ;
  assign n36468 = n36466 | n36467 ;
  assign n36469 = n77227 & n36468 ;
  assign n36470 = n36150 & n77221 ;
  assign n36471 = n36257 & n36470 ;
  assign n36472 = n36469 | n36471 ;
  assign n36473 = n65721 & n36472 ;
  assign n36474 = n3713 & n36143 ;
  assign n36475 = n77224 & n36474 ;
  assign n77264 = ~n36475 ;
  assign n36476 = n36263 & n77264 ;
  assign n36477 = n77227 & n36476 ;
  assign n36478 = n36146 & n77221 ;
  assign n36479 = n36257 & n36478 ;
  assign n36480 = n36477 | n36479 ;
  assign n36481 = n65686 & n36480 ;
  assign n36260 = n3713 & n77227 ;
  assign n36486 = x64 & n77227 ;
  assign n77265 = ~n36486 ;
  assign n36487 = x43 & n77265 ;
  assign n36488 = n36260 | n36487 ;
  assign n36490 = x65 & n36488 ;
  assign n36482 = n36256 | n36313 ;
  assign n36483 = n77221 & n36482 ;
  assign n77266 = ~n36483 ;
  assign n36484 = x64 & n77266 ;
  assign n77267 = ~n36484 ;
  assign n36485 = x43 & n77267 ;
  assign n36489 = x65 | n36260 ;
  assign n36491 = n36485 | n36489 ;
  assign n77268 = ~n36490 ;
  assign n36492 = n77268 & n36491 ;
  assign n36493 = n4058 | n36492 ;
  assign n36494 = n65670 & n36488 ;
  assign n77269 = ~n36494 ;
  assign n36495 = n36493 & n77269 ;
  assign n77270 = ~n36479 ;
  assign n36496 = x66 & n77270 ;
  assign n77271 = ~n36477 ;
  assign n36497 = n77271 & n36496 ;
  assign n36498 = n36481 | n36497 ;
  assign n36499 = n36495 | n36498 ;
  assign n77272 = ~n36481 ;
  assign n36500 = n77272 & n36499 ;
  assign n77273 = ~n36471 ;
  assign n36501 = x67 & n77273 ;
  assign n77274 = ~n36469 ;
  assign n36502 = n77274 & n36501 ;
  assign n36503 = n36500 | n36502 ;
  assign n77275 = ~n36473 ;
  assign n36504 = n77275 & n36503 ;
  assign n77276 = ~n36462 ;
  assign n36505 = x68 & n77276 ;
  assign n77277 = ~n36460 ;
  assign n36506 = n77277 & n36505 ;
  assign n36507 = n36464 | n36506 ;
  assign n36508 = n36504 | n36507 ;
  assign n77278 = ~n36464 ;
  assign n36509 = n77278 & n36508 ;
  assign n77279 = ~n36452 ;
  assign n36510 = x69 & n77279 ;
  assign n77280 = ~n36450 ;
  assign n36511 = n77280 & n36510 ;
  assign n36512 = n36509 | n36511 ;
  assign n77281 = ~n36454 ;
  assign n36513 = n77281 & n36512 ;
  assign n77282 = ~n36443 ;
  assign n36514 = x70 & n77282 ;
  assign n77283 = ~n36441 ;
  assign n36515 = n77283 & n36514 ;
  assign n36516 = n36445 | n36515 ;
  assign n36517 = n36513 | n36516 ;
  assign n77284 = ~n36445 ;
  assign n36518 = n77284 & n36517 ;
  assign n77285 = ~n36434 ;
  assign n36519 = x71 & n77285 ;
  assign n77286 = ~n36432 ;
  assign n36520 = n77286 & n36519 ;
  assign n36521 = n36436 | n36520 ;
  assign n36524 = n36518 | n36521 ;
  assign n77287 = ~n36436 ;
  assign n36525 = n77287 & n36524 ;
  assign n77288 = ~n36426 ;
  assign n36526 = x72 & n77288 ;
  assign n77289 = ~n36424 ;
  assign n36527 = n77289 & n36526 ;
  assign n36528 = n36428 | n36527 ;
  assign n36529 = n36525 | n36528 ;
  assign n77290 = ~n36428 ;
  assign n36530 = n77290 & n36529 ;
  assign n77291 = ~n36417 ;
  assign n36531 = x73 & n77291 ;
  assign n77292 = ~n36415 ;
  assign n36532 = n77292 & n36531 ;
  assign n36533 = n36419 | n36532 ;
  assign n36535 = n36530 | n36533 ;
  assign n77293 = ~n36419 ;
  assign n36536 = n77293 & n36535 ;
  assign n77294 = ~n36408 ;
  assign n36537 = x74 & n77294 ;
  assign n77295 = ~n36406 ;
  assign n36538 = n77295 & n36537 ;
  assign n36539 = n36410 | n36538 ;
  assign n36540 = n36536 | n36539 ;
  assign n77296 = ~n36410 ;
  assign n36541 = n77296 & n36540 ;
  assign n77297 = ~n36399 ;
  assign n36542 = x75 & n77297 ;
  assign n77298 = ~n36397 ;
  assign n36543 = n77298 & n36542 ;
  assign n36544 = n36401 | n36543 ;
  assign n36546 = n36541 | n36544 ;
  assign n77299 = ~n36401 ;
  assign n36547 = n77299 & n36546 ;
  assign n77300 = ~n36390 ;
  assign n36548 = x76 & n77300 ;
  assign n77301 = ~n36388 ;
  assign n36549 = n77301 & n36548 ;
  assign n36550 = n36392 | n36549 ;
  assign n36551 = n36547 | n36550 ;
  assign n77302 = ~n36392 ;
  assign n36552 = n77302 & n36551 ;
  assign n77303 = ~n36381 ;
  assign n36553 = x77 & n77303 ;
  assign n77304 = ~n36379 ;
  assign n36554 = n77304 & n36553 ;
  assign n36555 = n36383 | n36554 ;
  assign n36557 = n36552 | n36555 ;
  assign n77305 = ~n36383 ;
  assign n36558 = n77305 & n36557 ;
  assign n77306 = ~n36373 ;
  assign n36559 = x78 & n77306 ;
  assign n77307 = ~n36371 ;
  assign n36560 = n77307 & n36559 ;
  assign n36561 = n36375 | n36560 ;
  assign n36562 = n36558 | n36561 ;
  assign n77308 = ~n36375 ;
  assign n36563 = n77308 & n36562 ;
  assign n77309 = ~n36365 ;
  assign n36564 = x79 & n77309 ;
  assign n77310 = ~n36363 ;
  assign n36565 = n77310 & n36564 ;
  assign n36566 = n36367 | n36565 ;
  assign n36568 = n36563 | n36566 ;
  assign n77311 = ~n36367 ;
  assign n36569 = n77311 & n36568 ;
  assign n77312 = ~n36356 ;
  assign n36570 = x80 & n77312 ;
  assign n77313 = ~n36354 ;
  assign n36571 = n77313 & n36570 ;
  assign n36572 = n36358 | n36571 ;
  assign n36573 = n36569 | n36572 ;
  assign n77314 = ~n36358 ;
  assign n36574 = n77314 & n36573 ;
  assign n77315 = ~n36347 ;
  assign n36575 = x81 & n77315 ;
  assign n77316 = ~n36345 ;
  assign n36576 = n77316 & n36575 ;
  assign n36577 = n36349 | n36576 ;
  assign n36579 = n36574 | n36577 ;
  assign n77317 = ~n36349 ;
  assign n36580 = n77317 & n36579 ;
  assign n77318 = ~n36338 ;
  assign n36581 = x82 & n77318 ;
  assign n77319 = ~n36336 ;
  assign n36582 = n77319 & n36581 ;
  assign n36583 = n36340 | n36582 ;
  assign n36584 = n36580 | n36583 ;
  assign n77320 = ~n36340 ;
  assign n36585 = n77320 & n36584 ;
  assign n77321 = ~n36329 ;
  assign n36586 = x83 & n77321 ;
  assign n77322 = ~n36327 ;
  assign n36587 = n77322 & n36586 ;
  assign n36588 = n36331 | n36587 ;
  assign n36590 = n36585 | n36588 ;
  assign n77323 = ~n36331 ;
  assign n36591 = n77323 & n36590 ;
  assign n77324 = ~n36307 ;
  assign n36592 = x84 & n77324 ;
  assign n77325 = ~n36305 ;
  assign n36593 = n77325 & n36592 ;
  assign n36594 = n36322 | n36593 ;
  assign n36595 = n36591 | n36594 ;
  assign n77326 = ~n36322 ;
  assign n36596 = n77326 & n36595 ;
  assign n77327 = ~n36319 ;
  assign n36597 = x85 & n77327 ;
  assign n77328 = ~n36317 ;
  assign n36598 = n77328 & n36597 ;
  assign n36599 = n36321 | n36598 ;
  assign n36601 = n36596 | n36599 ;
  assign n77329 = ~n36321 ;
  assign n36602 = n77329 & n36601 ;
  assign n36603 = n4182 | n36602 ;
  assign n77330 = ~n36320 ;
  assign n36604 = n77330 & n36603 ;
  assign n77331 = ~n36596 ;
  assign n36600 = n77331 & n36599 ;
  assign n36611 = n36260 | n36485 ;
  assign n36612 = x65 & n36611 ;
  assign n77332 = ~n36612 ;
  assign n36613 = n36491 & n77332 ;
  assign n36614 = n4058 | n36613 ;
  assign n36615 = n77269 & n36614 ;
  assign n36616 = n36498 | n36615 ;
  assign n36617 = n77272 & n36616 ;
  assign n36618 = n36473 | n36502 ;
  assign n36620 = n36617 | n36618 ;
  assign n36621 = n77275 & n36620 ;
  assign n36622 = n36506 | n36621 ;
  assign n36624 = n77278 & n36622 ;
  assign n36625 = n36454 | n36511 ;
  assign n36627 = n36624 | n36625 ;
  assign n36628 = n77281 & n36627 ;
  assign n36629 = n36515 | n36628 ;
  assign n36631 = n77284 & n36629 ;
  assign n36632 = n36521 | n36631 ;
  assign n36633 = n77287 & n36632 ;
  assign n36634 = n36528 | n36633 ;
  assign n36636 = n77290 & n36634 ;
  assign n36637 = n36533 | n36636 ;
  assign n36638 = n77293 & n36637 ;
  assign n36639 = n36539 | n36638 ;
  assign n36641 = n77296 & n36639 ;
  assign n36642 = n36544 | n36641 ;
  assign n36643 = n77299 & n36642 ;
  assign n36644 = n36550 | n36643 ;
  assign n36646 = n77302 & n36644 ;
  assign n36647 = n36555 | n36646 ;
  assign n36648 = n77305 & n36647 ;
  assign n36649 = n36561 | n36648 ;
  assign n36651 = n77308 & n36649 ;
  assign n36652 = n36566 | n36651 ;
  assign n36653 = n77311 & n36652 ;
  assign n36654 = n36572 | n36653 ;
  assign n36656 = n77314 & n36654 ;
  assign n36657 = n36577 | n36656 ;
  assign n36658 = n77317 & n36657 ;
  assign n36659 = n36583 | n36658 ;
  assign n36661 = n77320 & n36659 ;
  assign n36662 = n36588 | n36661 ;
  assign n36663 = n77323 & n36662 ;
  assign n36665 = n36594 | n36663 ;
  assign n36672 = n36322 | n36599 ;
  assign n77333 = ~n36672 ;
  assign n36673 = n36665 & n77333 ;
  assign n36674 = n36600 | n36673 ;
  assign n36675 = n36603 | n36674 ;
  assign n77334 = ~n36604 ;
  assign n36676 = n77334 & n36675 ;
  assign n36677 = n66979 & n36676 ;
  assign n77335 = ~n36603 ;
  assign n36960 = n77335 & n36674 ;
  assign n36961 = n36320 & n36603 ;
  assign n77336 = ~n36961 ;
  assign n36962 = x86 & n77336 ;
  assign n77337 = ~n36960 ;
  assign n36963 = n77337 & n36962 ;
  assign n36964 = n36677 | n36963 ;
  assign n36609 = n36308 & n36603 ;
  assign n77338 = ~n36663 ;
  assign n36664 = n36594 & n77338 ;
  assign n36666 = n36331 | n36594 ;
  assign n77339 = ~n36666 ;
  assign n36667 = n36590 & n77339 ;
  assign n36668 = n36664 | n36667 ;
  assign n36669 = n66973 & n36668 ;
  assign n77340 = ~n36602 ;
  assign n36670 = n77340 & n36669 ;
  assign n36671 = n36609 | n36670 ;
  assign n36678 = n66868 & n36671 ;
  assign n36679 = n36330 & n36603 ;
  assign n77341 = ~n36585 ;
  assign n36589 = n77341 & n36588 ;
  assign n36680 = n36340 | n36588 ;
  assign n77342 = ~n36680 ;
  assign n36681 = n36659 & n77342 ;
  assign n36682 = n36589 | n36681 ;
  assign n36683 = n66973 & n36682 ;
  assign n36684 = n77340 & n36683 ;
  assign n36685 = n36679 | n36684 ;
  assign n36686 = n66797 & n36685 ;
  assign n77343 = ~n36684 ;
  assign n36948 = x84 & n77343 ;
  assign n77344 = ~n36679 ;
  assign n36949 = n77344 & n36948 ;
  assign n36950 = n36686 | n36949 ;
  assign n36687 = n36339 & n36603 ;
  assign n77345 = ~n36658 ;
  assign n36660 = n36583 & n77345 ;
  assign n36688 = n36349 | n36583 ;
  assign n77346 = ~n36688 ;
  assign n36689 = n36579 & n77346 ;
  assign n36690 = n36660 | n36689 ;
  assign n36691 = n66973 & n36690 ;
  assign n36692 = n77340 & n36691 ;
  assign n36693 = n36687 | n36692 ;
  assign n36694 = n66654 & n36693 ;
  assign n36695 = n36348 & n36603 ;
  assign n77347 = ~n36574 ;
  assign n36578 = n77347 & n36577 ;
  assign n36696 = n36358 | n36577 ;
  assign n77348 = ~n36696 ;
  assign n36697 = n36654 & n77348 ;
  assign n36698 = n36578 | n36697 ;
  assign n36699 = n66973 & n36698 ;
  assign n36700 = n77340 & n36699 ;
  assign n36701 = n36695 | n36700 ;
  assign n36702 = n66560 & n36701 ;
  assign n77349 = ~n36700 ;
  assign n36936 = x82 & n77349 ;
  assign n77350 = ~n36695 ;
  assign n36937 = n77350 & n36936 ;
  assign n36938 = n36702 | n36937 ;
  assign n36703 = n36357 & n36603 ;
  assign n77351 = ~n36653 ;
  assign n36655 = n36572 & n77351 ;
  assign n36704 = n36367 | n36572 ;
  assign n77352 = ~n36704 ;
  assign n36705 = n36568 & n77352 ;
  assign n36706 = n36655 | n36705 ;
  assign n36707 = n66973 & n36706 ;
  assign n36708 = n77340 & n36707 ;
  assign n36709 = n36703 | n36708 ;
  assign n36710 = n66505 & n36709 ;
  assign n36711 = n36366 & n36603 ;
  assign n77353 = ~n36563 ;
  assign n36567 = n77353 & n36566 ;
  assign n36712 = n36375 | n36566 ;
  assign n77354 = ~n36712 ;
  assign n36713 = n36649 & n77354 ;
  assign n36714 = n36567 | n36713 ;
  assign n36715 = n66973 & n36714 ;
  assign n36716 = n77340 & n36715 ;
  assign n36717 = n36711 | n36716 ;
  assign n36718 = n66379 & n36717 ;
  assign n77355 = ~n36716 ;
  assign n36924 = x80 & n77355 ;
  assign n77356 = ~n36711 ;
  assign n36925 = n77356 & n36924 ;
  assign n36926 = n36718 | n36925 ;
  assign n36719 = n36374 & n36603 ;
  assign n77357 = ~n36648 ;
  assign n36650 = n36561 & n77357 ;
  assign n36720 = n36383 | n36561 ;
  assign n77358 = ~n36720 ;
  assign n36721 = n36557 & n77358 ;
  assign n36722 = n36650 | n36721 ;
  assign n36723 = n66973 & n36722 ;
  assign n36724 = n77340 & n36723 ;
  assign n36725 = n36719 | n36724 ;
  assign n36726 = n66299 & n36725 ;
  assign n36727 = n36382 & n36603 ;
  assign n77359 = ~n36552 ;
  assign n36556 = n77359 & n36555 ;
  assign n36728 = n36392 | n36555 ;
  assign n77360 = ~n36728 ;
  assign n36729 = n36644 & n77360 ;
  assign n36730 = n36556 | n36729 ;
  assign n36731 = n66973 & n36730 ;
  assign n36732 = n77340 & n36731 ;
  assign n36733 = n36727 | n36732 ;
  assign n36734 = n66244 & n36733 ;
  assign n77361 = ~n36732 ;
  assign n36912 = x78 & n77361 ;
  assign n77362 = ~n36727 ;
  assign n36913 = n77362 & n36912 ;
  assign n36914 = n36734 | n36913 ;
  assign n36735 = n36391 & n36603 ;
  assign n77363 = ~n36643 ;
  assign n36645 = n36550 & n77363 ;
  assign n36736 = n36401 | n36550 ;
  assign n77364 = ~n36736 ;
  assign n36737 = n36546 & n77364 ;
  assign n36738 = n36645 | n36737 ;
  assign n36739 = n66973 & n36738 ;
  assign n36740 = n77340 & n36739 ;
  assign n36741 = n36735 | n36740 ;
  assign n36742 = n66145 & n36741 ;
  assign n36743 = n36400 & n36603 ;
  assign n77365 = ~n36541 ;
  assign n36545 = n77365 & n36544 ;
  assign n36744 = n36410 | n36544 ;
  assign n77366 = ~n36744 ;
  assign n36745 = n36639 & n77366 ;
  assign n36746 = n36545 | n36745 ;
  assign n36747 = n66973 & n36746 ;
  assign n36748 = n77340 & n36747 ;
  assign n36749 = n36743 | n36748 ;
  assign n36750 = n66081 & n36749 ;
  assign n77367 = ~n36748 ;
  assign n36900 = x76 & n77367 ;
  assign n77368 = ~n36743 ;
  assign n36901 = n77368 & n36900 ;
  assign n36902 = n36750 | n36901 ;
  assign n36751 = n36409 & n36603 ;
  assign n77369 = ~n36638 ;
  assign n36640 = n36539 & n77369 ;
  assign n36752 = n36419 | n36539 ;
  assign n77370 = ~n36752 ;
  assign n36753 = n36535 & n77370 ;
  assign n36754 = n36640 | n36753 ;
  assign n36755 = n66973 & n36754 ;
  assign n36756 = n77340 & n36755 ;
  assign n36757 = n36751 | n36756 ;
  assign n36758 = n66043 & n36757 ;
  assign n36759 = n36418 & n36603 ;
  assign n77371 = ~n36530 ;
  assign n36534 = n77371 & n36533 ;
  assign n36760 = n36428 | n36533 ;
  assign n77372 = ~n36760 ;
  assign n36761 = n36634 & n77372 ;
  assign n36762 = n36534 | n36761 ;
  assign n36763 = n66973 & n36762 ;
  assign n36764 = n77340 & n36763 ;
  assign n36765 = n36759 | n36764 ;
  assign n36766 = n65960 & n36765 ;
  assign n77373 = ~n36764 ;
  assign n36888 = x74 & n77373 ;
  assign n77374 = ~n36759 ;
  assign n36889 = n77374 & n36888 ;
  assign n36890 = n36766 | n36889 ;
  assign n36767 = n36427 & n36603 ;
  assign n77375 = ~n36633 ;
  assign n36635 = n36528 & n77375 ;
  assign n36768 = n36436 | n36528 ;
  assign n77376 = ~n36768 ;
  assign n36769 = n36524 & n77376 ;
  assign n36770 = n36635 | n36769 ;
  assign n36771 = n66973 & n36770 ;
  assign n36772 = n77340 & n36771 ;
  assign n36773 = n36767 | n36772 ;
  assign n36774 = n65909 & n36773 ;
  assign n36775 = n36435 & n36603 ;
  assign n77377 = ~n36518 ;
  assign n36522 = n77377 & n36521 ;
  assign n36523 = n36445 | n36521 ;
  assign n36776 = n36516 | n36628 ;
  assign n77378 = ~n36523 ;
  assign n36777 = n77378 & n36776 ;
  assign n36778 = n36522 | n36777 ;
  assign n36779 = n66973 & n36778 ;
  assign n36780 = n77340 & n36779 ;
  assign n36781 = n36775 | n36780 ;
  assign n36782 = n65877 & n36781 ;
  assign n77379 = ~n36780 ;
  assign n36876 = x72 & n77379 ;
  assign n77380 = ~n36775 ;
  assign n36877 = n77380 & n36876 ;
  assign n36878 = n36782 | n36877 ;
  assign n36606 = n36444 & n36603 ;
  assign n77381 = ~n36628 ;
  assign n36630 = n36516 & n77381 ;
  assign n36783 = n36509 | n36625 ;
  assign n36784 = n36454 | n36516 ;
  assign n77382 = ~n36784 ;
  assign n36785 = n36783 & n77382 ;
  assign n36786 = n36630 | n36785 ;
  assign n36787 = n66973 & n36786 ;
  assign n36788 = n77340 & n36787 ;
  assign n36789 = n36606 | n36788 ;
  assign n36790 = n65820 & n36789 ;
  assign n36607 = n36453 & n36603 ;
  assign n77383 = ~n36509 ;
  assign n36626 = n77383 & n36625 ;
  assign n36791 = n36507 | n36621 ;
  assign n36792 = n36464 | n36625 ;
  assign n77384 = ~n36792 ;
  assign n36793 = n36791 & n77384 ;
  assign n36794 = n36626 | n36793 ;
  assign n36795 = n66973 & n36794 ;
  assign n36796 = n77340 & n36795 ;
  assign n36797 = n36607 | n36796 ;
  assign n36798 = n65791 & n36797 ;
  assign n77385 = ~n36796 ;
  assign n36864 = x70 & n77385 ;
  assign n77386 = ~n36607 ;
  assign n36865 = n77386 & n36864 ;
  assign n36866 = n36798 | n36865 ;
  assign n36605 = n36463 & n36603 ;
  assign n77387 = ~n36621 ;
  assign n36623 = n36507 & n77387 ;
  assign n36799 = n36500 | n36618 ;
  assign n36800 = n36473 | n36507 ;
  assign n77388 = ~n36800 ;
  assign n36801 = n36799 & n77388 ;
  assign n36802 = n36623 | n36801 ;
  assign n36803 = n66973 & n36802 ;
  assign n36804 = n77340 & n36803 ;
  assign n36805 = n36605 | n36804 ;
  assign n36806 = n65772 & n36805 ;
  assign n36608 = n36472 & n36603 ;
  assign n77389 = ~n36500 ;
  assign n36619 = n77389 & n36618 ;
  assign n36807 = n36481 | n36618 ;
  assign n77390 = ~n36807 ;
  assign n36808 = n36499 & n77390 ;
  assign n36809 = n36619 | n36808 ;
  assign n36810 = n66973 & n36809 ;
  assign n36811 = n77340 & n36810 ;
  assign n36812 = n36608 | n36811 ;
  assign n36813 = n65746 & n36812 ;
  assign n77391 = ~n36811 ;
  assign n36854 = x68 & n77391 ;
  assign n77392 = ~n36608 ;
  assign n36855 = n77392 & n36854 ;
  assign n36856 = n36813 | n36855 ;
  assign n36610 = n36480 & n36603 ;
  assign n36814 = n36494 | n36498 ;
  assign n77393 = ~n36814 ;
  assign n36815 = n36614 & n77393 ;
  assign n77394 = ~n36615 ;
  assign n36816 = n36498 & n77394 ;
  assign n36817 = n36815 | n36816 ;
  assign n36818 = n66973 & n36817 ;
  assign n36819 = n77340 & n36818 ;
  assign n36820 = n36610 | n36819 ;
  assign n36821 = n65721 & n36820 ;
  assign n36822 = n36603 & n36611 ;
  assign n36823 = n4058 & n36491 ;
  assign n36824 = n77268 & n36823 ;
  assign n36825 = n4182 | n36824 ;
  assign n77395 = ~n36825 ;
  assign n36826 = n36614 & n77395 ;
  assign n36827 = n77340 & n36826 ;
  assign n36828 = n36822 | n36827 ;
  assign n36829 = n65686 & n36828 ;
  assign n77396 = ~n36827 ;
  assign n36844 = x66 & n77396 ;
  assign n77397 = ~n36822 ;
  assign n36845 = n77397 & n36844 ;
  assign n36846 = n36829 | n36845 ;
  assign n36830 = n77326 & n36665 ;
  assign n36831 = n36599 | n36830 ;
  assign n36832 = n77329 & n36831 ;
  assign n77398 = ~n36832 ;
  assign n36833 = n4403 & n77398 ;
  assign n77399 = ~n36833 ;
  assign n36834 = x42 & n77399 ;
  assign n36835 = n4410 & n77340 ;
  assign n36836 = n36834 | n36835 ;
  assign n36837 = x65 & n36836 ;
  assign n36838 = x65 | n36835 ;
  assign n36839 = n36834 | n36838 ;
  assign n77400 = ~n36837 ;
  assign n36840 = n77400 & n36839 ;
  assign n36842 = n4418 | n36840 ;
  assign n36843 = n65670 & n36836 ;
  assign n77401 = ~n36843 ;
  assign n36847 = n36842 & n77401 ;
  assign n36848 = n36846 | n36847 ;
  assign n77402 = ~n36829 ;
  assign n36849 = n77402 & n36848 ;
  assign n77403 = ~n36819 ;
  assign n36850 = x67 & n77403 ;
  assign n77404 = ~n36610 ;
  assign n36851 = n77404 & n36850 ;
  assign n36852 = n36821 | n36851 ;
  assign n36853 = n36849 | n36852 ;
  assign n77405 = ~n36821 ;
  assign n36857 = n77405 & n36853 ;
  assign n36858 = n36856 | n36857 ;
  assign n77406 = ~n36813 ;
  assign n36859 = n77406 & n36858 ;
  assign n77407 = ~n36804 ;
  assign n36860 = x69 & n77407 ;
  assign n77408 = ~n36605 ;
  assign n36861 = n77408 & n36860 ;
  assign n36862 = n36806 | n36861 ;
  assign n36863 = n36859 | n36862 ;
  assign n77409 = ~n36806 ;
  assign n36868 = n77409 & n36863 ;
  assign n36869 = n36866 | n36868 ;
  assign n77410 = ~n36798 ;
  assign n36870 = n77410 & n36869 ;
  assign n77411 = ~n36788 ;
  assign n36871 = x71 & n77411 ;
  assign n77412 = ~n36606 ;
  assign n36872 = n77412 & n36871 ;
  assign n36873 = n36790 | n36872 ;
  assign n36875 = n36870 | n36873 ;
  assign n77413 = ~n36790 ;
  assign n36880 = n77413 & n36875 ;
  assign n36881 = n36878 | n36880 ;
  assign n77414 = ~n36782 ;
  assign n36882 = n77414 & n36881 ;
  assign n77415 = ~n36772 ;
  assign n36883 = x73 & n77415 ;
  assign n77416 = ~n36767 ;
  assign n36884 = n77416 & n36883 ;
  assign n36885 = n36774 | n36884 ;
  assign n36887 = n36882 | n36885 ;
  assign n77417 = ~n36774 ;
  assign n36892 = n77417 & n36887 ;
  assign n36893 = n36890 | n36892 ;
  assign n77418 = ~n36766 ;
  assign n36894 = n77418 & n36893 ;
  assign n77419 = ~n36756 ;
  assign n36895 = x75 & n77419 ;
  assign n77420 = ~n36751 ;
  assign n36896 = n77420 & n36895 ;
  assign n36897 = n36758 | n36896 ;
  assign n36899 = n36894 | n36897 ;
  assign n77421 = ~n36758 ;
  assign n36904 = n77421 & n36899 ;
  assign n36905 = n36902 | n36904 ;
  assign n77422 = ~n36750 ;
  assign n36906 = n77422 & n36905 ;
  assign n77423 = ~n36740 ;
  assign n36907 = x77 & n77423 ;
  assign n77424 = ~n36735 ;
  assign n36908 = n77424 & n36907 ;
  assign n36909 = n36742 | n36908 ;
  assign n36911 = n36906 | n36909 ;
  assign n77425 = ~n36742 ;
  assign n36916 = n77425 & n36911 ;
  assign n36917 = n36914 | n36916 ;
  assign n77426 = ~n36734 ;
  assign n36918 = n77426 & n36917 ;
  assign n77427 = ~n36724 ;
  assign n36919 = x79 & n77427 ;
  assign n77428 = ~n36719 ;
  assign n36920 = n77428 & n36919 ;
  assign n36921 = n36726 | n36920 ;
  assign n36923 = n36918 | n36921 ;
  assign n77429 = ~n36726 ;
  assign n36928 = n77429 & n36923 ;
  assign n36929 = n36926 | n36928 ;
  assign n77430 = ~n36718 ;
  assign n36930 = n77430 & n36929 ;
  assign n77431 = ~n36708 ;
  assign n36931 = x81 & n77431 ;
  assign n77432 = ~n36703 ;
  assign n36932 = n77432 & n36931 ;
  assign n36933 = n36710 | n36932 ;
  assign n36935 = n36930 | n36933 ;
  assign n77433 = ~n36710 ;
  assign n36940 = n77433 & n36935 ;
  assign n36941 = n36938 | n36940 ;
  assign n77434 = ~n36702 ;
  assign n36942 = n77434 & n36941 ;
  assign n77435 = ~n36692 ;
  assign n36943 = x83 & n77435 ;
  assign n77436 = ~n36687 ;
  assign n36944 = n77436 & n36943 ;
  assign n36945 = n36694 | n36944 ;
  assign n36947 = n36942 | n36945 ;
  assign n77437 = ~n36694 ;
  assign n36952 = n77437 & n36947 ;
  assign n36953 = n36950 | n36952 ;
  assign n77438 = ~n36686 ;
  assign n36954 = n77438 & n36953 ;
  assign n77439 = ~n36670 ;
  assign n36955 = x85 & n77439 ;
  assign n77440 = ~n36609 ;
  assign n36956 = n77440 & n36955 ;
  assign n36957 = n36678 | n36956 ;
  assign n36959 = n36954 | n36957 ;
  assign n77441 = ~n36678 ;
  assign n36965 = n77441 & n36959 ;
  assign n36966 = n36964 | n36965 ;
  assign n77442 = ~n36677 ;
  assign n36967 = n77442 & n36966 ;
  assign n36968 = n4546 | n36967 ;
  assign n77443 = ~n36676 ;
  assign n36970 = n77443 & n36968 ;
  assign n77444 = ~n36965 ;
  assign n37317 = n36964 & n77444 ;
  assign n36972 = n4403 & n77340 ;
  assign n77445 = ~n36972 ;
  assign n36973 = x42 & n77445 ;
  assign n36974 = n36835 | n36973 ;
  assign n36975 = x65 & n36974 ;
  assign n77446 = ~n36975 ;
  assign n36976 = n36839 & n77446 ;
  assign n36977 = n4418 | n36976 ;
  assign n36978 = n77401 & n36977 ;
  assign n36979 = n36846 | n36978 ;
  assign n36980 = n77402 & n36979 ;
  assign n36981 = n36852 | n36980 ;
  assign n36982 = n77405 & n36981 ;
  assign n36983 = n36856 | n36982 ;
  assign n36984 = n77406 & n36983 ;
  assign n36985 = n36862 | n36984 ;
  assign n36986 = n77409 & n36985 ;
  assign n36987 = n36866 | n36986 ;
  assign n36988 = n77410 & n36987 ;
  assign n36989 = n36873 | n36988 ;
  assign n36990 = n77413 & n36989 ;
  assign n36991 = n36878 | n36990 ;
  assign n36992 = n77414 & n36991 ;
  assign n36993 = n36885 | n36992 ;
  assign n36994 = n77417 & n36993 ;
  assign n36995 = n36890 | n36994 ;
  assign n36996 = n77418 & n36995 ;
  assign n36997 = n36897 | n36996 ;
  assign n36998 = n77421 & n36997 ;
  assign n36999 = n36902 | n36998 ;
  assign n37000 = n77422 & n36999 ;
  assign n37001 = n36909 | n37000 ;
  assign n37002 = n77425 & n37001 ;
  assign n37003 = n36914 | n37002 ;
  assign n37004 = n77426 & n37003 ;
  assign n37005 = n36921 | n37004 ;
  assign n37006 = n77429 & n37005 ;
  assign n37007 = n36926 | n37006 ;
  assign n37008 = n77430 & n37007 ;
  assign n37009 = n36933 | n37008 ;
  assign n37010 = n77433 & n37009 ;
  assign n37011 = n36938 | n37010 ;
  assign n37012 = n77434 & n37011 ;
  assign n37013 = n36945 | n37012 ;
  assign n37014 = n77437 & n37013 ;
  assign n37015 = n36950 | n37014 ;
  assign n37017 = n77438 & n37015 ;
  assign n37187 = n36957 | n37017 ;
  assign n37318 = n36678 | n36964 ;
  assign n77447 = ~n37318 ;
  assign n37319 = n37187 & n77447 ;
  assign n37320 = n37317 | n37319 ;
  assign n37321 = n36968 | n37320 ;
  assign n77448 = ~n36970 ;
  assign n37322 = n77448 & n37321 ;
  assign n37330 = n67101 & n37322 ;
  assign n36971 = n36671 & n36968 ;
  assign n36958 = n36686 | n36957 ;
  assign n77449 = ~n36958 ;
  assign n37016 = n77449 & n37015 ;
  assign n77450 = ~n37017 ;
  assign n37018 = n36957 & n77450 ;
  assign n37019 = n37016 | n37018 ;
  assign n37020 = n67101 & n37019 ;
  assign n77451 = ~n36967 ;
  assign n37021 = n77451 & n37020 ;
  assign n37022 = n36971 | n37021 ;
  assign n37023 = n66979 & n37022 ;
  assign n37024 = n36685 & n36968 ;
  assign n36951 = n36694 | n36950 ;
  assign n77452 = ~n36951 ;
  assign n37025 = n36947 & n77452 ;
  assign n77453 = ~n36952 ;
  assign n37026 = n36950 & n77453 ;
  assign n37027 = n37025 | n37026 ;
  assign n37028 = n67101 & n37027 ;
  assign n37029 = n77451 & n37028 ;
  assign n37030 = n37024 | n37029 ;
  assign n37031 = n66868 & n37030 ;
  assign n37032 = n36693 & n36968 ;
  assign n36946 = n36702 | n36945 ;
  assign n77454 = ~n36946 ;
  assign n37033 = n77454 & n37011 ;
  assign n77455 = ~n37012 ;
  assign n37034 = n36945 & n77455 ;
  assign n37035 = n37033 | n37034 ;
  assign n37036 = n67101 & n37035 ;
  assign n37037 = n77451 & n37036 ;
  assign n37038 = n37032 | n37037 ;
  assign n37039 = n66797 & n37038 ;
  assign n37040 = n36701 & n36968 ;
  assign n36939 = n36710 | n36938 ;
  assign n77456 = ~n36939 ;
  assign n37041 = n36935 & n77456 ;
  assign n77457 = ~n36940 ;
  assign n37042 = n36938 & n77457 ;
  assign n37043 = n37041 | n37042 ;
  assign n37044 = n67101 & n37043 ;
  assign n37045 = n77451 & n37044 ;
  assign n37046 = n37040 | n37045 ;
  assign n37047 = n66654 & n37046 ;
  assign n37048 = n36709 & n36968 ;
  assign n36934 = n36718 | n36933 ;
  assign n77458 = ~n36934 ;
  assign n37049 = n77458 & n37007 ;
  assign n77459 = ~n37008 ;
  assign n37050 = n36933 & n77459 ;
  assign n37051 = n37049 | n37050 ;
  assign n37052 = n67101 & n37051 ;
  assign n37053 = n77451 & n37052 ;
  assign n37054 = n37048 | n37053 ;
  assign n37055 = n66560 & n37054 ;
  assign n37056 = n36717 & n36968 ;
  assign n36927 = n36726 | n36926 ;
  assign n77460 = ~n36927 ;
  assign n37057 = n36923 & n77460 ;
  assign n77461 = ~n36928 ;
  assign n37058 = n36926 & n77461 ;
  assign n37059 = n37057 | n37058 ;
  assign n37060 = n67101 & n37059 ;
  assign n37061 = n77451 & n37060 ;
  assign n37062 = n37056 | n37061 ;
  assign n37063 = n66505 & n37062 ;
  assign n37064 = n36725 & n36968 ;
  assign n36922 = n36734 | n36921 ;
  assign n77462 = ~n36922 ;
  assign n37065 = n77462 & n37003 ;
  assign n77463 = ~n37004 ;
  assign n37066 = n36921 & n77463 ;
  assign n37067 = n37065 | n37066 ;
  assign n37068 = n67101 & n37067 ;
  assign n37069 = n77451 & n37068 ;
  assign n37070 = n37064 | n37069 ;
  assign n37071 = n66379 & n37070 ;
  assign n37072 = n36733 & n36968 ;
  assign n36915 = n36742 | n36914 ;
  assign n77464 = ~n36915 ;
  assign n37073 = n36911 & n77464 ;
  assign n77465 = ~n36916 ;
  assign n37074 = n36914 & n77465 ;
  assign n37075 = n37073 | n37074 ;
  assign n37076 = n67101 & n37075 ;
  assign n37077 = n77451 & n37076 ;
  assign n37078 = n37072 | n37077 ;
  assign n37079 = n66299 & n37078 ;
  assign n37080 = n36741 & n36968 ;
  assign n36910 = n36750 | n36909 ;
  assign n77466 = ~n36910 ;
  assign n37081 = n77466 & n36999 ;
  assign n77467 = ~n37000 ;
  assign n37082 = n36909 & n77467 ;
  assign n37083 = n37081 | n37082 ;
  assign n37084 = n67101 & n37083 ;
  assign n37085 = n77451 & n37084 ;
  assign n37086 = n37080 | n37085 ;
  assign n37087 = n66244 & n37086 ;
  assign n37088 = n36749 & n36968 ;
  assign n36903 = n36758 | n36902 ;
  assign n77468 = ~n36903 ;
  assign n37089 = n36899 & n77468 ;
  assign n77469 = ~n36904 ;
  assign n37090 = n36902 & n77469 ;
  assign n37091 = n37089 | n37090 ;
  assign n37092 = n67101 & n37091 ;
  assign n37093 = n77451 & n37092 ;
  assign n37094 = n37088 | n37093 ;
  assign n37095 = n66145 & n37094 ;
  assign n37096 = n36757 & n36968 ;
  assign n36898 = n36766 | n36897 ;
  assign n77470 = ~n36898 ;
  assign n37097 = n77470 & n36995 ;
  assign n77471 = ~n36996 ;
  assign n37098 = n36897 & n77471 ;
  assign n37099 = n37097 | n37098 ;
  assign n37100 = n67101 & n37099 ;
  assign n37101 = n77451 & n37100 ;
  assign n37102 = n37096 | n37101 ;
  assign n37103 = n66081 & n37102 ;
  assign n37104 = n36765 & n36968 ;
  assign n36891 = n36774 | n36890 ;
  assign n77472 = ~n36891 ;
  assign n37105 = n36887 & n77472 ;
  assign n77473 = ~n36892 ;
  assign n37106 = n36890 & n77473 ;
  assign n37107 = n37105 | n37106 ;
  assign n37108 = n67101 & n37107 ;
  assign n37109 = n77451 & n37108 ;
  assign n37110 = n37104 | n37109 ;
  assign n37111 = n66043 & n37110 ;
  assign n37112 = n36773 & n36968 ;
  assign n36886 = n36782 | n36885 ;
  assign n77474 = ~n36886 ;
  assign n37113 = n77474 & n36991 ;
  assign n77475 = ~n36992 ;
  assign n37114 = n36885 & n77475 ;
  assign n37115 = n37113 | n37114 ;
  assign n37116 = n67101 & n37115 ;
  assign n37117 = n77451 & n37116 ;
  assign n37118 = n37112 | n37117 ;
  assign n37119 = n65960 & n37118 ;
  assign n37120 = n36781 & n36968 ;
  assign n36879 = n36790 | n36878 ;
  assign n77476 = ~n36879 ;
  assign n37121 = n36875 & n77476 ;
  assign n77477 = ~n36880 ;
  assign n37122 = n36878 & n77477 ;
  assign n37123 = n37121 | n37122 ;
  assign n37124 = n67101 & n37123 ;
  assign n37125 = n77451 & n37124 ;
  assign n37126 = n37120 | n37125 ;
  assign n37127 = n65909 & n37126 ;
  assign n37128 = n36789 & n36968 ;
  assign n36874 = n36798 | n36873 ;
  assign n77478 = ~n36874 ;
  assign n37129 = n77478 & n36987 ;
  assign n77479 = ~n36988 ;
  assign n37130 = n36873 & n77479 ;
  assign n37131 = n37129 | n37130 ;
  assign n37132 = n67101 & n37131 ;
  assign n37133 = n77451 & n37132 ;
  assign n37134 = n37128 | n37133 ;
  assign n37135 = n65877 & n37134 ;
  assign n37136 = n36797 & n36968 ;
  assign n36867 = n36806 | n36866 ;
  assign n77480 = ~n36867 ;
  assign n37137 = n77480 & n36985 ;
  assign n77481 = ~n36868 ;
  assign n37138 = n36866 & n77481 ;
  assign n37139 = n37137 | n37138 ;
  assign n37140 = n67101 & n37139 ;
  assign n37141 = n77451 & n37140 ;
  assign n37142 = n37136 | n37141 ;
  assign n37143 = n65820 & n37142 ;
  assign n37144 = n36805 & n36968 ;
  assign n37145 = n36813 | n36862 ;
  assign n77482 = ~n37145 ;
  assign n37146 = n36983 & n77482 ;
  assign n77483 = ~n36984 ;
  assign n37147 = n36862 & n77483 ;
  assign n37148 = n37146 | n37147 ;
  assign n37149 = n67101 & n37148 ;
  assign n37150 = n77451 & n37149 ;
  assign n37151 = n37144 | n37150 ;
  assign n37152 = n65791 & n37151 ;
  assign n37153 = n36812 & n36968 ;
  assign n37154 = n36821 | n36856 ;
  assign n77484 = ~n37154 ;
  assign n37155 = n36981 & n77484 ;
  assign n77485 = ~n36857 ;
  assign n37156 = n36856 & n77485 ;
  assign n37157 = n37155 | n37156 ;
  assign n37158 = n67101 & n37157 ;
  assign n37159 = n77451 & n37158 ;
  assign n37160 = n37153 | n37159 ;
  assign n37161 = n65772 & n37160 ;
  assign n37162 = n36820 & n36968 ;
  assign n37163 = n36829 | n36852 ;
  assign n77486 = ~n37163 ;
  assign n37164 = n36979 & n77486 ;
  assign n77487 = ~n36980 ;
  assign n37165 = n36852 & n77487 ;
  assign n37166 = n37164 | n37165 ;
  assign n37167 = n67101 & n37166 ;
  assign n37168 = n77451 & n37167 ;
  assign n37169 = n37162 | n37168 ;
  assign n37170 = n65746 & n37169 ;
  assign n37171 = n36828 & n36968 ;
  assign n77488 = ~n36978 ;
  assign n37172 = n36846 & n77488 ;
  assign n37173 = n36843 | n36846 ;
  assign n77489 = ~n37173 ;
  assign n37174 = n36977 & n77489 ;
  assign n37175 = n37172 | n37174 ;
  assign n37176 = n67101 & n37175 ;
  assign n37177 = n77451 & n37176 ;
  assign n37178 = n37171 | n37177 ;
  assign n37179 = n65721 & n37178 ;
  assign n36969 = n36836 & n36968 ;
  assign n36841 = n4418 & n36839 ;
  assign n37180 = n36841 & n77446 ;
  assign n37181 = n4546 | n37180 ;
  assign n77490 = ~n37181 ;
  assign n37182 = n36977 & n77490 ;
  assign n37183 = n77451 & n37182 ;
  assign n37184 = n36969 | n37183 ;
  assign n37185 = n65686 & n37184 ;
  assign n37186 = n4787 & n77451 ;
  assign n37188 = n77441 & n37187 ;
  assign n37189 = n36964 | n37188 ;
  assign n37190 = n77442 & n37189 ;
  assign n77491 = ~n37190 ;
  assign n37191 = n4780 & n77491 ;
  assign n77492 = ~n37191 ;
  assign n37192 = x41 & n77492 ;
  assign n37193 = n37186 | n37192 ;
  assign n37201 = n65670 & n37193 ;
  assign n37194 = n4780 & n77451 ;
  assign n77493 = ~n37194 ;
  assign n37195 = x41 & n77493 ;
  assign n37196 = n37186 | n37195 ;
  assign n37197 = x65 & n37196 ;
  assign n37198 = x65 | n37186 ;
  assign n37199 = n37195 | n37198 ;
  assign n77494 = ~n37197 ;
  assign n37200 = n77494 & n37199 ;
  assign n37202 = n4794 | n37200 ;
  assign n77495 = ~n37201 ;
  assign n37203 = n77495 & n37202 ;
  assign n77496 = ~n37183 ;
  assign n37204 = x66 & n77496 ;
  assign n77497 = ~n36969 ;
  assign n37205 = n77497 & n37204 ;
  assign n37206 = n37203 | n37205 ;
  assign n77498 = ~n37185 ;
  assign n37207 = n77498 & n37206 ;
  assign n77499 = ~n37177 ;
  assign n37208 = x67 & n77499 ;
  assign n77500 = ~n37171 ;
  assign n37209 = n77500 & n37208 ;
  assign n37210 = n37179 | n37209 ;
  assign n37211 = n37207 | n37210 ;
  assign n77501 = ~n37179 ;
  assign n37212 = n77501 & n37211 ;
  assign n77502 = ~n37168 ;
  assign n37213 = x68 & n77502 ;
  assign n77503 = ~n37162 ;
  assign n37214 = n77503 & n37213 ;
  assign n37215 = n37170 | n37214 ;
  assign n37216 = n37212 | n37215 ;
  assign n77504 = ~n37170 ;
  assign n37217 = n77504 & n37216 ;
  assign n77505 = ~n37159 ;
  assign n37218 = x69 & n77505 ;
  assign n77506 = ~n37153 ;
  assign n37219 = n77506 & n37218 ;
  assign n37220 = n37161 | n37219 ;
  assign n37221 = n37217 | n37220 ;
  assign n77507 = ~n37161 ;
  assign n37222 = n77507 & n37221 ;
  assign n77508 = ~n37150 ;
  assign n37223 = x70 & n77508 ;
  assign n77509 = ~n37144 ;
  assign n37224 = n77509 & n37223 ;
  assign n37225 = n37152 | n37224 ;
  assign n37227 = n37222 | n37225 ;
  assign n77510 = ~n37152 ;
  assign n37228 = n77510 & n37227 ;
  assign n77511 = ~n37141 ;
  assign n37229 = x71 & n77511 ;
  assign n77512 = ~n37136 ;
  assign n37230 = n77512 & n37229 ;
  assign n37231 = n37143 | n37230 ;
  assign n37232 = n37228 | n37231 ;
  assign n77513 = ~n37143 ;
  assign n37233 = n77513 & n37232 ;
  assign n77514 = ~n37133 ;
  assign n37234 = x72 & n77514 ;
  assign n77515 = ~n37128 ;
  assign n37235 = n77515 & n37234 ;
  assign n37236 = n37135 | n37235 ;
  assign n37238 = n37233 | n37236 ;
  assign n77516 = ~n37135 ;
  assign n37239 = n77516 & n37238 ;
  assign n77517 = ~n37125 ;
  assign n37240 = x73 & n77517 ;
  assign n77518 = ~n37120 ;
  assign n37241 = n77518 & n37240 ;
  assign n37242 = n37127 | n37241 ;
  assign n37243 = n37239 | n37242 ;
  assign n77519 = ~n37127 ;
  assign n37244 = n77519 & n37243 ;
  assign n77520 = ~n37117 ;
  assign n37245 = x74 & n77520 ;
  assign n77521 = ~n37112 ;
  assign n37246 = n77521 & n37245 ;
  assign n37247 = n37119 | n37246 ;
  assign n37249 = n37244 | n37247 ;
  assign n77522 = ~n37119 ;
  assign n37250 = n77522 & n37249 ;
  assign n77523 = ~n37109 ;
  assign n37251 = x75 & n77523 ;
  assign n77524 = ~n37104 ;
  assign n37252 = n77524 & n37251 ;
  assign n37253 = n37111 | n37252 ;
  assign n37254 = n37250 | n37253 ;
  assign n77525 = ~n37111 ;
  assign n37255 = n77525 & n37254 ;
  assign n77526 = ~n37101 ;
  assign n37256 = x76 & n77526 ;
  assign n77527 = ~n37096 ;
  assign n37257 = n77527 & n37256 ;
  assign n37258 = n37103 | n37257 ;
  assign n37260 = n37255 | n37258 ;
  assign n77528 = ~n37103 ;
  assign n37261 = n77528 & n37260 ;
  assign n77529 = ~n37093 ;
  assign n37262 = x77 & n77529 ;
  assign n77530 = ~n37088 ;
  assign n37263 = n77530 & n37262 ;
  assign n37264 = n37095 | n37263 ;
  assign n37265 = n37261 | n37264 ;
  assign n77531 = ~n37095 ;
  assign n37266 = n77531 & n37265 ;
  assign n77532 = ~n37085 ;
  assign n37267 = x78 & n77532 ;
  assign n77533 = ~n37080 ;
  assign n37268 = n77533 & n37267 ;
  assign n37269 = n37087 | n37268 ;
  assign n37271 = n37266 | n37269 ;
  assign n77534 = ~n37087 ;
  assign n37272 = n77534 & n37271 ;
  assign n77535 = ~n37077 ;
  assign n37273 = x79 & n77535 ;
  assign n77536 = ~n37072 ;
  assign n37274 = n77536 & n37273 ;
  assign n37275 = n37079 | n37274 ;
  assign n37276 = n37272 | n37275 ;
  assign n77537 = ~n37079 ;
  assign n37277 = n77537 & n37276 ;
  assign n77538 = ~n37069 ;
  assign n37278 = x80 & n77538 ;
  assign n77539 = ~n37064 ;
  assign n37279 = n77539 & n37278 ;
  assign n37280 = n37071 | n37279 ;
  assign n37282 = n37277 | n37280 ;
  assign n77540 = ~n37071 ;
  assign n37283 = n77540 & n37282 ;
  assign n77541 = ~n37061 ;
  assign n37284 = x81 & n77541 ;
  assign n77542 = ~n37056 ;
  assign n37285 = n77542 & n37284 ;
  assign n37286 = n37063 | n37285 ;
  assign n37287 = n37283 | n37286 ;
  assign n77543 = ~n37063 ;
  assign n37288 = n77543 & n37287 ;
  assign n77544 = ~n37053 ;
  assign n37289 = x82 & n77544 ;
  assign n77545 = ~n37048 ;
  assign n37290 = n77545 & n37289 ;
  assign n37291 = n37055 | n37290 ;
  assign n37293 = n37288 | n37291 ;
  assign n77546 = ~n37055 ;
  assign n37294 = n77546 & n37293 ;
  assign n77547 = ~n37045 ;
  assign n37295 = x83 & n77547 ;
  assign n77548 = ~n37040 ;
  assign n37296 = n77548 & n37295 ;
  assign n37297 = n37047 | n37296 ;
  assign n37298 = n37294 | n37297 ;
  assign n77549 = ~n37047 ;
  assign n37299 = n77549 & n37298 ;
  assign n77550 = ~n37037 ;
  assign n37300 = x84 & n77550 ;
  assign n77551 = ~n37032 ;
  assign n37301 = n77551 & n37300 ;
  assign n37302 = n37039 | n37301 ;
  assign n37304 = n37299 | n37302 ;
  assign n77552 = ~n37039 ;
  assign n37305 = n77552 & n37304 ;
  assign n77553 = ~n37029 ;
  assign n37306 = x85 & n77553 ;
  assign n77554 = ~n37024 ;
  assign n37307 = n77554 & n37306 ;
  assign n37308 = n37031 | n37307 ;
  assign n37309 = n37305 | n37308 ;
  assign n77555 = ~n37031 ;
  assign n37310 = n77555 & n37309 ;
  assign n77556 = ~n37021 ;
  assign n37311 = x86 & n77556 ;
  assign n77557 = ~n36971 ;
  assign n37312 = n77557 & n37311 ;
  assign n37313 = n37023 | n37312 ;
  assign n37315 = n37310 | n37313 ;
  assign n77558 = ~n37023 ;
  assign n37316 = n77558 & n37315 ;
  assign n37323 = n67164 & n37322 ;
  assign n77559 = ~n36968 ;
  assign n37324 = n77559 & n37320 ;
  assign n37325 = n36676 & n36968 ;
  assign n77560 = ~n37325 ;
  assign n37326 = x87 & n77560 ;
  assign n77561 = ~n37324 ;
  assign n37327 = n77561 & n37326 ;
  assign n37328 = n4915 | n37327 ;
  assign n37329 = n37323 | n37328 ;
  assign n37331 = n37316 | n37329 ;
  assign n77562 = ~n37330 ;
  assign n37332 = n77562 & n37331 ;
  assign n77563 = ~n37310 ;
  assign n37314 = n77563 & n37313 ;
  assign n37335 = x65 & n37193 ;
  assign n77564 = ~n37335 ;
  assign n37336 = n37199 & n77564 ;
  assign n37337 = n4794 | n37336 ;
  assign n37338 = n77495 & n37337 ;
  assign n37339 = n37185 | n37205 ;
  assign n37341 = n37338 | n37339 ;
  assign n37342 = n77498 & n37341 ;
  assign n37343 = n37209 | n37342 ;
  assign n37345 = n77501 & n37343 ;
  assign n37347 = n37215 | n37345 ;
  assign n37348 = n77504 & n37347 ;
  assign n37350 = n37220 | n37348 ;
  assign n37351 = n77507 & n37350 ;
  assign n37352 = n37225 | n37351 ;
  assign n37353 = n77510 & n37352 ;
  assign n37354 = n37231 | n37353 ;
  assign n37356 = n77513 & n37354 ;
  assign n37357 = n37236 | n37356 ;
  assign n37358 = n77516 & n37357 ;
  assign n37359 = n37242 | n37358 ;
  assign n37361 = n77519 & n37359 ;
  assign n37362 = n37247 | n37361 ;
  assign n37363 = n77522 & n37362 ;
  assign n37364 = n37253 | n37363 ;
  assign n37366 = n77525 & n37364 ;
  assign n37367 = n37258 | n37366 ;
  assign n37368 = n77528 & n37367 ;
  assign n37369 = n37264 | n37368 ;
  assign n37371 = n77531 & n37369 ;
  assign n37372 = n37269 | n37371 ;
  assign n37373 = n77534 & n37372 ;
  assign n37374 = n37275 | n37373 ;
  assign n37376 = n77537 & n37374 ;
  assign n37377 = n37280 | n37376 ;
  assign n37378 = n77540 & n37377 ;
  assign n37379 = n37286 | n37378 ;
  assign n37381 = n77543 & n37379 ;
  assign n37382 = n37291 | n37381 ;
  assign n37383 = n77546 & n37382 ;
  assign n37384 = n37297 | n37383 ;
  assign n37386 = n77549 & n37384 ;
  assign n37387 = n37302 | n37386 ;
  assign n37388 = n77552 & n37387 ;
  assign n37389 = n37308 | n37388 ;
  assign n37391 = n37031 | n37313 ;
  assign n77565 = ~n37391 ;
  assign n37392 = n37389 & n77565 ;
  assign n37393 = n37314 | n37392 ;
  assign n77566 = ~n37332 ;
  assign n37394 = n77566 & n37393 ;
  assign n37395 = n77555 & n37389 ;
  assign n37396 = n37313 | n37395 ;
  assign n37397 = n77558 & n37396 ;
  assign n37398 = n37329 | n37397 ;
  assign n37399 = n37022 & n77562 ;
  assign n37400 = n37398 & n37399 ;
  assign n37401 = n37394 | n37400 ;
  assign n37402 = n37023 | n37327 ;
  assign n37403 = n37323 | n37402 ;
  assign n77567 = ~n37403 ;
  assign n37404 = n37315 & n77567 ;
  assign n37405 = n37323 | n37327 ;
  assign n77568 = ~n37397 ;
  assign n37406 = n77568 & n37405 ;
  assign n37407 = n37404 | n37406 ;
  assign n37408 = n77566 & n37407 ;
  assign n37409 = n4546 & n36676 ;
  assign n37410 = n37398 & n37409 ;
  assign n37411 = n37408 | n37410 ;
  assign n37412 = n67222 & n37411 ;
  assign n77569 = ~n37410 ;
  assign n37723 = x88 & n77569 ;
  assign n77570 = ~n37408 ;
  assign n37724 = n77570 & n37723 ;
  assign n37725 = n37412 | n37724 ;
  assign n37413 = n67164 & n37401 ;
  assign n77571 = ~n37388 ;
  assign n37390 = n37308 & n77571 ;
  assign n37414 = n37039 | n37308 ;
  assign n77572 = ~n37414 ;
  assign n37415 = n37304 & n77572 ;
  assign n37416 = n37390 | n37415 ;
  assign n37417 = n77566 & n37416 ;
  assign n37418 = n37030 & n77562 ;
  assign n37419 = n37398 & n37418 ;
  assign n37420 = n37417 | n37419 ;
  assign n37421 = n66979 & n37420 ;
  assign n77573 = ~n37419 ;
  assign n37711 = x86 & n77573 ;
  assign n77574 = ~n37417 ;
  assign n37712 = n77574 & n37711 ;
  assign n37713 = n37421 | n37712 ;
  assign n77575 = ~n37299 ;
  assign n37303 = n77575 & n37302 ;
  assign n37422 = n37047 | n37302 ;
  assign n77576 = ~n37422 ;
  assign n37423 = n37384 & n77576 ;
  assign n37424 = n37303 | n37423 ;
  assign n37425 = n77566 & n37424 ;
  assign n37426 = n37038 & n77562 ;
  assign n37427 = n37398 & n37426 ;
  assign n37428 = n37425 | n37427 ;
  assign n37429 = n66868 & n37428 ;
  assign n77577 = ~n37383 ;
  assign n37385 = n37297 & n77577 ;
  assign n37430 = n37055 | n37297 ;
  assign n77578 = ~n37430 ;
  assign n37431 = n37293 & n77578 ;
  assign n37432 = n37385 | n37431 ;
  assign n37433 = n77566 & n37432 ;
  assign n37434 = n37046 & n77562 ;
  assign n37435 = n37398 & n37434 ;
  assign n37436 = n37433 | n37435 ;
  assign n37437 = n66797 & n37436 ;
  assign n77579 = ~n37435 ;
  assign n37699 = x84 & n77579 ;
  assign n77580 = ~n37433 ;
  assign n37700 = n77580 & n37699 ;
  assign n37701 = n37437 | n37700 ;
  assign n77581 = ~n37288 ;
  assign n37292 = n77581 & n37291 ;
  assign n37438 = n37063 | n37291 ;
  assign n77582 = ~n37438 ;
  assign n37439 = n37379 & n77582 ;
  assign n37440 = n37292 | n37439 ;
  assign n37441 = n77566 & n37440 ;
  assign n37442 = n37054 & n77562 ;
  assign n37443 = n37398 & n37442 ;
  assign n37444 = n37441 | n37443 ;
  assign n37445 = n66654 & n37444 ;
  assign n77583 = ~n37378 ;
  assign n37380 = n37286 & n77583 ;
  assign n37446 = n37071 | n37286 ;
  assign n77584 = ~n37446 ;
  assign n37447 = n37282 & n77584 ;
  assign n37448 = n37380 | n37447 ;
  assign n37449 = n77566 & n37448 ;
  assign n37450 = n37062 & n77562 ;
  assign n37451 = n37398 & n37450 ;
  assign n37452 = n37449 | n37451 ;
  assign n37453 = n66560 & n37452 ;
  assign n77585 = ~n37451 ;
  assign n37687 = x82 & n77585 ;
  assign n77586 = ~n37449 ;
  assign n37688 = n77586 & n37687 ;
  assign n37689 = n37453 | n37688 ;
  assign n77587 = ~n37277 ;
  assign n37281 = n77587 & n37280 ;
  assign n37454 = n37079 | n37280 ;
  assign n77588 = ~n37454 ;
  assign n37455 = n37374 & n77588 ;
  assign n37456 = n37281 | n37455 ;
  assign n37457 = n77566 & n37456 ;
  assign n37458 = n37070 & n77562 ;
  assign n37459 = n37398 & n37458 ;
  assign n37460 = n37457 | n37459 ;
  assign n37461 = n66505 & n37460 ;
  assign n77589 = ~n37373 ;
  assign n37375 = n37275 & n77589 ;
  assign n37462 = n37087 | n37275 ;
  assign n77590 = ~n37462 ;
  assign n37463 = n37271 & n77590 ;
  assign n37464 = n37375 | n37463 ;
  assign n37465 = n77566 & n37464 ;
  assign n37466 = n37078 & n77562 ;
  assign n37467 = n37398 & n37466 ;
  assign n37468 = n37465 | n37467 ;
  assign n37469 = n66379 & n37468 ;
  assign n77591 = ~n37467 ;
  assign n37675 = x80 & n77591 ;
  assign n77592 = ~n37465 ;
  assign n37676 = n77592 & n37675 ;
  assign n37677 = n37469 | n37676 ;
  assign n77593 = ~n37266 ;
  assign n37270 = n77593 & n37269 ;
  assign n37470 = n37095 | n37269 ;
  assign n77594 = ~n37470 ;
  assign n37471 = n37369 & n77594 ;
  assign n37472 = n37270 | n37471 ;
  assign n37473 = n77566 & n37472 ;
  assign n37474 = n37086 & n77562 ;
  assign n37475 = n37398 & n37474 ;
  assign n37476 = n37473 | n37475 ;
  assign n37477 = n66299 & n37476 ;
  assign n77595 = ~n37368 ;
  assign n37370 = n37264 & n77595 ;
  assign n37478 = n37103 | n37264 ;
  assign n77596 = ~n37478 ;
  assign n37479 = n37260 & n77596 ;
  assign n37480 = n37370 | n37479 ;
  assign n37481 = n77566 & n37480 ;
  assign n37482 = n37094 & n77562 ;
  assign n37483 = n37398 & n37482 ;
  assign n37484 = n37481 | n37483 ;
  assign n37485 = n66244 & n37484 ;
  assign n77597 = ~n37483 ;
  assign n37663 = x78 & n77597 ;
  assign n77598 = ~n37481 ;
  assign n37664 = n77598 & n37663 ;
  assign n37665 = n37485 | n37664 ;
  assign n77599 = ~n37255 ;
  assign n37259 = n77599 & n37258 ;
  assign n37486 = n37111 | n37258 ;
  assign n77600 = ~n37486 ;
  assign n37487 = n37364 & n77600 ;
  assign n37488 = n37259 | n37487 ;
  assign n37489 = n77566 & n37488 ;
  assign n37490 = n37102 & n77562 ;
  assign n37491 = n37398 & n37490 ;
  assign n37492 = n37489 | n37491 ;
  assign n37493 = n66145 & n37492 ;
  assign n77601 = ~n37363 ;
  assign n37365 = n37253 & n77601 ;
  assign n37494 = n37119 | n37253 ;
  assign n77602 = ~n37494 ;
  assign n37495 = n37249 & n77602 ;
  assign n37496 = n37365 | n37495 ;
  assign n37497 = n77566 & n37496 ;
  assign n37498 = n37110 & n77562 ;
  assign n37499 = n37398 & n37498 ;
  assign n37500 = n37497 | n37499 ;
  assign n37501 = n66081 & n37500 ;
  assign n77603 = ~n37499 ;
  assign n37651 = x76 & n77603 ;
  assign n77604 = ~n37497 ;
  assign n37652 = n77604 & n37651 ;
  assign n37653 = n37501 | n37652 ;
  assign n77605 = ~n37244 ;
  assign n37248 = n77605 & n37247 ;
  assign n37502 = n37127 | n37247 ;
  assign n77606 = ~n37502 ;
  assign n37503 = n37359 & n77606 ;
  assign n37504 = n37248 | n37503 ;
  assign n37505 = n77566 & n37504 ;
  assign n37506 = n37118 & n77562 ;
  assign n37507 = n37398 & n37506 ;
  assign n37508 = n37505 | n37507 ;
  assign n37509 = n66043 & n37508 ;
  assign n77607 = ~n37358 ;
  assign n37360 = n37242 & n77607 ;
  assign n37510 = n37135 | n37242 ;
  assign n77608 = ~n37510 ;
  assign n37511 = n37238 & n77608 ;
  assign n37512 = n37360 | n37511 ;
  assign n37513 = n77566 & n37512 ;
  assign n37514 = n37126 & n77562 ;
  assign n37515 = n37398 & n37514 ;
  assign n37516 = n37513 | n37515 ;
  assign n37517 = n65960 & n37516 ;
  assign n77609 = ~n37515 ;
  assign n37639 = x74 & n77609 ;
  assign n77610 = ~n37513 ;
  assign n37640 = n77610 & n37639 ;
  assign n37641 = n37517 | n37640 ;
  assign n77611 = ~n37233 ;
  assign n37237 = n77611 & n37236 ;
  assign n37518 = n37143 | n37236 ;
  assign n77612 = ~n37518 ;
  assign n37519 = n37354 & n77612 ;
  assign n37520 = n37237 | n37519 ;
  assign n37521 = n77566 & n37520 ;
  assign n37522 = n37134 & n77562 ;
  assign n37523 = n37398 & n37522 ;
  assign n37524 = n37521 | n37523 ;
  assign n37525 = n65909 & n37524 ;
  assign n77613 = ~n37353 ;
  assign n37355 = n37231 & n77613 ;
  assign n37526 = n37152 | n37231 ;
  assign n77614 = ~n37526 ;
  assign n37527 = n37227 & n77614 ;
  assign n37528 = n37355 | n37527 ;
  assign n37529 = n77566 & n37528 ;
  assign n37530 = n37142 & n77562 ;
  assign n37531 = n37398 & n37530 ;
  assign n37532 = n37529 | n37531 ;
  assign n37533 = n65877 & n37532 ;
  assign n77615 = ~n37531 ;
  assign n37627 = x72 & n77615 ;
  assign n77616 = ~n37529 ;
  assign n37628 = n77616 & n37627 ;
  assign n37629 = n37533 | n37628 ;
  assign n77617 = ~n37222 ;
  assign n37226 = n77617 & n37225 ;
  assign n37534 = n37161 | n37225 ;
  assign n77618 = ~n37534 ;
  assign n37535 = n37350 & n77618 ;
  assign n37536 = n37226 | n37535 ;
  assign n37537 = n77566 & n37536 ;
  assign n37538 = n37151 & n77562 ;
  assign n37539 = n37398 & n37538 ;
  assign n37540 = n37537 | n37539 ;
  assign n37541 = n65820 & n37540 ;
  assign n77619 = ~n37348 ;
  assign n37349 = n37220 & n77619 ;
  assign n37542 = n37170 | n37220 ;
  assign n77620 = ~n37542 ;
  assign n37543 = n37216 & n77620 ;
  assign n37544 = n37349 | n37543 ;
  assign n37545 = n77566 & n37544 ;
  assign n37546 = n37160 & n77562 ;
  assign n37547 = n37398 & n37546 ;
  assign n37548 = n37545 | n37547 ;
  assign n37549 = n65791 & n37548 ;
  assign n77621 = ~n37547 ;
  assign n37615 = x70 & n77621 ;
  assign n77622 = ~n37545 ;
  assign n37616 = n77622 & n37615 ;
  assign n37617 = n37549 | n37616 ;
  assign n77623 = ~n37212 ;
  assign n37346 = n77623 & n37215 ;
  assign n37550 = n37210 | n37342 ;
  assign n37551 = n37179 | n37215 ;
  assign n77624 = ~n37551 ;
  assign n37552 = n37550 & n77624 ;
  assign n37553 = n37346 | n37552 ;
  assign n37554 = n77566 & n37553 ;
  assign n37555 = n37169 & n77562 ;
  assign n37556 = n37398 & n37555 ;
  assign n37557 = n37554 | n37556 ;
  assign n37558 = n65772 & n37557 ;
  assign n77625 = ~n37342 ;
  assign n37344 = n37210 & n77625 ;
  assign n37559 = n37185 | n37210 ;
  assign n77626 = ~n37559 ;
  assign n37560 = n37341 & n77626 ;
  assign n37561 = n37344 | n37560 ;
  assign n37562 = n77566 & n37561 ;
  assign n37563 = n37178 & n77562 ;
  assign n37564 = n37398 & n37563 ;
  assign n37565 = n37562 | n37564 ;
  assign n37566 = n65746 & n37565 ;
  assign n77627 = ~n37564 ;
  assign n37604 = x68 & n77627 ;
  assign n77628 = ~n37562 ;
  assign n37605 = n77628 & n37604 ;
  assign n37606 = n37566 | n37605 ;
  assign n77629 = ~n37203 ;
  assign n37340 = n77629 & n37339 ;
  assign n37567 = n37201 | n37339 ;
  assign n77630 = ~n37567 ;
  assign n37568 = n37202 & n77630 ;
  assign n37569 = n37340 | n37568 ;
  assign n37570 = n77566 & n37569 ;
  assign n37571 = n37184 & n77562 ;
  assign n37572 = n37398 & n37571 ;
  assign n37573 = n37570 | n37572 ;
  assign n37574 = n65721 & n37573 ;
  assign n37575 = n4794 & n37199 ;
  assign n37576 = n77564 & n37575 ;
  assign n77631 = ~n37576 ;
  assign n37577 = n37202 & n77631 ;
  assign n37578 = n77566 & n37577 ;
  assign n37579 = n37193 & n77562 ;
  assign n37580 = n37398 & n37579 ;
  assign n37581 = n37578 | n37580 ;
  assign n37582 = n65686 & n37581 ;
  assign n77632 = ~n37580 ;
  assign n37594 = x66 & n77632 ;
  assign n77633 = ~n37578 ;
  assign n37595 = n77633 & n37594 ;
  assign n37596 = n37582 | n37595 ;
  assign n37334 = n4794 & n77566 ;
  assign n37333 = x64 & n77566 ;
  assign n77634 = ~n37333 ;
  assign n37583 = x40 & n77634 ;
  assign n37584 = n37334 | n37583 ;
  assign n37585 = x65 & n37584 ;
  assign n37586 = n77562 & n37398 ;
  assign n77635 = ~n37586 ;
  assign n37587 = n4794 & n77635 ;
  assign n37588 = x65 | n37587 ;
  assign n37589 = n37583 | n37588 ;
  assign n77636 = ~n37585 ;
  assign n37590 = n77636 & n37589 ;
  assign n37592 = n5190 | n37590 ;
  assign n37593 = n65670 & n37584 ;
  assign n77637 = ~n37593 ;
  assign n37597 = n37592 & n77637 ;
  assign n37598 = n37596 | n37597 ;
  assign n77638 = ~n37582 ;
  assign n37599 = n77638 & n37598 ;
  assign n77639 = ~n37572 ;
  assign n37600 = x67 & n77639 ;
  assign n77640 = ~n37570 ;
  assign n37601 = n77640 & n37600 ;
  assign n37602 = n37574 | n37601 ;
  assign n37603 = n37599 | n37602 ;
  assign n77641 = ~n37574 ;
  assign n37607 = n77641 & n37603 ;
  assign n37608 = n37606 | n37607 ;
  assign n77642 = ~n37566 ;
  assign n37609 = n77642 & n37608 ;
  assign n77643 = ~n37556 ;
  assign n37610 = x69 & n77643 ;
  assign n77644 = ~n37554 ;
  assign n37611 = n77644 & n37610 ;
  assign n37612 = n37558 | n37611 ;
  assign n37614 = n37609 | n37612 ;
  assign n77645 = ~n37558 ;
  assign n37619 = n77645 & n37614 ;
  assign n37620 = n37617 | n37619 ;
  assign n77646 = ~n37549 ;
  assign n37621 = n77646 & n37620 ;
  assign n77647 = ~n37539 ;
  assign n37622 = x71 & n77647 ;
  assign n77648 = ~n37537 ;
  assign n37623 = n77648 & n37622 ;
  assign n37624 = n37541 | n37623 ;
  assign n37626 = n37621 | n37624 ;
  assign n77649 = ~n37541 ;
  assign n37631 = n77649 & n37626 ;
  assign n37632 = n37629 | n37631 ;
  assign n77650 = ~n37533 ;
  assign n37633 = n77650 & n37632 ;
  assign n77651 = ~n37523 ;
  assign n37634 = x73 & n77651 ;
  assign n77652 = ~n37521 ;
  assign n37635 = n77652 & n37634 ;
  assign n37636 = n37525 | n37635 ;
  assign n37638 = n37633 | n37636 ;
  assign n77653 = ~n37525 ;
  assign n37643 = n77653 & n37638 ;
  assign n37644 = n37641 | n37643 ;
  assign n77654 = ~n37517 ;
  assign n37645 = n77654 & n37644 ;
  assign n77655 = ~n37507 ;
  assign n37646 = x75 & n77655 ;
  assign n77656 = ~n37505 ;
  assign n37647 = n77656 & n37646 ;
  assign n37648 = n37509 | n37647 ;
  assign n37650 = n37645 | n37648 ;
  assign n77657 = ~n37509 ;
  assign n37655 = n77657 & n37650 ;
  assign n37656 = n37653 | n37655 ;
  assign n77658 = ~n37501 ;
  assign n37657 = n77658 & n37656 ;
  assign n77659 = ~n37491 ;
  assign n37658 = x77 & n77659 ;
  assign n77660 = ~n37489 ;
  assign n37659 = n77660 & n37658 ;
  assign n37660 = n37493 | n37659 ;
  assign n37662 = n37657 | n37660 ;
  assign n77661 = ~n37493 ;
  assign n37667 = n77661 & n37662 ;
  assign n37668 = n37665 | n37667 ;
  assign n77662 = ~n37485 ;
  assign n37669 = n77662 & n37668 ;
  assign n77663 = ~n37475 ;
  assign n37670 = x79 & n77663 ;
  assign n77664 = ~n37473 ;
  assign n37671 = n77664 & n37670 ;
  assign n37672 = n37477 | n37671 ;
  assign n37674 = n37669 | n37672 ;
  assign n77665 = ~n37477 ;
  assign n37679 = n77665 & n37674 ;
  assign n37680 = n37677 | n37679 ;
  assign n77666 = ~n37469 ;
  assign n37681 = n77666 & n37680 ;
  assign n77667 = ~n37459 ;
  assign n37682 = x81 & n77667 ;
  assign n77668 = ~n37457 ;
  assign n37683 = n77668 & n37682 ;
  assign n37684 = n37461 | n37683 ;
  assign n37686 = n37681 | n37684 ;
  assign n77669 = ~n37461 ;
  assign n37691 = n77669 & n37686 ;
  assign n37692 = n37689 | n37691 ;
  assign n77670 = ~n37453 ;
  assign n37693 = n77670 & n37692 ;
  assign n77671 = ~n37443 ;
  assign n37694 = x83 & n77671 ;
  assign n77672 = ~n37441 ;
  assign n37695 = n77672 & n37694 ;
  assign n37696 = n37445 | n37695 ;
  assign n37698 = n37693 | n37696 ;
  assign n77673 = ~n37445 ;
  assign n37703 = n77673 & n37698 ;
  assign n37704 = n37701 | n37703 ;
  assign n77674 = ~n37437 ;
  assign n37705 = n77674 & n37704 ;
  assign n77675 = ~n37427 ;
  assign n37706 = x85 & n77675 ;
  assign n77676 = ~n37425 ;
  assign n37707 = n77676 & n37706 ;
  assign n37708 = n37429 | n37707 ;
  assign n37710 = n37705 | n37708 ;
  assign n77677 = ~n37429 ;
  assign n37715 = n77677 & n37710 ;
  assign n37716 = n37713 | n37715 ;
  assign n77678 = ~n37421 ;
  assign n37717 = n77678 & n37716 ;
  assign n77679 = ~n37400 ;
  assign n37718 = x87 & n77679 ;
  assign n77680 = ~n37394 ;
  assign n37719 = n77680 & n37718 ;
  assign n37720 = n37413 | n37719 ;
  assign n37722 = n37717 | n37720 ;
  assign n77681 = ~n37413 ;
  assign n37726 = n77681 & n37722 ;
  assign n37727 = n37725 | n37726 ;
  assign n77682 = ~n37412 ;
  assign n37728 = n77682 & n37727 ;
  assign n37729 = n5320 | n37728 ;
  assign n37732 = n37401 & n37729 ;
  assign n37721 = n37421 | n37720 ;
  assign n37733 = x64 & n77635 ;
  assign n77683 = ~n37733 ;
  assign n37734 = x40 & n77683 ;
  assign n37735 = n37334 | n37734 ;
  assign n37736 = x65 & n37735 ;
  assign n77684 = ~n37736 ;
  assign n37737 = n37589 & n77684 ;
  assign n37738 = n5190 | n37737 ;
  assign n37739 = n77637 & n37738 ;
  assign n37741 = n37596 | n37739 ;
  assign n37742 = n77638 & n37741 ;
  assign n37743 = n37602 | n37742 ;
  assign n37744 = n77641 & n37743 ;
  assign n37745 = n37606 | n37744 ;
  assign n37746 = n77642 & n37745 ;
  assign n37747 = n37612 | n37746 ;
  assign n37748 = n77645 & n37747 ;
  assign n37749 = n37617 | n37748 ;
  assign n37750 = n77646 & n37749 ;
  assign n37751 = n37624 | n37750 ;
  assign n37752 = n77649 & n37751 ;
  assign n37753 = n37629 | n37752 ;
  assign n37754 = n77650 & n37753 ;
  assign n37755 = n37636 | n37754 ;
  assign n37756 = n77653 & n37755 ;
  assign n37757 = n37641 | n37756 ;
  assign n37758 = n77654 & n37757 ;
  assign n37759 = n37648 | n37758 ;
  assign n37760 = n77657 & n37759 ;
  assign n37761 = n37653 | n37760 ;
  assign n37762 = n77658 & n37761 ;
  assign n37763 = n37660 | n37762 ;
  assign n37764 = n77661 & n37763 ;
  assign n37765 = n37665 | n37764 ;
  assign n37766 = n77662 & n37765 ;
  assign n37767 = n37672 | n37766 ;
  assign n37768 = n77665 & n37767 ;
  assign n37769 = n37677 | n37768 ;
  assign n37770 = n77666 & n37769 ;
  assign n37771 = n37684 | n37770 ;
  assign n37772 = n77669 & n37771 ;
  assign n37773 = n37689 | n37772 ;
  assign n37774 = n77670 & n37773 ;
  assign n37775 = n37696 | n37774 ;
  assign n37776 = n77673 & n37775 ;
  assign n37777 = n37701 | n37776 ;
  assign n37778 = n77674 & n37777 ;
  assign n37779 = n37708 | n37778 ;
  assign n37780 = n77677 & n37779 ;
  assign n37781 = n37713 | n37780 ;
  assign n77685 = ~n37721 ;
  assign n37782 = n77685 & n37781 ;
  assign n37783 = n77678 & n37781 ;
  assign n77686 = ~n37783 ;
  assign n37784 = n37720 & n77686 ;
  assign n37785 = n37782 | n37784 ;
  assign n37786 = n67354 & n37785 ;
  assign n77687 = ~n37728 ;
  assign n37787 = n77687 & n37786 ;
  assign n37788 = n37732 | n37787 ;
  assign n77688 = ~n37411 ;
  assign n37730 = n77688 & n37729 ;
  assign n77689 = ~n37726 ;
  assign n37791 = n37725 & n77689 ;
  assign n37789 = n37720 | n37783 ;
  assign n37792 = n37413 | n37725 ;
  assign n77690 = ~n37792 ;
  assign n37793 = n37789 & n77690 ;
  assign n37794 = n37791 | n37793 ;
  assign n37795 = n37729 | n37794 ;
  assign n77691 = ~n37730 ;
  assign n37796 = n77691 & n37795 ;
  assign n37797 = n67348 & n37796 ;
  assign n37798 = n67222 & n37788 ;
  assign n37799 = n37420 & n37729 ;
  assign n37714 = n37429 | n37713 ;
  assign n77692 = ~n37714 ;
  assign n37800 = n37710 & n77692 ;
  assign n77693 = ~n37715 ;
  assign n37801 = n37713 & n77693 ;
  assign n37802 = n37800 | n37801 ;
  assign n37803 = n67354 & n37802 ;
  assign n37804 = n77687 & n37803 ;
  assign n37805 = n37799 | n37804 ;
  assign n37806 = n67164 & n37805 ;
  assign n37807 = n37428 & n37729 ;
  assign n37709 = n37437 | n37708 ;
  assign n77694 = ~n37709 ;
  assign n37808 = n77694 & n37777 ;
  assign n77695 = ~n37778 ;
  assign n37809 = n37708 & n77695 ;
  assign n37810 = n37808 | n37809 ;
  assign n37811 = n67354 & n37810 ;
  assign n37812 = n77687 & n37811 ;
  assign n37813 = n37807 | n37812 ;
  assign n37814 = n66979 & n37813 ;
  assign n37815 = n37436 & n37729 ;
  assign n37702 = n37445 | n37701 ;
  assign n77696 = ~n37702 ;
  assign n37816 = n37698 & n77696 ;
  assign n77697 = ~n37703 ;
  assign n37817 = n37701 & n77697 ;
  assign n37818 = n37816 | n37817 ;
  assign n37819 = n67354 & n37818 ;
  assign n37820 = n77687 & n37819 ;
  assign n37821 = n37815 | n37820 ;
  assign n37822 = n66868 & n37821 ;
  assign n37823 = n37444 & n37729 ;
  assign n37697 = n37453 | n37696 ;
  assign n77698 = ~n37697 ;
  assign n37824 = n77698 & n37773 ;
  assign n77699 = ~n37774 ;
  assign n37825 = n37696 & n77699 ;
  assign n37826 = n37824 | n37825 ;
  assign n37827 = n67354 & n37826 ;
  assign n37828 = n77687 & n37827 ;
  assign n37829 = n37823 | n37828 ;
  assign n37830 = n66797 & n37829 ;
  assign n37831 = n37452 & n37729 ;
  assign n37690 = n37461 | n37689 ;
  assign n77700 = ~n37690 ;
  assign n37832 = n37686 & n77700 ;
  assign n77701 = ~n37691 ;
  assign n37833 = n37689 & n77701 ;
  assign n37834 = n37832 | n37833 ;
  assign n37835 = n67354 & n37834 ;
  assign n37836 = n77687 & n37835 ;
  assign n37837 = n37831 | n37836 ;
  assign n37838 = n66654 & n37837 ;
  assign n37839 = n37460 & n37729 ;
  assign n37685 = n37469 | n37684 ;
  assign n77702 = ~n37685 ;
  assign n37840 = n77702 & n37769 ;
  assign n77703 = ~n37770 ;
  assign n37841 = n37684 & n77703 ;
  assign n37842 = n37840 | n37841 ;
  assign n37843 = n67354 & n37842 ;
  assign n37844 = n77687 & n37843 ;
  assign n37845 = n37839 | n37844 ;
  assign n37846 = n66560 & n37845 ;
  assign n37847 = n37468 & n37729 ;
  assign n37678 = n37477 | n37677 ;
  assign n77704 = ~n37678 ;
  assign n37848 = n37674 & n77704 ;
  assign n77705 = ~n37679 ;
  assign n37849 = n37677 & n77705 ;
  assign n37850 = n37848 | n37849 ;
  assign n37851 = n67354 & n37850 ;
  assign n37852 = n77687 & n37851 ;
  assign n37853 = n37847 | n37852 ;
  assign n37854 = n66505 & n37853 ;
  assign n37855 = n37476 & n37729 ;
  assign n37673 = n37485 | n37672 ;
  assign n77706 = ~n37673 ;
  assign n37856 = n77706 & n37765 ;
  assign n77707 = ~n37766 ;
  assign n37857 = n37672 & n77707 ;
  assign n37858 = n37856 | n37857 ;
  assign n37859 = n67354 & n37858 ;
  assign n37860 = n77687 & n37859 ;
  assign n37861 = n37855 | n37860 ;
  assign n37862 = n66379 & n37861 ;
  assign n37863 = n37484 & n37729 ;
  assign n37666 = n37493 | n37665 ;
  assign n77708 = ~n37666 ;
  assign n37864 = n37662 & n77708 ;
  assign n77709 = ~n37667 ;
  assign n37865 = n37665 & n77709 ;
  assign n37866 = n37864 | n37865 ;
  assign n37867 = n67354 & n37866 ;
  assign n37868 = n77687 & n37867 ;
  assign n37869 = n37863 | n37868 ;
  assign n37870 = n66299 & n37869 ;
  assign n37871 = n37492 & n37729 ;
  assign n37661 = n37501 | n37660 ;
  assign n77710 = ~n37661 ;
  assign n37872 = n77710 & n37761 ;
  assign n77711 = ~n37762 ;
  assign n37873 = n37660 & n77711 ;
  assign n37874 = n37872 | n37873 ;
  assign n37875 = n67354 & n37874 ;
  assign n37876 = n77687 & n37875 ;
  assign n37877 = n37871 | n37876 ;
  assign n37878 = n66244 & n37877 ;
  assign n37879 = n37500 & n37729 ;
  assign n37654 = n37509 | n37653 ;
  assign n77712 = ~n37654 ;
  assign n37880 = n37650 & n77712 ;
  assign n77713 = ~n37655 ;
  assign n37881 = n37653 & n77713 ;
  assign n37882 = n37880 | n37881 ;
  assign n37883 = n67354 & n37882 ;
  assign n37884 = n77687 & n37883 ;
  assign n37885 = n37879 | n37884 ;
  assign n37886 = n66145 & n37885 ;
  assign n37887 = n37508 & n37729 ;
  assign n37649 = n37517 | n37648 ;
  assign n77714 = ~n37649 ;
  assign n37888 = n77714 & n37757 ;
  assign n77715 = ~n37758 ;
  assign n37889 = n37648 & n77715 ;
  assign n37890 = n37888 | n37889 ;
  assign n37891 = n67354 & n37890 ;
  assign n37892 = n77687 & n37891 ;
  assign n37893 = n37887 | n37892 ;
  assign n37894 = n66081 & n37893 ;
  assign n37895 = n37516 & n37729 ;
  assign n37642 = n37525 | n37641 ;
  assign n77716 = ~n37642 ;
  assign n37896 = n37638 & n77716 ;
  assign n77717 = ~n37643 ;
  assign n37897 = n37641 & n77717 ;
  assign n37898 = n37896 | n37897 ;
  assign n37899 = n67354 & n37898 ;
  assign n37900 = n77687 & n37899 ;
  assign n37901 = n37895 | n37900 ;
  assign n37902 = n66043 & n37901 ;
  assign n37903 = n37524 & n37729 ;
  assign n37637 = n37533 | n37636 ;
  assign n77718 = ~n37637 ;
  assign n37904 = n77718 & n37753 ;
  assign n77719 = ~n37754 ;
  assign n37905 = n37636 & n77719 ;
  assign n37906 = n37904 | n37905 ;
  assign n37907 = n67354 & n37906 ;
  assign n37908 = n77687 & n37907 ;
  assign n37909 = n37903 | n37908 ;
  assign n37910 = n65960 & n37909 ;
  assign n37911 = n37532 & n37729 ;
  assign n37630 = n37541 | n37629 ;
  assign n77720 = ~n37630 ;
  assign n37912 = n37626 & n77720 ;
  assign n77721 = ~n37631 ;
  assign n37913 = n37629 & n77721 ;
  assign n37914 = n37912 | n37913 ;
  assign n37915 = n67354 & n37914 ;
  assign n37916 = n77687 & n37915 ;
  assign n37917 = n37911 | n37916 ;
  assign n37918 = n65909 & n37917 ;
  assign n37919 = n37540 & n37729 ;
  assign n37625 = n37549 | n37624 ;
  assign n77722 = ~n37625 ;
  assign n37920 = n77722 & n37749 ;
  assign n77723 = ~n37750 ;
  assign n37921 = n37624 & n77723 ;
  assign n37922 = n37920 | n37921 ;
  assign n37923 = n67354 & n37922 ;
  assign n37924 = n77687 & n37923 ;
  assign n37925 = n37919 | n37924 ;
  assign n37926 = n65877 & n37925 ;
  assign n37927 = n37548 & n37729 ;
  assign n37618 = n37558 | n37617 ;
  assign n77724 = ~n37618 ;
  assign n37928 = n37614 & n77724 ;
  assign n77725 = ~n37619 ;
  assign n37929 = n37617 & n77725 ;
  assign n37930 = n37928 | n37929 ;
  assign n37931 = n67354 & n37930 ;
  assign n37932 = n77687 & n37931 ;
  assign n37933 = n37927 | n37932 ;
  assign n37934 = n65820 & n37933 ;
  assign n37935 = n37557 & n37729 ;
  assign n37613 = n37566 | n37612 ;
  assign n77726 = ~n37613 ;
  assign n37936 = n77726 & n37745 ;
  assign n77727 = ~n37746 ;
  assign n37937 = n37612 & n77727 ;
  assign n37938 = n37936 | n37937 ;
  assign n37939 = n67354 & n37938 ;
  assign n37940 = n77687 & n37939 ;
  assign n37941 = n37935 | n37940 ;
  assign n37942 = n65791 & n37941 ;
  assign n37943 = n37565 & n37729 ;
  assign n37944 = n37574 | n37606 ;
  assign n77728 = ~n37944 ;
  assign n37945 = n37603 & n77728 ;
  assign n77729 = ~n37607 ;
  assign n37946 = n37606 & n77729 ;
  assign n37947 = n37945 | n37946 ;
  assign n37948 = n67354 & n37947 ;
  assign n37949 = n77687 & n37948 ;
  assign n37950 = n37943 | n37949 ;
  assign n37951 = n65772 & n37950 ;
  assign n37952 = n37573 & n37729 ;
  assign n37953 = n37582 | n37602 ;
  assign n77730 = ~n37953 ;
  assign n37954 = n37598 & n77730 ;
  assign n77731 = ~n37742 ;
  assign n37955 = n37602 & n77731 ;
  assign n37956 = n37954 | n37955 ;
  assign n37957 = n67354 & n37956 ;
  assign n37958 = n77687 & n37957 ;
  assign n37959 = n37952 | n37958 ;
  assign n37960 = n65746 & n37959 ;
  assign n37961 = n37581 & n37729 ;
  assign n37740 = n37593 | n37596 ;
  assign n77732 = ~n37740 ;
  assign n37962 = n37738 & n77732 ;
  assign n77733 = ~n37597 ;
  assign n37963 = n37596 & n77733 ;
  assign n37964 = n37962 | n37963 ;
  assign n37965 = n67354 & n37964 ;
  assign n37966 = n77687 & n37965 ;
  assign n37967 = n37961 | n37966 ;
  assign n37968 = n65721 & n37967 ;
  assign n37731 = n37584 & n37729 ;
  assign n37591 = n5190 & n37589 ;
  assign n37970 = n37591 & n77684 ;
  assign n37971 = n5320 | n37970 ;
  assign n77734 = ~n37971 ;
  assign n37972 = n37738 & n77734 ;
  assign n37973 = n77687 & n37972 ;
  assign n37974 = n37731 | n37973 ;
  assign n37975 = n65686 & n37974 ;
  assign n37969 = n5583 & n77687 ;
  assign n37976 = n5577 & n77687 ;
  assign n77735 = ~n37976 ;
  assign n37977 = x39 & n77735 ;
  assign n37978 = n37969 | n37977 ;
  assign n37979 = n65670 & n37978 ;
  assign n37790 = n77681 & n37789 ;
  assign n37981 = n37725 | n37790 ;
  assign n37982 = n77682 & n37981 ;
  assign n77736 = ~n37982 ;
  assign n37983 = n5577 & n77736 ;
  assign n77737 = ~n37983 ;
  assign n37984 = x39 & n77737 ;
  assign n37985 = n37969 | n37984 ;
  assign n37987 = x65 & n37985 ;
  assign n37986 = x65 | n37969 ;
  assign n37988 = n37977 | n37986 ;
  assign n77738 = ~n37987 ;
  assign n37989 = n77738 & n37988 ;
  assign n37990 = n5594 | n37989 ;
  assign n77739 = ~n37979 ;
  assign n37991 = n77739 & n37990 ;
  assign n77740 = ~n37973 ;
  assign n37992 = x66 & n77740 ;
  assign n77741 = ~n37731 ;
  assign n37993 = n77741 & n37992 ;
  assign n37994 = n37975 | n37993 ;
  assign n37995 = n37991 | n37994 ;
  assign n77742 = ~n37975 ;
  assign n37996 = n77742 & n37995 ;
  assign n77743 = ~n37966 ;
  assign n37997 = x67 & n77743 ;
  assign n77744 = ~n37961 ;
  assign n37998 = n77744 & n37997 ;
  assign n37999 = n37996 | n37998 ;
  assign n77745 = ~n37968 ;
  assign n38000 = n77745 & n37999 ;
  assign n77746 = ~n37958 ;
  assign n38001 = x68 & n77746 ;
  assign n77747 = ~n37952 ;
  assign n38002 = n77747 & n38001 ;
  assign n38003 = n37960 | n38002 ;
  assign n38004 = n38000 | n38003 ;
  assign n77748 = ~n37960 ;
  assign n38005 = n77748 & n38004 ;
  assign n77749 = ~n37949 ;
  assign n38006 = x69 & n77749 ;
  assign n77750 = ~n37943 ;
  assign n38007 = n77750 & n38006 ;
  assign n38008 = n37951 | n38007 ;
  assign n38009 = n38005 | n38008 ;
  assign n77751 = ~n37951 ;
  assign n38010 = n77751 & n38009 ;
  assign n77752 = ~n37940 ;
  assign n38011 = x70 & n77752 ;
  assign n77753 = ~n37935 ;
  assign n38012 = n77753 & n38011 ;
  assign n38013 = n37942 | n38012 ;
  assign n38014 = n38010 | n38013 ;
  assign n77754 = ~n37942 ;
  assign n38015 = n77754 & n38014 ;
  assign n77755 = ~n37932 ;
  assign n38016 = x71 & n77755 ;
  assign n77756 = ~n37927 ;
  assign n38017 = n77756 & n38016 ;
  assign n38018 = n37934 | n38017 ;
  assign n38020 = n38015 | n38018 ;
  assign n77757 = ~n37934 ;
  assign n38021 = n77757 & n38020 ;
  assign n77758 = ~n37924 ;
  assign n38022 = x72 & n77758 ;
  assign n77759 = ~n37919 ;
  assign n38023 = n77759 & n38022 ;
  assign n38024 = n37926 | n38023 ;
  assign n38025 = n38021 | n38024 ;
  assign n77760 = ~n37926 ;
  assign n38026 = n77760 & n38025 ;
  assign n77761 = ~n37916 ;
  assign n38027 = x73 & n77761 ;
  assign n77762 = ~n37911 ;
  assign n38028 = n77762 & n38027 ;
  assign n38029 = n37918 | n38028 ;
  assign n38031 = n38026 | n38029 ;
  assign n77763 = ~n37918 ;
  assign n38032 = n77763 & n38031 ;
  assign n77764 = ~n37908 ;
  assign n38033 = x74 & n77764 ;
  assign n77765 = ~n37903 ;
  assign n38034 = n77765 & n38033 ;
  assign n38035 = n37910 | n38034 ;
  assign n38036 = n38032 | n38035 ;
  assign n77766 = ~n37910 ;
  assign n38037 = n77766 & n38036 ;
  assign n77767 = ~n37900 ;
  assign n38038 = x75 & n77767 ;
  assign n77768 = ~n37895 ;
  assign n38039 = n77768 & n38038 ;
  assign n38040 = n37902 | n38039 ;
  assign n38042 = n38037 | n38040 ;
  assign n77769 = ~n37902 ;
  assign n38043 = n77769 & n38042 ;
  assign n77770 = ~n37892 ;
  assign n38044 = x76 & n77770 ;
  assign n77771 = ~n37887 ;
  assign n38045 = n77771 & n38044 ;
  assign n38046 = n37894 | n38045 ;
  assign n38047 = n38043 | n38046 ;
  assign n77772 = ~n37894 ;
  assign n38048 = n77772 & n38047 ;
  assign n77773 = ~n37884 ;
  assign n38049 = x77 & n77773 ;
  assign n77774 = ~n37879 ;
  assign n38050 = n77774 & n38049 ;
  assign n38051 = n37886 | n38050 ;
  assign n38053 = n38048 | n38051 ;
  assign n77775 = ~n37886 ;
  assign n38054 = n77775 & n38053 ;
  assign n77776 = ~n37876 ;
  assign n38055 = x78 & n77776 ;
  assign n77777 = ~n37871 ;
  assign n38056 = n77777 & n38055 ;
  assign n38057 = n37878 | n38056 ;
  assign n38058 = n38054 | n38057 ;
  assign n77778 = ~n37878 ;
  assign n38059 = n77778 & n38058 ;
  assign n77779 = ~n37868 ;
  assign n38060 = x79 & n77779 ;
  assign n77780 = ~n37863 ;
  assign n38061 = n77780 & n38060 ;
  assign n38062 = n37870 | n38061 ;
  assign n38064 = n38059 | n38062 ;
  assign n77781 = ~n37870 ;
  assign n38065 = n77781 & n38064 ;
  assign n77782 = ~n37860 ;
  assign n38066 = x80 & n77782 ;
  assign n77783 = ~n37855 ;
  assign n38067 = n77783 & n38066 ;
  assign n38068 = n37862 | n38067 ;
  assign n38069 = n38065 | n38068 ;
  assign n77784 = ~n37862 ;
  assign n38070 = n77784 & n38069 ;
  assign n77785 = ~n37852 ;
  assign n38071 = x81 & n77785 ;
  assign n77786 = ~n37847 ;
  assign n38072 = n77786 & n38071 ;
  assign n38073 = n37854 | n38072 ;
  assign n38075 = n38070 | n38073 ;
  assign n77787 = ~n37854 ;
  assign n38076 = n77787 & n38075 ;
  assign n77788 = ~n37844 ;
  assign n38077 = x82 & n77788 ;
  assign n77789 = ~n37839 ;
  assign n38078 = n77789 & n38077 ;
  assign n38079 = n37846 | n38078 ;
  assign n38080 = n38076 | n38079 ;
  assign n77790 = ~n37846 ;
  assign n38081 = n77790 & n38080 ;
  assign n77791 = ~n37836 ;
  assign n38082 = x83 & n77791 ;
  assign n77792 = ~n37831 ;
  assign n38083 = n77792 & n38082 ;
  assign n38084 = n37838 | n38083 ;
  assign n38086 = n38081 | n38084 ;
  assign n77793 = ~n37838 ;
  assign n38087 = n77793 & n38086 ;
  assign n77794 = ~n37828 ;
  assign n38088 = x84 & n77794 ;
  assign n77795 = ~n37823 ;
  assign n38089 = n77795 & n38088 ;
  assign n38090 = n37830 | n38089 ;
  assign n38091 = n38087 | n38090 ;
  assign n77796 = ~n37830 ;
  assign n38092 = n77796 & n38091 ;
  assign n77797 = ~n37820 ;
  assign n38093 = x85 & n77797 ;
  assign n77798 = ~n37815 ;
  assign n38094 = n77798 & n38093 ;
  assign n38095 = n37822 | n38094 ;
  assign n38097 = n38092 | n38095 ;
  assign n77799 = ~n37822 ;
  assign n38098 = n77799 & n38097 ;
  assign n77800 = ~n37812 ;
  assign n38099 = x86 & n77800 ;
  assign n77801 = ~n37807 ;
  assign n38100 = n77801 & n38099 ;
  assign n38101 = n37814 | n38100 ;
  assign n38102 = n38098 | n38101 ;
  assign n77802 = ~n37814 ;
  assign n38103 = n77802 & n38102 ;
  assign n77803 = ~n37804 ;
  assign n38104 = x87 & n77803 ;
  assign n77804 = ~n37799 ;
  assign n38105 = n77804 & n38104 ;
  assign n38106 = n37806 | n38105 ;
  assign n38108 = n38103 | n38106 ;
  assign n77805 = ~n37806 ;
  assign n38109 = n77805 & n38108 ;
  assign n77806 = ~n37787 ;
  assign n38110 = x88 & n77806 ;
  assign n77807 = ~n37732 ;
  assign n38111 = n77807 & n38110 ;
  assign n38112 = n37798 | n38111 ;
  assign n38113 = n38109 | n38112 ;
  assign n77808 = ~n37798 ;
  assign n38114 = n77808 & n38113 ;
  assign n77809 = ~n37729 ;
  assign n38115 = n77809 & n37794 ;
  assign n38116 = n37411 & n37729 ;
  assign n77810 = ~n38116 ;
  assign n38117 = x89 & n77810 ;
  assign n77811 = ~n38115 ;
  assign n38118 = n77811 & n38117 ;
  assign n38119 = n37797 | n38118 ;
  assign n38121 = n38114 | n38119 ;
  assign n77812 = ~n37797 ;
  assign n38122 = n77812 & n38121 ;
  assign n38123 = n5743 | n38122 ;
  assign n38124 = n37788 & n38123 ;
  assign n38126 = n65670 & n37985 ;
  assign n37980 = x65 & n37978 ;
  assign n77813 = ~n37980 ;
  assign n38125 = n77813 & n37988 ;
  assign n38127 = n5594 | n38125 ;
  assign n77814 = ~n38126 ;
  assign n38128 = n77814 & n38127 ;
  assign n38129 = n37994 | n38128 ;
  assign n38130 = n77742 & n38129 ;
  assign n38131 = n37968 | n37998 ;
  assign n38133 = n38130 | n38131 ;
  assign n38134 = n77745 & n38133 ;
  assign n38136 = n38003 | n38134 ;
  assign n38137 = n77748 & n38136 ;
  assign n38139 = n38008 | n38137 ;
  assign n38140 = n77751 & n38139 ;
  assign n38141 = n38013 | n38140 ;
  assign n38143 = n77754 & n38141 ;
  assign n38144 = n38018 | n38143 ;
  assign n38145 = n77757 & n38144 ;
  assign n38146 = n38024 | n38145 ;
  assign n38148 = n77760 & n38146 ;
  assign n38149 = n38029 | n38148 ;
  assign n38150 = n77763 & n38149 ;
  assign n38151 = n38035 | n38150 ;
  assign n38153 = n77766 & n38151 ;
  assign n38154 = n38040 | n38153 ;
  assign n38155 = n77769 & n38154 ;
  assign n38156 = n38046 | n38155 ;
  assign n38158 = n77772 & n38156 ;
  assign n38159 = n38051 | n38158 ;
  assign n38160 = n77775 & n38159 ;
  assign n38161 = n38057 | n38160 ;
  assign n38163 = n77778 & n38161 ;
  assign n38164 = n38062 | n38163 ;
  assign n38165 = n77781 & n38164 ;
  assign n38166 = n38068 | n38165 ;
  assign n38168 = n77784 & n38166 ;
  assign n38169 = n38073 | n38168 ;
  assign n38170 = n77787 & n38169 ;
  assign n38171 = n38079 | n38170 ;
  assign n38173 = n77790 & n38171 ;
  assign n38174 = n38084 | n38173 ;
  assign n38175 = n77793 & n38174 ;
  assign n38176 = n38090 | n38175 ;
  assign n38178 = n77796 & n38176 ;
  assign n38179 = n38095 | n38178 ;
  assign n38180 = n77799 & n38179 ;
  assign n38181 = n38101 | n38180 ;
  assign n38183 = n77802 & n38181 ;
  assign n38184 = n38106 | n38183 ;
  assign n38185 = n77805 & n38184 ;
  assign n77815 = ~n38185 ;
  assign n38186 = n38112 & n77815 ;
  assign n38188 = n37806 | n38112 ;
  assign n77816 = ~n38188 ;
  assign n38189 = n38108 & n77816 ;
  assign n38190 = n38186 | n38189 ;
  assign n38191 = n67482 & n38190 ;
  assign n77817 = ~n38122 ;
  assign n38192 = n77817 & n38191 ;
  assign n38193 = n38124 | n38192 ;
  assign n38194 = n67348 & n38193 ;
  assign n77818 = ~n38192 ;
  assign n38516 = x89 & n77818 ;
  assign n77819 = ~n38124 ;
  assign n38517 = n77819 & n38516 ;
  assign n38518 = n38194 | n38517 ;
  assign n38195 = n37805 & n38123 ;
  assign n77820 = ~n38103 ;
  assign n38107 = n77820 & n38106 ;
  assign n38196 = n37814 | n38106 ;
  assign n77821 = ~n38196 ;
  assign n38197 = n38181 & n77821 ;
  assign n38198 = n38107 | n38197 ;
  assign n38199 = n67482 & n38198 ;
  assign n38200 = n77817 & n38199 ;
  assign n38201 = n38195 | n38200 ;
  assign n38202 = n67222 & n38201 ;
  assign n38203 = n37813 & n38123 ;
  assign n77822 = ~n38180 ;
  assign n38182 = n38101 & n77822 ;
  assign n38204 = n37822 | n38101 ;
  assign n77823 = ~n38204 ;
  assign n38205 = n38097 & n77823 ;
  assign n38206 = n38182 | n38205 ;
  assign n38207 = n67482 & n38206 ;
  assign n38208 = n77817 & n38207 ;
  assign n38209 = n38203 | n38208 ;
  assign n38210 = n67164 & n38209 ;
  assign n77824 = ~n38208 ;
  assign n38506 = x87 & n77824 ;
  assign n77825 = ~n38203 ;
  assign n38507 = n77825 & n38506 ;
  assign n38508 = n38210 | n38507 ;
  assign n38211 = n37821 & n38123 ;
  assign n77826 = ~n38092 ;
  assign n38096 = n77826 & n38095 ;
  assign n38212 = n37830 | n38095 ;
  assign n77827 = ~n38212 ;
  assign n38213 = n38176 & n77827 ;
  assign n38214 = n38096 | n38213 ;
  assign n38215 = n67482 & n38214 ;
  assign n38216 = n77817 & n38215 ;
  assign n38217 = n38211 | n38216 ;
  assign n38218 = n66979 & n38217 ;
  assign n38219 = n37829 & n38123 ;
  assign n77828 = ~n38175 ;
  assign n38177 = n38090 & n77828 ;
  assign n38220 = n37838 | n38090 ;
  assign n77829 = ~n38220 ;
  assign n38221 = n38086 & n77829 ;
  assign n38222 = n38177 | n38221 ;
  assign n38223 = n67482 & n38222 ;
  assign n38224 = n77817 & n38223 ;
  assign n38225 = n38219 | n38224 ;
  assign n38226 = n66868 & n38225 ;
  assign n77830 = ~n38224 ;
  assign n38496 = x85 & n77830 ;
  assign n77831 = ~n38219 ;
  assign n38497 = n77831 & n38496 ;
  assign n38498 = n38226 | n38497 ;
  assign n38227 = n37837 & n38123 ;
  assign n77832 = ~n38081 ;
  assign n38085 = n77832 & n38084 ;
  assign n38228 = n37846 | n38084 ;
  assign n77833 = ~n38228 ;
  assign n38229 = n38171 & n77833 ;
  assign n38230 = n38085 | n38229 ;
  assign n38231 = n67482 & n38230 ;
  assign n38232 = n77817 & n38231 ;
  assign n38233 = n38227 | n38232 ;
  assign n38234 = n66797 & n38233 ;
  assign n38235 = n37845 & n38123 ;
  assign n77834 = ~n38170 ;
  assign n38172 = n38079 & n77834 ;
  assign n38236 = n37854 | n38079 ;
  assign n77835 = ~n38236 ;
  assign n38237 = n38075 & n77835 ;
  assign n38238 = n38172 | n38237 ;
  assign n38239 = n67482 & n38238 ;
  assign n38240 = n77817 & n38239 ;
  assign n38241 = n38235 | n38240 ;
  assign n38242 = n66654 & n38241 ;
  assign n77836 = ~n38240 ;
  assign n38486 = x83 & n77836 ;
  assign n77837 = ~n38235 ;
  assign n38487 = n77837 & n38486 ;
  assign n38488 = n38242 | n38487 ;
  assign n38243 = n37853 & n38123 ;
  assign n77838 = ~n38070 ;
  assign n38074 = n77838 & n38073 ;
  assign n38244 = n37862 | n38073 ;
  assign n77839 = ~n38244 ;
  assign n38245 = n38166 & n77839 ;
  assign n38246 = n38074 | n38245 ;
  assign n38247 = n67482 & n38246 ;
  assign n38248 = n77817 & n38247 ;
  assign n38249 = n38243 | n38248 ;
  assign n38250 = n66560 & n38249 ;
  assign n38251 = n37861 & n38123 ;
  assign n77840 = ~n38165 ;
  assign n38167 = n38068 & n77840 ;
  assign n38252 = n37870 | n38068 ;
  assign n77841 = ~n38252 ;
  assign n38253 = n38064 & n77841 ;
  assign n38254 = n38167 | n38253 ;
  assign n38255 = n67482 & n38254 ;
  assign n38256 = n77817 & n38255 ;
  assign n38257 = n38251 | n38256 ;
  assign n38258 = n66505 & n38257 ;
  assign n77842 = ~n38256 ;
  assign n38476 = x81 & n77842 ;
  assign n77843 = ~n38251 ;
  assign n38477 = n77843 & n38476 ;
  assign n38478 = n38258 | n38477 ;
  assign n38259 = n37869 & n38123 ;
  assign n77844 = ~n38059 ;
  assign n38063 = n77844 & n38062 ;
  assign n38260 = n37878 | n38062 ;
  assign n77845 = ~n38260 ;
  assign n38261 = n38161 & n77845 ;
  assign n38262 = n38063 | n38261 ;
  assign n38263 = n67482 & n38262 ;
  assign n38264 = n77817 & n38263 ;
  assign n38265 = n38259 | n38264 ;
  assign n38266 = n66379 & n38265 ;
  assign n38267 = n37877 & n38123 ;
  assign n77846 = ~n38160 ;
  assign n38162 = n38057 & n77846 ;
  assign n38268 = n37886 | n38057 ;
  assign n77847 = ~n38268 ;
  assign n38269 = n38053 & n77847 ;
  assign n38270 = n38162 | n38269 ;
  assign n38271 = n67482 & n38270 ;
  assign n38272 = n77817 & n38271 ;
  assign n38273 = n38267 | n38272 ;
  assign n38274 = n66299 & n38273 ;
  assign n77848 = ~n38272 ;
  assign n38466 = x79 & n77848 ;
  assign n77849 = ~n38267 ;
  assign n38467 = n77849 & n38466 ;
  assign n38468 = n38274 | n38467 ;
  assign n38275 = n37885 & n38123 ;
  assign n77850 = ~n38048 ;
  assign n38052 = n77850 & n38051 ;
  assign n38276 = n37894 | n38051 ;
  assign n77851 = ~n38276 ;
  assign n38277 = n38156 & n77851 ;
  assign n38278 = n38052 | n38277 ;
  assign n38279 = n67482 & n38278 ;
  assign n38280 = n77817 & n38279 ;
  assign n38281 = n38275 | n38280 ;
  assign n38282 = n66244 & n38281 ;
  assign n38283 = n37893 & n38123 ;
  assign n77852 = ~n38155 ;
  assign n38157 = n38046 & n77852 ;
  assign n38284 = n37902 | n38046 ;
  assign n77853 = ~n38284 ;
  assign n38285 = n38042 & n77853 ;
  assign n38286 = n38157 | n38285 ;
  assign n38287 = n67482 & n38286 ;
  assign n38288 = n77817 & n38287 ;
  assign n38289 = n38283 | n38288 ;
  assign n38290 = n66145 & n38289 ;
  assign n77854 = ~n38288 ;
  assign n38455 = x77 & n77854 ;
  assign n77855 = ~n38283 ;
  assign n38456 = n77855 & n38455 ;
  assign n38457 = n38290 | n38456 ;
  assign n38291 = n37901 & n38123 ;
  assign n77856 = ~n38037 ;
  assign n38041 = n77856 & n38040 ;
  assign n38292 = n37910 | n38040 ;
  assign n77857 = ~n38292 ;
  assign n38293 = n38151 & n77857 ;
  assign n38294 = n38041 | n38293 ;
  assign n38295 = n67482 & n38294 ;
  assign n38296 = n77817 & n38295 ;
  assign n38297 = n38291 | n38296 ;
  assign n38298 = n66081 & n38297 ;
  assign n38299 = n37909 & n38123 ;
  assign n77858 = ~n38150 ;
  assign n38152 = n38035 & n77858 ;
  assign n38300 = n37918 | n38035 ;
  assign n77859 = ~n38300 ;
  assign n38301 = n38031 & n77859 ;
  assign n38302 = n38152 | n38301 ;
  assign n38303 = n67482 & n38302 ;
  assign n38304 = n77817 & n38303 ;
  assign n38305 = n38299 | n38304 ;
  assign n38306 = n66043 & n38305 ;
  assign n77860 = ~n38304 ;
  assign n38445 = x75 & n77860 ;
  assign n77861 = ~n38299 ;
  assign n38446 = n77861 & n38445 ;
  assign n38447 = n38306 | n38446 ;
  assign n38307 = n37917 & n38123 ;
  assign n77862 = ~n38026 ;
  assign n38030 = n77862 & n38029 ;
  assign n38308 = n37926 | n38029 ;
  assign n77863 = ~n38308 ;
  assign n38309 = n38146 & n77863 ;
  assign n38310 = n38030 | n38309 ;
  assign n38311 = n67482 & n38310 ;
  assign n38312 = n77817 & n38311 ;
  assign n38313 = n38307 | n38312 ;
  assign n38314 = n65960 & n38313 ;
  assign n38315 = n37925 & n38123 ;
  assign n77864 = ~n38145 ;
  assign n38147 = n38024 & n77864 ;
  assign n38316 = n37934 | n38024 ;
  assign n77865 = ~n38316 ;
  assign n38317 = n38020 & n77865 ;
  assign n38318 = n38147 | n38317 ;
  assign n38319 = n67482 & n38318 ;
  assign n38320 = n77817 & n38319 ;
  assign n38321 = n38315 | n38320 ;
  assign n38322 = n65909 & n38321 ;
  assign n77866 = ~n38320 ;
  assign n38434 = x73 & n77866 ;
  assign n77867 = ~n38315 ;
  assign n38435 = n77867 & n38434 ;
  assign n38436 = n38322 | n38435 ;
  assign n38323 = n37933 & n38123 ;
  assign n77868 = ~n38015 ;
  assign n38019 = n77868 & n38018 ;
  assign n38324 = n37942 | n38018 ;
  assign n77869 = ~n38324 ;
  assign n38325 = n38141 & n77869 ;
  assign n38326 = n38019 | n38325 ;
  assign n38327 = n67482 & n38326 ;
  assign n38328 = n77817 & n38327 ;
  assign n38329 = n38323 | n38328 ;
  assign n38330 = n65877 & n38329 ;
  assign n38331 = n37941 & n38123 ;
  assign n77870 = ~n38140 ;
  assign n38142 = n38013 & n77870 ;
  assign n38332 = n37951 | n38013 ;
  assign n77871 = ~n38332 ;
  assign n38333 = n38009 & n77871 ;
  assign n38334 = n38142 | n38333 ;
  assign n38335 = n67482 & n38334 ;
  assign n38336 = n77817 & n38335 ;
  assign n38337 = n38331 | n38336 ;
  assign n38338 = n65820 & n38337 ;
  assign n77872 = ~n38336 ;
  assign n38423 = x71 & n77872 ;
  assign n77873 = ~n38331 ;
  assign n38424 = n77873 & n38423 ;
  assign n38425 = n38338 | n38424 ;
  assign n38339 = n37950 & n38123 ;
  assign n77874 = ~n38005 ;
  assign n38138 = n77874 & n38008 ;
  assign n38340 = n37960 | n38008 ;
  assign n77875 = ~n38340 ;
  assign n38341 = n38004 & n77875 ;
  assign n38342 = n38138 | n38341 ;
  assign n38343 = n67482 & n38342 ;
  assign n38344 = n77817 & n38343 ;
  assign n38345 = n38339 | n38344 ;
  assign n38346 = n65791 & n38345 ;
  assign n38347 = n37959 & n38123 ;
  assign n77876 = ~n38134 ;
  assign n38135 = n38003 & n77876 ;
  assign n38348 = n37996 | n38131 ;
  assign n38349 = n37968 | n38003 ;
  assign n77877 = ~n38349 ;
  assign n38350 = n38348 & n77877 ;
  assign n38351 = n38135 | n38350 ;
  assign n38352 = n67482 & n38351 ;
  assign n38353 = n77817 & n38352 ;
  assign n38354 = n38347 | n38353 ;
  assign n38355 = n65772 & n38354 ;
  assign n77878 = ~n38353 ;
  assign n38412 = x69 & n77878 ;
  assign n77879 = ~n38347 ;
  assign n38413 = n77879 & n38412 ;
  assign n38414 = n38355 | n38413 ;
  assign n38356 = n37967 & n38123 ;
  assign n77880 = ~n37996 ;
  assign n38132 = n77880 & n38131 ;
  assign n38357 = n37975 | n38131 ;
  assign n77881 = ~n38357 ;
  assign n38358 = n37995 & n77881 ;
  assign n38359 = n38132 | n38358 ;
  assign n38360 = n67482 & n38359 ;
  assign n38361 = n77817 & n38360 ;
  assign n38362 = n38356 | n38361 ;
  assign n38363 = n65746 & n38362 ;
  assign n38364 = n37974 & n38123 ;
  assign n38365 = n37994 | n38126 ;
  assign n77882 = ~n38365 ;
  assign n38366 = n38127 & n77882 ;
  assign n77883 = ~n38128 ;
  assign n38367 = n37994 & n77883 ;
  assign n38368 = n38366 | n38367 ;
  assign n38369 = n67482 & n38368 ;
  assign n38370 = n77817 & n38369 ;
  assign n38371 = n38364 | n38370 ;
  assign n38373 = n65721 & n38371 ;
  assign n77884 = ~n38370 ;
  assign n38372 = x67 & n77884 ;
  assign n77885 = ~n38364 ;
  assign n38403 = n77885 & n38372 ;
  assign n38404 = n38373 | n38403 ;
  assign n38374 = n37978 & n38123 ;
  assign n38375 = n5594 & n37988 ;
  assign n38376 = n77738 & n38375 ;
  assign n38377 = n5743 | n38376 ;
  assign n77886 = ~n38377 ;
  assign n38378 = n38127 & n77886 ;
  assign n38379 = n77817 & n38378 ;
  assign n38380 = n38374 | n38379 ;
  assign n38381 = n65686 & n38380 ;
  assign n38382 = n5994 & n77817 ;
  assign n77887 = ~n38382 ;
  assign n38383 = x38 & n77887 ;
  assign n38384 = n6006 & n77817 ;
  assign n38385 = n38383 | n38384 ;
  assign n38386 = x65 & n38385 ;
  assign n38187 = n38112 | n38185 ;
  assign n38387 = n77808 & n38187 ;
  assign n38388 = n38119 | n38387 ;
  assign n38389 = n77812 & n38388 ;
  assign n77888 = ~n38389 ;
  assign n38390 = n5994 & n77888 ;
  assign n77889 = ~n38390 ;
  assign n38391 = x38 & n77889 ;
  assign n38392 = x65 | n38384 ;
  assign n38393 = n38391 | n38392 ;
  assign n77890 = ~n38386 ;
  assign n38394 = n77890 & n38393 ;
  assign n38395 = n6013 | n38394 ;
  assign n38396 = n38384 | n38391 ;
  assign n38397 = n65670 & n38396 ;
  assign n77891 = ~n38397 ;
  assign n38398 = n38395 & n77891 ;
  assign n77892 = ~n38379 ;
  assign n38399 = x66 & n77892 ;
  assign n77893 = ~n38374 ;
  assign n38400 = n77893 & n38399 ;
  assign n38401 = n38381 | n38400 ;
  assign n38402 = n38398 | n38401 ;
  assign n77894 = ~n38381 ;
  assign n38405 = n77894 & n38402 ;
  assign n38406 = n38404 | n38405 ;
  assign n77895 = ~n38373 ;
  assign n38407 = n77895 & n38406 ;
  assign n77896 = ~n38361 ;
  assign n38408 = x68 & n77896 ;
  assign n77897 = ~n38356 ;
  assign n38409 = n77897 & n38408 ;
  assign n38410 = n38363 | n38409 ;
  assign n38411 = n38407 | n38410 ;
  assign n77898 = ~n38363 ;
  assign n38415 = n77898 & n38411 ;
  assign n38416 = n38414 | n38415 ;
  assign n77899 = ~n38355 ;
  assign n38417 = n77899 & n38416 ;
  assign n77900 = ~n38344 ;
  assign n38418 = x70 & n77900 ;
  assign n77901 = ~n38339 ;
  assign n38419 = n77901 & n38418 ;
  assign n38420 = n38346 | n38419 ;
  assign n38422 = n38417 | n38420 ;
  assign n77902 = ~n38346 ;
  assign n38427 = n77902 & n38422 ;
  assign n38428 = n38425 | n38427 ;
  assign n77903 = ~n38338 ;
  assign n38429 = n77903 & n38428 ;
  assign n77904 = ~n38328 ;
  assign n38430 = x72 & n77904 ;
  assign n77905 = ~n38323 ;
  assign n38431 = n77905 & n38430 ;
  assign n38432 = n38330 | n38431 ;
  assign n38433 = n38429 | n38432 ;
  assign n77906 = ~n38330 ;
  assign n38437 = n77906 & n38433 ;
  assign n38438 = n38436 | n38437 ;
  assign n77907 = ~n38322 ;
  assign n38439 = n77907 & n38438 ;
  assign n77908 = ~n38312 ;
  assign n38440 = x74 & n77908 ;
  assign n77909 = ~n38307 ;
  assign n38441 = n77909 & n38440 ;
  assign n38442 = n38314 | n38441 ;
  assign n38444 = n38439 | n38442 ;
  assign n77910 = ~n38314 ;
  assign n38448 = n77910 & n38444 ;
  assign n38449 = n38447 | n38448 ;
  assign n77911 = ~n38306 ;
  assign n38450 = n77911 & n38449 ;
  assign n77912 = ~n38296 ;
  assign n38451 = x76 & n77912 ;
  assign n77913 = ~n38291 ;
  assign n38452 = n77913 & n38451 ;
  assign n38453 = n38298 | n38452 ;
  assign n38454 = n38450 | n38453 ;
  assign n77914 = ~n38298 ;
  assign n38459 = n77914 & n38454 ;
  assign n38460 = n38457 | n38459 ;
  assign n77915 = ~n38290 ;
  assign n38461 = n77915 & n38460 ;
  assign n77916 = ~n38280 ;
  assign n38462 = x78 & n77916 ;
  assign n77917 = ~n38275 ;
  assign n38463 = n77917 & n38462 ;
  assign n38464 = n38282 | n38463 ;
  assign n38465 = n38461 | n38464 ;
  assign n77918 = ~n38282 ;
  assign n38469 = n77918 & n38465 ;
  assign n38470 = n38468 | n38469 ;
  assign n77919 = ~n38274 ;
  assign n38471 = n77919 & n38470 ;
  assign n77920 = ~n38264 ;
  assign n38472 = x80 & n77920 ;
  assign n77921 = ~n38259 ;
  assign n38473 = n77921 & n38472 ;
  assign n38474 = n38266 | n38473 ;
  assign n38475 = n38471 | n38474 ;
  assign n77922 = ~n38266 ;
  assign n38479 = n77922 & n38475 ;
  assign n38480 = n38478 | n38479 ;
  assign n77923 = ~n38258 ;
  assign n38481 = n77923 & n38480 ;
  assign n77924 = ~n38248 ;
  assign n38482 = x82 & n77924 ;
  assign n77925 = ~n38243 ;
  assign n38483 = n77925 & n38482 ;
  assign n38484 = n38250 | n38483 ;
  assign n38485 = n38481 | n38484 ;
  assign n77926 = ~n38250 ;
  assign n38489 = n77926 & n38485 ;
  assign n38490 = n38488 | n38489 ;
  assign n77927 = ~n38242 ;
  assign n38491 = n77927 & n38490 ;
  assign n77928 = ~n38232 ;
  assign n38492 = x84 & n77928 ;
  assign n77929 = ~n38227 ;
  assign n38493 = n77929 & n38492 ;
  assign n38494 = n38234 | n38493 ;
  assign n38495 = n38491 | n38494 ;
  assign n77930 = ~n38234 ;
  assign n38499 = n77930 & n38495 ;
  assign n38500 = n38498 | n38499 ;
  assign n77931 = ~n38226 ;
  assign n38501 = n77931 & n38500 ;
  assign n77932 = ~n38216 ;
  assign n38502 = x86 & n77932 ;
  assign n77933 = ~n38211 ;
  assign n38503 = n77933 & n38502 ;
  assign n38504 = n38218 | n38503 ;
  assign n38505 = n38501 | n38504 ;
  assign n77934 = ~n38218 ;
  assign n38509 = n77934 & n38505 ;
  assign n38510 = n38508 | n38509 ;
  assign n77935 = ~n38210 ;
  assign n38511 = n77935 & n38510 ;
  assign n77936 = ~n38200 ;
  assign n38512 = x88 & n77936 ;
  assign n77937 = ~n38195 ;
  assign n38513 = n77937 & n38512 ;
  assign n38514 = n38202 | n38513 ;
  assign n38515 = n38511 | n38514 ;
  assign n77938 = ~n38202 ;
  assign n38519 = n77938 & n38515 ;
  assign n38520 = n38518 | n38519 ;
  assign n77939 = ~n38194 ;
  assign n38521 = n77939 & n38520 ;
  assign n77940 = ~n38114 ;
  assign n38120 = n77940 & n38119 ;
  assign n38522 = n37798 | n38119 ;
  assign n77941 = ~n38522 ;
  assign n38523 = n38187 & n77941 ;
  assign n38524 = n38120 | n38523 ;
  assign n38525 = n38123 | n38524 ;
  assign n77942 = ~n37796 ;
  assign n38526 = n77942 & n38123 ;
  assign n77943 = ~n38526 ;
  assign n38527 = n38525 & n77943 ;
  assign n38528 = n67531 & n38527 ;
  assign n77944 = ~n38123 ;
  assign n38529 = n77944 & n38524 ;
  assign n38530 = n37796 & n38123 ;
  assign n77945 = ~n38530 ;
  assign n38531 = x90 & n77945 ;
  assign n77946 = ~n38529 ;
  assign n38532 = n77946 & n38531 ;
  assign n38533 = n6159 | n38532 ;
  assign n38534 = n38528 | n38533 ;
  assign n38535 = n38521 | n38534 ;
  assign n38536 = n67482 & n38527 ;
  assign n77947 = ~n38536 ;
  assign n38537 = n38535 & n77947 ;
  assign n38597 = n38194 | n38532 ;
  assign n38598 = n38528 | n38597 ;
  assign n77948 = ~n38598 ;
  assign n38599 = n38520 & n77948 ;
  assign n38600 = n38528 | n38532 ;
  assign n77949 = ~n38521 ;
  assign n38601 = n77949 & n38600 ;
  assign n38602 = n38599 | n38601 ;
  assign n77950 = ~n38537 ;
  assign n38603 = n77950 & n38602 ;
  assign n38604 = n5743 & n37796 ;
  assign n38605 = n38535 & n38604 ;
  assign n38606 = n38603 | n38605 ;
  assign n38607 = n67622 & n38606 ;
  assign n77951 = ~n38519 ;
  assign n38589 = n38518 & n77951 ;
  assign n38539 = x65 & n38396 ;
  assign n77952 = ~n38539 ;
  assign n38540 = n38393 & n77952 ;
  assign n38541 = n6013 | n38540 ;
  assign n38542 = n77891 & n38541 ;
  assign n38543 = n38401 | n38542 ;
  assign n38544 = n77894 & n38543 ;
  assign n38545 = n38404 | n38544 ;
  assign n38546 = n77895 & n38545 ;
  assign n38547 = n38410 | n38546 ;
  assign n38548 = n77898 & n38547 ;
  assign n38549 = n38414 | n38548 ;
  assign n38550 = n77899 & n38549 ;
  assign n38551 = n38420 | n38550 ;
  assign n38552 = n77902 & n38551 ;
  assign n38553 = n38425 | n38552 ;
  assign n38554 = n77903 & n38553 ;
  assign n38555 = n38432 | n38554 ;
  assign n38556 = n77906 & n38555 ;
  assign n38557 = n38436 | n38556 ;
  assign n38558 = n77907 & n38557 ;
  assign n38559 = n38442 | n38558 ;
  assign n38560 = n77910 & n38559 ;
  assign n38561 = n38447 | n38560 ;
  assign n38562 = n77911 & n38561 ;
  assign n38563 = n38453 | n38562 ;
  assign n38564 = n77914 & n38563 ;
  assign n38565 = n38457 | n38564 ;
  assign n38566 = n77915 & n38565 ;
  assign n38567 = n38464 | n38566 ;
  assign n38568 = n77918 & n38567 ;
  assign n38569 = n38468 | n38568 ;
  assign n38570 = n77919 & n38569 ;
  assign n38571 = n38474 | n38570 ;
  assign n38572 = n77922 & n38571 ;
  assign n38573 = n38478 | n38572 ;
  assign n38574 = n77923 & n38573 ;
  assign n38575 = n38484 | n38574 ;
  assign n38576 = n77926 & n38575 ;
  assign n38577 = n38488 | n38576 ;
  assign n38578 = n77927 & n38577 ;
  assign n38579 = n38494 | n38578 ;
  assign n38580 = n77930 & n38579 ;
  assign n38581 = n38498 | n38580 ;
  assign n38582 = n77931 & n38581 ;
  assign n38583 = n38504 | n38582 ;
  assign n38584 = n77934 & n38583 ;
  assign n38585 = n38508 | n38584 ;
  assign n38586 = n77935 & n38585 ;
  assign n38587 = n38514 | n38586 ;
  assign n38590 = n38202 | n38518 ;
  assign n77953 = ~n38590 ;
  assign n38591 = n38587 & n77953 ;
  assign n38592 = n38589 | n38591 ;
  assign n38593 = n77950 & n38592 ;
  assign n38594 = n38193 & n77947 ;
  assign n38595 = n38535 & n38594 ;
  assign n38596 = n38593 | n38595 ;
  assign n38608 = n67531 & n38596 ;
  assign n77954 = ~n38586 ;
  assign n38609 = n38514 & n77954 ;
  assign n38610 = n38210 | n38514 ;
  assign n77955 = ~n38610 ;
  assign n38611 = n38510 & n77955 ;
  assign n38612 = n38609 | n38611 ;
  assign n38613 = n77950 & n38612 ;
  assign n38614 = n38201 & n77947 ;
  assign n38615 = n38535 & n38614 ;
  assign n38616 = n38613 | n38615 ;
  assign n38617 = n67348 & n38616 ;
  assign n77956 = ~n38509 ;
  assign n38618 = n38508 & n77956 ;
  assign n38619 = n38218 | n38508 ;
  assign n77957 = ~n38619 ;
  assign n38620 = n38583 & n77957 ;
  assign n38621 = n38618 | n38620 ;
  assign n38622 = n77950 & n38621 ;
  assign n38623 = n38209 & n77947 ;
  assign n38624 = n38535 & n38623 ;
  assign n38625 = n38622 | n38624 ;
  assign n38626 = n67222 & n38625 ;
  assign n77958 = ~n38582 ;
  assign n38627 = n38504 & n77958 ;
  assign n38628 = n38226 | n38504 ;
  assign n77959 = ~n38628 ;
  assign n38629 = n38500 & n77959 ;
  assign n38630 = n38627 | n38629 ;
  assign n38631 = n77950 & n38630 ;
  assign n38632 = n38217 & n77947 ;
  assign n38633 = n38535 & n38632 ;
  assign n38634 = n38631 | n38633 ;
  assign n38635 = n67164 & n38634 ;
  assign n77960 = ~n38499 ;
  assign n38636 = n38498 & n77960 ;
  assign n38637 = n38234 | n38498 ;
  assign n77961 = ~n38637 ;
  assign n38638 = n38579 & n77961 ;
  assign n38639 = n38636 | n38638 ;
  assign n38640 = n77950 & n38639 ;
  assign n38641 = n38225 & n77947 ;
  assign n38642 = n38535 & n38641 ;
  assign n38643 = n38640 | n38642 ;
  assign n38644 = n66979 & n38643 ;
  assign n77962 = ~n38578 ;
  assign n38645 = n38494 & n77962 ;
  assign n38646 = n38242 | n38494 ;
  assign n77963 = ~n38646 ;
  assign n38647 = n38490 & n77963 ;
  assign n38648 = n38645 | n38647 ;
  assign n38649 = n77950 & n38648 ;
  assign n38650 = n38233 & n77947 ;
  assign n38651 = n38535 & n38650 ;
  assign n38652 = n38649 | n38651 ;
  assign n38653 = n66868 & n38652 ;
  assign n77964 = ~n38489 ;
  assign n38654 = n38488 & n77964 ;
  assign n38655 = n38250 | n38488 ;
  assign n77965 = ~n38655 ;
  assign n38656 = n38575 & n77965 ;
  assign n38657 = n38654 | n38656 ;
  assign n38658 = n77950 & n38657 ;
  assign n38659 = n38241 & n77947 ;
  assign n38660 = n38535 & n38659 ;
  assign n38661 = n38658 | n38660 ;
  assign n38662 = n66797 & n38661 ;
  assign n77966 = ~n38574 ;
  assign n38663 = n38484 & n77966 ;
  assign n38664 = n38258 | n38484 ;
  assign n77967 = ~n38664 ;
  assign n38665 = n38480 & n77967 ;
  assign n38666 = n38663 | n38665 ;
  assign n38667 = n77950 & n38666 ;
  assign n38668 = n38249 & n77947 ;
  assign n38669 = n38535 & n38668 ;
  assign n38670 = n38667 | n38669 ;
  assign n38671 = n66654 & n38670 ;
  assign n77968 = ~n38479 ;
  assign n38672 = n38478 & n77968 ;
  assign n38673 = n38266 | n38478 ;
  assign n77969 = ~n38673 ;
  assign n38674 = n38571 & n77969 ;
  assign n38675 = n38672 | n38674 ;
  assign n38676 = n77950 & n38675 ;
  assign n38677 = n38257 & n77947 ;
  assign n38678 = n38535 & n38677 ;
  assign n38679 = n38676 | n38678 ;
  assign n38680 = n66560 & n38679 ;
  assign n77970 = ~n38570 ;
  assign n38681 = n38474 & n77970 ;
  assign n38682 = n38274 | n38474 ;
  assign n77971 = ~n38682 ;
  assign n38683 = n38470 & n77971 ;
  assign n38684 = n38681 | n38683 ;
  assign n38685 = n77950 & n38684 ;
  assign n38686 = n38265 & n77947 ;
  assign n38687 = n38535 & n38686 ;
  assign n38688 = n38685 | n38687 ;
  assign n38689 = n66505 & n38688 ;
  assign n77972 = ~n38469 ;
  assign n38690 = n38468 & n77972 ;
  assign n38691 = n38282 | n38468 ;
  assign n77973 = ~n38691 ;
  assign n38692 = n38567 & n77973 ;
  assign n38693 = n38690 | n38692 ;
  assign n38694 = n77950 & n38693 ;
  assign n38695 = n38273 & n77947 ;
  assign n38696 = n38535 & n38695 ;
  assign n38697 = n38694 | n38696 ;
  assign n38698 = n66379 & n38697 ;
  assign n77974 = ~n38566 ;
  assign n38699 = n38464 & n77974 ;
  assign n38700 = n38290 | n38464 ;
  assign n77975 = ~n38700 ;
  assign n38701 = n38460 & n77975 ;
  assign n38702 = n38699 | n38701 ;
  assign n38703 = n77950 & n38702 ;
  assign n38704 = n38281 & n77947 ;
  assign n38705 = n38535 & n38704 ;
  assign n38706 = n38703 | n38705 ;
  assign n38707 = n66299 & n38706 ;
  assign n77976 = ~n38459 ;
  assign n38708 = n38457 & n77976 ;
  assign n38458 = n38298 | n38457 ;
  assign n77977 = ~n38458 ;
  assign n38709 = n38454 & n77977 ;
  assign n38710 = n38708 | n38709 ;
  assign n38711 = n77950 & n38710 ;
  assign n38712 = n38289 & n77947 ;
  assign n38713 = n38535 & n38712 ;
  assign n38714 = n38711 | n38713 ;
  assign n38715 = n66244 & n38714 ;
  assign n77978 = ~n38562 ;
  assign n38716 = n38453 & n77978 ;
  assign n38717 = n38306 | n38453 ;
  assign n77979 = ~n38717 ;
  assign n38718 = n38449 & n77979 ;
  assign n38719 = n38716 | n38718 ;
  assign n38720 = n77950 & n38719 ;
  assign n38721 = n38297 & n77947 ;
  assign n38722 = n38535 & n38721 ;
  assign n38723 = n38720 | n38722 ;
  assign n38724 = n66145 & n38723 ;
  assign n77980 = ~n38448 ;
  assign n38725 = n38447 & n77980 ;
  assign n38726 = n38314 | n38447 ;
  assign n77981 = ~n38726 ;
  assign n38727 = n38559 & n77981 ;
  assign n38728 = n38725 | n38727 ;
  assign n38729 = n77950 & n38728 ;
  assign n38730 = n38305 & n77947 ;
  assign n38731 = n38535 & n38730 ;
  assign n38732 = n38729 | n38731 ;
  assign n38733 = n66081 & n38732 ;
  assign n77982 = ~n38558 ;
  assign n38734 = n38442 & n77982 ;
  assign n38443 = n38322 | n38442 ;
  assign n77983 = ~n38443 ;
  assign n38735 = n77983 & n38557 ;
  assign n38736 = n38734 | n38735 ;
  assign n38737 = n77950 & n38736 ;
  assign n38738 = n38313 & n77947 ;
  assign n38739 = n38535 & n38738 ;
  assign n38740 = n38737 | n38739 ;
  assign n38741 = n66043 & n38740 ;
  assign n77984 = ~n38437 ;
  assign n38742 = n38436 & n77984 ;
  assign n38743 = n38330 | n38436 ;
  assign n77985 = ~n38743 ;
  assign n38744 = n38555 & n77985 ;
  assign n38745 = n38742 | n38744 ;
  assign n38746 = n77950 & n38745 ;
  assign n38747 = n38321 & n77947 ;
  assign n38748 = n38535 & n38747 ;
  assign n38749 = n38746 | n38748 ;
  assign n38750 = n65960 & n38749 ;
  assign n77986 = ~n38554 ;
  assign n38751 = n38432 & n77986 ;
  assign n38752 = n38338 | n38432 ;
  assign n77987 = ~n38752 ;
  assign n38753 = n38428 & n77987 ;
  assign n38754 = n38751 | n38753 ;
  assign n38755 = n77950 & n38754 ;
  assign n38756 = n38329 & n77947 ;
  assign n38757 = n38535 & n38756 ;
  assign n38758 = n38755 | n38757 ;
  assign n38759 = n65909 & n38758 ;
  assign n77988 = ~n38427 ;
  assign n38760 = n38425 & n77988 ;
  assign n38426 = n38346 | n38425 ;
  assign n77989 = ~n38426 ;
  assign n38761 = n38422 & n77989 ;
  assign n38762 = n38760 | n38761 ;
  assign n38763 = n77950 & n38762 ;
  assign n38764 = n38337 & n77947 ;
  assign n38765 = n38535 & n38764 ;
  assign n38766 = n38763 | n38765 ;
  assign n38767 = n65877 & n38766 ;
  assign n77990 = ~n38550 ;
  assign n38768 = n38420 & n77990 ;
  assign n38421 = n38355 | n38420 ;
  assign n77991 = ~n38421 ;
  assign n38769 = n77991 & n38549 ;
  assign n38770 = n38768 | n38769 ;
  assign n38771 = n77950 & n38770 ;
  assign n38772 = n38345 & n77947 ;
  assign n38773 = n38535 & n38772 ;
  assign n38774 = n38771 | n38773 ;
  assign n38775 = n65820 & n38774 ;
  assign n77992 = ~n38415 ;
  assign n38776 = n38414 & n77992 ;
  assign n38777 = n38363 | n38414 ;
  assign n77993 = ~n38777 ;
  assign n38778 = n38547 & n77993 ;
  assign n38779 = n38776 | n38778 ;
  assign n38780 = n77950 & n38779 ;
  assign n38781 = n38354 & n77947 ;
  assign n38782 = n38535 & n38781 ;
  assign n38783 = n38780 | n38782 ;
  assign n38784 = n65791 & n38783 ;
  assign n77994 = ~n38546 ;
  assign n38785 = n38410 & n77994 ;
  assign n38786 = n38373 | n38410 ;
  assign n77995 = ~n38786 ;
  assign n38787 = n38406 & n77995 ;
  assign n38788 = n38785 | n38787 ;
  assign n38789 = n77950 & n38788 ;
  assign n38790 = n38362 & n77947 ;
  assign n38791 = n38535 & n38790 ;
  assign n38792 = n38789 | n38791 ;
  assign n38793 = n65772 & n38792 ;
  assign n77996 = ~n38405 ;
  assign n38795 = n38404 & n77996 ;
  assign n38794 = n38381 | n38404 ;
  assign n77997 = ~n38794 ;
  assign n38796 = n38402 & n77997 ;
  assign n38797 = n38795 | n38796 ;
  assign n38798 = n77950 & n38797 ;
  assign n38799 = n38371 & n77947 ;
  assign n38800 = n38535 & n38799 ;
  assign n38801 = n38798 | n38800 ;
  assign n38802 = n65746 & n38801 ;
  assign n77998 = ~n38542 ;
  assign n38804 = n38401 & n77998 ;
  assign n38803 = n38397 | n38401 ;
  assign n77999 = ~n38803 ;
  assign n38805 = n38541 & n77999 ;
  assign n38806 = n38804 | n38805 ;
  assign n38807 = n77950 & n38806 ;
  assign n38808 = n38380 & n77947 ;
  assign n38809 = n38535 & n38808 ;
  assign n38810 = n38807 | n38809 ;
  assign n38811 = n65721 & n38810 ;
  assign n38812 = n6013 & n38393 ;
  assign n38813 = n77952 & n38812 ;
  assign n78000 = ~n38813 ;
  assign n38814 = n38541 & n78000 ;
  assign n38815 = n77950 & n38814 ;
  assign n38816 = n38396 & n77947 ;
  assign n38817 = n38535 & n38816 ;
  assign n38818 = n38815 | n38817 ;
  assign n38819 = n65686 & n38818 ;
  assign n38538 = n6013 & n77950 ;
  assign n38826 = x64 & n77950 ;
  assign n78001 = ~n38826 ;
  assign n38827 = x37 & n78001 ;
  assign n38828 = n38538 | n38827 ;
  assign n38830 = x65 & n38828 ;
  assign n38588 = n77938 & n38587 ;
  assign n38820 = n38518 | n38588 ;
  assign n38821 = n77939 & n38820 ;
  assign n38822 = n38534 | n38821 ;
  assign n38823 = n77947 & n38822 ;
  assign n78002 = ~n38823 ;
  assign n38824 = x64 & n78002 ;
  assign n78003 = ~n38824 ;
  assign n38825 = x37 & n78003 ;
  assign n38829 = x65 | n38538 ;
  assign n38831 = n38825 | n38829 ;
  assign n78004 = ~n38830 ;
  assign n38832 = n78004 & n38831 ;
  assign n38833 = n6457 | n38832 ;
  assign n38834 = n65670 & n38828 ;
  assign n78005 = ~n38834 ;
  assign n38835 = n38833 & n78005 ;
  assign n78006 = ~n38817 ;
  assign n38836 = x66 & n78006 ;
  assign n78007 = ~n38815 ;
  assign n38837 = n78007 & n38836 ;
  assign n38838 = n38819 | n38837 ;
  assign n38839 = n38835 | n38838 ;
  assign n78008 = ~n38819 ;
  assign n38840 = n78008 & n38839 ;
  assign n78009 = ~n38809 ;
  assign n38841 = x67 & n78009 ;
  assign n78010 = ~n38807 ;
  assign n38842 = n78010 & n38841 ;
  assign n38843 = n38840 | n38842 ;
  assign n78011 = ~n38811 ;
  assign n38844 = n78011 & n38843 ;
  assign n78012 = ~n38800 ;
  assign n38845 = x68 & n78012 ;
  assign n78013 = ~n38798 ;
  assign n38846 = n78013 & n38845 ;
  assign n38847 = n38802 | n38846 ;
  assign n38848 = n38844 | n38847 ;
  assign n78014 = ~n38802 ;
  assign n38849 = n78014 & n38848 ;
  assign n78015 = ~n38791 ;
  assign n38850 = x69 & n78015 ;
  assign n78016 = ~n38789 ;
  assign n38851 = n78016 & n38850 ;
  assign n38852 = n38793 | n38851 ;
  assign n38855 = n38849 | n38852 ;
  assign n78017 = ~n38793 ;
  assign n38856 = n78017 & n38855 ;
  assign n78018 = ~n38782 ;
  assign n38857 = x70 & n78018 ;
  assign n78019 = ~n38780 ;
  assign n38858 = n78019 & n38857 ;
  assign n38859 = n38784 | n38858 ;
  assign n38860 = n38856 | n38859 ;
  assign n78020 = ~n38784 ;
  assign n38861 = n78020 & n38860 ;
  assign n78021 = ~n38773 ;
  assign n38862 = x71 & n78021 ;
  assign n78022 = ~n38771 ;
  assign n38863 = n78022 & n38862 ;
  assign n38864 = n38775 | n38863 ;
  assign n38867 = n38861 | n38864 ;
  assign n78023 = ~n38775 ;
  assign n38868 = n78023 & n38867 ;
  assign n78024 = ~n38765 ;
  assign n38869 = x72 & n78024 ;
  assign n78025 = ~n38763 ;
  assign n38870 = n78025 & n38869 ;
  assign n38871 = n38767 | n38870 ;
  assign n38872 = n38868 | n38871 ;
  assign n78026 = ~n38767 ;
  assign n38873 = n78026 & n38872 ;
  assign n78027 = ~n38757 ;
  assign n38874 = x73 & n78027 ;
  assign n78028 = ~n38755 ;
  assign n38875 = n78028 & n38874 ;
  assign n38876 = n38759 | n38875 ;
  assign n38878 = n38873 | n38876 ;
  assign n78029 = ~n38759 ;
  assign n38879 = n78029 & n38878 ;
  assign n78030 = ~n38748 ;
  assign n38880 = x74 & n78030 ;
  assign n78031 = ~n38746 ;
  assign n38881 = n78031 & n38880 ;
  assign n38882 = n38750 | n38881 ;
  assign n38883 = n38879 | n38882 ;
  assign n78032 = ~n38750 ;
  assign n38884 = n78032 & n38883 ;
  assign n78033 = ~n38739 ;
  assign n38885 = x75 & n78033 ;
  assign n78034 = ~n38737 ;
  assign n38886 = n78034 & n38885 ;
  assign n38887 = n38741 | n38886 ;
  assign n38889 = n38884 | n38887 ;
  assign n78035 = ~n38741 ;
  assign n38890 = n78035 & n38889 ;
  assign n78036 = ~n38731 ;
  assign n38891 = x76 & n78036 ;
  assign n78037 = ~n38729 ;
  assign n38892 = n78037 & n38891 ;
  assign n38893 = n38733 | n38892 ;
  assign n38894 = n38890 | n38893 ;
  assign n78038 = ~n38733 ;
  assign n38895 = n78038 & n38894 ;
  assign n78039 = ~n38722 ;
  assign n38896 = x77 & n78039 ;
  assign n78040 = ~n38720 ;
  assign n38897 = n78040 & n38896 ;
  assign n38898 = n38724 | n38897 ;
  assign n38900 = n38895 | n38898 ;
  assign n78041 = ~n38724 ;
  assign n38901 = n78041 & n38900 ;
  assign n78042 = ~n38713 ;
  assign n38902 = x78 & n78042 ;
  assign n78043 = ~n38711 ;
  assign n38903 = n78043 & n38902 ;
  assign n38904 = n38715 | n38903 ;
  assign n38905 = n38901 | n38904 ;
  assign n78044 = ~n38715 ;
  assign n38906 = n78044 & n38905 ;
  assign n78045 = ~n38705 ;
  assign n38907 = x79 & n78045 ;
  assign n78046 = ~n38703 ;
  assign n38908 = n78046 & n38907 ;
  assign n38909 = n38707 | n38908 ;
  assign n38911 = n38906 | n38909 ;
  assign n78047 = ~n38707 ;
  assign n38912 = n78047 & n38911 ;
  assign n78048 = ~n38696 ;
  assign n38913 = x80 & n78048 ;
  assign n78049 = ~n38694 ;
  assign n38914 = n78049 & n38913 ;
  assign n38915 = n38698 | n38914 ;
  assign n38916 = n38912 | n38915 ;
  assign n78050 = ~n38698 ;
  assign n38917 = n78050 & n38916 ;
  assign n78051 = ~n38687 ;
  assign n38918 = x81 & n78051 ;
  assign n78052 = ~n38685 ;
  assign n38919 = n78052 & n38918 ;
  assign n38920 = n38689 | n38919 ;
  assign n38922 = n38917 | n38920 ;
  assign n78053 = ~n38689 ;
  assign n38923 = n78053 & n38922 ;
  assign n78054 = ~n38678 ;
  assign n38924 = x82 & n78054 ;
  assign n78055 = ~n38676 ;
  assign n38925 = n78055 & n38924 ;
  assign n38926 = n38680 | n38925 ;
  assign n38927 = n38923 | n38926 ;
  assign n78056 = ~n38680 ;
  assign n38928 = n78056 & n38927 ;
  assign n78057 = ~n38669 ;
  assign n38929 = x83 & n78057 ;
  assign n78058 = ~n38667 ;
  assign n38930 = n78058 & n38929 ;
  assign n38931 = n38671 | n38930 ;
  assign n38933 = n38928 | n38931 ;
  assign n78059 = ~n38671 ;
  assign n38934 = n78059 & n38933 ;
  assign n78060 = ~n38660 ;
  assign n38935 = x84 & n78060 ;
  assign n78061 = ~n38658 ;
  assign n38936 = n78061 & n38935 ;
  assign n38937 = n38662 | n38936 ;
  assign n38938 = n38934 | n38937 ;
  assign n78062 = ~n38662 ;
  assign n38939 = n78062 & n38938 ;
  assign n78063 = ~n38651 ;
  assign n38940 = x85 & n78063 ;
  assign n78064 = ~n38649 ;
  assign n38941 = n78064 & n38940 ;
  assign n38942 = n38653 | n38941 ;
  assign n38944 = n38939 | n38942 ;
  assign n78065 = ~n38653 ;
  assign n38945 = n78065 & n38944 ;
  assign n78066 = ~n38642 ;
  assign n38946 = x86 & n78066 ;
  assign n78067 = ~n38640 ;
  assign n38947 = n78067 & n38946 ;
  assign n38948 = n38644 | n38947 ;
  assign n38949 = n38945 | n38948 ;
  assign n78068 = ~n38644 ;
  assign n38950 = n78068 & n38949 ;
  assign n78069 = ~n38633 ;
  assign n38951 = x87 & n78069 ;
  assign n78070 = ~n38631 ;
  assign n38952 = n78070 & n38951 ;
  assign n38953 = n38635 | n38952 ;
  assign n38955 = n38950 | n38953 ;
  assign n78071 = ~n38635 ;
  assign n38956 = n78071 & n38955 ;
  assign n78072 = ~n38624 ;
  assign n38957 = x88 & n78072 ;
  assign n78073 = ~n38622 ;
  assign n38958 = n78073 & n38957 ;
  assign n38959 = n38626 | n38958 ;
  assign n38960 = n38956 | n38959 ;
  assign n78074 = ~n38626 ;
  assign n38961 = n78074 & n38960 ;
  assign n78075 = ~n38615 ;
  assign n38962 = x89 & n78075 ;
  assign n78076 = ~n38613 ;
  assign n38963 = n78076 & n38962 ;
  assign n38964 = n38617 | n38963 ;
  assign n38966 = n38961 | n38964 ;
  assign n78077 = ~n38617 ;
  assign n38967 = n78077 & n38966 ;
  assign n78078 = ~n38595 ;
  assign n38968 = x90 & n78078 ;
  assign n78079 = ~n38593 ;
  assign n38969 = n78079 & n38968 ;
  assign n38970 = n38608 | n38969 ;
  assign n38971 = n38967 | n38970 ;
  assign n78080 = ~n38608 ;
  assign n38972 = n78080 & n38971 ;
  assign n78081 = ~n38605 ;
  assign n38973 = x91 & n78081 ;
  assign n78082 = ~n38603 ;
  assign n38974 = n78082 & n38973 ;
  assign n38975 = n38607 | n38974 ;
  assign n38977 = n38972 | n38975 ;
  assign n78083 = ~n38607 ;
  assign n38978 = n78083 & n38977 ;
  assign n38979 = n6615 | n38978 ;
  assign n78084 = ~n38606 ;
  assign n38980 = n78084 & n38979 ;
  assign n78085 = ~n38972 ;
  assign n38976 = n78085 & n38975 ;
  assign n38986 = n38538 | n38825 ;
  assign n38987 = x65 & n38986 ;
  assign n78086 = ~n38987 ;
  assign n38988 = n38831 & n78086 ;
  assign n38989 = n6457 | n38988 ;
  assign n38990 = n78005 & n38989 ;
  assign n38991 = n38838 | n38990 ;
  assign n38992 = n78008 & n38991 ;
  assign n38993 = n38811 | n38842 ;
  assign n38995 = n38992 | n38993 ;
  assign n38996 = n78011 & n38995 ;
  assign n38997 = n38846 | n38996 ;
  assign n38999 = n78014 & n38997 ;
  assign n39000 = n38852 | n38999 ;
  assign n39001 = n78017 & n39000 ;
  assign n39002 = n38858 | n39001 ;
  assign n39004 = n78020 & n39002 ;
  assign n39005 = n38864 | n39004 ;
  assign n39006 = n78023 & n39005 ;
  assign n39007 = n38871 | n39006 ;
  assign n39009 = n78026 & n39007 ;
  assign n39010 = n38876 | n39009 ;
  assign n39011 = n78029 & n39010 ;
  assign n39012 = n38882 | n39011 ;
  assign n39014 = n78032 & n39012 ;
  assign n39015 = n38887 | n39014 ;
  assign n39016 = n78035 & n39015 ;
  assign n39017 = n38893 | n39016 ;
  assign n39019 = n78038 & n39017 ;
  assign n39020 = n38898 | n39019 ;
  assign n39021 = n78041 & n39020 ;
  assign n39022 = n38904 | n39021 ;
  assign n39024 = n78044 & n39022 ;
  assign n39025 = n38909 | n39024 ;
  assign n39026 = n78047 & n39025 ;
  assign n39027 = n38915 | n39026 ;
  assign n39029 = n78050 & n39027 ;
  assign n39030 = n38920 | n39029 ;
  assign n39031 = n78053 & n39030 ;
  assign n39032 = n38926 | n39031 ;
  assign n39034 = n78056 & n39032 ;
  assign n39035 = n38931 | n39034 ;
  assign n39036 = n78059 & n39035 ;
  assign n39037 = n38937 | n39036 ;
  assign n39039 = n78062 & n39037 ;
  assign n39040 = n38942 | n39039 ;
  assign n39041 = n78065 & n39040 ;
  assign n39042 = n38948 | n39041 ;
  assign n39044 = n78068 & n39042 ;
  assign n39045 = n38953 | n39044 ;
  assign n39046 = n78071 & n39045 ;
  assign n39047 = n38959 | n39046 ;
  assign n39049 = n78074 & n39047 ;
  assign n39050 = n38964 | n39049 ;
  assign n39051 = n78077 & n39050 ;
  assign n39053 = n38970 | n39051 ;
  assign n39060 = n38608 | n38975 ;
  assign n78087 = ~n39060 ;
  assign n39061 = n39053 & n78087 ;
  assign n39062 = n38976 | n39061 ;
  assign n39063 = n38979 | n39062 ;
  assign n78088 = ~n38980 ;
  assign n39064 = n78088 & n39063 ;
  assign n39065 = n67763 & n39064 ;
  assign n78089 = ~n38979 ;
  assign n39431 = n78089 & n39062 ;
  assign n39432 = n38606 & n38979 ;
  assign n78090 = ~n39432 ;
  assign n39433 = x92 & n78090 ;
  assign n78091 = ~n39431 ;
  assign n39434 = n78091 & n39433 ;
  assign n39435 = n39065 | n39434 ;
  assign n38984 = n38596 & n38979 ;
  assign n78092 = ~n39051 ;
  assign n39052 = n38970 & n78092 ;
  assign n39054 = n38617 | n38970 ;
  assign n78093 = ~n39054 ;
  assign n39055 = n38966 & n78093 ;
  assign n39056 = n39052 | n39055 ;
  assign n39057 = n67757 & n39056 ;
  assign n78094 = ~n38978 ;
  assign n39058 = n78094 & n39057 ;
  assign n39059 = n38984 | n39058 ;
  assign n39066 = n67622 & n39059 ;
  assign n39067 = n38616 & n38979 ;
  assign n78095 = ~n38961 ;
  assign n38965 = n78095 & n38964 ;
  assign n39068 = n38626 | n38964 ;
  assign n78096 = ~n39068 ;
  assign n39069 = n39047 & n78096 ;
  assign n39070 = n38965 | n39069 ;
  assign n39071 = n67757 & n39070 ;
  assign n39072 = n78094 & n39071 ;
  assign n39073 = n39067 | n39072 ;
  assign n39074 = n67531 & n39073 ;
  assign n78097 = ~n39072 ;
  assign n39419 = x90 & n78097 ;
  assign n78098 = ~n39067 ;
  assign n39420 = n78098 & n39419 ;
  assign n39421 = n39074 | n39420 ;
  assign n39075 = n38625 & n38979 ;
  assign n78099 = ~n39046 ;
  assign n39048 = n38959 & n78099 ;
  assign n39076 = n38635 | n38959 ;
  assign n78100 = ~n39076 ;
  assign n39077 = n38955 & n78100 ;
  assign n39078 = n39048 | n39077 ;
  assign n39079 = n67757 & n39078 ;
  assign n39080 = n78094 & n39079 ;
  assign n39081 = n39075 | n39080 ;
  assign n39082 = n67348 & n39081 ;
  assign n39083 = n38634 & n38979 ;
  assign n78101 = ~n38950 ;
  assign n38954 = n78101 & n38953 ;
  assign n39084 = n38644 | n38953 ;
  assign n78102 = ~n39084 ;
  assign n39085 = n39042 & n78102 ;
  assign n39086 = n38954 | n39085 ;
  assign n39087 = n67757 & n39086 ;
  assign n39088 = n78094 & n39087 ;
  assign n39089 = n39083 | n39088 ;
  assign n39090 = n67222 & n39089 ;
  assign n78103 = ~n39088 ;
  assign n39407 = x88 & n78103 ;
  assign n78104 = ~n39083 ;
  assign n39408 = n78104 & n39407 ;
  assign n39409 = n39090 | n39408 ;
  assign n39091 = n38643 & n38979 ;
  assign n78105 = ~n39041 ;
  assign n39043 = n38948 & n78105 ;
  assign n39092 = n38653 | n38948 ;
  assign n78106 = ~n39092 ;
  assign n39093 = n38944 & n78106 ;
  assign n39094 = n39043 | n39093 ;
  assign n39095 = n67757 & n39094 ;
  assign n39096 = n78094 & n39095 ;
  assign n39097 = n39091 | n39096 ;
  assign n39098 = n67164 & n39097 ;
  assign n39099 = n38652 & n38979 ;
  assign n78107 = ~n38939 ;
  assign n38943 = n78107 & n38942 ;
  assign n39100 = n38662 | n38942 ;
  assign n78108 = ~n39100 ;
  assign n39101 = n39037 & n78108 ;
  assign n39102 = n38943 | n39101 ;
  assign n39103 = n67757 & n39102 ;
  assign n39104 = n78094 & n39103 ;
  assign n39105 = n39099 | n39104 ;
  assign n39106 = n66979 & n39105 ;
  assign n78109 = ~n39104 ;
  assign n39395 = x86 & n78109 ;
  assign n78110 = ~n39099 ;
  assign n39396 = n78110 & n39395 ;
  assign n39397 = n39106 | n39396 ;
  assign n39107 = n38661 & n38979 ;
  assign n78111 = ~n39036 ;
  assign n39038 = n38937 & n78111 ;
  assign n39108 = n38671 | n38937 ;
  assign n78112 = ~n39108 ;
  assign n39109 = n38933 & n78112 ;
  assign n39110 = n39038 | n39109 ;
  assign n39111 = n67757 & n39110 ;
  assign n39112 = n78094 & n39111 ;
  assign n39113 = n39107 | n39112 ;
  assign n39114 = n66868 & n39113 ;
  assign n39115 = n38670 & n38979 ;
  assign n78113 = ~n38928 ;
  assign n38932 = n78113 & n38931 ;
  assign n39116 = n38680 | n38931 ;
  assign n78114 = ~n39116 ;
  assign n39117 = n39032 & n78114 ;
  assign n39118 = n38932 | n39117 ;
  assign n39119 = n67757 & n39118 ;
  assign n39120 = n78094 & n39119 ;
  assign n39121 = n39115 | n39120 ;
  assign n39122 = n66797 & n39121 ;
  assign n78115 = ~n39120 ;
  assign n39383 = x84 & n78115 ;
  assign n78116 = ~n39115 ;
  assign n39384 = n78116 & n39383 ;
  assign n39385 = n39122 | n39384 ;
  assign n39123 = n38679 & n38979 ;
  assign n78117 = ~n39031 ;
  assign n39033 = n38926 & n78117 ;
  assign n39124 = n38689 | n38926 ;
  assign n78118 = ~n39124 ;
  assign n39125 = n38922 & n78118 ;
  assign n39126 = n39033 | n39125 ;
  assign n39127 = n67757 & n39126 ;
  assign n39128 = n78094 & n39127 ;
  assign n39129 = n39123 | n39128 ;
  assign n39130 = n66654 & n39129 ;
  assign n39131 = n38688 & n38979 ;
  assign n78119 = ~n38917 ;
  assign n38921 = n78119 & n38920 ;
  assign n39132 = n38698 | n38920 ;
  assign n78120 = ~n39132 ;
  assign n39133 = n39027 & n78120 ;
  assign n39134 = n38921 | n39133 ;
  assign n39135 = n67757 & n39134 ;
  assign n39136 = n78094 & n39135 ;
  assign n39137 = n39131 | n39136 ;
  assign n39138 = n66560 & n39137 ;
  assign n78121 = ~n39136 ;
  assign n39371 = x82 & n78121 ;
  assign n78122 = ~n39131 ;
  assign n39372 = n78122 & n39371 ;
  assign n39373 = n39138 | n39372 ;
  assign n39139 = n38697 & n38979 ;
  assign n78123 = ~n39026 ;
  assign n39028 = n38915 & n78123 ;
  assign n39140 = n38707 | n38915 ;
  assign n78124 = ~n39140 ;
  assign n39141 = n38911 & n78124 ;
  assign n39142 = n39028 | n39141 ;
  assign n39143 = n67757 & n39142 ;
  assign n39144 = n78094 & n39143 ;
  assign n39145 = n39139 | n39144 ;
  assign n39146 = n66505 & n39145 ;
  assign n39147 = n38706 & n38979 ;
  assign n78125 = ~n38906 ;
  assign n38910 = n78125 & n38909 ;
  assign n39148 = n38715 | n38909 ;
  assign n78126 = ~n39148 ;
  assign n39149 = n39022 & n78126 ;
  assign n39150 = n38910 | n39149 ;
  assign n39151 = n67757 & n39150 ;
  assign n39152 = n78094 & n39151 ;
  assign n39153 = n39147 | n39152 ;
  assign n39154 = n66379 & n39153 ;
  assign n78127 = ~n39152 ;
  assign n39359 = x80 & n78127 ;
  assign n78128 = ~n39147 ;
  assign n39360 = n78128 & n39359 ;
  assign n39361 = n39154 | n39360 ;
  assign n39155 = n38714 & n38979 ;
  assign n78129 = ~n39021 ;
  assign n39023 = n38904 & n78129 ;
  assign n39156 = n38724 | n38904 ;
  assign n78130 = ~n39156 ;
  assign n39157 = n38900 & n78130 ;
  assign n39158 = n39023 | n39157 ;
  assign n39159 = n67757 & n39158 ;
  assign n39160 = n78094 & n39159 ;
  assign n39161 = n39155 | n39160 ;
  assign n39162 = n66299 & n39161 ;
  assign n39163 = n38723 & n38979 ;
  assign n78131 = ~n38895 ;
  assign n38899 = n78131 & n38898 ;
  assign n39164 = n38733 | n38898 ;
  assign n78132 = ~n39164 ;
  assign n39165 = n39017 & n78132 ;
  assign n39166 = n38899 | n39165 ;
  assign n39167 = n67757 & n39166 ;
  assign n39168 = n78094 & n39167 ;
  assign n39169 = n39163 | n39168 ;
  assign n39170 = n66244 & n39169 ;
  assign n78133 = ~n39168 ;
  assign n39347 = x78 & n78133 ;
  assign n78134 = ~n39163 ;
  assign n39348 = n78134 & n39347 ;
  assign n39349 = n39170 | n39348 ;
  assign n39171 = n38732 & n38979 ;
  assign n78135 = ~n39016 ;
  assign n39018 = n38893 & n78135 ;
  assign n39172 = n38741 | n38893 ;
  assign n78136 = ~n39172 ;
  assign n39173 = n38889 & n78136 ;
  assign n39174 = n39018 | n39173 ;
  assign n39175 = n67757 & n39174 ;
  assign n39176 = n78094 & n39175 ;
  assign n39177 = n39171 | n39176 ;
  assign n39178 = n66145 & n39177 ;
  assign n39179 = n38740 & n38979 ;
  assign n78137 = ~n38884 ;
  assign n38888 = n78137 & n38887 ;
  assign n39180 = n38750 | n38887 ;
  assign n78138 = ~n39180 ;
  assign n39181 = n39012 & n78138 ;
  assign n39182 = n38888 | n39181 ;
  assign n39183 = n67757 & n39182 ;
  assign n39184 = n78094 & n39183 ;
  assign n39185 = n39179 | n39184 ;
  assign n39186 = n66081 & n39185 ;
  assign n78139 = ~n39184 ;
  assign n39335 = x76 & n78139 ;
  assign n78140 = ~n39179 ;
  assign n39336 = n78140 & n39335 ;
  assign n39337 = n39186 | n39336 ;
  assign n39187 = n38749 & n38979 ;
  assign n78141 = ~n39011 ;
  assign n39013 = n38882 & n78141 ;
  assign n39188 = n38759 | n38882 ;
  assign n78142 = ~n39188 ;
  assign n39189 = n38878 & n78142 ;
  assign n39190 = n39013 | n39189 ;
  assign n39191 = n67757 & n39190 ;
  assign n39192 = n78094 & n39191 ;
  assign n39193 = n39187 | n39192 ;
  assign n39194 = n66043 & n39193 ;
  assign n39195 = n38758 & n38979 ;
  assign n78143 = ~n38873 ;
  assign n38877 = n78143 & n38876 ;
  assign n39196 = n38767 | n38876 ;
  assign n78144 = ~n39196 ;
  assign n39197 = n39007 & n78144 ;
  assign n39198 = n38877 | n39197 ;
  assign n39199 = n67757 & n39198 ;
  assign n39200 = n78094 & n39199 ;
  assign n39201 = n39195 | n39200 ;
  assign n39202 = n65960 & n39201 ;
  assign n78145 = ~n39200 ;
  assign n39323 = x74 & n78145 ;
  assign n78146 = ~n39195 ;
  assign n39324 = n78146 & n39323 ;
  assign n39325 = n39202 | n39324 ;
  assign n39203 = n38766 & n38979 ;
  assign n78147 = ~n39006 ;
  assign n39008 = n38871 & n78147 ;
  assign n39204 = n38775 | n38871 ;
  assign n78148 = ~n39204 ;
  assign n39205 = n38867 & n78148 ;
  assign n39206 = n39008 | n39205 ;
  assign n39207 = n67757 & n39206 ;
  assign n39208 = n78094 & n39207 ;
  assign n39209 = n39203 | n39208 ;
  assign n39210 = n65909 & n39209 ;
  assign n39211 = n38774 & n38979 ;
  assign n78149 = ~n38861 ;
  assign n38865 = n78149 & n38864 ;
  assign n38866 = n38784 | n38864 ;
  assign n39212 = n38859 | n39001 ;
  assign n78150 = ~n38866 ;
  assign n39213 = n78150 & n39212 ;
  assign n39214 = n38865 | n39213 ;
  assign n39215 = n67757 & n39214 ;
  assign n39216 = n78094 & n39215 ;
  assign n39217 = n39211 | n39216 ;
  assign n39218 = n65877 & n39217 ;
  assign n78151 = ~n39216 ;
  assign n39311 = x72 & n78151 ;
  assign n78152 = ~n39211 ;
  assign n39312 = n78152 & n39311 ;
  assign n39313 = n39218 | n39312 ;
  assign n38981 = n38783 & n38979 ;
  assign n78153 = ~n39001 ;
  assign n39003 = n38859 & n78153 ;
  assign n39219 = n38793 | n38859 ;
  assign n78154 = ~n39219 ;
  assign n39220 = n38855 & n78154 ;
  assign n39221 = n39003 | n39220 ;
  assign n39222 = n67757 & n39221 ;
  assign n39223 = n78094 & n39222 ;
  assign n39224 = n38981 | n39223 ;
  assign n39225 = n65820 & n39224 ;
  assign n39226 = n38792 & n38979 ;
  assign n78155 = ~n38849 ;
  assign n38853 = n78155 & n38852 ;
  assign n38854 = n38802 | n38852 ;
  assign n39227 = n38847 | n38996 ;
  assign n78156 = ~n38854 ;
  assign n39228 = n78156 & n39227 ;
  assign n39229 = n38853 | n39228 ;
  assign n39230 = n67757 & n39229 ;
  assign n39231 = n78094 & n39230 ;
  assign n39232 = n39226 | n39231 ;
  assign n39233 = n65791 & n39232 ;
  assign n78157 = ~n39231 ;
  assign n39299 = x70 & n78157 ;
  assign n78158 = ~n39226 ;
  assign n39300 = n78158 & n39299 ;
  assign n39301 = n39233 | n39300 ;
  assign n38983 = n38801 & n38979 ;
  assign n78159 = ~n38996 ;
  assign n38998 = n38847 & n78159 ;
  assign n39234 = n38840 | n38993 ;
  assign n39235 = n38811 | n38847 ;
  assign n78160 = ~n39235 ;
  assign n39236 = n39234 & n78160 ;
  assign n39237 = n38998 | n39236 ;
  assign n39238 = n67757 & n39237 ;
  assign n39239 = n78094 & n39238 ;
  assign n39240 = n38983 | n39239 ;
  assign n39241 = n65772 & n39240 ;
  assign n38982 = n38810 & n38979 ;
  assign n78161 = ~n38840 ;
  assign n38994 = n78161 & n38993 ;
  assign n39242 = n38819 | n38993 ;
  assign n78162 = ~n39242 ;
  assign n39243 = n38839 & n78162 ;
  assign n39244 = n38994 | n39243 ;
  assign n39245 = n67757 & n39244 ;
  assign n39246 = n78094 & n39245 ;
  assign n39247 = n38982 | n39246 ;
  assign n39248 = n65746 & n39247 ;
  assign n78163 = ~n39246 ;
  assign n39289 = x68 & n78163 ;
  assign n78164 = ~n38982 ;
  assign n39290 = n78164 & n39289 ;
  assign n39291 = n39248 | n39290 ;
  assign n38985 = n38818 & n38979 ;
  assign n39249 = n38834 | n38838 ;
  assign n78165 = ~n39249 ;
  assign n39250 = n38989 & n78165 ;
  assign n78166 = ~n38990 ;
  assign n39251 = n38838 & n78166 ;
  assign n39252 = n39250 | n39251 ;
  assign n39253 = n67757 & n39252 ;
  assign n39254 = n78094 & n39253 ;
  assign n39255 = n38985 | n39254 ;
  assign n39256 = n65721 & n39255 ;
  assign n39257 = n38979 & n38986 ;
  assign n39258 = n6457 & n38831 ;
  assign n39259 = n78004 & n39258 ;
  assign n39260 = n6615 | n39259 ;
  assign n78167 = ~n39260 ;
  assign n39261 = n38989 & n78167 ;
  assign n39262 = n78094 & n39261 ;
  assign n39263 = n39257 | n39262 ;
  assign n39264 = n65686 & n39263 ;
  assign n78168 = ~n39262 ;
  assign n39279 = x66 & n78168 ;
  assign n78169 = ~n39257 ;
  assign n39280 = n78169 & n39279 ;
  assign n39281 = n39264 | n39280 ;
  assign n39265 = n78080 & n39053 ;
  assign n39266 = n38975 | n39265 ;
  assign n39267 = n78083 & n39266 ;
  assign n78170 = ~n39267 ;
  assign n39268 = n6894 & n78170 ;
  assign n78171 = ~n39268 ;
  assign n39269 = x36 & n78171 ;
  assign n39270 = n6899 & n78094 ;
  assign n39271 = n39269 | n39270 ;
  assign n39272 = x65 & n39271 ;
  assign n39273 = x65 | n39270 ;
  assign n39274 = n39269 | n39273 ;
  assign n78172 = ~n39272 ;
  assign n39275 = n78172 & n39274 ;
  assign n39277 = n6907 | n39275 ;
  assign n39278 = n65670 & n39271 ;
  assign n78173 = ~n39278 ;
  assign n39282 = n39277 & n78173 ;
  assign n39283 = n39281 | n39282 ;
  assign n78174 = ~n39264 ;
  assign n39284 = n78174 & n39283 ;
  assign n78175 = ~n39254 ;
  assign n39285 = x67 & n78175 ;
  assign n78176 = ~n38985 ;
  assign n39286 = n78176 & n39285 ;
  assign n39287 = n39256 | n39286 ;
  assign n39288 = n39284 | n39287 ;
  assign n78177 = ~n39256 ;
  assign n39292 = n78177 & n39288 ;
  assign n39293 = n39291 | n39292 ;
  assign n78178 = ~n39248 ;
  assign n39294 = n78178 & n39293 ;
  assign n78179 = ~n39239 ;
  assign n39295 = x69 & n78179 ;
  assign n78180 = ~n38983 ;
  assign n39296 = n78180 & n39295 ;
  assign n39297 = n39241 | n39296 ;
  assign n39298 = n39294 | n39297 ;
  assign n78181 = ~n39241 ;
  assign n39303 = n78181 & n39298 ;
  assign n39304 = n39301 | n39303 ;
  assign n78182 = ~n39233 ;
  assign n39305 = n78182 & n39304 ;
  assign n78183 = ~n39223 ;
  assign n39306 = x71 & n78183 ;
  assign n78184 = ~n38981 ;
  assign n39307 = n78184 & n39306 ;
  assign n39308 = n39225 | n39307 ;
  assign n39310 = n39305 | n39308 ;
  assign n78185 = ~n39225 ;
  assign n39315 = n78185 & n39310 ;
  assign n39316 = n39313 | n39315 ;
  assign n78186 = ~n39218 ;
  assign n39317 = n78186 & n39316 ;
  assign n78187 = ~n39208 ;
  assign n39318 = x73 & n78187 ;
  assign n78188 = ~n39203 ;
  assign n39319 = n78188 & n39318 ;
  assign n39320 = n39210 | n39319 ;
  assign n39322 = n39317 | n39320 ;
  assign n78189 = ~n39210 ;
  assign n39327 = n78189 & n39322 ;
  assign n39328 = n39325 | n39327 ;
  assign n78190 = ~n39202 ;
  assign n39329 = n78190 & n39328 ;
  assign n78191 = ~n39192 ;
  assign n39330 = x75 & n78191 ;
  assign n78192 = ~n39187 ;
  assign n39331 = n78192 & n39330 ;
  assign n39332 = n39194 | n39331 ;
  assign n39334 = n39329 | n39332 ;
  assign n78193 = ~n39194 ;
  assign n39339 = n78193 & n39334 ;
  assign n39340 = n39337 | n39339 ;
  assign n78194 = ~n39186 ;
  assign n39341 = n78194 & n39340 ;
  assign n78195 = ~n39176 ;
  assign n39342 = x77 & n78195 ;
  assign n78196 = ~n39171 ;
  assign n39343 = n78196 & n39342 ;
  assign n39344 = n39178 | n39343 ;
  assign n39346 = n39341 | n39344 ;
  assign n78197 = ~n39178 ;
  assign n39351 = n78197 & n39346 ;
  assign n39352 = n39349 | n39351 ;
  assign n78198 = ~n39170 ;
  assign n39353 = n78198 & n39352 ;
  assign n78199 = ~n39160 ;
  assign n39354 = x79 & n78199 ;
  assign n78200 = ~n39155 ;
  assign n39355 = n78200 & n39354 ;
  assign n39356 = n39162 | n39355 ;
  assign n39358 = n39353 | n39356 ;
  assign n78201 = ~n39162 ;
  assign n39363 = n78201 & n39358 ;
  assign n39364 = n39361 | n39363 ;
  assign n78202 = ~n39154 ;
  assign n39365 = n78202 & n39364 ;
  assign n78203 = ~n39144 ;
  assign n39366 = x81 & n78203 ;
  assign n78204 = ~n39139 ;
  assign n39367 = n78204 & n39366 ;
  assign n39368 = n39146 | n39367 ;
  assign n39370 = n39365 | n39368 ;
  assign n78205 = ~n39146 ;
  assign n39375 = n78205 & n39370 ;
  assign n39376 = n39373 | n39375 ;
  assign n78206 = ~n39138 ;
  assign n39377 = n78206 & n39376 ;
  assign n78207 = ~n39128 ;
  assign n39378 = x83 & n78207 ;
  assign n78208 = ~n39123 ;
  assign n39379 = n78208 & n39378 ;
  assign n39380 = n39130 | n39379 ;
  assign n39382 = n39377 | n39380 ;
  assign n78209 = ~n39130 ;
  assign n39387 = n78209 & n39382 ;
  assign n39388 = n39385 | n39387 ;
  assign n78210 = ~n39122 ;
  assign n39389 = n78210 & n39388 ;
  assign n78211 = ~n39112 ;
  assign n39390 = x85 & n78211 ;
  assign n78212 = ~n39107 ;
  assign n39391 = n78212 & n39390 ;
  assign n39392 = n39114 | n39391 ;
  assign n39394 = n39389 | n39392 ;
  assign n78213 = ~n39114 ;
  assign n39399 = n78213 & n39394 ;
  assign n39400 = n39397 | n39399 ;
  assign n78214 = ~n39106 ;
  assign n39401 = n78214 & n39400 ;
  assign n78215 = ~n39096 ;
  assign n39402 = x87 & n78215 ;
  assign n78216 = ~n39091 ;
  assign n39403 = n78216 & n39402 ;
  assign n39404 = n39098 | n39403 ;
  assign n39406 = n39401 | n39404 ;
  assign n78217 = ~n39098 ;
  assign n39411 = n78217 & n39406 ;
  assign n39412 = n39409 | n39411 ;
  assign n78218 = ~n39090 ;
  assign n39413 = n78218 & n39412 ;
  assign n78219 = ~n39080 ;
  assign n39414 = x89 & n78219 ;
  assign n78220 = ~n39075 ;
  assign n39415 = n78220 & n39414 ;
  assign n39416 = n39082 | n39415 ;
  assign n39418 = n39413 | n39416 ;
  assign n78221 = ~n39082 ;
  assign n39423 = n78221 & n39418 ;
  assign n39424 = n39421 | n39423 ;
  assign n78222 = ~n39074 ;
  assign n39425 = n78222 & n39424 ;
  assign n78223 = ~n39058 ;
  assign n39426 = x91 & n78223 ;
  assign n78224 = ~n38984 ;
  assign n39427 = n78224 & n39426 ;
  assign n39428 = n39066 | n39427 ;
  assign n39430 = n39425 | n39428 ;
  assign n78225 = ~n39066 ;
  assign n39436 = n78225 & n39430 ;
  assign n39437 = n39435 | n39436 ;
  assign n78226 = ~n39065 ;
  assign n39438 = n78226 & n39437 ;
  assign n39439 = n7066 | n39438 ;
  assign n78227 = ~n39064 ;
  assign n39441 = n78227 & n39439 ;
  assign n78228 = ~n39436 ;
  assign n39881 = n39435 & n78228 ;
  assign n39443 = n6894 & n78094 ;
  assign n78229 = ~n39443 ;
  assign n39444 = x36 & n78229 ;
  assign n39445 = n39270 | n39444 ;
  assign n39446 = x65 & n39445 ;
  assign n78230 = ~n39446 ;
  assign n39447 = n39274 & n78230 ;
  assign n39448 = n6907 | n39447 ;
  assign n39449 = n78173 & n39448 ;
  assign n39450 = n39281 | n39449 ;
  assign n39451 = n78174 & n39450 ;
  assign n39452 = n39287 | n39451 ;
  assign n39453 = n78177 & n39452 ;
  assign n39454 = n39291 | n39453 ;
  assign n39455 = n78178 & n39454 ;
  assign n39456 = n39297 | n39455 ;
  assign n39457 = n78181 & n39456 ;
  assign n39458 = n39301 | n39457 ;
  assign n39459 = n78182 & n39458 ;
  assign n39460 = n39308 | n39459 ;
  assign n39461 = n78185 & n39460 ;
  assign n39462 = n39313 | n39461 ;
  assign n39463 = n78186 & n39462 ;
  assign n39464 = n39320 | n39463 ;
  assign n39465 = n78189 & n39464 ;
  assign n39466 = n39325 | n39465 ;
  assign n39467 = n78190 & n39466 ;
  assign n39468 = n39332 | n39467 ;
  assign n39469 = n78193 & n39468 ;
  assign n39470 = n39337 | n39469 ;
  assign n39471 = n78194 & n39470 ;
  assign n39472 = n39344 | n39471 ;
  assign n39473 = n78197 & n39472 ;
  assign n39474 = n39349 | n39473 ;
  assign n39475 = n78198 & n39474 ;
  assign n39476 = n39356 | n39475 ;
  assign n39477 = n78201 & n39476 ;
  assign n39478 = n39361 | n39477 ;
  assign n39479 = n78202 & n39478 ;
  assign n39480 = n39368 | n39479 ;
  assign n39481 = n78205 & n39480 ;
  assign n39482 = n39373 | n39481 ;
  assign n39483 = n78206 & n39482 ;
  assign n39484 = n39380 | n39483 ;
  assign n39485 = n78209 & n39484 ;
  assign n39486 = n39385 | n39485 ;
  assign n39487 = n78210 & n39486 ;
  assign n39488 = n39392 | n39487 ;
  assign n39489 = n78213 & n39488 ;
  assign n39490 = n39397 | n39489 ;
  assign n39491 = n78214 & n39490 ;
  assign n39492 = n39404 | n39491 ;
  assign n39493 = n78217 & n39492 ;
  assign n39494 = n39409 | n39493 ;
  assign n39495 = n78218 & n39494 ;
  assign n39496 = n39416 | n39495 ;
  assign n39497 = n78221 & n39496 ;
  assign n39498 = n39421 | n39497 ;
  assign n39500 = n78222 & n39498 ;
  assign n39718 = n39428 | n39500 ;
  assign n39882 = n39066 | n39435 ;
  assign n78231 = ~n39882 ;
  assign n39883 = n39718 & n78231 ;
  assign n39884 = n39881 | n39883 ;
  assign n39885 = n39439 | n39884 ;
  assign n78232 = ~n39441 ;
  assign n39886 = n78232 & n39885 ;
  assign n39894 = n67905 & n39886 ;
  assign n39442 = n39059 & n39439 ;
  assign n39429 = n39074 | n39428 ;
  assign n78233 = ~n39429 ;
  assign n39499 = n78233 & n39498 ;
  assign n78234 = ~n39500 ;
  assign n39501 = n39428 & n78234 ;
  assign n39502 = n39499 | n39501 ;
  assign n39503 = n67905 & n39502 ;
  assign n78235 = ~n39438 ;
  assign n39504 = n78235 & n39503 ;
  assign n39505 = n39442 | n39504 ;
  assign n39506 = n67763 & n39505 ;
  assign n39507 = n39073 & n39439 ;
  assign n39422 = n39082 | n39421 ;
  assign n78236 = ~n39422 ;
  assign n39508 = n39418 & n78236 ;
  assign n78237 = ~n39423 ;
  assign n39509 = n39421 & n78237 ;
  assign n39510 = n39508 | n39509 ;
  assign n39511 = n67905 & n39510 ;
  assign n39512 = n78235 & n39511 ;
  assign n39513 = n39507 | n39512 ;
  assign n39514 = n67622 & n39513 ;
  assign n39515 = n39081 & n39439 ;
  assign n39417 = n39090 | n39416 ;
  assign n78238 = ~n39417 ;
  assign n39516 = n78238 & n39494 ;
  assign n78239 = ~n39495 ;
  assign n39517 = n39416 & n78239 ;
  assign n39518 = n39516 | n39517 ;
  assign n39519 = n67905 & n39518 ;
  assign n39520 = n78235 & n39519 ;
  assign n39521 = n39515 | n39520 ;
  assign n39522 = n67531 & n39521 ;
  assign n39523 = n39089 & n39439 ;
  assign n39410 = n39098 | n39409 ;
  assign n78240 = ~n39410 ;
  assign n39524 = n39406 & n78240 ;
  assign n78241 = ~n39411 ;
  assign n39525 = n39409 & n78241 ;
  assign n39526 = n39524 | n39525 ;
  assign n39527 = n67905 & n39526 ;
  assign n39528 = n78235 & n39527 ;
  assign n39529 = n39523 | n39528 ;
  assign n39530 = n67348 & n39529 ;
  assign n39531 = n39097 & n39439 ;
  assign n39405 = n39106 | n39404 ;
  assign n78242 = ~n39405 ;
  assign n39532 = n78242 & n39490 ;
  assign n78243 = ~n39491 ;
  assign n39533 = n39404 & n78243 ;
  assign n39534 = n39532 | n39533 ;
  assign n39535 = n67905 & n39534 ;
  assign n39536 = n78235 & n39535 ;
  assign n39537 = n39531 | n39536 ;
  assign n39538 = n67222 & n39537 ;
  assign n39539 = n39105 & n39439 ;
  assign n39398 = n39114 | n39397 ;
  assign n78244 = ~n39398 ;
  assign n39540 = n39394 & n78244 ;
  assign n78245 = ~n39399 ;
  assign n39541 = n39397 & n78245 ;
  assign n39542 = n39540 | n39541 ;
  assign n39543 = n67905 & n39542 ;
  assign n39544 = n78235 & n39543 ;
  assign n39545 = n39539 | n39544 ;
  assign n39546 = n67164 & n39545 ;
  assign n39547 = n39113 & n39439 ;
  assign n39393 = n39122 | n39392 ;
  assign n78246 = ~n39393 ;
  assign n39548 = n78246 & n39486 ;
  assign n78247 = ~n39487 ;
  assign n39549 = n39392 & n78247 ;
  assign n39550 = n39548 | n39549 ;
  assign n39551 = n67905 & n39550 ;
  assign n39552 = n78235 & n39551 ;
  assign n39553 = n39547 | n39552 ;
  assign n39554 = n66979 & n39553 ;
  assign n39555 = n39121 & n39439 ;
  assign n39386 = n39130 | n39385 ;
  assign n78248 = ~n39386 ;
  assign n39556 = n39382 & n78248 ;
  assign n78249 = ~n39387 ;
  assign n39557 = n39385 & n78249 ;
  assign n39558 = n39556 | n39557 ;
  assign n39559 = n67905 & n39558 ;
  assign n39560 = n78235 & n39559 ;
  assign n39561 = n39555 | n39560 ;
  assign n39562 = n66868 & n39561 ;
  assign n39563 = n39129 & n39439 ;
  assign n39381 = n39138 | n39380 ;
  assign n78250 = ~n39381 ;
  assign n39564 = n78250 & n39482 ;
  assign n78251 = ~n39483 ;
  assign n39565 = n39380 & n78251 ;
  assign n39566 = n39564 | n39565 ;
  assign n39567 = n67905 & n39566 ;
  assign n39568 = n78235 & n39567 ;
  assign n39569 = n39563 | n39568 ;
  assign n39570 = n66797 & n39569 ;
  assign n39571 = n39137 & n39439 ;
  assign n39374 = n39146 | n39373 ;
  assign n78252 = ~n39374 ;
  assign n39572 = n39370 & n78252 ;
  assign n78253 = ~n39375 ;
  assign n39573 = n39373 & n78253 ;
  assign n39574 = n39572 | n39573 ;
  assign n39575 = n67905 & n39574 ;
  assign n39576 = n78235 & n39575 ;
  assign n39577 = n39571 | n39576 ;
  assign n39578 = n66654 & n39577 ;
  assign n39579 = n39145 & n39439 ;
  assign n39369 = n39154 | n39368 ;
  assign n78254 = ~n39369 ;
  assign n39580 = n78254 & n39478 ;
  assign n78255 = ~n39479 ;
  assign n39581 = n39368 & n78255 ;
  assign n39582 = n39580 | n39581 ;
  assign n39583 = n67905 & n39582 ;
  assign n39584 = n78235 & n39583 ;
  assign n39585 = n39579 | n39584 ;
  assign n39586 = n66560 & n39585 ;
  assign n39587 = n39153 & n39439 ;
  assign n39362 = n39162 | n39361 ;
  assign n78256 = ~n39362 ;
  assign n39588 = n39358 & n78256 ;
  assign n78257 = ~n39363 ;
  assign n39589 = n39361 & n78257 ;
  assign n39590 = n39588 | n39589 ;
  assign n39591 = n67905 & n39590 ;
  assign n39592 = n78235 & n39591 ;
  assign n39593 = n39587 | n39592 ;
  assign n39594 = n66505 & n39593 ;
  assign n39595 = n39161 & n39439 ;
  assign n39357 = n39170 | n39356 ;
  assign n78258 = ~n39357 ;
  assign n39596 = n78258 & n39474 ;
  assign n78259 = ~n39475 ;
  assign n39597 = n39356 & n78259 ;
  assign n39598 = n39596 | n39597 ;
  assign n39599 = n67905 & n39598 ;
  assign n39600 = n78235 & n39599 ;
  assign n39601 = n39595 | n39600 ;
  assign n39602 = n66379 & n39601 ;
  assign n39603 = n39169 & n39439 ;
  assign n39350 = n39178 | n39349 ;
  assign n78260 = ~n39350 ;
  assign n39604 = n39346 & n78260 ;
  assign n78261 = ~n39351 ;
  assign n39605 = n39349 & n78261 ;
  assign n39606 = n39604 | n39605 ;
  assign n39607 = n67905 & n39606 ;
  assign n39608 = n78235 & n39607 ;
  assign n39609 = n39603 | n39608 ;
  assign n39610 = n66299 & n39609 ;
  assign n39611 = n39177 & n39439 ;
  assign n39345 = n39186 | n39344 ;
  assign n78262 = ~n39345 ;
  assign n39612 = n78262 & n39470 ;
  assign n78263 = ~n39471 ;
  assign n39613 = n39344 & n78263 ;
  assign n39614 = n39612 | n39613 ;
  assign n39615 = n67905 & n39614 ;
  assign n39616 = n78235 & n39615 ;
  assign n39617 = n39611 | n39616 ;
  assign n39618 = n66244 & n39617 ;
  assign n39619 = n39185 & n39439 ;
  assign n39338 = n39194 | n39337 ;
  assign n78264 = ~n39338 ;
  assign n39620 = n39334 & n78264 ;
  assign n78265 = ~n39339 ;
  assign n39621 = n39337 & n78265 ;
  assign n39622 = n39620 | n39621 ;
  assign n39623 = n67905 & n39622 ;
  assign n39624 = n78235 & n39623 ;
  assign n39625 = n39619 | n39624 ;
  assign n39626 = n66145 & n39625 ;
  assign n39627 = n39193 & n39439 ;
  assign n39333 = n39202 | n39332 ;
  assign n78266 = ~n39333 ;
  assign n39628 = n78266 & n39466 ;
  assign n78267 = ~n39467 ;
  assign n39629 = n39332 & n78267 ;
  assign n39630 = n39628 | n39629 ;
  assign n39631 = n67905 & n39630 ;
  assign n39632 = n78235 & n39631 ;
  assign n39633 = n39627 | n39632 ;
  assign n39634 = n66081 & n39633 ;
  assign n39635 = n39201 & n39439 ;
  assign n39326 = n39210 | n39325 ;
  assign n78268 = ~n39326 ;
  assign n39636 = n39322 & n78268 ;
  assign n78269 = ~n39327 ;
  assign n39637 = n39325 & n78269 ;
  assign n39638 = n39636 | n39637 ;
  assign n39639 = n67905 & n39638 ;
  assign n39640 = n78235 & n39639 ;
  assign n39641 = n39635 | n39640 ;
  assign n39642 = n66043 & n39641 ;
  assign n39643 = n39209 & n39439 ;
  assign n39321 = n39218 | n39320 ;
  assign n78270 = ~n39321 ;
  assign n39644 = n78270 & n39462 ;
  assign n78271 = ~n39463 ;
  assign n39645 = n39320 & n78271 ;
  assign n39646 = n39644 | n39645 ;
  assign n39647 = n67905 & n39646 ;
  assign n39648 = n78235 & n39647 ;
  assign n39649 = n39643 | n39648 ;
  assign n39650 = n65960 & n39649 ;
  assign n39651 = n39217 & n39439 ;
  assign n39314 = n39225 | n39313 ;
  assign n78272 = ~n39314 ;
  assign n39652 = n39310 & n78272 ;
  assign n78273 = ~n39315 ;
  assign n39653 = n39313 & n78273 ;
  assign n39654 = n39652 | n39653 ;
  assign n39655 = n67905 & n39654 ;
  assign n39656 = n78235 & n39655 ;
  assign n39657 = n39651 | n39656 ;
  assign n39658 = n65909 & n39657 ;
  assign n39659 = n39224 & n39439 ;
  assign n39309 = n39233 | n39308 ;
  assign n78274 = ~n39309 ;
  assign n39660 = n78274 & n39458 ;
  assign n78275 = ~n39459 ;
  assign n39661 = n39308 & n78275 ;
  assign n39662 = n39660 | n39661 ;
  assign n39663 = n67905 & n39662 ;
  assign n39664 = n78235 & n39663 ;
  assign n39665 = n39659 | n39664 ;
  assign n39666 = n65877 & n39665 ;
  assign n39667 = n39232 & n39439 ;
  assign n39302 = n39241 | n39301 ;
  assign n78276 = ~n39302 ;
  assign n39668 = n78276 & n39456 ;
  assign n78277 = ~n39303 ;
  assign n39669 = n39301 & n78277 ;
  assign n39670 = n39668 | n39669 ;
  assign n39671 = n67905 & n39670 ;
  assign n39672 = n78235 & n39671 ;
  assign n39673 = n39667 | n39672 ;
  assign n39674 = n65820 & n39673 ;
  assign n39675 = n39240 & n39439 ;
  assign n39676 = n39248 | n39297 ;
  assign n78278 = ~n39676 ;
  assign n39677 = n39454 & n78278 ;
  assign n78279 = ~n39455 ;
  assign n39678 = n39297 & n78279 ;
  assign n39679 = n39677 | n39678 ;
  assign n39680 = n67905 & n39679 ;
  assign n39681 = n78235 & n39680 ;
  assign n39682 = n39675 | n39681 ;
  assign n39683 = n65791 & n39682 ;
  assign n39684 = n39247 & n39439 ;
  assign n39685 = n39256 | n39291 ;
  assign n78280 = ~n39685 ;
  assign n39686 = n39452 & n78280 ;
  assign n78281 = ~n39292 ;
  assign n39687 = n39291 & n78281 ;
  assign n39688 = n39686 | n39687 ;
  assign n39689 = n67905 & n39688 ;
  assign n39690 = n78235 & n39689 ;
  assign n39691 = n39684 | n39690 ;
  assign n39692 = n65772 & n39691 ;
  assign n39693 = n39255 & n39439 ;
  assign n39694 = n39264 | n39287 ;
  assign n78282 = ~n39694 ;
  assign n39695 = n39450 & n78282 ;
  assign n78283 = ~n39451 ;
  assign n39696 = n39287 & n78283 ;
  assign n39697 = n39695 | n39696 ;
  assign n39698 = n67905 & n39697 ;
  assign n39699 = n78235 & n39698 ;
  assign n39700 = n39693 | n39699 ;
  assign n39701 = n65746 & n39700 ;
  assign n39702 = n39263 & n39439 ;
  assign n78284 = ~n39449 ;
  assign n39703 = n39281 & n78284 ;
  assign n39704 = n39278 | n39281 ;
  assign n78285 = ~n39704 ;
  assign n39705 = n39448 & n78285 ;
  assign n39706 = n39703 | n39705 ;
  assign n39707 = n67905 & n39706 ;
  assign n39708 = n78235 & n39707 ;
  assign n39709 = n39702 | n39708 ;
  assign n39710 = n65721 & n39709 ;
  assign n39440 = n39271 & n39439 ;
  assign n39276 = n6907 & n39274 ;
  assign n39711 = n39276 & n78230 ;
  assign n39712 = n7066 | n39711 ;
  assign n78286 = ~n39712 ;
  assign n39713 = n39448 & n78286 ;
  assign n39714 = n78235 & n39713 ;
  assign n39715 = n39440 | n39714 ;
  assign n39716 = n65686 & n39715 ;
  assign n39717 = n7368 & n78235 ;
  assign n39719 = n78225 & n39718 ;
  assign n39720 = n39435 | n39719 ;
  assign n39721 = n78226 & n39720 ;
  assign n78287 = ~n39721 ;
  assign n39722 = n7363 & n78287 ;
  assign n78288 = ~n39722 ;
  assign n39723 = x35 & n78288 ;
  assign n39724 = n39717 | n39723 ;
  assign n39732 = n65670 & n39724 ;
  assign n39725 = n7363 & n78235 ;
  assign n78289 = ~n39725 ;
  assign n39726 = x35 & n78289 ;
  assign n39727 = n39717 | n39726 ;
  assign n39728 = x65 & n39727 ;
  assign n39729 = x65 | n39717 ;
  assign n39730 = n39726 | n39729 ;
  assign n78290 = ~n39728 ;
  assign n39731 = n78290 & n39730 ;
  assign n39733 = n7375 | n39731 ;
  assign n78291 = ~n39732 ;
  assign n39734 = n78291 & n39733 ;
  assign n78292 = ~n39714 ;
  assign n39735 = x66 & n78292 ;
  assign n78293 = ~n39440 ;
  assign n39736 = n78293 & n39735 ;
  assign n39737 = n39734 | n39736 ;
  assign n78294 = ~n39716 ;
  assign n39738 = n78294 & n39737 ;
  assign n78295 = ~n39708 ;
  assign n39739 = x67 & n78295 ;
  assign n78296 = ~n39702 ;
  assign n39740 = n78296 & n39739 ;
  assign n39741 = n39710 | n39740 ;
  assign n39742 = n39738 | n39741 ;
  assign n78297 = ~n39710 ;
  assign n39743 = n78297 & n39742 ;
  assign n78298 = ~n39699 ;
  assign n39744 = x68 & n78298 ;
  assign n78299 = ~n39693 ;
  assign n39745 = n78299 & n39744 ;
  assign n39746 = n39701 | n39745 ;
  assign n39747 = n39743 | n39746 ;
  assign n78300 = ~n39701 ;
  assign n39748 = n78300 & n39747 ;
  assign n78301 = ~n39690 ;
  assign n39749 = x69 & n78301 ;
  assign n78302 = ~n39684 ;
  assign n39750 = n78302 & n39749 ;
  assign n39751 = n39692 | n39750 ;
  assign n39752 = n39748 | n39751 ;
  assign n78303 = ~n39692 ;
  assign n39753 = n78303 & n39752 ;
  assign n78304 = ~n39681 ;
  assign n39754 = x70 & n78304 ;
  assign n78305 = ~n39675 ;
  assign n39755 = n78305 & n39754 ;
  assign n39756 = n39683 | n39755 ;
  assign n39758 = n39753 | n39756 ;
  assign n78306 = ~n39683 ;
  assign n39759 = n78306 & n39758 ;
  assign n78307 = ~n39672 ;
  assign n39760 = x71 & n78307 ;
  assign n78308 = ~n39667 ;
  assign n39761 = n78308 & n39760 ;
  assign n39762 = n39674 | n39761 ;
  assign n39763 = n39759 | n39762 ;
  assign n78309 = ~n39674 ;
  assign n39764 = n78309 & n39763 ;
  assign n78310 = ~n39664 ;
  assign n39765 = x72 & n78310 ;
  assign n78311 = ~n39659 ;
  assign n39766 = n78311 & n39765 ;
  assign n39767 = n39666 | n39766 ;
  assign n39769 = n39764 | n39767 ;
  assign n78312 = ~n39666 ;
  assign n39770 = n78312 & n39769 ;
  assign n78313 = ~n39656 ;
  assign n39771 = x73 & n78313 ;
  assign n78314 = ~n39651 ;
  assign n39772 = n78314 & n39771 ;
  assign n39773 = n39658 | n39772 ;
  assign n39774 = n39770 | n39773 ;
  assign n78315 = ~n39658 ;
  assign n39775 = n78315 & n39774 ;
  assign n78316 = ~n39648 ;
  assign n39776 = x74 & n78316 ;
  assign n78317 = ~n39643 ;
  assign n39777 = n78317 & n39776 ;
  assign n39778 = n39650 | n39777 ;
  assign n39780 = n39775 | n39778 ;
  assign n78318 = ~n39650 ;
  assign n39781 = n78318 & n39780 ;
  assign n78319 = ~n39640 ;
  assign n39782 = x75 & n78319 ;
  assign n78320 = ~n39635 ;
  assign n39783 = n78320 & n39782 ;
  assign n39784 = n39642 | n39783 ;
  assign n39785 = n39781 | n39784 ;
  assign n78321 = ~n39642 ;
  assign n39786 = n78321 & n39785 ;
  assign n78322 = ~n39632 ;
  assign n39787 = x76 & n78322 ;
  assign n78323 = ~n39627 ;
  assign n39788 = n78323 & n39787 ;
  assign n39789 = n39634 | n39788 ;
  assign n39791 = n39786 | n39789 ;
  assign n78324 = ~n39634 ;
  assign n39792 = n78324 & n39791 ;
  assign n78325 = ~n39624 ;
  assign n39793 = x77 & n78325 ;
  assign n78326 = ~n39619 ;
  assign n39794 = n78326 & n39793 ;
  assign n39795 = n39626 | n39794 ;
  assign n39796 = n39792 | n39795 ;
  assign n78327 = ~n39626 ;
  assign n39797 = n78327 & n39796 ;
  assign n78328 = ~n39616 ;
  assign n39798 = x78 & n78328 ;
  assign n78329 = ~n39611 ;
  assign n39799 = n78329 & n39798 ;
  assign n39800 = n39618 | n39799 ;
  assign n39802 = n39797 | n39800 ;
  assign n78330 = ~n39618 ;
  assign n39803 = n78330 & n39802 ;
  assign n78331 = ~n39608 ;
  assign n39804 = x79 & n78331 ;
  assign n78332 = ~n39603 ;
  assign n39805 = n78332 & n39804 ;
  assign n39806 = n39610 | n39805 ;
  assign n39807 = n39803 | n39806 ;
  assign n78333 = ~n39610 ;
  assign n39808 = n78333 & n39807 ;
  assign n78334 = ~n39600 ;
  assign n39809 = x80 & n78334 ;
  assign n78335 = ~n39595 ;
  assign n39810 = n78335 & n39809 ;
  assign n39811 = n39602 | n39810 ;
  assign n39813 = n39808 | n39811 ;
  assign n78336 = ~n39602 ;
  assign n39814 = n78336 & n39813 ;
  assign n78337 = ~n39592 ;
  assign n39815 = x81 & n78337 ;
  assign n78338 = ~n39587 ;
  assign n39816 = n78338 & n39815 ;
  assign n39817 = n39594 | n39816 ;
  assign n39818 = n39814 | n39817 ;
  assign n78339 = ~n39594 ;
  assign n39819 = n78339 & n39818 ;
  assign n78340 = ~n39584 ;
  assign n39820 = x82 & n78340 ;
  assign n78341 = ~n39579 ;
  assign n39821 = n78341 & n39820 ;
  assign n39822 = n39586 | n39821 ;
  assign n39824 = n39819 | n39822 ;
  assign n78342 = ~n39586 ;
  assign n39825 = n78342 & n39824 ;
  assign n78343 = ~n39576 ;
  assign n39826 = x83 & n78343 ;
  assign n78344 = ~n39571 ;
  assign n39827 = n78344 & n39826 ;
  assign n39828 = n39578 | n39827 ;
  assign n39829 = n39825 | n39828 ;
  assign n78345 = ~n39578 ;
  assign n39830 = n78345 & n39829 ;
  assign n78346 = ~n39568 ;
  assign n39831 = x84 & n78346 ;
  assign n78347 = ~n39563 ;
  assign n39832 = n78347 & n39831 ;
  assign n39833 = n39570 | n39832 ;
  assign n39835 = n39830 | n39833 ;
  assign n78348 = ~n39570 ;
  assign n39836 = n78348 & n39835 ;
  assign n78349 = ~n39560 ;
  assign n39837 = x85 & n78349 ;
  assign n78350 = ~n39555 ;
  assign n39838 = n78350 & n39837 ;
  assign n39839 = n39562 | n39838 ;
  assign n39840 = n39836 | n39839 ;
  assign n78351 = ~n39562 ;
  assign n39841 = n78351 & n39840 ;
  assign n78352 = ~n39552 ;
  assign n39842 = x86 & n78352 ;
  assign n78353 = ~n39547 ;
  assign n39843 = n78353 & n39842 ;
  assign n39844 = n39554 | n39843 ;
  assign n39846 = n39841 | n39844 ;
  assign n78354 = ~n39554 ;
  assign n39847 = n78354 & n39846 ;
  assign n78355 = ~n39544 ;
  assign n39848 = x87 & n78355 ;
  assign n78356 = ~n39539 ;
  assign n39849 = n78356 & n39848 ;
  assign n39850 = n39546 | n39849 ;
  assign n39851 = n39847 | n39850 ;
  assign n78357 = ~n39546 ;
  assign n39852 = n78357 & n39851 ;
  assign n78358 = ~n39536 ;
  assign n39853 = x88 & n78358 ;
  assign n78359 = ~n39531 ;
  assign n39854 = n78359 & n39853 ;
  assign n39855 = n39538 | n39854 ;
  assign n39857 = n39852 | n39855 ;
  assign n78360 = ~n39538 ;
  assign n39858 = n78360 & n39857 ;
  assign n78361 = ~n39528 ;
  assign n39859 = x89 & n78361 ;
  assign n78362 = ~n39523 ;
  assign n39860 = n78362 & n39859 ;
  assign n39861 = n39530 | n39860 ;
  assign n39862 = n39858 | n39861 ;
  assign n78363 = ~n39530 ;
  assign n39863 = n78363 & n39862 ;
  assign n78364 = ~n39520 ;
  assign n39864 = x90 & n78364 ;
  assign n78365 = ~n39515 ;
  assign n39865 = n78365 & n39864 ;
  assign n39866 = n39522 | n39865 ;
  assign n39868 = n39863 | n39866 ;
  assign n78366 = ~n39522 ;
  assign n39869 = n78366 & n39868 ;
  assign n78367 = ~n39512 ;
  assign n39870 = x91 & n78367 ;
  assign n78368 = ~n39507 ;
  assign n39871 = n78368 & n39870 ;
  assign n39872 = n39514 | n39871 ;
  assign n39873 = n39869 | n39872 ;
  assign n78369 = ~n39514 ;
  assign n39874 = n78369 & n39873 ;
  assign n78370 = ~n39504 ;
  assign n39875 = x92 & n78370 ;
  assign n78371 = ~n39442 ;
  assign n39876 = n78371 & n39875 ;
  assign n39877 = n39506 | n39876 ;
  assign n39879 = n39874 | n39877 ;
  assign n78372 = ~n39506 ;
  assign n39880 = n78372 & n39879 ;
  assign n39887 = n67986 & n39886 ;
  assign n78373 = ~n39439 ;
  assign n39888 = n78373 & n39884 ;
  assign n39889 = n39064 & n39439 ;
  assign n78374 = ~n39889 ;
  assign n39890 = x93 & n78374 ;
  assign n78375 = ~n39888 ;
  assign n39891 = n78375 & n39890 ;
  assign n39892 = n7527 | n39891 ;
  assign n39893 = n39887 | n39892 ;
  assign n39895 = n39880 | n39893 ;
  assign n78376 = ~n39894 ;
  assign n39896 = n78376 & n39895 ;
  assign n78377 = ~n39874 ;
  assign n39878 = n78377 & n39877 ;
  assign n39899 = x65 & n39724 ;
  assign n78378 = ~n39899 ;
  assign n39900 = n39730 & n78378 ;
  assign n39901 = n7375 | n39900 ;
  assign n39902 = n78291 & n39901 ;
  assign n39903 = n39716 | n39736 ;
  assign n39905 = n39902 | n39903 ;
  assign n39906 = n78294 & n39905 ;
  assign n39907 = n39740 | n39906 ;
  assign n39909 = n78297 & n39907 ;
  assign n39911 = n39746 | n39909 ;
  assign n39912 = n78300 & n39911 ;
  assign n39914 = n39751 | n39912 ;
  assign n39915 = n78303 & n39914 ;
  assign n39916 = n39756 | n39915 ;
  assign n39917 = n78306 & n39916 ;
  assign n39918 = n39762 | n39917 ;
  assign n39920 = n78309 & n39918 ;
  assign n39921 = n39767 | n39920 ;
  assign n39922 = n78312 & n39921 ;
  assign n39923 = n39773 | n39922 ;
  assign n39925 = n78315 & n39923 ;
  assign n39926 = n39778 | n39925 ;
  assign n39927 = n78318 & n39926 ;
  assign n39928 = n39784 | n39927 ;
  assign n39930 = n78321 & n39928 ;
  assign n39931 = n39789 | n39930 ;
  assign n39932 = n78324 & n39931 ;
  assign n39933 = n39795 | n39932 ;
  assign n39935 = n78327 & n39933 ;
  assign n39936 = n39800 | n39935 ;
  assign n39937 = n78330 & n39936 ;
  assign n39938 = n39806 | n39937 ;
  assign n39940 = n78333 & n39938 ;
  assign n39941 = n39811 | n39940 ;
  assign n39942 = n78336 & n39941 ;
  assign n39943 = n39817 | n39942 ;
  assign n39945 = n78339 & n39943 ;
  assign n39946 = n39822 | n39945 ;
  assign n39947 = n78342 & n39946 ;
  assign n39948 = n39828 | n39947 ;
  assign n39950 = n78345 & n39948 ;
  assign n39951 = n39833 | n39950 ;
  assign n39952 = n78348 & n39951 ;
  assign n39953 = n39839 | n39952 ;
  assign n39955 = n78351 & n39953 ;
  assign n39956 = n39844 | n39955 ;
  assign n39957 = n78354 & n39956 ;
  assign n39958 = n39850 | n39957 ;
  assign n39960 = n78357 & n39958 ;
  assign n39961 = n39855 | n39960 ;
  assign n39962 = n78360 & n39961 ;
  assign n39963 = n39861 | n39962 ;
  assign n39965 = n78363 & n39963 ;
  assign n39966 = n39866 | n39965 ;
  assign n39967 = n78366 & n39966 ;
  assign n39968 = n39872 | n39967 ;
  assign n39970 = n39514 | n39877 ;
  assign n78379 = ~n39970 ;
  assign n39971 = n39968 & n78379 ;
  assign n39972 = n39878 | n39971 ;
  assign n78380 = ~n39896 ;
  assign n39973 = n78380 & n39972 ;
  assign n39974 = n78369 & n39968 ;
  assign n39975 = n39877 | n39974 ;
  assign n39976 = n78372 & n39975 ;
  assign n39977 = n39893 | n39976 ;
  assign n39978 = n39505 & n78376 ;
  assign n39979 = n39977 & n39978 ;
  assign n39980 = n39973 | n39979 ;
  assign n39981 = n39506 | n39891 ;
  assign n39982 = n39887 | n39981 ;
  assign n78381 = ~n39982 ;
  assign n39983 = n39879 & n78381 ;
  assign n39984 = n39887 | n39891 ;
  assign n78382 = ~n39976 ;
  assign n39985 = n78382 & n39984 ;
  assign n39986 = n39983 | n39985 ;
  assign n39987 = n78380 & n39986 ;
  assign n39988 = n7066 & n39064 ;
  assign n39989 = n39977 & n39988 ;
  assign n39990 = n39987 | n39989 ;
  assign n39991 = n68058 & n39990 ;
  assign n78383 = ~n39989 ;
  assign n40386 = x94 & n78383 ;
  assign n78384 = ~n39987 ;
  assign n40387 = n78384 & n40386 ;
  assign n40388 = n39991 | n40387 ;
  assign n39992 = n67986 & n39980 ;
  assign n78385 = ~n39967 ;
  assign n39969 = n39872 & n78385 ;
  assign n39993 = n39522 | n39872 ;
  assign n78386 = ~n39993 ;
  assign n39994 = n39868 & n78386 ;
  assign n39995 = n39969 | n39994 ;
  assign n39996 = n78380 & n39995 ;
  assign n39997 = n39513 & n78376 ;
  assign n39998 = n39977 & n39997 ;
  assign n39999 = n39996 | n39998 ;
  assign n40000 = n67763 & n39999 ;
  assign n78387 = ~n39998 ;
  assign n40374 = x92 & n78387 ;
  assign n78388 = ~n39996 ;
  assign n40375 = n78388 & n40374 ;
  assign n40376 = n40000 | n40375 ;
  assign n78389 = ~n39863 ;
  assign n39867 = n78389 & n39866 ;
  assign n40001 = n39530 | n39866 ;
  assign n78390 = ~n40001 ;
  assign n40002 = n39963 & n78390 ;
  assign n40003 = n39867 | n40002 ;
  assign n40004 = n78380 & n40003 ;
  assign n40005 = n39521 & n78376 ;
  assign n40006 = n39977 & n40005 ;
  assign n40007 = n40004 | n40006 ;
  assign n40008 = n67622 & n40007 ;
  assign n78391 = ~n39962 ;
  assign n39964 = n39861 & n78391 ;
  assign n40009 = n39538 | n39861 ;
  assign n78392 = ~n40009 ;
  assign n40010 = n39857 & n78392 ;
  assign n40011 = n39964 | n40010 ;
  assign n40012 = n78380 & n40011 ;
  assign n40013 = n39529 & n78376 ;
  assign n40014 = n39977 & n40013 ;
  assign n40015 = n40012 | n40014 ;
  assign n40016 = n67531 & n40015 ;
  assign n78393 = ~n40014 ;
  assign n40362 = x90 & n78393 ;
  assign n78394 = ~n40012 ;
  assign n40363 = n78394 & n40362 ;
  assign n40364 = n40016 | n40363 ;
  assign n78395 = ~n39852 ;
  assign n39856 = n78395 & n39855 ;
  assign n40017 = n39546 | n39855 ;
  assign n78396 = ~n40017 ;
  assign n40018 = n39958 & n78396 ;
  assign n40019 = n39856 | n40018 ;
  assign n40020 = n78380 & n40019 ;
  assign n40021 = n39537 & n78376 ;
  assign n40022 = n39977 & n40021 ;
  assign n40023 = n40020 | n40022 ;
  assign n40024 = n67348 & n40023 ;
  assign n78397 = ~n39957 ;
  assign n39959 = n39850 & n78397 ;
  assign n40025 = n39554 | n39850 ;
  assign n78398 = ~n40025 ;
  assign n40026 = n39846 & n78398 ;
  assign n40027 = n39959 | n40026 ;
  assign n40028 = n78380 & n40027 ;
  assign n40029 = n39545 & n78376 ;
  assign n40030 = n39977 & n40029 ;
  assign n40031 = n40028 | n40030 ;
  assign n40032 = n67222 & n40031 ;
  assign n78399 = ~n40030 ;
  assign n40350 = x88 & n78399 ;
  assign n78400 = ~n40028 ;
  assign n40351 = n78400 & n40350 ;
  assign n40352 = n40032 | n40351 ;
  assign n78401 = ~n39841 ;
  assign n39845 = n78401 & n39844 ;
  assign n40033 = n39562 | n39844 ;
  assign n78402 = ~n40033 ;
  assign n40034 = n39953 & n78402 ;
  assign n40035 = n39845 | n40034 ;
  assign n40036 = n78380 & n40035 ;
  assign n40037 = n39553 & n78376 ;
  assign n40038 = n39977 & n40037 ;
  assign n40039 = n40036 | n40038 ;
  assign n40040 = n67164 & n40039 ;
  assign n78403 = ~n39952 ;
  assign n39954 = n39839 & n78403 ;
  assign n40041 = n39570 | n39839 ;
  assign n78404 = ~n40041 ;
  assign n40042 = n39835 & n78404 ;
  assign n40043 = n39954 | n40042 ;
  assign n40044 = n78380 & n40043 ;
  assign n40045 = n39561 & n78376 ;
  assign n40046 = n39977 & n40045 ;
  assign n40047 = n40044 | n40046 ;
  assign n40048 = n66979 & n40047 ;
  assign n78405 = ~n40046 ;
  assign n40338 = x86 & n78405 ;
  assign n78406 = ~n40044 ;
  assign n40339 = n78406 & n40338 ;
  assign n40340 = n40048 | n40339 ;
  assign n78407 = ~n39830 ;
  assign n39834 = n78407 & n39833 ;
  assign n40049 = n39578 | n39833 ;
  assign n78408 = ~n40049 ;
  assign n40050 = n39948 & n78408 ;
  assign n40051 = n39834 | n40050 ;
  assign n40052 = n78380 & n40051 ;
  assign n40053 = n39569 & n78376 ;
  assign n40054 = n39977 & n40053 ;
  assign n40055 = n40052 | n40054 ;
  assign n40056 = n66868 & n40055 ;
  assign n78409 = ~n39947 ;
  assign n39949 = n39828 & n78409 ;
  assign n40057 = n39586 | n39828 ;
  assign n78410 = ~n40057 ;
  assign n40058 = n39824 & n78410 ;
  assign n40059 = n39949 | n40058 ;
  assign n40060 = n78380 & n40059 ;
  assign n40061 = n39577 & n78376 ;
  assign n40062 = n39977 & n40061 ;
  assign n40063 = n40060 | n40062 ;
  assign n40064 = n66797 & n40063 ;
  assign n78411 = ~n40062 ;
  assign n40326 = x84 & n78411 ;
  assign n78412 = ~n40060 ;
  assign n40327 = n78412 & n40326 ;
  assign n40328 = n40064 | n40327 ;
  assign n78413 = ~n39819 ;
  assign n39823 = n78413 & n39822 ;
  assign n40065 = n39594 | n39822 ;
  assign n78414 = ~n40065 ;
  assign n40066 = n39943 & n78414 ;
  assign n40067 = n39823 | n40066 ;
  assign n40068 = n78380 & n40067 ;
  assign n40069 = n39585 & n78376 ;
  assign n40070 = n39977 & n40069 ;
  assign n40071 = n40068 | n40070 ;
  assign n40072 = n66654 & n40071 ;
  assign n78415 = ~n39942 ;
  assign n39944 = n39817 & n78415 ;
  assign n40073 = n39602 | n39817 ;
  assign n78416 = ~n40073 ;
  assign n40074 = n39813 & n78416 ;
  assign n40075 = n39944 | n40074 ;
  assign n40076 = n78380 & n40075 ;
  assign n40077 = n39593 & n78376 ;
  assign n40078 = n39977 & n40077 ;
  assign n40079 = n40076 | n40078 ;
  assign n40080 = n66560 & n40079 ;
  assign n78417 = ~n40078 ;
  assign n40314 = x82 & n78417 ;
  assign n78418 = ~n40076 ;
  assign n40315 = n78418 & n40314 ;
  assign n40316 = n40080 | n40315 ;
  assign n78419 = ~n39808 ;
  assign n39812 = n78419 & n39811 ;
  assign n40081 = n39610 | n39811 ;
  assign n78420 = ~n40081 ;
  assign n40082 = n39938 & n78420 ;
  assign n40083 = n39812 | n40082 ;
  assign n40084 = n78380 & n40083 ;
  assign n40085 = n39601 & n78376 ;
  assign n40086 = n39977 & n40085 ;
  assign n40087 = n40084 | n40086 ;
  assign n40088 = n66505 & n40087 ;
  assign n78421 = ~n39937 ;
  assign n39939 = n39806 & n78421 ;
  assign n40089 = n39618 | n39806 ;
  assign n78422 = ~n40089 ;
  assign n40090 = n39802 & n78422 ;
  assign n40091 = n39939 | n40090 ;
  assign n40092 = n78380 & n40091 ;
  assign n40093 = n39609 & n78376 ;
  assign n40094 = n39977 & n40093 ;
  assign n40095 = n40092 | n40094 ;
  assign n40096 = n66379 & n40095 ;
  assign n78423 = ~n40094 ;
  assign n40302 = x80 & n78423 ;
  assign n78424 = ~n40092 ;
  assign n40303 = n78424 & n40302 ;
  assign n40304 = n40096 | n40303 ;
  assign n78425 = ~n39797 ;
  assign n39801 = n78425 & n39800 ;
  assign n40097 = n39626 | n39800 ;
  assign n78426 = ~n40097 ;
  assign n40098 = n39933 & n78426 ;
  assign n40099 = n39801 | n40098 ;
  assign n40100 = n78380 & n40099 ;
  assign n40101 = n39617 & n78376 ;
  assign n40102 = n39977 & n40101 ;
  assign n40103 = n40100 | n40102 ;
  assign n40104 = n66299 & n40103 ;
  assign n78427 = ~n39932 ;
  assign n39934 = n39795 & n78427 ;
  assign n40105 = n39634 | n39795 ;
  assign n78428 = ~n40105 ;
  assign n40106 = n39791 & n78428 ;
  assign n40107 = n39934 | n40106 ;
  assign n40108 = n78380 & n40107 ;
  assign n40109 = n39625 & n78376 ;
  assign n40110 = n39977 & n40109 ;
  assign n40111 = n40108 | n40110 ;
  assign n40112 = n66244 & n40111 ;
  assign n78429 = ~n40110 ;
  assign n40290 = x78 & n78429 ;
  assign n78430 = ~n40108 ;
  assign n40291 = n78430 & n40290 ;
  assign n40292 = n40112 | n40291 ;
  assign n78431 = ~n39786 ;
  assign n39790 = n78431 & n39789 ;
  assign n40113 = n39642 | n39789 ;
  assign n78432 = ~n40113 ;
  assign n40114 = n39928 & n78432 ;
  assign n40115 = n39790 | n40114 ;
  assign n40116 = n78380 & n40115 ;
  assign n40117 = n39633 & n78376 ;
  assign n40118 = n39977 & n40117 ;
  assign n40119 = n40116 | n40118 ;
  assign n40120 = n66145 & n40119 ;
  assign n78433 = ~n39927 ;
  assign n39929 = n39784 & n78433 ;
  assign n40121 = n39650 | n39784 ;
  assign n78434 = ~n40121 ;
  assign n40122 = n39780 & n78434 ;
  assign n40123 = n39929 | n40122 ;
  assign n40124 = n78380 & n40123 ;
  assign n40125 = n39641 & n78376 ;
  assign n40126 = n39977 & n40125 ;
  assign n40127 = n40124 | n40126 ;
  assign n40128 = n66081 & n40127 ;
  assign n78435 = ~n40126 ;
  assign n40278 = x76 & n78435 ;
  assign n78436 = ~n40124 ;
  assign n40279 = n78436 & n40278 ;
  assign n40280 = n40128 | n40279 ;
  assign n78437 = ~n39775 ;
  assign n39779 = n78437 & n39778 ;
  assign n40129 = n39658 | n39778 ;
  assign n78438 = ~n40129 ;
  assign n40130 = n39923 & n78438 ;
  assign n40131 = n39779 | n40130 ;
  assign n40132 = n78380 & n40131 ;
  assign n40133 = n39649 & n78376 ;
  assign n40134 = n39977 & n40133 ;
  assign n40135 = n40132 | n40134 ;
  assign n40136 = n66043 & n40135 ;
  assign n78439 = ~n39922 ;
  assign n39924 = n39773 & n78439 ;
  assign n40137 = n39666 | n39773 ;
  assign n78440 = ~n40137 ;
  assign n40138 = n39769 & n78440 ;
  assign n40139 = n39924 | n40138 ;
  assign n40140 = n78380 & n40139 ;
  assign n40141 = n39657 & n78376 ;
  assign n40142 = n39977 & n40141 ;
  assign n40143 = n40140 | n40142 ;
  assign n40144 = n65960 & n40143 ;
  assign n78441 = ~n40142 ;
  assign n40266 = x74 & n78441 ;
  assign n78442 = ~n40140 ;
  assign n40267 = n78442 & n40266 ;
  assign n40268 = n40144 | n40267 ;
  assign n78443 = ~n39764 ;
  assign n39768 = n78443 & n39767 ;
  assign n40145 = n39674 | n39767 ;
  assign n78444 = ~n40145 ;
  assign n40146 = n39918 & n78444 ;
  assign n40147 = n39768 | n40146 ;
  assign n40148 = n78380 & n40147 ;
  assign n40149 = n39665 & n78376 ;
  assign n40150 = n39977 & n40149 ;
  assign n40151 = n40148 | n40150 ;
  assign n40152 = n65909 & n40151 ;
  assign n78445 = ~n39917 ;
  assign n39919 = n39762 & n78445 ;
  assign n40153 = n39683 | n39762 ;
  assign n78446 = ~n40153 ;
  assign n40154 = n39758 & n78446 ;
  assign n40155 = n39919 | n40154 ;
  assign n40156 = n78380 & n40155 ;
  assign n40157 = n39673 & n78376 ;
  assign n40158 = n39977 & n40157 ;
  assign n40159 = n40156 | n40158 ;
  assign n40160 = n65877 & n40159 ;
  assign n78447 = ~n40158 ;
  assign n40254 = x72 & n78447 ;
  assign n78448 = ~n40156 ;
  assign n40255 = n78448 & n40254 ;
  assign n40256 = n40160 | n40255 ;
  assign n78449 = ~n39753 ;
  assign n39757 = n78449 & n39756 ;
  assign n40161 = n39692 | n39756 ;
  assign n78450 = ~n40161 ;
  assign n40162 = n39914 & n78450 ;
  assign n40163 = n39757 | n40162 ;
  assign n40164 = n78380 & n40163 ;
  assign n40165 = n39682 & n78376 ;
  assign n40166 = n39977 & n40165 ;
  assign n40167 = n40164 | n40166 ;
  assign n40168 = n65820 & n40167 ;
  assign n78451 = ~n39912 ;
  assign n39913 = n39751 & n78451 ;
  assign n40169 = n39701 | n39751 ;
  assign n78452 = ~n40169 ;
  assign n40170 = n39747 & n78452 ;
  assign n40171 = n39913 | n40170 ;
  assign n40172 = n78380 & n40171 ;
  assign n40173 = n39691 & n78376 ;
  assign n40174 = n39977 & n40173 ;
  assign n40175 = n40172 | n40174 ;
  assign n40176 = n65791 & n40175 ;
  assign n78453 = ~n40174 ;
  assign n40242 = x70 & n78453 ;
  assign n78454 = ~n40172 ;
  assign n40243 = n78454 & n40242 ;
  assign n40244 = n40176 | n40243 ;
  assign n78455 = ~n39743 ;
  assign n39910 = n78455 & n39746 ;
  assign n40177 = n39741 | n39906 ;
  assign n40178 = n39710 | n39746 ;
  assign n78456 = ~n40178 ;
  assign n40179 = n40177 & n78456 ;
  assign n40180 = n39910 | n40179 ;
  assign n40181 = n78380 & n40180 ;
  assign n40182 = n39700 & n78376 ;
  assign n40183 = n39977 & n40182 ;
  assign n40184 = n40181 | n40183 ;
  assign n40185 = n65772 & n40184 ;
  assign n78457 = ~n39906 ;
  assign n39908 = n39741 & n78457 ;
  assign n40186 = n39716 | n39741 ;
  assign n78458 = ~n40186 ;
  assign n40187 = n39905 & n78458 ;
  assign n40188 = n39908 | n40187 ;
  assign n40189 = n78380 & n40188 ;
  assign n40190 = n39709 & n78376 ;
  assign n40191 = n39977 & n40190 ;
  assign n40192 = n40189 | n40191 ;
  assign n40193 = n65746 & n40192 ;
  assign n78459 = ~n40191 ;
  assign n40231 = x68 & n78459 ;
  assign n78460 = ~n40189 ;
  assign n40232 = n78460 & n40231 ;
  assign n40233 = n40193 | n40232 ;
  assign n78461 = ~n39734 ;
  assign n39904 = n78461 & n39903 ;
  assign n40194 = n39732 | n39903 ;
  assign n78462 = ~n40194 ;
  assign n40195 = n39733 & n78462 ;
  assign n40196 = n39904 | n40195 ;
  assign n40197 = n78380 & n40196 ;
  assign n40198 = n39715 & n78376 ;
  assign n40199 = n39977 & n40198 ;
  assign n40200 = n40197 | n40199 ;
  assign n40201 = n65721 & n40200 ;
  assign n40202 = n7375 & n39730 ;
  assign n40203 = n78378 & n40202 ;
  assign n78463 = ~n40203 ;
  assign n40204 = n39733 & n78463 ;
  assign n40205 = n78380 & n40204 ;
  assign n40206 = n39724 & n78376 ;
  assign n40207 = n39977 & n40206 ;
  assign n40208 = n40205 | n40207 ;
  assign n40209 = n65686 & n40208 ;
  assign n78464 = ~n40207 ;
  assign n40221 = x66 & n78464 ;
  assign n78465 = ~n40205 ;
  assign n40222 = n78465 & n40221 ;
  assign n40223 = n40209 | n40222 ;
  assign n39897 = n7375 & n78380 ;
  assign n39898 = x64 & n78380 ;
  assign n78466 = ~n39898 ;
  assign n40210 = x34 & n78466 ;
  assign n40211 = n39897 | n40210 ;
  assign n40212 = x65 & n40211 ;
  assign n40213 = n78376 & n39977 ;
  assign n78467 = ~n40213 ;
  assign n40214 = n7375 & n78467 ;
  assign n40215 = x65 | n40214 ;
  assign n40216 = n40210 | n40215 ;
  assign n78468 = ~n40212 ;
  assign n40217 = n78468 & n40216 ;
  assign n40219 = n7868 | n40217 ;
  assign n40220 = n65670 & n40211 ;
  assign n78469 = ~n40220 ;
  assign n40224 = n40219 & n78469 ;
  assign n40225 = n40223 | n40224 ;
  assign n78470 = ~n40209 ;
  assign n40226 = n78470 & n40225 ;
  assign n78471 = ~n40199 ;
  assign n40227 = x67 & n78471 ;
  assign n78472 = ~n40197 ;
  assign n40228 = n78472 & n40227 ;
  assign n40229 = n40201 | n40228 ;
  assign n40230 = n40226 | n40229 ;
  assign n78473 = ~n40201 ;
  assign n40234 = n78473 & n40230 ;
  assign n40235 = n40233 | n40234 ;
  assign n78474 = ~n40193 ;
  assign n40236 = n78474 & n40235 ;
  assign n78475 = ~n40183 ;
  assign n40237 = x69 & n78475 ;
  assign n78476 = ~n40181 ;
  assign n40238 = n78476 & n40237 ;
  assign n40239 = n40185 | n40238 ;
  assign n40241 = n40236 | n40239 ;
  assign n78477 = ~n40185 ;
  assign n40246 = n78477 & n40241 ;
  assign n40247 = n40244 | n40246 ;
  assign n78478 = ~n40176 ;
  assign n40248 = n78478 & n40247 ;
  assign n78479 = ~n40166 ;
  assign n40249 = x71 & n78479 ;
  assign n78480 = ~n40164 ;
  assign n40250 = n78480 & n40249 ;
  assign n40251 = n40168 | n40250 ;
  assign n40253 = n40248 | n40251 ;
  assign n78481 = ~n40168 ;
  assign n40258 = n78481 & n40253 ;
  assign n40259 = n40256 | n40258 ;
  assign n78482 = ~n40160 ;
  assign n40260 = n78482 & n40259 ;
  assign n78483 = ~n40150 ;
  assign n40261 = x73 & n78483 ;
  assign n78484 = ~n40148 ;
  assign n40262 = n78484 & n40261 ;
  assign n40263 = n40152 | n40262 ;
  assign n40265 = n40260 | n40263 ;
  assign n78485 = ~n40152 ;
  assign n40270 = n78485 & n40265 ;
  assign n40271 = n40268 | n40270 ;
  assign n78486 = ~n40144 ;
  assign n40272 = n78486 & n40271 ;
  assign n78487 = ~n40134 ;
  assign n40273 = x75 & n78487 ;
  assign n78488 = ~n40132 ;
  assign n40274 = n78488 & n40273 ;
  assign n40275 = n40136 | n40274 ;
  assign n40277 = n40272 | n40275 ;
  assign n78489 = ~n40136 ;
  assign n40282 = n78489 & n40277 ;
  assign n40283 = n40280 | n40282 ;
  assign n78490 = ~n40128 ;
  assign n40284 = n78490 & n40283 ;
  assign n78491 = ~n40118 ;
  assign n40285 = x77 & n78491 ;
  assign n78492 = ~n40116 ;
  assign n40286 = n78492 & n40285 ;
  assign n40287 = n40120 | n40286 ;
  assign n40289 = n40284 | n40287 ;
  assign n78493 = ~n40120 ;
  assign n40294 = n78493 & n40289 ;
  assign n40295 = n40292 | n40294 ;
  assign n78494 = ~n40112 ;
  assign n40296 = n78494 & n40295 ;
  assign n78495 = ~n40102 ;
  assign n40297 = x79 & n78495 ;
  assign n78496 = ~n40100 ;
  assign n40298 = n78496 & n40297 ;
  assign n40299 = n40104 | n40298 ;
  assign n40301 = n40296 | n40299 ;
  assign n78497 = ~n40104 ;
  assign n40306 = n78497 & n40301 ;
  assign n40307 = n40304 | n40306 ;
  assign n78498 = ~n40096 ;
  assign n40308 = n78498 & n40307 ;
  assign n78499 = ~n40086 ;
  assign n40309 = x81 & n78499 ;
  assign n78500 = ~n40084 ;
  assign n40310 = n78500 & n40309 ;
  assign n40311 = n40088 | n40310 ;
  assign n40313 = n40308 | n40311 ;
  assign n78501 = ~n40088 ;
  assign n40318 = n78501 & n40313 ;
  assign n40319 = n40316 | n40318 ;
  assign n78502 = ~n40080 ;
  assign n40320 = n78502 & n40319 ;
  assign n78503 = ~n40070 ;
  assign n40321 = x83 & n78503 ;
  assign n78504 = ~n40068 ;
  assign n40322 = n78504 & n40321 ;
  assign n40323 = n40072 | n40322 ;
  assign n40325 = n40320 | n40323 ;
  assign n78505 = ~n40072 ;
  assign n40330 = n78505 & n40325 ;
  assign n40331 = n40328 | n40330 ;
  assign n78506 = ~n40064 ;
  assign n40332 = n78506 & n40331 ;
  assign n78507 = ~n40054 ;
  assign n40333 = x85 & n78507 ;
  assign n78508 = ~n40052 ;
  assign n40334 = n78508 & n40333 ;
  assign n40335 = n40056 | n40334 ;
  assign n40337 = n40332 | n40335 ;
  assign n78509 = ~n40056 ;
  assign n40342 = n78509 & n40337 ;
  assign n40343 = n40340 | n40342 ;
  assign n78510 = ~n40048 ;
  assign n40344 = n78510 & n40343 ;
  assign n78511 = ~n40038 ;
  assign n40345 = x87 & n78511 ;
  assign n78512 = ~n40036 ;
  assign n40346 = n78512 & n40345 ;
  assign n40347 = n40040 | n40346 ;
  assign n40349 = n40344 | n40347 ;
  assign n78513 = ~n40040 ;
  assign n40354 = n78513 & n40349 ;
  assign n40355 = n40352 | n40354 ;
  assign n78514 = ~n40032 ;
  assign n40356 = n78514 & n40355 ;
  assign n78515 = ~n40022 ;
  assign n40357 = x89 & n78515 ;
  assign n78516 = ~n40020 ;
  assign n40358 = n78516 & n40357 ;
  assign n40359 = n40024 | n40358 ;
  assign n40361 = n40356 | n40359 ;
  assign n78517 = ~n40024 ;
  assign n40366 = n78517 & n40361 ;
  assign n40367 = n40364 | n40366 ;
  assign n78518 = ~n40016 ;
  assign n40368 = n78518 & n40367 ;
  assign n78519 = ~n40006 ;
  assign n40369 = x91 & n78519 ;
  assign n78520 = ~n40004 ;
  assign n40370 = n78520 & n40369 ;
  assign n40371 = n40008 | n40370 ;
  assign n40373 = n40368 | n40371 ;
  assign n78521 = ~n40008 ;
  assign n40378 = n78521 & n40373 ;
  assign n40379 = n40376 | n40378 ;
  assign n78522 = ~n40000 ;
  assign n40380 = n78522 & n40379 ;
  assign n78523 = ~n39979 ;
  assign n40381 = x93 & n78523 ;
  assign n78524 = ~n39973 ;
  assign n40382 = n78524 & n40381 ;
  assign n40383 = n39992 | n40382 ;
  assign n40385 = n40380 | n40383 ;
  assign n78525 = ~n39992 ;
  assign n40389 = n78525 & n40385 ;
  assign n40390 = n40388 | n40389 ;
  assign n78526 = ~n39991 ;
  assign n40391 = n78526 & n40390 ;
  assign n40392 = n8032 | n40391 ;
  assign n40395 = n39980 & n40392 ;
  assign n40384 = n40000 | n40383 ;
  assign n40396 = x64 & n78467 ;
  assign n78527 = ~n40396 ;
  assign n40397 = x34 & n78527 ;
  assign n40398 = n39897 | n40397 ;
  assign n40399 = x65 & n40398 ;
  assign n78528 = ~n40399 ;
  assign n40400 = n40216 & n78528 ;
  assign n40401 = n7868 | n40400 ;
  assign n40402 = n78469 & n40401 ;
  assign n40404 = n40223 | n40402 ;
  assign n40405 = n78470 & n40404 ;
  assign n40406 = n40229 | n40405 ;
  assign n40407 = n78473 & n40406 ;
  assign n40408 = n40233 | n40407 ;
  assign n40409 = n78474 & n40408 ;
  assign n40410 = n40239 | n40409 ;
  assign n40411 = n78477 & n40410 ;
  assign n40412 = n40244 | n40411 ;
  assign n40413 = n78478 & n40412 ;
  assign n40414 = n40251 | n40413 ;
  assign n40415 = n78481 & n40414 ;
  assign n40416 = n40256 | n40415 ;
  assign n40417 = n78482 & n40416 ;
  assign n40418 = n40263 | n40417 ;
  assign n40419 = n78485 & n40418 ;
  assign n40420 = n40268 | n40419 ;
  assign n40421 = n78486 & n40420 ;
  assign n40422 = n40275 | n40421 ;
  assign n40423 = n78489 & n40422 ;
  assign n40424 = n40280 | n40423 ;
  assign n40425 = n78490 & n40424 ;
  assign n40426 = n40287 | n40425 ;
  assign n40427 = n78493 & n40426 ;
  assign n40428 = n40292 | n40427 ;
  assign n40429 = n78494 & n40428 ;
  assign n40430 = n40299 | n40429 ;
  assign n40431 = n78497 & n40430 ;
  assign n40432 = n40304 | n40431 ;
  assign n40433 = n78498 & n40432 ;
  assign n40434 = n40311 | n40433 ;
  assign n40435 = n78501 & n40434 ;
  assign n40436 = n40316 | n40435 ;
  assign n40437 = n78502 & n40436 ;
  assign n40438 = n40323 | n40437 ;
  assign n40439 = n78505 & n40438 ;
  assign n40440 = n40328 | n40439 ;
  assign n40441 = n78506 & n40440 ;
  assign n40442 = n40335 | n40441 ;
  assign n40443 = n78509 & n40442 ;
  assign n40444 = n40340 | n40443 ;
  assign n40445 = n78510 & n40444 ;
  assign n40446 = n40347 | n40445 ;
  assign n40447 = n78513 & n40446 ;
  assign n40448 = n40352 | n40447 ;
  assign n40449 = n78514 & n40448 ;
  assign n40450 = n40359 | n40449 ;
  assign n40451 = n78517 & n40450 ;
  assign n40452 = n40364 | n40451 ;
  assign n40453 = n78518 & n40452 ;
  assign n40454 = n40371 | n40453 ;
  assign n40455 = n78521 & n40454 ;
  assign n40456 = n40376 | n40455 ;
  assign n78529 = ~n40384 ;
  assign n40457 = n78529 & n40456 ;
  assign n40458 = n78522 & n40456 ;
  assign n78530 = ~n40458 ;
  assign n40459 = n40383 & n78530 ;
  assign n40460 = n40457 | n40459 ;
  assign n40461 = n68220 & n40460 ;
  assign n78531 = ~n40391 ;
  assign n40462 = n78531 & n40461 ;
  assign n40463 = n40395 | n40462 ;
  assign n78532 = ~n39990 ;
  assign n40393 = n78532 & n40392 ;
  assign n78533 = ~n40389 ;
  assign n40466 = n40388 & n78533 ;
  assign n40464 = n40383 | n40458 ;
  assign n40467 = n39992 | n40388 ;
  assign n78534 = ~n40467 ;
  assign n40468 = n40464 & n78534 ;
  assign n40469 = n40466 | n40468 ;
  assign n40470 = n40392 | n40469 ;
  assign n78535 = ~n40393 ;
  assign n40471 = n78535 & n40470 ;
  assign n40472 = n68214 & n40471 ;
  assign n40473 = n68058 & n40463 ;
  assign n40474 = n39999 & n40392 ;
  assign n40377 = n40008 | n40376 ;
  assign n78536 = ~n40377 ;
  assign n40475 = n40373 & n78536 ;
  assign n78537 = ~n40378 ;
  assign n40476 = n40376 & n78537 ;
  assign n40477 = n40475 | n40476 ;
  assign n40478 = n68220 & n40477 ;
  assign n40479 = n78531 & n40478 ;
  assign n40480 = n40474 | n40479 ;
  assign n40481 = n67986 & n40480 ;
  assign n40482 = n40007 & n40392 ;
  assign n40372 = n40016 | n40371 ;
  assign n78538 = ~n40372 ;
  assign n40483 = n78538 & n40452 ;
  assign n78539 = ~n40453 ;
  assign n40484 = n40371 & n78539 ;
  assign n40485 = n40483 | n40484 ;
  assign n40486 = n68220 & n40485 ;
  assign n40487 = n78531 & n40486 ;
  assign n40488 = n40482 | n40487 ;
  assign n40489 = n67763 & n40488 ;
  assign n40490 = n40015 & n40392 ;
  assign n40365 = n40024 | n40364 ;
  assign n78540 = ~n40365 ;
  assign n40491 = n40361 & n78540 ;
  assign n78541 = ~n40366 ;
  assign n40492 = n40364 & n78541 ;
  assign n40493 = n40491 | n40492 ;
  assign n40494 = n68220 & n40493 ;
  assign n40495 = n78531 & n40494 ;
  assign n40496 = n40490 | n40495 ;
  assign n40497 = n67622 & n40496 ;
  assign n40498 = n40023 & n40392 ;
  assign n40360 = n40032 | n40359 ;
  assign n78542 = ~n40360 ;
  assign n40499 = n78542 & n40448 ;
  assign n78543 = ~n40449 ;
  assign n40500 = n40359 & n78543 ;
  assign n40501 = n40499 | n40500 ;
  assign n40502 = n68220 & n40501 ;
  assign n40503 = n78531 & n40502 ;
  assign n40504 = n40498 | n40503 ;
  assign n40505 = n67531 & n40504 ;
  assign n40506 = n40031 & n40392 ;
  assign n40353 = n40040 | n40352 ;
  assign n78544 = ~n40353 ;
  assign n40507 = n40349 & n78544 ;
  assign n78545 = ~n40354 ;
  assign n40508 = n40352 & n78545 ;
  assign n40509 = n40507 | n40508 ;
  assign n40510 = n68220 & n40509 ;
  assign n40511 = n78531 & n40510 ;
  assign n40512 = n40506 | n40511 ;
  assign n40513 = n67348 & n40512 ;
  assign n40514 = n40039 & n40392 ;
  assign n40348 = n40048 | n40347 ;
  assign n78546 = ~n40348 ;
  assign n40515 = n78546 & n40444 ;
  assign n78547 = ~n40445 ;
  assign n40516 = n40347 & n78547 ;
  assign n40517 = n40515 | n40516 ;
  assign n40518 = n68220 & n40517 ;
  assign n40519 = n78531 & n40518 ;
  assign n40520 = n40514 | n40519 ;
  assign n40521 = n67222 & n40520 ;
  assign n40522 = n40047 & n40392 ;
  assign n40341 = n40056 | n40340 ;
  assign n78548 = ~n40341 ;
  assign n40523 = n40337 & n78548 ;
  assign n78549 = ~n40342 ;
  assign n40524 = n40340 & n78549 ;
  assign n40525 = n40523 | n40524 ;
  assign n40526 = n68220 & n40525 ;
  assign n40527 = n78531 & n40526 ;
  assign n40528 = n40522 | n40527 ;
  assign n40529 = n67164 & n40528 ;
  assign n40530 = n40055 & n40392 ;
  assign n40336 = n40064 | n40335 ;
  assign n78550 = ~n40336 ;
  assign n40531 = n78550 & n40440 ;
  assign n78551 = ~n40441 ;
  assign n40532 = n40335 & n78551 ;
  assign n40533 = n40531 | n40532 ;
  assign n40534 = n68220 & n40533 ;
  assign n40535 = n78531 & n40534 ;
  assign n40536 = n40530 | n40535 ;
  assign n40537 = n66979 & n40536 ;
  assign n40538 = n40063 & n40392 ;
  assign n40329 = n40072 | n40328 ;
  assign n78552 = ~n40329 ;
  assign n40539 = n40325 & n78552 ;
  assign n78553 = ~n40330 ;
  assign n40540 = n40328 & n78553 ;
  assign n40541 = n40539 | n40540 ;
  assign n40542 = n68220 & n40541 ;
  assign n40543 = n78531 & n40542 ;
  assign n40544 = n40538 | n40543 ;
  assign n40545 = n66868 & n40544 ;
  assign n40546 = n40071 & n40392 ;
  assign n40324 = n40080 | n40323 ;
  assign n78554 = ~n40324 ;
  assign n40547 = n78554 & n40436 ;
  assign n78555 = ~n40437 ;
  assign n40548 = n40323 & n78555 ;
  assign n40549 = n40547 | n40548 ;
  assign n40550 = n68220 & n40549 ;
  assign n40551 = n78531 & n40550 ;
  assign n40552 = n40546 | n40551 ;
  assign n40553 = n66797 & n40552 ;
  assign n40554 = n40079 & n40392 ;
  assign n40317 = n40088 | n40316 ;
  assign n78556 = ~n40317 ;
  assign n40555 = n40313 & n78556 ;
  assign n78557 = ~n40318 ;
  assign n40556 = n40316 & n78557 ;
  assign n40557 = n40555 | n40556 ;
  assign n40558 = n68220 & n40557 ;
  assign n40559 = n78531 & n40558 ;
  assign n40560 = n40554 | n40559 ;
  assign n40561 = n66654 & n40560 ;
  assign n40562 = n40087 & n40392 ;
  assign n40312 = n40096 | n40311 ;
  assign n78558 = ~n40312 ;
  assign n40563 = n78558 & n40432 ;
  assign n78559 = ~n40433 ;
  assign n40564 = n40311 & n78559 ;
  assign n40565 = n40563 | n40564 ;
  assign n40566 = n68220 & n40565 ;
  assign n40567 = n78531 & n40566 ;
  assign n40568 = n40562 | n40567 ;
  assign n40569 = n66560 & n40568 ;
  assign n40570 = n40095 & n40392 ;
  assign n40305 = n40104 | n40304 ;
  assign n78560 = ~n40305 ;
  assign n40571 = n40301 & n78560 ;
  assign n78561 = ~n40306 ;
  assign n40572 = n40304 & n78561 ;
  assign n40573 = n40571 | n40572 ;
  assign n40574 = n68220 & n40573 ;
  assign n40575 = n78531 & n40574 ;
  assign n40576 = n40570 | n40575 ;
  assign n40577 = n66505 & n40576 ;
  assign n40578 = n40103 & n40392 ;
  assign n40300 = n40112 | n40299 ;
  assign n78562 = ~n40300 ;
  assign n40579 = n78562 & n40428 ;
  assign n78563 = ~n40429 ;
  assign n40580 = n40299 & n78563 ;
  assign n40581 = n40579 | n40580 ;
  assign n40582 = n68220 & n40581 ;
  assign n40583 = n78531 & n40582 ;
  assign n40584 = n40578 | n40583 ;
  assign n40585 = n66379 & n40584 ;
  assign n40586 = n40111 & n40392 ;
  assign n40293 = n40120 | n40292 ;
  assign n78564 = ~n40293 ;
  assign n40587 = n40289 & n78564 ;
  assign n78565 = ~n40294 ;
  assign n40588 = n40292 & n78565 ;
  assign n40589 = n40587 | n40588 ;
  assign n40590 = n68220 & n40589 ;
  assign n40591 = n78531 & n40590 ;
  assign n40592 = n40586 | n40591 ;
  assign n40593 = n66299 & n40592 ;
  assign n40594 = n40119 & n40392 ;
  assign n40288 = n40128 | n40287 ;
  assign n78566 = ~n40288 ;
  assign n40595 = n78566 & n40424 ;
  assign n78567 = ~n40425 ;
  assign n40596 = n40287 & n78567 ;
  assign n40597 = n40595 | n40596 ;
  assign n40598 = n68220 & n40597 ;
  assign n40599 = n78531 & n40598 ;
  assign n40600 = n40594 | n40599 ;
  assign n40601 = n66244 & n40600 ;
  assign n40602 = n40127 & n40392 ;
  assign n40281 = n40136 | n40280 ;
  assign n78568 = ~n40281 ;
  assign n40603 = n40277 & n78568 ;
  assign n78569 = ~n40282 ;
  assign n40604 = n40280 & n78569 ;
  assign n40605 = n40603 | n40604 ;
  assign n40606 = n68220 & n40605 ;
  assign n40607 = n78531 & n40606 ;
  assign n40608 = n40602 | n40607 ;
  assign n40609 = n66145 & n40608 ;
  assign n40610 = n40135 & n40392 ;
  assign n40276 = n40144 | n40275 ;
  assign n78570 = ~n40276 ;
  assign n40611 = n78570 & n40420 ;
  assign n78571 = ~n40421 ;
  assign n40612 = n40275 & n78571 ;
  assign n40613 = n40611 | n40612 ;
  assign n40614 = n68220 & n40613 ;
  assign n40615 = n78531 & n40614 ;
  assign n40616 = n40610 | n40615 ;
  assign n40617 = n66081 & n40616 ;
  assign n40618 = n40143 & n40392 ;
  assign n40269 = n40152 | n40268 ;
  assign n78572 = ~n40269 ;
  assign n40619 = n40265 & n78572 ;
  assign n78573 = ~n40270 ;
  assign n40620 = n40268 & n78573 ;
  assign n40621 = n40619 | n40620 ;
  assign n40622 = n68220 & n40621 ;
  assign n40623 = n78531 & n40622 ;
  assign n40624 = n40618 | n40623 ;
  assign n40625 = n66043 & n40624 ;
  assign n40626 = n40151 & n40392 ;
  assign n40264 = n40160 | n40263 ;
  assign n78574 = ~n40264 ;
  assign n40627 = n78574 & n40416 ;
  assign n78575 = ~n40417 ;
  assign n40628 = n40263 & n78575 ;
  assign n40629 = n40627 | n40628 ;
  assign n40630 = n68220 & n40629 ;
  assign n40631 = n78531 & n40630 ;
  assign n40632 = n40626 | n40631 ;
  assign n40633 = n65960 & n40632 ;
  assign n40634 = n40159 & n40392 ;
  assign n40257 = n40168 | n40256 ;
  assign n78576 = ~n40257 ;
  assign n40635 = n40253 & n78576 ;
  assign n78577 = ~n40258 ;
  assign n40636 = n40256 & n78577 ;
  assign n40637 = n40635 | n40636 ;
  assign n40638 = n68220 & n40637 ;
  assign n40639 = n78531 & n40638 ;
  assign n40640 = n40634 | n40639 ;
  assign n40641 = n65909 & n40640 ;
  assign n40642 = n40167 & n40392 ;
  assign n40252 = n40176 | n40251 ;
  assign n78578 = ~n40252 ;
  assign n40643 = n78578 & n40412 ;
  assign n78579 = ~n40413 ;
  assign n40644 = n40251 & n78579 ;
  assign n40645 = n40643 | n40644 ;
  assign n40646 = n68220 & n40645 ;
  assign n40647 = n78531 & n40646 ;
  assign n40648 = n40642 | n40647 ;
  assign n40649 = n65877 & n40648 ;
  assign n40650 = n40175 & n40392 ;
  assign n40245 = n40185 | n40244 ;
  assign n78580 = ~n40245 ;
  assign n40651 = n40241 & n78580 ;
  assign n78581 = ~n40246 ;
  assign n40652 = n40244 & n78581 ;
  assign n40653 = n40651 | n40652 ;
  assign n40654 = n68220 & n40653 ;
  assign n40655 = n78531 & n40654 ;
  assign n40656 = n40650 | n40655 ;
  assign n40657 = n65820 & n40656 ;
  assign n40658 = n40184 & n40392 ;
  assign n40240 = n40193 | n40239 ;
  assign n78582 = ~n40240 ;
  assign n40659 = n78582 & n40408 ;
  assign n78583 = ~n40409 ;
  assign n40660 = n40239 & n78583 ;
  assign n40661 = n40659 | n40660 ;
  assign n40662 = n68220 & n40661 ;
  assign n40663 = n78531 & n40662 ;
  assign n40664 = n40658 | n40663 ;
  assign n40665 = n65791 & n40664 ;
  assign n40666 = n40192 & n40392 ;
  assign n40667 = n40201 | n40233 ;
  assign n78584 = ~n40667 ;
  assign n40668 = n40230 & n78584 ;
  assign n78585 = ~n40234 ;
  assign n40669 = n40233 & n78585 ;
  assign n40670 = n40668 | n40669 ;
  assign n40671 = n68220 & n40670 ;
  assign n40672 = n78531 & n40671 ;
  assign n40673 = n40666 | n40672 ;
  assign n40674 = n65772 & n40673 ;
  assign n40675 = n40200 & n40392 ;
  assign n40676 = n40209 | n40229 ;
  assign n78586 = ~n40676 ;
  assign n40677 = n40225 & n78586 ;
  assign n78587 = ~n40405 ;
  assign n40678 = n40229 & n78587 ;
  assign n40679 = n40677 | n40678 ;
  assign n40680 = n68220 & n40679 ;
  assign n40681 = n78531 & n40680 ;
  assign n40682 = n40675 | n40681 ;
  assign n40683 = n65746 & n40682 ;
  assign n40684 = n40208 & n40392 ;
  assign n40403 = n40220 | n40223 ;
  assign n78588 = ~n40403 ;
  assign n40685 = n40401 & n78588 ;
  assign n78589 = ~n40224 ;
  assign n40686 = n40223 & n78589 ;
  assign n40687 = n40685 | n40686 ;
  assign n40688 = n68220 & n40687 ;
  assign n40689 = n78531 & n40688 ;
  assign n40690 = n40684 | n40689 ;
  assign n40691 = n65721 & n40690 ;
  assign n40394 = n40211 & n40392 ;
  assign n40218 = n7868 & n40216 ;
  assign n40693 = n40218 & n78528 ;
  assign n40694 = n8032 | n40693 ;
  assign n78590 = ~n40694 ;
  assign n40695 = n40401 & n78590 ;
  assign n40696 = n78531 & n40695 ;
  assign n40697 = n40394 | n40696 ;
  assign n40698 = n65686 & n40697 ;
  assign n40692 = n8357 & n78531 ;
  assign n40699 = n8351 & n78531 ;
  assign n78591 = ~n40699 ;
  assign n40700 = x33 & n78591 ;
  assign n40701 = n40692 | n40700 ;
  assign n40702 = n65670 & n40701 ;
  assign n40465 = n78525 & n40464 ;
  assign n40704 = n40388 | n40465 ;
  assign n40705 = n78526 & n40704 ;
  assign n78592 = ~n40705 ;
  assign n40706 = n8351 & n78592 ;
  assign n78593 = ~n40706 ;
  assign n40707 = x33 & n78593 ;
  assign n40708 = n40692 | n40707 ;
  assign n40710 = x65 & n40708 ;
  assign n40709 = x65 | n40692 ;
  assign n40711 = n40700 | n40709 ;
  assign n78594 = ~n40710 ;
  assign n40712 = n78594 & n40711 ;
  assign n40713 = n8368 | n40712 ;
  assign n78595 = ~n40702 ;
  assign n40714 = n78595 & n40713 ;
  assign n78596 = ~n40696 ;
  assign n40715 = x66 & n78596 ;
  assign n78597 = ~n40394 ;
  assign n40716 = n78597 & n40715 ;
  assign n40717 = n40698 | n40716 ;
  assign n40718 = n40714 | n40717 ;
  assign n78598 = ~n40698 ;
  assign n40719 = n78598 & n40718 ;
  assign n78599 = ~n40689 ;
  assign n40720 = x67 & n78599 ;
  assign n78600 = ~n40684 ;
  assign n40721 = n78600 & n40720 ;
  assign n40722 = n40719 | n40721 ;
  assign n78601 = ~n40691 ;
  assign n40723 = n78601 & n40722 ;
  assign n78602 = ~n40681 ;
  assign n40724 = x68 & n78602 ;
  assign n78603 = ~n40675 ;
  assign n40725 = n78603 & n40724 ;
  assign n40726 = n40683 | n40725 ;
  assign n40727 = n40723 | n40726 ;
  assign n78604 = ~n40683 ;
  assign n40728 = n78604 & n40727 ;
  assign n78605 = ~n40672 ;
  assign n40729 = x69 & n78605 ;
  assign n78606 = ~n40666 ;
  assign n40730 = n78606 & n40729 ;
  assign n40731 = n40674 | n40730 ;
  assign n40732 = n40728 | n40731 ;
  assign n78607 = ~n40674 ;
  assign n40733 = n78607 & n40732 ;
  assign n78608 = ~n40663 ;
  assign n40734 = x70 & n78608 ;
  assign n78609 = ~n40658 ;
  assign n40735 = n78609 & n40734 ;
  assign n40736 = n40665 | n40735 ;
  assign n40737 = n40733 | n40736 ;
  assign n78610 = ~n40665 ;
  assign n40738 = n78610 & n40737 ;
  assign n78611 = ~n40655 ;
  assign n40739 = x71 & n78611 ;
  assign n78612 = ~n40650 ;
  assign n40740 = n78612 & n40739 ;
  assign n40741 = n40657 | n40740 ;
  assign n40743 = n40738 | n40741 ;
  assign n78613 = ~n40657 ;
  assign n40744 = n78613 & n40743 ;
  assign n78614 = ~n40647 ;
  assign n40745 = x72 & n78614 ;
  assign n78615 = ~n40642 ;
  assign n40746 = n78615 & n40745 ;
  assign n40747 = n40649 | n40746 ;
  assign n40748 = n40744 | n40747 ;
  assign n78616 = ~n40649 ;
  assign n40749 = n78616 & n40748 ;
  assign n78617 = ~n40639 ;
  assign n40750 = x73 & n78617 ;
  assign n78618 = ~n40634 ;
  assign n40751 = n78618 & n40750 ;
  assign n40752 = n40641 | n40751 ;
  assign n40754 = n40749 | n40752 ;
  assign n78619 = ~n40641 ;
  assign n40755 = n78619 & n40754 ;
  assign n78620 = ~n40631 ;
  assign n40756 = x74 & n78620 ;
  assign n78621 = ~n40626 ;
  assign n40757 = n78621 & n40756 ;
  assign n40758 = n40633 | n40757 ;
  assign n40759 = n40755 | n40758 ;
  assign n78622 = ~n40633 ;
  assign n40760 = n78622 & n40759 ;
  assign n78623 = ~n40623 ;
  assign n40761 = x75 & n78623 ;
  assign n78624 = ~n40618 ;
  assign n40762 = n78624 & n40761 ;
  assign n40763 = n40625 | n40762 ;
  assign n40765 = n40760 | n40763 ;
  assign n78625 = ~n40625 ;
  assign n40766 = n78625 & n40765 ;
  assign n78626 = ~n40615 ;
  assign n40767 = x76 & n78626 ;
  assign n78627 = ~n40610 ;
  assign n40768 = n78627 & n40767 ;
  assign n40769 = n40617 | n40768 ;
  assign n40770 = n40766 | n40769 ;
  assign n78628 = ~n40617 ;
  assign n40771 = n78628 & n40770 ;
  assign n78629 = ~n40607 ;
  assign n40772 = x77 & n78629 ;
  assign n78630 = ~n40602 ;
  assign n40773 = n78630 & n40772 ;
  assign n40774 = n40609 | n40773 ;
  assign n40776 = n40771 | n40774 ;
  assign n78631 = ~n40609 ;
  assign n40777 = n78631 & n40776 ;
  assign n78632 = ~n40599 ;
  assign n40778 = x78 & n78632 ;
  assign n78633 = ~n40594 ;
  assign n40779 = n78633 & n40778 ;
  assign n40780 = n40601 | n40779 ;
  assign n40781 = n40777 | n40780 ;
  assign n78634 = ~n40601 ;
  assign n40782 = n78634 & n40781 ;
  assign n78635 = ~n40591 ;
  assign n40783 = x79 & n78635 ;
  assign n78636 = ~n40586 ;
  assign n40784 = n78636 & n40783 ;
  assign n40785 = n40593 | n40784 ;
  assign n40787 = n40782 | n40785 ;
  assign n78637 = ~n40593 ;
  assign n40788 = n78637 & n40787 ;
  assign n78638 = ~n40583 ;
  assign n40789 = x80 & n78638 ;
  assign n78639 = ~n40578 ;
  assign n40790 = n78639 & n40789 ;
  assign n40791 = n40585 | n40790 ;
  assign n40792 = n40788 | n40791 ;
  assign n78640 = ~n40585 ;
  assign n40793 = n78640 & n40792 ;
  assign n78641 = ~n40575 ;
  assign n40794 = x81 & n78641 ;
  assign n78642 = ~n40570 ;
  assign n40795 = n78642 & n40794 ;
  assign n40796 = n40577 | n40795 ;
  assign n40798 = n40793 | n40796 ;
  assign n78643 = ~n40577 ;
  assign n40799 = n78643 & n40798 ;
  assign n78644 = ~n40567 ;
  assign n40800 = x82 & n78644 ;
  assign n78645 = ~n40562 ;
  assign n40801 = n78645 & n40800 ;
  assign n40802 = n40569 | n40801 ;
  assign n40803 = n40799 | n40802 ;
  assign n78646 = ~n40569 ;
  assign n40804 = n78646 & n40803 ;
  assign n78647 = ~n40559 ;
  assign n40805 = x83 & n78647 ;
  assign n78648 = ~n40554 ;
  assign n40806 = n78648 & n40805 ;
  assign n40807 = n40561 | n40806 ;
  assign n40809 = n40804 | n40807 ;
  assign n78649 = ~n40561 ;
  assign n40810 = n78649 & n40809 ;
  assign n78650 = ~n40551 ;
  assign n40811 = x84 & n78650 ;
  assign n78651 = ~n40546 ;
  assign n40812 = n78651 & n40811 ;
  assign n40813 = n40553 | n40812 ;
  assign n40814 = n40810 | n40813 ;
  assign n78652 = ~n40553 ;
  assign n40815 = n78652 & n40814 ;
  assign n78653 = ~n40543 ;
  assign n40816 = x85 & n78653 ;
  assign n78654 = ~n40538 ;
  assign n40817 = n78654 & n40816 ;
  assign n40818 = n40545 | n40817 ;
  assign n40820 = n40815 | n40818 ;
  assign n78655 = ~n40545 ;
  assign n40821 = n78655 & n40820 ;
  assign n78656 = ~n40535 ;
  assign n40822 = x86 & n78656 ;
  assign n78657 = ~n40530 ;
  assign n40823 = n78657 & n40822 ;
  assign n40824 = n40537 | n40823 ;
  assign n40825 = n40821 | n40824 ;
  assign n78658 = ~n40537 ;
  assign n40826 = n78658 & n40825 ;
  assign n78659 = ~n40527 ;
  assign n40827 = x87 & n78659 ;
  assign n78660 = ~n40522 ;
  assign n40828 = n78660 & n40827 ;
  assign n40829 = n40529 | n40828 ;
  assign n40831 = n40826 | n40829 ;
  assign n78661 = ~n40529 ;
  assign n40832 = n78661 & n40831 ;
  assign n78662 = ~n40519 ;
  assign n40833 = x88 & n78662 ;
  assign n78663 = ~n40514 ;
  assign n40834 = n78663 & n40833 ;
  assign n40835 = n40521 | n40834 ;
  assign n40836 = n40832 | n40835 ;
  assign n78664 = ~n40521 ;
  assign n40837 = n78664 & n40836 ;
  assign n78665 = ~n40511 ;
  assign n40838 = x89 & n78665 ;
  assign n78666 = ~n40506 ;
  assign n40839 = n78666 & n40838 ;
  assign n40840 = n40513 | n40839 ;
  assign n40842 = n40837 | n40840 ;
  assign n78667 = ~n40513 ;
  assign n40843 = n78667 & n40842 ;
  assign n78668 = ~n40503 ;
  assign n40844 = x90 & n78668 ;
  assign n78669 = ~n40498 ;
  assign n40845 = n78669 & n40844 ;
  assign n40846 = n40505 | n40845 ;
  assign n40847 = n40843 | n40846 ;
  assign n78670 = ~n40505 ;
  assign n40848 = n78670 & n40847 ;
  assign n78671 = ~n40495 ;
  assign n40849 = x91 & n78671 ;
  assign n78672 = ~n40490 ;
  assign n40850 = n78672 & n40849 ;
  assign n40851 = n40497 | n40850 ;
  assign n40853 = n40848 | n40851 ;
  assign n78673 = ~n40497 ;
  assign n40854 = n78673 & n40853 ;
  assign n78674 = ~n40487 ;
  assign n40855 = x92 & n78674 ;
  assign n78675 = ~n40482 ;
  assign n40856 = n78675 & n40855 ;
  assign n40857 = n40489 | n40856 ;
  assign n40858 = n40854 | n40857 ;
  assign n78676 = ~n40489 ;
  assign n40859 = n78676 & n40858 ;
  assign n78677 = ~n40479 ;
  assign n40860 = x93 & n78677 ;
  assign n78678 = ~n40474 ;
  assign n40861 = n78678 & n40860 ;
  assign n40862 = n40481 | n40861 ;
  assign n40864 = n40859 | n40862 ;
  assign n78679 = ~n40481 ;
  assign n40865 = n78679 & n40864 ;
  assign n78680 = ~n40462 ;
  assign n40866 = x94 & n78680 ;
  assign n78681 = ~n40395 ;
  assign n40867 = n78681 & n40866 ;
  assign n40868 = n40473 | n40867 ;
  assign n40869 = n40865 | n40868 ;
  assign n78682 = ~n40473 ;
  assign n40870 = n78682 & n40869 ;
  assign n78683 = ~n40392 ;
  assign n40871 = n78683 & n40469 ;
  assign n40872 = n39990 & n40392 ;
  assign n78684 = ~n40872 ;
  assign n40873 = x95 & n78684 ;
  assign n78685 = ~n40871 ;
  assign n40874 = n78685 & n40873 ;
  assign n40875 = n40472 | n40874 ;
  assign n40877 = n40870 | n40875 ;
  assign n78686 = ~n40472 ;
  assign n40878 = n78686 & n40877 ;
  assign n40879 = n303 | n40878 ;
  assign n40880 = n40463 & n40879 ;
  assign n40882 = n65670 & n40708 ;
  assign n40703 = x65 & n40701 ;
  assign n78687 = ~n40703 ;
  assign n40881 = n78687 & n40711 ;
  assign n40883 = n8368 | n40881 ;
  assign n78688 = ~n40882 ;
  assign n40884 = n78688 & n40883 ;
  assign n40885 = n40717 | n40884 ;
  assign n40886 = n78598 & n40885 ;
  assign n40887 = n40691 | n40721 ;
  assign n40889 = n40886 | n40887 ;
  assign n40890 = n78601 & n40889 ;
  assign n40892 = n40726 | n40890 ;
  assign n40893 = n78604 & n40892 ;
  assign n40895 = n40731 | n40893 ;
  assign n40896 = n78607 & n40895 ;
  assign n40897 = n40736 | n40896 ;
  assign n40899 = n78610 & n40897 ;
  assign n40900 = n40741 | n40899 ;
  assign n40901 = n78613 & n40900 ;
  assign n40902 = n40747 | n40901 ;
  assign n40904 = n78616 & n40902 ;
  assign n40905 = n40752 | n40904 ;
  assign n40906 = n78619 & n40905 ;
  assign n40907 = n40758 | n40906 ;
  assign n40909 = n78622 & n40907 ;
  assign n40910 = n40763 | n40909 ;
  assign n40911 = n78625 & n40910 ;
  assign n40912 = n40769 | n40911 ;
  assign n40914 = n78628 & n40912 ;
  assign n40915 = n40774 | n40914 ;
  assign n40916 = n78631 & n40915 ;
  assign n40917 = n40780 | n40916 ;
  assign n40919 = n78634 & n40917 ;
  assign n40920 = n40785 | n40919 ;
  assign n40921 = n78637 & n40920 ;
  assign n40922 = n40791 | n40921 ;
  assign n40924 = n78640 & n40922 ;
  assign n40925 = n40796 | n40924 ;
  assign n40926 = n78643 & n40925 ;
  assign n40927 = n40802 | n40926 ;
  assign n40929 = n78646 & n40927 ;
  assign n40930 = n40807 | n40929 ;
  assign n40931 = n78649 & n40930 ;
  assign n40932 = n40813 | n40931 ;
  assign n40934 = n78652 & n40932 ;
  assign n40935 = n40818 | n40934 ;
  assign n40936 = n78655 & n40935 ;
  assign n40937 = n40824 | n40936 ;
  assign n40939 = n78658 & n40937 ;
  assign n40940 = n40829 | n40939 ;
  assign n40941 = n78661 & n40940 ;
  assign n40942 = n40835 | n40941 ;
  assign n40944 = n78664 & n40942 ;
  assign n40945 = n40840 | n40944 ;
  assign n40946 = n78667 & n40945 ;
  assign n40947 = n40846 | n40946 ;
  assign n40949 = n78670 & n40947 ;
  assign n40950 = n40851 | n40949 ;
  assign n40951 = n78673 & n40950 ;
  assign n40952 = n40857 | n40951 ;
  assign n40954 = n78676 & n40952 ;
  assign n40955 = n40862 | n40954 ;
  assign n40956 = n78679 & n40955 ;
  assign n78689 = ~n40956 ;
  assign n40957 = n40868 & n78689 ;
  assign n40959 = n40481 | n40868 ;
  assign n78690 = ~n40959 ;
  assign n40960 = n40864 & n78690 ;
  assign n40961 = n40957 | n40960 ;
  assign n40962 = n65696 & n40961 ;
  assign n78691 = ~n40878 ;
  assign n40963 = n78691 & n40962 ;
  assign n40964 = n40880 | n40963 ;
  assign n40965 = n68214 & n40964 ;
  assign n78692 = ~n40963 ;
  assign n41365 = x95 & n78692 ;
  assign n78693 = ~n40880 ;
  assign n41366 = n78693 & n41365 ;
  assign n41367 = n40965 | n41366 ;
  assign n40966 = n40480 & n40879 ;
  assign n78694 = ~n40859 ;
  assign n40863 = n78694 & n40862 ;
  assign n40967 = n40489 | n40862 ;
  assign n78695 = ~n40967 ;
  assign n40968 = n40952 & n78695 ;
  assign n40969 = n40863 | n40968 ;
  assign n40970 = n65696 & n40969 ;
  assign n40971 = n78691 & n40970 ;
  assign n40972 = n40966 | n40971 ;
  assign n40973 = n68058 & n40972 ;
  assign n40974 = n40488 & n40879 ;
  assign n78696 = ~n40951 ;
  assign n40953 = n40857 & n78696 ;
  assign n40975 = n40497 | n40857 ;
  assign n78697 = ~n40975 ;
  assign n40976 = n40853 & n78697 ;
  assign n40977 = n40953 | n40976 ;
  assign n40978 = n65696 & n40977 ;
  assign n40979 = n78691 & n40978 ;
  assign n40980 = n40974 | n40979 ;
  assign n40981 = n67986 & n40980 ;
  assign n78698 = ~n40979 ;
  assign n41355 = x93 & n78698 ;
  assign n78699 = ~n40974 ;
  assign n41356 = n78699 & n41355 ;
  assign n41357 = n40981 | n41356 ;
  assign n40982 = n40496 & n40879 ;
  assign n78700 = ~n40848 ;
  assign n40852 = n78700 & n40851 ;
  assign n40983 = n40505 | n40851 ;
  assign n78701 = ~n40983 ;
  assign n40984 = n40947 & n78701 ;
  assign n40985 = n40852 | n40984 ;
  assign n40986 = n65696 & n40985 ;
  assign n40987 = n78691 & n40986 ;
  assign n40988 = n40982 | n40987 ;
  assign n40989 = n67763 & n40988 ;
  assign n40990 = n40504 & n40879 ;
  assign n78702 = ~n40946 ;
  assign n40948 = n40846 & n78702 ;
  assign n40991 = n40513 | n40846 ;
  assign n78703 = ~n40991 ;
  assign n40992 = n40842 & n78703 ;
  assign n40993 = n40948 | n40992 ;
  assign n40994 = n65696 & n40993 ;
  assign n40995 = n78691 & n40994 ;
  assign n40996 = n40990 | n40995 ;
  assign n40997 = n67622 & n40996 ;
  assign n78704 = ~n40995 ;
  assign n41345 = x91 & n78704 ;
  assign n78705 = ~n40990 ;
  assign n41346 = n78705 & n41345 ;
  assign n41347 = n40997 | n41346 ;
  assign n40998 = n40512 & n40879 ;
  assign n78706 = ~n40837 ;
  assign n40841 = n78706 & n40840 ;
  assign n40999 = n40521 | n40840 ;
  assign n78707 = ~n40999 ;
  assign n41000 = n40942 & n78707 ;
  assign n41001 = n40841 | n41000 ;
  assign n41002 = n65696 & n41001 ;
  assign n41003 = n78691 & n41002 ;
  assign n41004 = n40998 | n41003 ;
  assign n41005 = n67531 & n41004 ;
  assign n41006 = n40520 & n40879 ;
  assign n78708 = ~n40941 ;
  assign n40943 = n40835 & n78708 ;
  assign n41007 = n40529 | n40835 ;
  assign n78709 = ~n41007 ;
  assign n41008 = n40831 & n78709 ;
  assign n41009 = n40943 | n41008 ;
  assign n41010 = n65696 & n41009 ;
  assign n41011 = n78691 & n41010 ;
  assign n41012 = n41006 | n41011 ;
  assign n41013 = n67348 & n41012 ;
  assign n78710 = ~n41011 ;
  assign n41335 = x89 & n78710 ;
  assign n78711 = ~n41006 ;
  assign n41336 = n78711 & n41335 ;
  assign n41337 = n41013 | n41336 ;
  assign n41014 = n40528 & n40879 ;
  assign n78712 = ~n40826 ;
  assign n40830 = n78712 & n40829 ;
  assign n41015 = n40537 | n40829 ;
  assign n78713 = ~n41015 ;
  assign n41016 = n40937 & n78713 ;
  assign n41017 = n40830 | n41016 ;
  assign n41018 = n65696 & n41017 ;
  assign n41019 = n78691 & n41018 ;
  assign n41020 = n41014 | n41019 ;
  assign n41021 = n67222 & n41020 ;
  assign n41022 = n40536 & n40879 ;
  assign n78714 = ~n40936 ;
  assign n40938 = n40824 & n78714 ;
  assign n41023 = n40545 | n40824 ;
  assign n78715 = ~n41023 ;
  assign n41024 = n40820 & n78715 ;
  assign n41025 = n40938 | n41024 ;
  assign n41026 = n65696 & n41025 ;
  assign n41027 = n78691 & n41026 ;
  assign n41028 = n41022 | n41027 ;
  assign n41029 = n67164 & n41028 ;
  assign n78716 = ~n41027 ;
  assign n41325 = x87 & n78716 ;
  assign n78717 = ~n41022 ;
  assign n41326 = n78717 & n41325 ;
  assign n41327 = n41029 | n41326 ;
  assign n41030 = n40544 & n40879 ;
  assign n78718 = ~n40815 ;
  assign n40819 = n78718 & n40818 ;
  assign n41031 = n40553 | n40818 ;
  assign n78719 = ~n41031 ;
  assign n41032 = n40932 & n78719 ;
  assign n41033 = n40819 | n41032 ;
  assign n41034 = n65696 & n41033 ;
  assign n41035 = n78691 & n41034 ;
  assign n41036 = n41030 | n41035 ;
  assign n41037 = n66979 & n41036 ;
  assign n41038 = n40552 & n40879 ;
  assign n78720 = ~n40931 ;
  assign n40933 = n40813 & n78720 ;
  assign n41039 = n40561 | n40813 ;
  assign n78721 = ~n41039 ;
  assign n41040 = n40809 & n78721 ;
  assign n41041 = n40933 | n41040 ;
  assign n41042 = n65696 & n41041 ;
  assign n41043 = n78691 & n41042 ;
  assign n41044 = n41038 | n41043 ;
  assign n41045 = n66868 & n41044 ;
  assign n78722 = ~n41043 ;
  assign n41314 = x85 & n78722 ;
  assign n78723 = ~n41038 ;
  assign n41315 = n78723 & n41314 ;
  assign n41316 = n41045 | n41315 ;
  assign n41046 = n40560 & n40879 ;
  assign n78724 = ~n40804 ;
  assign n40808 = n78724 & n40807 ;
  assign n41047 = n40569 | n40807 ;
  assign n78725 = ~n41047 ;
  assign n41048 = n40927 & n78725 ;
  assign n41049 = n40808 | n41048 ;
  assign n41050 = n65696 & n41049 ;
  assign n41051 = n78691 & n41050 ;
  assign n41052 = n41046 | n41051 ;
  assign n41053 = n66797 & n41052 ;
  assign n41054 = n40568 & n40879 ;
  assign n78726 = ~n40926 ;
  assign n40928 = n40802 & n78726 ;
  assign n41055 = n40577 | n40802 ;
  assign n78727 = ~n41055 ;
  assign n41056 = n40798 & n78727 ;
  assign n41057 = n40928 | n41056 ;
  assign n41058 = n65696 & n41057 ;
  assign n41059 = n78691 & n41058 ;
  assign n41060 = n41054 | n41059 ;
  assign n41061 = n66654 & n41060 ;
  assign n78728 = ~n41059 ;
  assign n41304 = x83 & n78728 ;
  assign n78729 = ~n41054 ;
  assign n41305 = n78729 & n41304 ;
  assign n41306 = n41061 | n41305 ;
  assign n41062 = n40576 & n40879 ;
  assign n78730 = ~n40793 ;
  assign n40797 = n78730 & n40796 ;
  assign n41063 = n40585 | n40796 ;
  assign n78731 = ~n41063 ;
  assign n41064 = n40922 & n78731 ;
  assign n41065 = n40797 | n41064 ;
  assign n41066 = n65696 & n41065 ;
  assign n41067 = n78691 & n41066 ;
  assign n41068 = n41062 | n41067 ;
  assign n41069 = n66560 & n41068 ;
  assign n41070 = n40584 & n40879 ;
  assign n78732 = ~n40921 ;
  assign n40923 = n40791 & n78732 ;
  assign n41071 = n40593 | n40791 ;
  assign n78733 = ~n41071 ;
  assign n41072 = n40787 & n78733 ;
  assign n41073 = n40923 | n41072 ;
  assign n41074 = n65696 & n41073 ;
  assign n41075 = n78691 & n41074 ;
  assign n41076 = n41070 | n41075 ;
  assign n41077 = n66505 & n41076 ;
  assign n78734 = ~n41075 ;
  assign n41294 = x81 & n78734 ;
  assign n78735 = ~n41070 ;
  assign n41295 = n78735 & n41294 ;
  assign n41296 = n41077 | n41295 ;
  assign n41078 = n40592 & n40879 ;
  assign n78736 = ~n40782 ;
  assign n40786 = n78736 & n40785 ;
  assign n41079 = n40601 | n40785 ;
  assign n78737 = ~n41079 ;
  assign n41080 = n40917 & n78737 ;
  assign n41081 = n40786 | n41080 ;
  assign n41082 = n65696 & n41081 ;
  assign n41083 = n78691 & n41082 ;
  assign n41084 = n41078 | n41083 ;
  assign n41085 = n66379 & n41084 ;
  assign n41086 = n40600 & n40879 ;
  assign n78738 = ~n40916 ;
  assign n40918 = n40780 & n78738 ;
  assign n41087 = n40609 | n40780 ;
  assign n78739 = ~n41087 ;
  assign n41088 = n40776 & n78739 ;
  assign n41089 = n40918 | n41088 ;
  assign n41090 = n65696 & n41089 ;
  assign n41091 = n78691 & n41090 ;
  assign n41092 = n41086 | n41091 ;
  assign n41093 = n66299 & n41092 ;
  assign n78740 = ~n41091 ;
  assign n41284 = x79 & n78740 ;
  assign n78741 = ~n41086 ;
  assign n41285 = n78741 & n41284 ;
  assign n41286 = n41093 | n41285 ;
  assign n41094 = n40608 & n40879 ;
  assign n78742 = ~n40771 ;
  assign n40775 = n78742 & n40774 ;
  assign n41095 = n40617 | n40774 ;
  assign n78743 = ~n41095 ;
  assign n41096 = n40912 & n78743 ;
  assign n41097 = n40775 | n41096 ;
  assign n41098 = n65696 & n41097 ;
  assign n41099 = n78691 & n41098 ;
  assign n41100 = n41094 | n41099 ;
  assign n41101 = n66244 & n41100 ;
  assign n41102 = n40616 & n40879 ;
  assign n78744 = ~n40911 ;
  assign n40913 = n40769 & n78744 ;
  assign n41103 = n40625 | n40769 ;
  assign n78745 = ~n41103 ;
  assign n41104 = n40765 & n78745 ;
  assign n41105 = n40913 | n41104 ;
  assign n41106 = n65696 & n41105 ;
  assign n41107 = n78691 & n41106 ;
  assign n41108 = n41102 | n41107 ;
  assign n41109 = n66145 & n41108 ;
  assign n78746 = ~n41107 ;
  assign n41273 = x77 & n78746 ;
  assign n78747 = ~n41102 ;
  assign n41274 = n78747 & n41273 ;
  assign n41275 = n41109 | n41274 ;
  assign n41110 = n40624 & n40879 ;
  assign n78748 = ~n40760 ;
  assign n40764 = n78748 & n40763 ;
  assign n41111 = n40633 | n40763 ;
  assign n78749 = ~n41111 ;
  assign n41112 = n40907 & n78749 ;
  assign n41113 = n40764 | n41112 ;
  assign n41114 = n65696 & n41113 ;
  assign n41115 = n78691 & n41114 ;
  assign n41116 = n41110 | n41115 ;
  assign n41117 = n66081 & n41116 ;
  assign n41118 = n40632 & n40879 ;
  assign n78750 = ~n40906 ;
  assign n40908 = n40758 & n78750 ;
  assign n41119 = n40641 | n40758 ;
  assign n78751 = ~n41119 ;
  assign n41120 = n40754 & n78751 ;
  assign n41121 = n40908 | n41120 ;
  assign n41122 = n65696 & n41121 ;
  assign n41123 = n78691 & n41122 ;
  assign n41124 = n41118 | n41123 ;
  assign n41125 = n66043 & n41124 ;
  assign n78752 = ~n41123 ;
  assign n41261 = x75 & n78752 ;
  assign n78753 = ~n41118 ;
  assign n41262 = n78753 & n41261 ;
  assign n41263 = n41125 | n41262 ;
  assign n41126 = n40640 & n40879 ;
  assign n78754 = ~n40749 ;
  assign n40753 = n78754 & n40752 ;
  assign n41127 = n40649 | n40752 ;
  assign n78755 = ~n41127 ;
  assign n41128 = n40902 & n78755 ;
  assign n41129 = n40753 | n41128 ;
  assign n41130 = n65696 & n41129 ;
  assign n41131 = n78691 & n41130 ;
  assign n41132 = n41126 | n41131 ;
  assign n41133 = n65960 & n41132 ;
  assign n41134 = n40648 & n40879 ;
  assign n78756 = ~n40901 ;
  assign n40903 = n40747 & n78756 ;
  assign n41135 = n40657 | n40747 ;
  assign n78757 = ~n41135 ;
  assign n41136 = n40743 & n78757 ;
  assign n41137 = n40903 | n41136 ;
  assign n41138 = n65696 & n41137 ;
  assign n41139 = n78691 & n41138 ;
  assign n41140 = n41134 | n41139 ;
  assign n41141 = n65909 & n41140 ;
  assign n78758 = ~n41139 ;
  assign n41251 = x73 & n78758 ;
  assign n78759 = ~n41134 ;
  assign n41252 = n78759 & n41251 ;
  assign n41253 = n41141 | n41252 ;
  assign n41142 = n40656 & n40879 ;
  assign n78760 = ~n40738 ;
  assign n40742 = n78760 & n40741 ;
  assign n41143 = n40665 | n40741 ;
  assign n78761 = ~n41143 ;
  assign n41144 = n40897 & n78761 ;
  assign n41145 = n40742 | n41144 ;
  assign n41146 = n65696 & n41145 ;
  assign n41147 = n78691 & n41146 ;
  assign n41148 = n41142 | n41147 ;
  assign n41149 = n65877 & n41148 ;
  assign n41150 = n40664 & n40879 ;
  assign n78762 = ~n40896 ;
  assign n40898 = n40736 & n78762 ;
  assign n41151 = n40674 | n40736 ;
  assign n78763 = ~n41151 ;
  assign n41152 = n40732 & n78763 ;
  assign n41153 = n40898 | n41152 ;
  assign n41154 = n65696 & n41153 ;
  assign n41155 = n78691 & n41154 ;
  assign n41156 = n41150 | n41155 ;
  assign n41157 = n65820 & n41156 ;
  assign n78764 = ~n41155 ;
  assign n41241 = x71 & n78764 ;
  assign n78765 = ~n41150 ;
  assign n41242 = n78765 & n41241 ;
  assign n41243 = n41157 | n41242 ;
  assign n41158 = n40673 & n40879 ;
  assign n78766 = ~n40728 ;
  assign n40894 = n78766 & n40731 ;
  assign n41159 = n40683 | n40731 ;
  assign n78767 = ~n41159 ;
  assign n41160 = n40727 & n78767 ;
  assign n41161 = n40894 | n41160 ;
  assign n41162 = n65696 & n41161 ;
  assign n41163 = n78691 & n41162 ;
  assign n41164 = n41158 | n41163 ;
  assign n41165 = n65791 & n41164 ;
  assign n41166 = n40682 & n40879 ;
  assign n78768 = ~n40890 ;
  assign n40891 = n40726 & n78768 ;
  assign n41167 = n40719 | n40887 ;
  assign n41168 = n40691 | n40726 ;
  assign n78769 = ~n41168 ;
  assign n41169 = n41167 & n78769 ;
  assign n41170 = n40891 | n41169 ;
  assign n41171 = n65696 & n41170 ;
  assign n41172 = n78691 & n41171 ;
  assign n41173 = n41166 | n41172 ;
  assign n41174 = n65772 & n41173 ;
  assign n78770 = ~n41172 ;
  assign n41231 = x69 & n78770 ;
  assign n78771 = ~n41166 ;
  assign n41232 = n78771 & n41231 ;
  assign n41233 = n41174 | n41232 ;
  assign n41175 = n40690 & n40879 ;
  assign n78772 = ~n40719 ;
  assign n40888 = n78772 & n40887 ;
  assign n41176 = n40698 | n40887 ;
  assign n78773 = ~n41176 ;
  assign n41177 = n40718 & n78773 ;
  assign n41178 = n40888 | n41177 ;
  assign n41179 = n65696 & n41178 ;
  assign n41180 = n78691 & n41179 ;
  assign n41181 = n41175 | n41180 ;
  assign n41182 = n65746 & n41181 ;
  assign n41183 = n40697 & n40879 ;
  assign n41184 = n40717 | n40882 ;
  assign n78774 = ~n41184 ;
  assign n41185 = n40883 & n78774 ;
  assign n78775 = ~n40884 ;
  assign n41186 = n40717 & n78775 ;
  assign n41187 = n41185 | n41186 ;
  assign n41188 = n65696 & n41187 ;
  assign n41189 = n78691 & n41188 ;
  assign n41190 = n41183 | n41189 ;
  assign n41192 = n65721 & n41190 ;
  assign n78776 = ~n41189 ;
  assign n41191 = x67 & n78776 ;
  assign n78777 = ~n41183 ;
  assign n41222 = n78777 & n41191 ;
  assign n41223 = n41192 | n41222 ;
  assign n41193 = n40701 & n40879 ;
  assign n41194 = n8368 & n40711 ;
  assign n41195 = n78594 & n41194 ;
  assign n41196 = n303 | n41195 ;
  assign n78778 = ~n41196 ;
  assign n41197 = n40883 & n78778 ;
  assign n41198 = n78691 & n41197 ;
  assign n41199 = n41193 | n41198 ;
  assign n41200 = n65686 & n41199 ;
  assign n41201 = n8860 & n78691 ;
  assign n78779 = ~n41201 ;
  assign n41202 = x32 & n78779 ;
  assign n41203 = n8871 & n78691 ;
  assign n41204 = n41202 | n41203 ;
  assign n41205 = x65 & n41204 ;
  assign n40958 = n40868 | n40956 ;
  assign n41206 = n78682 & n40958 ;
  assign n41207 = n40875 | n41206 ;
  assign n41208 = n78686 & n41207 ;
  assign n78780 = ~n41208 ;
  assign n41209 = n8860 & n78780 ;
  assign n78781 = ~n41209 ;
  assign n41210 = x32 & n78781 ;
  assign n41211 = x65 | n41203 ;
  assign n41212 = n41210 | n41211 ;
  assign n78782 = ~n41205 ;
  assign n41213 = n78782 & n41212 ;
  assign n41214 = n8878 | n41213 ;
  assign n41215 = n41203 | n41210 ;
  assign n41216 = n65670 & n41215 ;
  assign n78783 = ~n41216 ;
  assign n41217 = n41214 & n78783 ;
  assign n78784 = ~n41198 ;
  assign n41218 = x66 & n78784 ;
  assign n78785 = ~n41193 ;
  assign n41219 = n78785 & n41218 ;
  assign n41220 = n41200 | n41219 ;
  assign n41221 = n41217 | n41220 ;
  assign n78786 = ~n41200 ;
  assign n41224 = n78786 & n41221 ;
  assign n41225 = n41223 | n41224 ;
  assign n78787 = ~n41192 ;
  assign n41226 = n78787 & n41225 ;
  assign n78788 = ~n41180 ;
  assign n41227 = x68 & n78788 ;
  assign n78789 = ~n41175 ;
  assign n41228 = n78789 & n41227 ;
  assign n41229 = n41182 | n41228 ;
  assign n41230 = n41226 | n41229 ;
  assign n78790 = ~n41182 ;
  assign n41234 = n78790 & n41230 ;
  assign n41235 = n41233 | n41234 ;
  assign n78791 = ~n41174 ;
  assign n41236 = n78791 & n41235 ;
  assign n78792 = ~n41163 ;
  assign n41237 = x70 & n78792 ;
  assign n78793 = ~n41158 ;
  assign n41238 = n78793 & n41237 ;
  assign n41239 = n41165 | n41238 ;
  assign n41240 = n41236 | n41239 ;
  assign n78794 = ~n41165 ;
  assign n41244 = n78794 & n41240 ;
  assign n41245 = n41243 | n41244 ;
  assign n78795 = ~n41157 ;
  assign n41246 = n78795 & n41245 ;
  assign n78796 = ~n41147 ;
  assign n41247 = x72 & n78796 ;
  assign n78797 = ~n41142 ;
  assign n41248 = n78797 & n41247 ;
  assign n41249 = n41149 | n41248 ;
  assign n41250 = n41246 | n41249 ;
  assign n78798 = ~n41149 ;
  assign n41254 = n78798 & n41250 ;
  assign n41255 = n41253 | n41254 ;
  assign n78799 = ~n41141 ;
  assign n41256 = n78799 & n41255 ;
  assign n78800 = ~n41131 ;
  assign n41257 = x74 & n78800 ;
  assign n78801 = ~n41126 ;
  assign n41258 = n78801 & n41257 ;
  assign n41259 = n41133 | n41258 ;
  assign n41260 = n41256 | n41259 ;
  assign n78802 = ~n41133 ;
  assign n41265 = n78802 & n41260 ;
  assign n41266 = n41263 | n41265 ;
  assign n78803 = ~n41125 ;
  assign n41267 = n78803 & n41266 ;
  assign n78804 = ~n41115 ;
  assign n41268 = x76 & n78804 ;
  assign n78805 = ~n41110 ;
  assign n41269 = n78805 & n41268 ;
  assign n41270 = n41117 | n41269 ;
  assign n41272 = n41267 | n41270 ;
  assign n78806 = ~n41117 ;
  assign n41276 = n78806 & n41272 ;
  assign n41277 = n41275 | n41276 ;
  assign n78807 = ~n41109 ;
  assign n41278 = n78807 & n41277 ;
  assign n78808 = ~n41099 ;
  assign n41279 = x78 & n78808 ;
  assign n78809 = ~n41094 ;
  assign n41280 = n78809 & n41279 ;
  assign n41281 = n41101 | n41280 ;
  assign n41283 = n41278 | n41281 ;
  assign n78810 = ~n41101 ;
  assign n41287 = n78810 & n41283 ;
  assign n41288 = n41286 | n41287 ;
  assign n78811 = ~n41093 ;
  assign n41289 = n78811 & n41288 ;
  assign n78812 = ~n41083 ;
  assign n41290 = x80 & n78812 ;
  assign n78813 = ~n41078 ;
  assign n41291 = n78813 & n41290 ;
  assign n41292 = n41085 | n41291 ;
  assign n41293 = n41289 | n41292 ;
  assign n78814 = ~n41085 ;
  assign n41297 = n78814 & n41293 ;
  assign n41298 = n41296 | n41297 ;
  assign n78815 = ~n41077 ;
  assign n41299 = n78815 & n41298 ;
  assign n78816 = ~n41067 ;
  assign n41300 = x82 & n78816 ;
  assign n78817 = ~n41062 ;
  assign n41301 = n78817 & n41300 ;
  assign n41302 = n41069 | n41301 ;
  assign n41303 = n41299 | n41302 ;
  assign n78818 = ~n41069 ;
  assign n41307 = n78818 & n41303 ;
  assign n41308 = n41306 | n41307 ;
  assign n78819 = ~n41061 ;
  assign n41309 = n78819 & n41308 ;
  assign n78820 = ~n41051 ;
  assign n41310 = x84 & n78820 ;
  assign n78821 = ~n41046 ;
  assign n41311 = n78821 & n41310 ;
  assign n41312 = n41053 | n41311 ;
  assign n41313 = n41309 | n41312 ;
  assign n78822 = ~n41053 ;
  assign n41318 = n78822 & n41313 ;
  assign n41319 = n41316 | n41318 ;
  assign n78823 = ~n41045 ;
  assign n41320 = n78823 & n41319 ;
  assign n78824 = ~n41035 ;
  assign n41321 = x86 & n78824 ;
  assign n78825 = ~n41030 ;
  assign n41322 = n78825 & n41321 ;
  assign n41323 = n41037 | n41322 ;
  assign n41324 = n41320 | n41323 ;
  assign n78826 = ~n41037 ;
  assign n41328 = n78826 & n41324 ;
  assign n41329 = n41327 | n41328 ;
  assign n78827 = ~n41029 ;
  assign n41330 = n78827 & n41329 ;
  assign n78828 = ~n41019 ;
  assign n41331 = x88 & n78828 ;
  assign n78829 = ~n41014 ;
  assign n41332 = n78829 & n41331 ;
  assign n41333 = n41021 | n41332 ;
  assign n41334 = n41330 | n41333 ;
  assign n78830 = ~n41021 ;
  assign n41338 = n78830 & n41334 ;
  assign n41339 = n41337 | n41338 ;
  assign n78831 = ~n41013 ;
  assign n41340 = n78831 & n41339 ;
  assign n78832 = ~n41003 ;
  assign n41341 = x90 & n78832 ;
  assign n78833 = ~n40998 ;
  assign n41342 = n78833 & n41341 ;
  assign n41343 = n41005 | n41342 ;
  assign n41344 = n41340 | n41343 ;
  assign n78834 = ~n41005 ;
  assign n41348 = n78834 & n41344 ;
  assign n41349 = n41347 | n41348 ;
  assign n78835 = ~n40997 ;
  assign n41350 = n78835 & n41349 ;
  assign n78836 = ~n40987 ;
  assign n41351 = x92 & n78836 ;
  assign n78837 = ~n40982 ;
  assign n41352 = n78837 & n41351 ;
  assign n41353 = n40989 | n41352 ;
  assign n41354 = n41350 | n41353 ;
  assign n78838 = ~n40989 ;
  assign n41358 = n78838 & n41354 ;
  assign n41359 = n41357 | n41358 ;
  assign n78839 = ~n40981 ;
  assign n41360 = n78839 & n41359 ;
  assign n78840 = ~n40971 ;
  assign n41361 = x94 & n78840 ;
  assign n78841 = ~n40966 ;
  assign n41362 = n78841 & n41361 ;
  assign n41363 = n40973 | n41362 ;
  assign n41364 = n41360 | n41363 ;
  assign n78842 = ~n40973 ;
  assign n41368 = n78842 & n41364 ;
  assign n41369 = n41367 | n41368 ;
  assign n78843 = ~n40965 ;
  assign n41370 = n78843 & n41369 ;
  assign n78844 = ~n40870 ;
  assign n40876 = n78844 & n40875 ;
  assign n41371 = n40473 | n40875 ;
  assign n78845 = ~n41371 ;
  assign n41372 = n40958 & n78845 ;
  assign n41373 = n40876 | n41372 ;
  assign n41374 = n40879 | n41373 ;
  assign n78846 = ~n40471 ;
  assign n41375 = n78846 & n40879 ;
  assign n78847 = ~n41375 ;
  assign n41376 = n41374 & n78847 ;
  assign n41377 = n68438 & n41376 ;
  assign n78848 = ~n40879 ;
  assign n41378 = n78848 & n41373 ;
  assign n41379 = n40471 & n40879 ;
  assign n78849 = ~n41379 ;
  assign n41380 = x96 & n78849 ;
  assign n78850 = ~n41378 ;
  assign n41381 = n78850 & n41380 ;
  assign n41382 = n295 | n41381 ;
  assign n41383 = n41377 | n41382 ;
  assign n41384 = n41370 | n41383 ;
  assign n41385 = n65696 & n41376 ;
  assign n78851 = ~n41385 ;
  assign n41386 = n41384 & n78851 ;
  assign n41458 = n40965 | n41381 ;
  assign n41459 = n41377 | n41458 ;
  assign n78852 = ~n41459 ;
  assign n41460 = n41369 & n78852 ;
  assign n41388 = x65 & n41215 ;
  assign n78853 = ~n41388 ;
  assign n41389 = n41212 & n78853 ;
  assign n41390 = n8878 | n41389 ;
  assign n41391 = n78783 & n41390 ;
  assign n41392 = n41220 | n41391 ;
  assign n41393 = n78786 & n41392 ;
  assign n41394 = n41223 | n41393 ;
  assign n41395 = n78787 & n41394 ;
  assign n41396 = n41229 | n41395 ;
  assign n41397 = n78790 & n41396 ;
  assign n41398 = n41233 | n41397 ;
  assign n41399 = n78791 & n41398 ;
  assign n41400 = n41239 | n41399 ;
  assign n41401 = n78794 & n41400 ;
  assign n41402 = n41243 | n41401 ;
  assign n41403 = n78795 & n41402 ;
  assign n41404 = n41249 | n41403 ;
  assign n41405 = n78798 & n41404 ;
  assign n41406 = n41253 | n41405 ;
  assign n41407 = n78799 & n41406 ;
  assign n41408 = n41259 | n41407 ;
  assign n41409 = n78802 & n41408 ;
  assign n41410 = n41263 | n41409 ;
  assign n41411 = n78803 & n41410 ;
  assign n41412 = n41270 | n41411 ;
  assign n41413 = n78806 & n41412 ;
  assign n41414 = n41275 | n41413 ;
  assign n41415 = n78807 & n41414 ;
  assign n41416 = n41281 | n41415 ;
  assign n41417 = n78810 & n41416 ;
  assign n41418 = n41286 | n41417 ;
  assign n41419 = n78811 & n41418 ;
  assign n41420 = n41292 | n41419 ;
  assign n41421 = n78814 & n41420 ;
  assign n41422 = n41296 | n41421 ;
  assign n41423 = n78815 & n41422 ;
  assign n41424 = n41302 | n41423 ;
  assign n41425 = n78818 & n41424 ;
  assign n41426 = n41306 | n41425 ;
  assign n41427 = n78819 & n41426 ;
  assign n41428 = n41312 | n41427 ;
  assign n41429 = n78822 & n41428 ;
  assign n41430 = n41316 | n41429 ;
  assign n41431 = n78823 & n41430 ;
  assign n41432 = n41323 | n41431 ;
  assign n41433 = n78826 & n41432 ;
  assign n41434 = n41327 | n41433 ;
  assign n41435 = n78827 & n41434 ;
  assign n41436 = n41333 | n41435 ;
  assign n41437 = n78830 & n41436 ;
  assign n41438 = n41337 | n41437 ;
  assign n41439 = n78831 & n41438 ;
  assign n41440 = n41343 | n41439 ;
  assign n41441 = n78834 & n41440 ;
  assign n41442 = n41347 | n41441 ;
  assign n41443 = n78835 & n41442 ;
  assign n41444 = n41353 | n41443 ;
  assign n41445 = n78838 & n41444 ;
  assign n41446 = n41357 | n41445 ;
  assign n41447 = n78839 & n41446 ;
  assign n41448 = n41363 | n41447 ;
  assign n41449 = n78842 & n41448 ;
  assign n41461 = n41367 | n41449 ;
  assign n41462 = n78843 & n41461 ;
  assign n41463 = n41377 | n41381 ;
  assign n78854 = ~n41462 ;
  assign n41464 = n78854 & n41463 ;
  assign n41465 = n41460 | n41464 ;
  assign n78855 = ~n41386 ;
  assign n41466 = n78855 & n41465 ;
  assign n41467 = n303 & n40471 ;
  assign n41468 = n41384 & n41467 ;
  assign n41469 = n41466 | n41468 ;
  assign n41470 = n68545 & n41469 ;
  assign n78856 = ~n41368 ;
  assign n41450 = n41367 & n78856 ;
  assign n41451 = n40973 | n41367 ;
  assign n78857 = ~n41451 ;
  assign n41452 = n41448 & n78857 ;
  assign n41453 = n41450 | n41452 ;
  assign n41454 = n78855 & n41453 ;
  assign n41455 = n40964 & n78851 ;
  assign n41456 = n41384 & n41455 ;
  assign n41457 = n41454 | n41456 ;
  assign n41471 = n68438 & n41457 ;
  assign n78858 = ~n41447 ;
  assign n41472 = n41363 & n78858 ;
  assign n41473 = n40981 | n41363 ;
  assign n78859 = ~n41473 ;
  assign n41474 = n41359 & n78859 ;
  assign n41475 = n41472 | n41474 ;
  assign n41476 = n78855 & n41475 ;
  assign n41477 = n40972 & n78851 ;
  assign n41478 = n41384 & n41477 ;
  assign n41479 = n41476 | n41478 ;
  assign n41480 = n68214 & n41479 ;
  assign n78860 = ~n41358 ;
  assign n41481 = n41357 & n78860 ;
  assign n41482 = n40989 | n41357 ;
  assign n78861 = ~n41482 ;
  assign n41483 = n41444 & n78861 ;
  assign n41484 = n41481 | n41483 ;
  assign n41485 = n78855 & n41484 ;
  assign n41486 = n40980 & n78851 ;
  assign n41487 = n41384 & n41486 ;
  assign n41488 = n41485 | n41487 ;
  assign n41489 = n68058 & n41488 ;
  assign n78862 = ~n41443 ;
  assign n41490 = n41353 & n78862 ;
  assign n41491 = n40997 | n41353 ;
  assign n78863 = ~n41491 ;
  assign n41492 = n41349 & n78863 ;
  assign n41493 = n41490 | n41492 ;
  assign n41494 = n78855 & n41493 ;
  assign n41495 = n40988 & n78851 ;
  assign n41496 = n41384 & n41495 ;
  assign n41497 = n41494 | n41496 ;
  assign n41498 = n67986 & n41497 ;
  assign n78864 = ~n41348 ;
  assign n41499 = n41347 & n78864 ;
  assign n41500 = n41005 | n41347 ;
  assign n78865 = ~n41500 ;
  assign n41501 = n41440 & n78865 ;
  assign n41502 = n41499 | n41501 ;
  assign n41503 = n78855 & n41502 ;
  assign n41504 = n40996 & n78851 ;
  assign n41505 = n41384 & n41504 ;
  assign n41506 = n41503 | n41505 ;
  assign n41507 = n67763 & n41506 ;
  assign n78866 = ~n41439 ;
  assign n41508 = n41343 & n78866 ;
  assign n41509 = n41013 | n41343 ;
  assign n78867 = ~n41509 ;
  assign n41510 = n41339 & n78867 ;
  assign n41511 = n41508 | n41510 ;
  assign n41512 = n78855 & n41511 ;
  assign n41513 = n41004 & n78851 ;
  assign n41514 = n41384 & n41513 ;
  assign n41515 = n41512 | n41514 ;
  assign n41516 = n67622 & n41515 ;
  assign n78868 = ~n41338 ;
  assign n41517 = n41337 & n78868 ;
  assign n41518 = n41021 | n41337 ;
  assign n78869 = ~n41518 ;
  assign n41519 = n41436 & n78869 ;
  assign n41520 = n41517 | n41519 ;
  assign n41521 = n78855 & n41520 ;
  assign n41522 = n41012 & n78851 ;
  assign n41523 = n41384 & n41522 ;
  assign n41524 = n41521 | n41523 ;
  assign n41525 = n67531 & n41524 ;
  assign n78870 = ~n41435 ;
  assign n41526 = n41333 & n78870 ;
  assign n41527 = n41029 | n41333 ;
  assign n78871 = ~n41527 ;
  assign n41528 = n41329 & n78871 ;
  assign n41529 = n41526 | n41528 ;
  assign n41530 = n78855 & n41529 ;
  assign n41531 = n41020 & n78851 ;
  assign n41532 = n41384 & n41531 ;
  assign n41533 = n41530 | n41532 ;
  assign n41534 = n67348 & n41533 ;
  assign n78872 = ~n41328 ;
  assign n41535 = n41327 & n78872 ;
  assign n41536 = n41037 | n41327 ;
  assign n78873 = ~n41536 ;
  assign n41537 = n41432 & n78873 ;
  assign n41538 = n41535 | n41537 ;
  assign n41539 = n78855 & n41538 ;
  assign n41540 = n41028 & n78851 ;
  assign n41541 = n41384 & n41540 ;
  assign n41542 = n41539 | n41541 ;
  assign n41543 = n67222 & n41542 ;
  assign n78874 = ~n41431 ;
  assign n41544 = n41323 & n78874 ;
  assign n41545 = n41045 | n41323 ;
  assign n78875 = ~n41545 ;
  assign n41546 = n41319 & n78875 ;
  assign n41547 = n41544 | n41546 ;
  assign n41548 = n78855 & n41547 ;
  assign n41549 = n41036 & n78851 ;
  assign n41550 = n41384 & n41549 ;
  assign n41551 = n41548 | n41550 ;
  assign n41552 = n67164 & n41551 ;
  assign n78876 = ~n41318 ;
  assign n41553 = n41316 & n78876 ;
  assign n41317 = n41053 | n41316 ;
  assign n78877 = ~n41317 ;
  assign n41554 = n41313 & n78877 ;
  assign n41555 = n41553 | n41554 ;
  assign n41556 = n78855 & n41555 ;
  assign n41557 = n41044 & n78851 ;
  assign n41558 = n41384 & n41557 ;
  assign n41559 = n41556 | n41558 ;
  assign n41560 = n66979 & n41559 ;
  assign n78878 = ~n41427 ;
  assign n41561 = n41312 & n78878 ;
  assign n41562 = n41061 | n41312 ;
  assign n78879 = ~n41562 ;
  assign n41563 = n41308 & n78879 ;
  assign n41564 = n41561 | n41563 ;
  assign n41565 = n78855 & n41564 ;
  assign n41566 = n41052 & n78851 ;
  assign n41567 = n41384 & n41566 ;
  assign n41568 = n41565 | n41567 ;
  assign n41569 = n66868 & n41568 ;
  assign n78880 = ~n41307 ;
  assign n41570 = n41306 & n78880 ;
  assign n41571 = n41069 | n41306 ;
  assign n78881 = ~n41571 ;
  assign n41572 = n41424 & n78881 ;
  assign n41573 = n41570 | n41572 ;
  assign n41574 = n78855 & n41573 ;
  assign n41575 = n41060 & n78851 ;
  assign n41576 = n41384 & n41575 ;
  assign n41577 = n41574 | n41576 ;
  assign n41578 = n66797 & n41577 ;
  assign n78882 = ~n41423 ;
  assign n41579 = n41302 & n78882 ;
  assign n41580 = n41077 | n41302 ;
  assign n78883 = ~n41580 ;
  assign n41581 = n41298 & n78883 ;
  assign n41582 = n41579 | n41581 ;
  assign n41583 = n78855 & n41582 ;
  assign n41584 = n41068 & n78851 ;
  assign n41585 = n41384 & n41584 ;
  assign n41586 = n41583 | n41585 ;
  assign n41587 = n66654 & n41586 ;
  assign n78884 = ~n41297 ;
  assign n41588 = n41296 & n78884 ;
  assign n41589 = n41085 | n41296 ;
  assign n78885 = ~n41589 ;
  assign n41590 = n41420 & n78885 ;
  assign n41591 = n41588 | n41590 ;
  assign n41592 = n78855 & n41591 ;
  assign n41593 = n41076 & n78851 ;
  assign n41594 = n41384 & n41593 ;
  assign n41595 = n41592 | n41594 ;
  assign n41596 = n66560 & n41595 ;
  assign n78886 = ~n41419 ;
  assign n41597 = n41292 & n78886 ;
  assign n41598 = n41093 | n41292 ;
  assign n78887 = ~n41598 ;
  assign n41599 = n41288 & n78887 ;
  assign n41600 = n41597 | n41599 ;
  assign n41601 = n78855 & n41600 ;
  assign n41602 = n41084 & n78851 ;
  assign n41603 = n41384 & n41602 ;
  assign n41604 = n41601 | n41603 ;
  assign n41605 = n66505 & n41604 ;
  assign n78888 = ~n41287 ;
  assign n41606 = n41286 & n78888 ;
  assign n41607 = n41101 | n41286 ;
  assign n78889 = ~n41607 ;
  assign n41608 = n41416 & n78889 ;
  assign n41609 = n41606 | n41608 ;
  assign n41610 = n78855 & n41609 ;
  assign n41611 = n41092 & n78851 ;
  assign n41612 = n41384 & n41611 ;
  assign n41613 = n41610 | n41612 ;
  assign n41614 = n66379 & n41613 ;
  assign n78890 = ~n41415 ;
  assign n41615 = n41281 & n78890 ;
  assign n41282 = n41109 | n41281 ;
  assign n78891 = ~n41282 ;
  assign n41616 = n78891 & n41414 ;
  assign n41617 = n41615 | n41616 ;
  assign n41618 = n78855 & n41617 ;
  assign n41619 = n41100 & n78851 ;
  assign n41620 = n41384 & n41619 ;
  assign n41621 = n41618 | n41620 ;
  assign n41622 = n66299 & n41621 ;
  assign n78892 = ~n41276 ;
  assign n41623 = n41275 & n78892 ;
  assign n41624 = n41117 | n41275 ;
  assign n78893 = ~n41624 ;
  assign n41625 = n41412 & n78893 ;
  assign n41626 = n41623 | n41625 ;
  assign n41627 = n78855 & n41626 ;
  assign n41628 = n41108 & n78851 ;
  assign n41629 = n41384 & n41628 ;
  assign n41630 = n41627 | n41629 ;
  assign n41631 = n66244 & n41630 ;
  assign n78894 = ~n41411 ;
  assign n41632 = n41270 & n78894 ;
  assign n41271 = n41125 | n41270 ;
  assign n78895 = ~n41271 ;
  assign n41633 = n78895 & n41410 ;
  assign n41634 = n41632 | n41633 ;
  assign n41635 = n78855 & n41634 ;
  assign n41636 = n41116 & n78851 ;
  assign n41637 = n41384 & n41636 ;
  assign n41638 = n41635 | n41637 ;
  assign n41639 = n66145 & n41638 ;
  assign n78896 = ~n41265 ;
  assign n41640 = n41263 & n78896 ;
  assign n41264 = n41133 | n41263 ;
  assign n78897 = ~n41264 ;
  assign n41641 = n41260 & n78897 ;
  assign n41642 = n41640 | n41641 ;
  assign n41643 = n78855 & n41642 ;
  assign n41644 = n41124 & n78851 ;
  assign n41645 = n41384 & n41644 ;
  assign n41646 = n41643 | n41645 ;
  assign n41647 = n66081 & n41646 ;
  assign n78898 = ~n41407 ;
  assign n41648 = n41259 & n78898 ;
  assign n41649 = n41141 | n41259 ;
  assign n78899 = ~n41649 ;
  assign n41650 = n41255 & n78899 ;
  assign n41651 = n41648 | n41650 ;
  assign n41652 = n78855 & n41651 ;
  assign n41653 = n41132 & n78851 ;
  assign n41654 = n41384 & n41653 ;
  assign n41655 = n41652 | n41654 ;
  assign n41656 = n66043 & n41655 ;
  assign n78900 = ~n41254 ;
  assign n41657 = n41253 & n78900 ;
  assign n41658 = n41149 | n41253 ;
  assign n78901 = ~n41658 ;
  assign n41659 = n41404 & n78901 ;
  assign n41660 = n41657 | n41659 ;
  assign n41661 = n78855 & n41660 ;
  assign n41662 = n41140 & n78851 ;
  assign n41663 = n41384 & n41662 ;
  assign n41664 = n41661 | n41663 ;
  assign n41665 = n65960 & n41664 ;
  assign n78902 = ~n41403 ;
  assign n41666 = n41249 & n78902 ;
  assign n41667 = n41157 | n41249 ;
  assign n78903 = ~n41667 ;
  assign n41668 = n41245 & n78903 ;
  assign n41669 = n41666 | n41668 ;
  assign n41670 = n78855 & n41669 ;
  assign n41671 = n41148 & n78851 ;
  assign n41672 = n41384 & n41671 ;
  assign n41673 = n41670 | n41672 ;
  assign n41674 = n65909 & n41673 ;
  assign n78904 = ~n41244 ;
  assign n41675 = n41243 & n78904 ;
  assign n41676 = n41165 | n41243 ;
  assign n78905 = ~n41676 ;
  assign n41677 = n41400 & n78905 ;
  assign n41678 = n41675 | n41677 ;
  assign n41679 = n78855 & n41678 ;
  assign n41680 = n41156 & n78851 ;
  assign n41681 = n41384 & n41680 ;
  assign n41682 = n41679 | n41681 ;
  assign n41683 = n65877 & n41682 ;
  assign n78906 = ~n41399 ;
  assign n41684 = n41239 & n78906 ;
  assign n41685 = n41174 | n41239 ;
  assign n78907 = ~n41685 ;
  assign n41686 = n41235 & n78907 ;
  assign n41687 = n41684 | n41686 ;
  assign n41688 = n78855 & n41687 ;
  assign n41689 = n41164 & n78851 ;
  assign n41690 = n41384 & n41689 ;
  assign n41691 = n41688 | n41690 ;
  assign n41692 = n65820 & n41691 ;
  assign n78908 = ~n41234 ;
  assign n41694 = n41233 & n78908 ;
  assign n41693 = n41182 | n41233 ;
  assign n78909 = ~n41693 ;
  assign n41695 = n41230 & n78909 ;
  assign n41696 = n41694 | n41695 ;
  assign n41697 = n78855 & n41696 ;
  assign n41698 = n41173 & n78851 ;
  assign n41699 = n41384 & n41698 ;
  assign n41700 = n41697 | n41699 ;
  assign n41701 = n65791 & n41700 ;
  assign n78910 = ~n41395 ;
  assign n41702 = n41229 & n78910 ;
  assign n41703 = n41192 | n41229 ;
  assign n78911 = ~n41703 ;
  assign n41704 = n41225 & n78911 ;
  assign n41705 = n41702 | n41704 ;
  assign n41706 = n78855 & n41705 ;
  assign n41707 = n41181 & n78851 ;
  assign n41708 = n41384 & n41707 ;
  assign n41709 = n41706 | n41708 ;
  assign n41710 = n65772 & n41709 ;
  assign n78912 = ~n41224 ;
  assign n41712 = n41223 & n78912 ;
  assign n41711 = n41200 | n41223 ;
  assign n78913 = ~n41711 ;
  assign n41713 = n41221 & n78913 ;
  assign n41714 = n41712 | n41713 ;
  assign n41715 = n78855 & n41714 ;
  assign n41716 = n41190 & n78851 ;
  assign n41717 = n41384 & n41716 ;
  assign n41718 = n41715 | n41717 ;
  assign n41719 = n65746 & n41718 ;
  assign n78914 = ~n41391 ;
  assign n41721 = n41220 & n78914 ;
  assign n41720 = n41216 | n41220 ;
  assign n78915 = ~n41720 ;
  assign n41722 = n41390 & n78915 ;
  assign n41723 = n41721 | n41722 ;
  assign n41724 = n78855 & n41723 ;
  assign n41725 = n41199 & n78851 ;
  assign n41726 = n41384 & n41725 ;
  assign n41727 = n41724 | n41726 ;
  assign n41728 = n65721 & n41727 ;
  assign n41729 = n8878 & n41212 ;
  assign n41730 = n78853 & n41729 ;
  assign n78916 = ~n41730 ;
  assign n41731 = n41390 & n78916 ;
  assign n41732 = n78855 & n41731 ;
  assign n41733 = n41215 & n78851 ;
  assign n41734 = n41384 & n41733 ;
  assign n41735 = n41732 | n41734 ;
  assign n41736 = n65686 & n41735 ;
  assign n41387 = n8878 & n78855 ;
  assign n41741 = x64 & n78855 ;
  assign n78917 = ~n41741 ;
  assign n41742 = x31 & n78917 ;
  assign n41743 = n41387 | n41742 ;
  assign n41745 = x65 & n41743 ;
  assign n41737 = n41383 | n41462 ;
  assign n41738 = n78851 & n41737 ;
  assign n78918 = ~n41738 ;
  assign n41739 = x64 & n78918 ;
  assign n78919 = ~n41739 ;
  assign n41740 = x31 & n78919 ;
  assign n41744 = x65 | n41387 ;
  assign n41746 = n41740 | n41744 ;
  assign n78920 = ~n41745 ;
  assign n41747 = n78920 & n41746 ;
  assign n41748 = n9415 | n41747 ;
  assign n41749 = n65670 & n41743 ;
  assign n78921 = ~n41749 ;
  assign n41750 = n41748 & n78921 ;
  assign n78922 = ~n41734 ;
  assign n41751 = x66 & n78922 ;
  assign n78923 = ~n41732 ;
  assign n41752 = n78923 & n41751 ;
  assign n41753 = n41736 | n41752 ;
  assign n41754 = n41750 | n41753 ;
  assign n78924 = ~n41736 ;
  assign n41755 = n78924 & n41754 ;
  assign n78925 = ~n41726 ;
  assign n41756 = x67 & n78925 ;
  assign n78926 = ~n41724 ;
  assign n41757 = n78926 & n41756 ;
  assign n41758 = n41755 | n41757 ;
  assign n78927 = ~n41728 ;
  assign n41759 = n78927 & n41758 ;
  assign n78928 = ~n41717 ;
  assign n41760 = x68 & n78928 ;
  assign n78929 = ~n41715 ;
  assign n41761 = n78929 & n41760 ;
  assign n41762 = n41719 | n41761 ;
  assign n41763 = n41759 | n41762 ;
  assign n78930 = ~n41719 ;
  assign n41764 = n78930 & n41763 ;
  assign n78931 = ~n41708 ;
  assign n41765 = x69 & n78931 ;
  assign n78932 = ~n41706 ;
  assign n41766 = n78932 & n41765 ;
  assign n41767 = n41764 | n41766 ;
  assign n78933 = ~n41710 ;
  assign n41768 = n78933 & n41767 ;
  assign n78934 = ~n41699 ;
  assign n41769 = x70 & n78934 ;
  assign n78935 = ~n41697 ;
  assign n41770 = n78935 & n41769 ;
  assign n41771 = n41701 | n41770 ;
  assign n41772 = n41768 | n41771 ;
  assign n78936 = ~n41701 ;
  assign n41773 = n78936 & n41772 ;
  assign n78937 = ~n41690 ;
  assign n41774 = x71 & n78937 ;
  assign n78938 = ~n41688 ;
  assign n41775 = n78938 & n41774 ;
  assign n41776 = n41692 | n41775 ;
  assign n41779 = n41773 | n41776 ;
  assign n78939 = ~n41692 ;
  assign n41780 = n78939 & n41779 ;
  assign n78940 = ~n41681 ;
  assign n41781 = x72 & n78940 ;
  assign n78941 = ~n41679 ;
  assign n41782 = n78941 & n41781 ;
  assign n41783 = n41683 | n41782 ;
  assign n41784 = n41780 | n41783 ;
  assign n78942 = ~n41683 ;
  assign n41785 = n78942 & n41784 ;
  assign n78943 = ~n41672 ;
  assign n41786 = x73 & n78943 ;
  assign n78944 = ~n41670 ;
  assign n41787 = n78944 & n41786 ;
  assign n41788 = n41674 | n41787 ;
  assign n41790 = n41785 | n41788 ;
  assign n78945 = ~n41674 ;
  assign n41791 = n78945 & n41790 ;
  assign n78946 = ~n41663 ;
  assign n41792 = x74 & n78946 ;
  assign n78947 = ~n41661 ;
  assign n41793 = n78947 & n41792 ;
  assign n41794 = n41665 | n41793 ;
  assign n41795 = n41791 | n41794 ;
  assign n78948 = ~n41665 ;
  assign n41796 = n78948 & n41795 ;
  assign n78949 = ~n41654 ;
  assign n41797 = x75 & n78949 ;
  assign n78950 = ~n41652 ;
  assign n41798 = n78950 & n41797 ;
  assign n41799 = n41656 | n41798 ;
  assign n41801 = n41796 | n41799 ;
  assign n78951 = ~n41656 ;
  assign n41802 = n78951 & n41801 ;
  assign n78952 = ~n41645 ;
  assign n41803 = x76 & n78952 ;
  assign n78953 = ~n41643 ;
  assign n41804 = n78953 & n41803 ;
  assign n41805 = n41647 | n41804 ;
  assign n41806 = n41802 | n41805 ;
  assign n78954 = ~n41647 ;
  assign n41807 = n78954 & n41806 ;
  assign n78955 = ~n41637 ;
  assign n41808 = x77 & n78955 ;
  assign n78956 = ~n41635 ;
  assign n41809 = n78956 & n41808 ;
  assign n41810 = n41639 | n41809 ;
  assign n41812 = n41807 | n41810 ;
  assign n78957 = ~n41639 ;
  assign n41813 = n78957 & n41812 ;
  assign n78958 = ~n41629 ;
  assign n41814 = x78 & n78958 ;
  assign n78959 = ~n41627 ;
  assign n41815 = n78959 & n41814 ;
  assign n41816 = n41631 | n41815 ;
  assign n41817 = n41813 | n41816 ;
  assign n78960 = ~n41631 ;
  assign n41818 = n78960 & n41817 ;
  assign n78961 = ~n41620 ;
  assign n41819 = x79 & n78961 ;
  assign n78962 = ~n41618 ;
  assign n41820 = n78962 & n41819 ;
  assign n41821 = n41622 | n41820 ;
  assign n41823 = n41818 | n41821 ;
  assign n78963 = ~n41622 ;
  assign n41824 = n78963 & n41823 ;
  assign n78964 = ~n41612 ;
  assign n41825 = x80 & n78964 ;
  assign n78965 = ~n41610 ;
  assign n41826 = n78965 & n41825 ;
  assign n41827 = n41614 | n41826 ;
  assign n41828 = n41824 | n41827 ;
  assign n78966 = ~n41614 ;
  assign n41829 = n78966 & n41828 ;
  assign n78967 = ~n41603 ;
  assign n41830 = x81 & n78967 ;
  assign n78968 = ~n41601 ;
  assign n41831 = n78968 & n41830 ;
  assign n41832 = n41605 | n41831 ;
  assign n41834 = n41829 | n41832 ;
  assign n78969 = ~n41605 ;
  assign n41835 = n78969 & n41834 ;
  assign n78970 = ~n41594 ;
  assign n41836 = x82 & n78970 ;
  assign n78971 = ~n41592 ;
  assign n41837 = n78971 & n41836 ;
  assign n41838 = n41596 | n41837 ;
  assign n41839 = n41835 | n41838 ;
  assign n78972 = ~n41596 ;
  assign n41840 = n78972 & n41839 ;
  assign n78973 = ~n41585 ;
  assign n41841 = x83 & n78973 ;
  assign n78974 = ~n41583 ;
  assign n41842 = n78974 & n41841 ;
  assign n41843 = n41587 | n41842 ;
  assign n41845 = n41840 | n41843 ;
  assign n78975 = ~n41587 ;
  assign n41846 = n78975 & n41845 ;
  assign n78976 = ~n41576 ;
  assign n41847 = x84 & n78976 ;
  assign n78977 = ~n41574 ;
  assign n41848 = n78977 & n41847 ;
  assign n41849 = n41578 | n41848 ;
  assign n41850 = n41846 | n41849 ;
  assign n78978 = ~n41578 ;
  assign n41851 = n78978 & n41850 ;
  assign n78979 = ~n41567 ;
  assign n41852 = x85 & n78979 ;
  assign n78980 = ~n41565 ;
  assign n41853 = n78980 & n41852 ;
  assign n41854 = n41569 | n41853 ;
  assign n41856 = n41851 | n41854 ;
  assign n78981 = ~n41569 ;
  assign n41857 = n78981 & n41856 ;
  assign n78982 = ~n41558 ;
  assign n41858 = x86 & n78982 ;
  assign n78983 = ~n41556 ;
  assign n41859 = n78983 & n41858 ;
  assign n41860 = n41560 | n41859 ;
  assign n41861 = n41857 | n41860 ;
  assign n78984 = ~n41560 ;
  assign n41862 = n78984 & n41861 ;
  assign n78985 = ~n41550 ;
  assign n41863 = x87 & n78985 ;
  assign n78986 = ~n41548 ;
  assign n41864 = n78986 & n41863 ;
  assign n41865 = n41552 | n41864 ;
  assign n41867 = n41862 | n41865 ;
  assign n78987 = ~n41552 ;
  assign n41868 = n78987 & n41867 ;
  assign n78988 = ~n41541 ;
  assign n41869 = x88 & n78988 ;
  assign n78989 = ~n41539 ;
  assign n41870 = n78989 & n41869 ;
  assign n41871 = n41543 | n41870 ;
  assign n41872 = n41868 | n41871 ;
  assign n78990 = ~n41543 ;
  assign n41873 = n78990 & n41872 ;
  assign n78991 = ~n41532 ;
  assign n41874 = x89 & n78991 ;
  assign n78992 = ~n41530 ;
  assign n41875 = n78992 & n41874 ;
  assign n41876 = n41534 | n41875 ;
  assign n41878 = n41873 | n41876 ;
  assign n78993 = ~n41534 ;
  assign n41879 = n78993 & n41878 ;
  assign n78994 = ~n41523 ;
  assign n41880 = x90 & n78994 ;
  assign n78995 = ~n41521 ;
  assign n41881 = n78995 & n41880 ;
  assign n41882 = n41525 | n41881 ;
  assign n41883 = n41879 | n41882 ;
  assign n78996 = ~n41525 ;
  assign n41884 = n78996 & n41883 ;
  assign n78997 = ~n41514 ;
  assign n41885 = x91 & n78997 ;
  assign n78998 = ~n41512 ;
  assign n41886 = n78998 & n41885 ;
  assign n41887 = n41516 | n41886 ;
  assign n41889 = n41884 | n41887 ;
  assign n78999 = ~n41516 ;
  assign n41890 = n78999 & n41889 ;
  assign n79000 = ~n41505 ;
  assign n41891 = x92 & n79000 ;
  assign n79001 = ~n41503 ;
  assign n41892 = n79001 & n41891 ;
  assign n41893 = n41507 | n41892 ;
  assign n41894 = n41890 | n41893 ;
  assign n79002 = ~n41507 ;
  assign n41895 = n79002 & n41894 ;
  assign n79003 = ~n41496 ;
  assign n41896 = x93 & n79003 ;
  assign n79004 = ~n41494 ;
  assign n41897 = n79004 & n41896 ;
  assign n41898 = n41498 | n41897 ;
  assign n41900 = n41895 | n41898 ;
  assign n79005 = ~n41498 ;
  assign n41901 = n79005 & n41900 ;
  assign n79006 = ~n41487 ;
  assign n41902 = x94 & n79006 ;
  assign n79007 = ~n41485 ;
  assign n41903 = n79007 & n41902 ;
  assign n41904 = n41489 | n41903 ;
  assign n41905 = n41901 | n41904 ;
  assign n79008 = ~n41489 ;
  assign n41906 = n79008 & n41905 ;
  assign n79009 = ~n41478 ;
  assign n41907 = x95 & n79009 ;
  assign n79010 = ~n41476 ;
  assign n41908 = n79010 & n41907 ;
  assign n41909 = n41480 | n41908 ;
  assign n41911 = n41906 | n41909 ;
  assign n79011 = ~n41480 ;
  assign n41912 = n79011 & n41911 ;
  assign n79012 = ~n41456 ;
  assign n41913 = x96 & n79012 ;
  assign n79013 = ~n41454 ;
  assign n41914 = n79013 & n41913 ;
  assign n41915 = n41471 | n41914 ;
  assign n41916 = n41912 | n41915 ;
  assign n79014 = ~n41471 ;
  assign n41917 = n79014 & n41916 ;
  assign n79015 = ~n41468 ;
  assign n41918 = x97 & n79015 ;
  assign n79016 = ~n41466 ;
  assign n41919 = n79016 & n41918 ;
  assign n41920 = n41470 | n41919 ;
  assign n41922 = n41917 | n41920 ;
  assign n79017 = ~n41470 ;
  assign n41923 = n79017 & n41922 ;
  assign n41924 = n9610 | n41923 ;
  assign n79018 = ~n41469 ;
  assign n41928 = n79018 & n41924 ;
  assign n79019 = ~n41917 ;
  assign n41921 = n79019 & n41920 ;
  assign n41932 = n41387 | n41740 ;
  assign n41933 = x65 & n41932 ;
  assign n79020 = ~n41933 ;
  assign n41934 = n41746 & n79020 ;
  assign n41935 = n9415 | n41934 ;
  assign n41936 = n78921 & n41935 ;
  assign n41937 = n41753 | n41936 ;
  assign n41938 = n78924 & n41937 ;
  assign n41939 = n41728 | n41757 ;
  assign n41941 = n41938 | n41939 ;
  assign n41942 = n78927 & n41941 ;
  assign n41943 = n41761 | n41942 ;
  assign n41945 = n78930 & n41943 ;
  assign n41946 = n41710 | n41766 ;
  assign n41948 = n41945 | n41946 ;
  assign n41949 = n78933 & n41948 ;
  assign n41950 = n41770 | n41949 ;
  assign n41952 = n78936 & n41950 ;
  assign n41953 = n41776 | n41952 ;
  assign n41954 = n78939 & n41953 ;
  assign n41955 = n41783 | n41954 ;
  assign n41957 = n78942 & n41955 ;
  assign n41958 = n41788 | n41957 ;
  assign n41959 = n78945 & n41958 ;
  assign n41960 = n41794 | n41959 ;
  assign n41962 = n78948 & n41960 ;
  assign n41963 = n41799 | n41962 ;
  assign n41964 = n78951 & n41963 ;
  assign n41965 = n41805 | n41964 ;
  assign n41967 = n78954 & n41965 ;
  assign n41968 = n41810 | n41967 ;
  assign n41969 = n78957 & n41968 ;
  assign n41970 = n41816 | n41969 ;
  assign n41972 = n78960 & n41970 ;
  assign n41973 = n41821 | n41972 ;
  assign n41974 = n78963 & n41973 ;
  assign n41975 = n41827 | n41974 ;
  assign n41977 = n78966 & n41975 ;
  assign n41978 = n41832 | n41977 ;
  assign n41979 = n78969 & n41978 ;
  assign n41980 = n41838 | n41979 ;
  assign n41982 = n78972 & n41980 ;
  assign n41983 = n41843 | n41982 ;
  assign n41984 = n78975 & n41983 ;
  assign n41985 = n41849 | n41984 ;
  assign n41987 = n78978 & n41985 ;
  assign n41988 = n41854 | n41987 ;
  assign n41989 = n78981 & n41988 ;
  assign n41990 = n41860 | n41989 ;
  assign n41992 = n78984 & n41990 ;
  assign n41993 = n41865 | n41992 ;
  assign n41994 = n78987 & n41993 ;
  assign n41995 = n41871 | n41994 ;
  assign n41997 = n78990 & n41995 ;
  assign n41998 = n41876 | n41997 ;
  assign n41999 = n78993 & n41998 ;
  assign n42000 = n41882 | n41999 ;
  assign n42002 = n78996 & n42000 ;
  assign n42003 = n41887 | n42002 ;
  assign n42004 = n78999 & n42003 ;
  assign n42005 = n41893 | n42004 ;
  assign n42007 = n79002 & n42005 ;
  assign n42008 = n41898 | n42007 ;
  assign n42009 = n79005 & n42008 ;
  assign n42010 = n41904 | n42009 ;
  assign n42012 = n79008 & n42010 ;
  assign n42013 = n41909 | n42012 ;
  assign n42014 = n79011 & n42013 ;
  assign n42016 = n41915 | n42014 ;
  assign n42023 = n41471 | n41920 ;
  assign n79021 = ~n42023 ;
  assign n42024 = n42016 & n79021 ;
  assign n42025 = n41921 | n42024 ;
  assign n42026 = n41924 | n42025 ;
  assign n79022 = ~n41928 ;
  assign n42027 = n79022 & n42026 ;
  assign n42028 = n68716 & n42027 ;
  assign n79023 = ~n41924 ;
  assign n42479 = n79023 & n42025 ;
  assign n42480 = n41469 & n41924 ;
  assign n79024 = ~n42480 ;
  assign n42481 = x98 & n79024 ;
  assign n79025 = ~n42479 ;
  assign n42482 = n79025 & n42481 ;
  assign n42483 = n42028 | n42482 ;
  assign n41930 = n41457 & n41924 ;
  assign n79026 = ~n42014 ;
  assign n42015 = n41915 & n79026 ;
  assign n42017 = n41480 | n41915 ;
  assign n79027 = ~n42017 ;
  assign n42018 = n41911 & n79027 ;
  assign n42019 = n42015 | n42018 ;
  assign n42020 = n68710 & n42019 ;
  assign n79028 = ~n41923 ;
  assign n42021 = n79028 & n42020 ;
  assign n42022 = n41930 | n42021 ;
  assign n42029 = n68545 & n42022 ;
  assign n42030 = n41479 & n41924 ;
  assign n79029 = ~n41906 ;
  assign n41910 = n79029 & n41909 ;
  assign n42031 = n41489 | n41909 ;
  assign n79030 = ~n42031 ;
  assign n42032 = n42010 & n79030 ;
  assign n42033 = n41910 | n42032 ;
  assign n42034 = n68710 & n42033 ;
  assign n42035 = n79028 & n42034 ;
  assign n42036 = n42030 | n42035 ;
  assign n42037 = n68438 & n42036 ;
  assign n79031 = ~n42035 ;
  assign n42467 = x96 & n79031 ;
  assign n79032 = ~n42030 ;
  assign n42468 = n79032 & n42467 ;
  assign n42469 = n42037 | n42468 ;
  assign n42038 = n41488 & n41924 ;
  assign n79033 = ~n42009 ;
  assign n42011 = n41904 & n79033 ;
  assign n42039 = n41498 | n41904 ;
  assign n79034 = ~n42039 ;
  assign n42040 = n41900 & n79034 ;
  assign n42041 = n42011 | n42040 ;
  assign n42042 = n68710 & n42041 ;
  assign n42043 = n79028 & n42042 ;
  assign n42044 = n42038 | n42043 ;
  assign n42045 = n68214 & n42044 ;
  assign n42046 = n41497 & n41924 ;
  assign n79035 = ~n41895 ;
  assign n41899 = n79035 & n41898 ;
  assign n42047 = n41507 | n41898 ;
  assign n79036 = ~n42047 ;
  assign n42048 = n42005 & n79036 ;
  assign n42049 = n41899 | n42048 ;
  assign n42050 = n68710 & n42049 ;
  assign n42051 = n79028 & n42050 ;
  assign n42052 = n42046 | n42051 ;
  assign n42053 = n68058 & n42052 ;
  assign n79037 = ~n42051 ;
  assign n42455 = x94 & n79037 ;
  assign n79038 = ~n42046 ;
  assign n42456 = n79038 & n42455 ;
  assign n42457 = n42053 | n42456 ;
  assign n42054 = n41506 & n41924 ;
  assign n79039 = ~n42004 ;
  assign n42006 = n41893 & n79039 ;
  assign n42055 = n41516 | n41893 ;
  assign n79040 = ~n42055 ;
  assign n42056 = n41889 & n79040 ;
  assign n42057 = n42006 | n42056 ;
  assign n42058 = n68710 & n42057 ;
  assign n42059 = n79028 & n42058 ;
  assign n42060 = n42054 | n42059 ;
  assign n42061 = n67986 & n42060 ;
  assign n42062 = n41515 & n41924 ;
  assign n79041 = ~n41884 ;
  assign n41888 = n79041 & n41887 ;
  assign n42063 = n41525 | n41887 ;
  assign n79042 = ~n42063 ;
  assign n42064 = n42000 & n79042 ;
  assign n42065 = n41888 | n42064 ;
  assign n42066 = n68710 & n42065 ;
  assign n42067 = n79028 & n42066 ;
  assign n42068 = n42062 | n42067 ;
  assign n42069 = n67763 & n42068 ;
  assign n79043 = ~n42067 ;
  assign n42443 = x92 & n79043 ;
  assign n79044 = ~n42062 ;
  assign n42444 = n79044 & n42443 ;
  assign n42445 = n42069 | n42444 ;
  assign n42070 = n41524 & n41924 ;
  assign n79045 = ~n41999 ;
  assign n42001 = n41882 & n79045 ;
  assign n42071 = n41534 | n41882 ;
  assign n79046 = ~n42071 ;
  assign n42072 = n41878 & n79046 ;
  assign n42073 = n42001 | n42072 ;
  assign n42074 = n68710 & n42073 ;
  assign n42075 = n79028 & n42074 ;
  assign n42076 = n42070 | n42075 ;
  assign n42077 = n67622 & n42076 ;
  assign n42078 = n41533 & n41924 ;
  assign n79047 = ~n41873 ;
  assign n41877 = n79047 & n41876 ;
  assign n42079 = n41543 | n41876 ;
  assign n79048 = ~n42079 ;
  assign n42080 = n41995 & n79048 ;
  assign n42081 = n41877 | n42080 ;
  assign n42082 = n68710 & n42081 ;
  assign n42083 = n79028 & n42082 ;
  assign n42084 = n42078 | n42083 ;
  assign n42085 = n67531 & n42084 ;
  assign n79049 = ~n42083 ;
  assign n42431 = x90 & n79049 ;
  assign n79050 = ~n42078 ;
  assign n42432 = n79050 & n42431 ;
  assign n42433 = n42085 | n42432 ;
  assign n42086 = n41542 & n41924 ;
  assign n79051 = ~n41994 ;
  assign n41996 = n41871 & n79051 ;
  assign n42087 = n41552 | n41871 ;
  assign n79052 = ~n42087 ;
  assign n42088 = n41867 & n79052 ;
  assign n42089 = n41996 | n42088 ;
  assign n42090 = n68710 & n42089 ;
  assign n42091 = n79028 & n42090 ;
  assign n42092 = n42086 | n42091 ;
  assign n42093 = n67348 & n42092 ;
  assign n42094 = n41551 & n41924 ;
  assign n79053 = ~n41862 ;
  assign n41866 = n79053 & n41865 ;
  assign n42095 = n41560 | n41865 ;
  assign n79054 = ~n42095 ;
  assign n42096 = n41990 & n79054 ;
  assign n42097 = n41866 | n42096 ;
  assign n42098 = n68710 & n42097 ;
  assign n42099 = n79028 & n42098 ;
  assign n42100 = n42094 | n42099 ;
  assign n42101 = n67222 & n42100 ;
  assign n79055 = ~n42099 ;
  assign n42419 = x88 & n79055 ;
  assign n79056 = ~n42094 ;
  assign n42420 = n79056 & n42419 ;
  assign n42421 = n42101 | n42420 ;
  assign n42102 = n41559 & n41924 ;
  assign n79057 = ~n41989 ;
  assign n41991 = n41860 & n79057 ;
  assign n42103 = n41569 | n41860 ;
  assign n79058 = ~n42103 ;
  assign n42104 = n41856 & n79058 ;
  assign n42105 = n41991 | n42104 ;
  assign n42106 = n68710 & n42105 ;
  assign n42107 = n79028 & n42106 ;
  assign n42108 = n42102 | n42107 ;
  assign n42109 = n67164 & n42108 ;
  assign n42110 = n41568 & n41924 ;
  assign n79059 = ~n41851 ;
  assign n41855 = n79059 & n41854 ;
  assign n42111 = n41578 | n41854 ;
  assign n79060 = ~n42111 ;
  assign n42112 = n41985 & n79060 ;
  assign n42113 = n41855 | n42112 ;
  assign n42114 = n68710 & n42113 ;
  assign n42115 = n79028 & n42114 ;
  assign n42116 = n42110 | n42115 ;
  assign n42117 = n66979 & n42116 ;
  assign n79061 = ~n42115 ;
  assign n42407 = x86 & n79061 ;
  assign n79062 = ~n42110 ;
  assign n42408 = n79062 & n42407 ;
  assign n42409 = n42117 | n42408 ;
  assign n42118 = n41577 & n41924 ;
  assign n79063 = ~n41984 ;
  assign n41986 = n41849 & n79063 ;
  assign n42119 = n41587 | n41849 ;
  assign n79064 = ~n42119 ;
  assign n42120 = n41845 & n79064 ;
  assign n42121 = n41986 | n42120 ;
  assign n42122 = n68710 & n42121 ;
  assign n42123 = n79028 & n42122 ;
  assign n42124 = n42118 | n42123 ;
  assign n42125 = n66868 & n42124 ;
  assign n42126 = n41586 & n41924 ;
  assign n79065 = ~n41840 ;
  assign n41844 = n79065 & n41843 ;
  assign n42127 = n41596 | n41843 ;
  assign n79066 = ~n42127 ;
  assign n42128 = n41980 & n79066 ;
  assign n42129 = n41844 | n42128 ;
  assign n42130 = n68710 & n42129 ;
  assign n42131 = n79028 & n42130 ;
  assign n42132 = n42126 | n42131 ;
  assign n42133 = n66797 & n42132 ;
  assign n79067 = ~n42131 ;
  assign n42395 = x84 & n79067 ;
  assign n79068 = ~n42126 ;
  assign n42396 = n79068 & n42395 ;
  assign n42397 = n42133 | n42396 ;
  assign n42134 = n41595 & n41924 ;
  assign n79069 = ~n41979 ;
  assign n41981 = n41838 & n79069 ;
  assign n42135 = n41605 | n41838 ;
  assign n79070 = ~n42135 ;
  assign n42136 = n41834 & n79070 ;
  assign n42137 = n41981 | n42136 ;
  assign n42138 = n68710 & n42137 ;
  assign n42139 = n79028 & n42138 ;
  assign n42140 = n42134 | n42139 ;
  assign n42141 = n66654 & n42140 ;
  assign n42142 = n41604 & n41924 ;
  assign n79071 = ~n41829 ;
  assign n41833 = n79071 & n41832 ;
  assign n42143 = n41614 | n41832 ;
  assign n79072 = ~n42143 ;
  assign n42144 = n41975 & n79072 ;
  assign n42145 = n41833 | n42144 ;
  assign n42146 = n68710 & n42145 ;
  assign n42147 = n79028 & n42146 ;
  assign n42148 = n42142 | n42147 ;
  assign n42149 = n66560 & n42148 ;
  assign n79073 = ~n42147 ;
  assign n42383 = x82 & n79073 ;
  assign n79074 = ~n42142 ;
  assign n42384 = n79074 & n42383 ;
  assign n42385 = n42149 | n42384 ;
  assign n42150 = n41613 & n41924 ;
  assign n79075 = ~n41974 ;
  assign n41976 = n41827 & n79075 ;
  assign n42151 = n41622 | n41827 ;
  assign n79076 = ~n42151 ;
  assign n42152 = n41823 & n79076 ;
  assign n42153 = n41976 | n42152 ;
  assign n42154 = n68710 & n42153 ;
  assign n42155 = n79028 & n42154 ;
  assign n42156 = n42150 | n42155 ;
  assign n42157 = n66505 & n42156 ;
  assign n42158 = n41621 & n41924 ;
  assign n79077 = ~n41818 ;
  assign n41822 = n79077 & n41821 ;
  assign n42159 = n41631 | n41821 ;
  assign n79078 = ~n42159 ;
  assign n42160 = n41970 & n79078 ;
  assign n42161 = n41822 | n42160 ;
  assign n42162 = n68710 & n42161 ;
  assign n42163 = n79028 & n42162 ;
  assign n42164 = n42158 | n42163 ;
  assign n42165 = n66379 & n42164 ;
  assign n79079 = ~n42163 ;
  assign n42371 = x80 & n79079 ;
  assign n79080 = ~n42158 ;
  assign n42372 = n79080 & n42371 ;
  assign n42373 = n42165 | n42372 ;
  assign n42166 = n41630 & n41924 ;
  assign n79081 = ~n41969 ;
  assign n41971 = n41816 & n79081 ;
  assign n42167 = n41639 | n41816 ;
  assign n79082 = ~n42167 ;
  assign n42168 = n41812 & n79082 ;
  assign n42169 = n41971 | n42168 ;
  assign n42170 = n68710 & n42169 ;
  assign n42171 = n79028 & n42170 ;
  assign n42172 = n42166 | n42171 ;
  assign n42173 = n66299 & n42172 ;
  assign n42174 = n41638 & n41924 ;
  assign n79083 = ~n41807 ;
  assign n41811 = n79083 & n41810 ;
  assign n42175 = n41647 | n41810 ;
  assign n79084 = ~n42175 ;
  assign n42176 = n41965 & n79084 ;
  assign n42177 = n41811 | n42176 ;
  assign n42178 = n68710 & n42177 ;
  assign n42179 = n79028 & n42178 ;
  assign n42180 = n42174 | n42179 ;
  assign n42181 = n66244 & n42180 ;
  assign n79085 = ~n42179 ;
  assign n42359 = x78 & n79085 ;
  assign n79086 = ~n42174 ;
  assign n42360 = n79086 & n42359 ;
  assign n42361 = n42181 | n42360 ;
  assign n42182 = n41646 & n41924 ;
  assign n79087 = ~n41964 ;
  assign n41966 = n41805 & n79087 ;
  assign n42183 = n41656 | n41805 ;
  assign n79088 = ~n42183 ;
  assign n42184 = n41801 & n79088 ;
  assign n42185 = n41966 | n42184 ;
  assign n42186 = n68710 & n42185 ;
  assign n42187 = n79028 & n42186 ;
  assign n42188 = n42182 | n42187 ;
  assign n42189 = n66145 & n42188 ;
  assign n42190 = n41655 & n41924 ;
  assign n79089 = ~n41796 ;
  assign n41800 = n79089 & n41799 ;
  assign n42191 = n41665 | n41799 ;
  assign n79090 = ~n42191 ;
  assign n42192 = n41960 & n79090 ;
  assign n42193 = n41800 | n42192 ;
  assign n42194 = n68710 & n42193 ;
  assign n42195 = n79028 & n42194 ;
  assign n42196 = n42190 | n42195 ;
  assign n42197 = n66081 & n42196 ;
  assign n79091 = ~n42195 ;
  assign n42347 = x76 & n79091 ;
  assign n79092 = ~n42190 ;
  assign n42348 = n79092 & n42347 ;
  assign n42349 = n42197 | n42348 ;
  assign n42198 = n41664 & n41924 ;
  assign n79093 = ~n41959 ;
  assign n41961 = n41794 & n79093 ;
  assign n42199 = n41674 | n41794 ;
  assign n79094 = ~n42199 ;
  assign n42200 = n41790 & n79094 ;
  assign n42201 = n41961 | n42200 ;
  assign n42202 = n68710 & n42201 ;
  assign n42203 = n79028 & n42202 ;
  assign n42204 = n42198 | n42203 ;
  assign n42205 = n66043 & n42204 ;
  assign n42206 = n41673 & n41924 ;
  assign n79095 = ~n41785 ;
  assign n41789 = n79095 & n41788 ;
  assign n42207 = n41683 | n41788 ;
  assign n79096 = ~n42207 ;
  assign n42208 = n41955 & n79096 ;
  assign n42209 = n41789 | n42208 ;
  assign n42210 = n68710 & n42209 ;
  assign n42211 = n79028 & n42210 ;
  assign n42212 = n42206 | n42211 ;
  assign n42213 = n65960 & n42212 ;
  assign n79097 = ~n42211 ;
  assign n42335 = x74 & n79097 ;
  assign n79098 = ~n42206 ;
  assign n42336 = n79098 & n42335 ;
  assign n42337 = n42213 | n42336 ;
  assign n42214 = n41682 & n41924 ;
  assign n79099 = ~n41954 ;
  assign n41956 = n41783 & n79099 ;
  assign n42215 = n41692 | n41783 ;
  assign n79100 = ~n42215 ;
  assign n42216 = n41779 & n79100 ;
  assign n42217 = n41956 | n42216 ;
  assign n42218 = n68710 & n42217 ;
  assign n42219 = n79028 & n42218 ;
  assign n42220 = n42214 | n42219 ;
  assign n42221 = n65909 & n42220 ;
  assign n42222 = n41691 & n41924 ;
  assign n79101 = ~n41773 ;
  assign n41777 = n79101 & n41776 ;
  assign n41778 = n41701 | n41776 ;
  assign n42223 = n41771 | n41949 ;
  assign n79102 = ~n41778 ;
  assign n42224 = n79102 & n42223 ;
  assign n42225 = n41777 | n42224 ;
  assign n42226 = n68710 & n42225 ;
  assign n42227 = n79028 & n42226 ;
  assign n42228 = n42222 | n42227 ;
  assign n42229 = n65877 & n42228 ;
  assign n79103 = ~n42227 ;
  assign n42323 = x72 & n79103 ;
  assign n79104 = ~n42222 ;
  assign n42324 = n79104 & n42323 ;
  assign n42325 = n42229 | n42324 ;
  assign n41927 = n41700 & n41924 ;
  assign n79105 = ~n41949 ;
  assign n41951 = n41771 & n79105 ;
  assign n42230 = n41764 | n41946 ;
  assign n42231 = n41710 | n41771 ;
  assign n79106 = ~n42231 ;
  assign n42232 = n42230 & n79106 ;
  assign n42233 = n41951 | n42232 ;
  assign n42234 = n68710 & n42233 ;
  assign n42235 = n79028 & n42234 ;
  assign n42236 = n41927 | n42235 ;
  assign n42237 = n65820 & n42236 ;
  assign n41926 = n41709 & n41924 ;
  assign n79107 = ~n41764 ;
  assign n41947 = n79107 & n41946 ;
  assign n42238 = n41762 | n41942 ;
  assign n42239 = n41719 | n41946 ;
  assign n79108 = ~n42239 ;
  assign n42240 = n42238 & n79108 ;
  assign n42241 = n41947 | n42240 ;
  assign n42242 = n68710 & n42241 ;
  assign n42243 = n79028 & n42242 ;
  assign n42244 = n41926 | n42243 ;
  assign n42245 = n65791 & n42244 ;
  assign n79109 = ~n42243 ;
  assign n42311 = x70 & n79109 ;
  assign n79110 = ~n41926 ;
  assign n42312 = n79110 & n42311 ;
  assign n42313 = n42245 | n42312 ;
  assign n41925 = n41718 & n41924 ;
  assign n79111 = ~n41942 ;
  assign n41944 = n41762 & n79111 ;
  assign n42246 = n41755 | n41939 ;
  assign n42247 = n41728 | n41762 ;
  assign n79112 = ~n42247 ;
  assign n42248 = n42246 & n79112 ;
  assign n42249 = n41944 | n42248 ;
  assign n42250 = n68710 & n42249 ;
  assign n42251 = n79028 & n42250 ;
  assign n42252 = n41925 | n42251 ;
  assign n42253 = n65772 & n42252 ;
  assign n41929 = n41727 & n41924 ;
  assign n79113 = ~n41755 ;
  assign n41940 = n79113 & n41939 ;
  assign n42254 = n41736 | n41939 ;
  assign n79114 = ~n42254 ;
  assign n42255 = n41754 & n79114 ;
  assign n42256 = n41940 | n42255 ;
  assign n42257 = n68710 & n42256 ;
  assign n42258 = n79028 & n42257 ;
  assign n42259 = n41929 | n42258 ;
  assign n42260 = n65746 & n42259 ;
  assign n79115 = ~n42258 ;
  assign n42301 = x68 & n79115 ;
  assign n79116 = ~n41929 ;
  assign n42302 = n79116 & n42301 ;
  assign n42303 = n42260 | n42302 ;
  assign n41931 = n41735 & n41924 ;
  assign n42261 = n41749 | n41753 ;
  assign n79117 = ~n42261 ;
  assign n42262 = n41935 & n79117 ;
  assign n79118 = ~n41936 ;
  assign n42263 = n41753 & n79118 ;
  assign n42264 = n42262 | n42263 ;
  assign n42265 = n68710 & n42264 ;
  assign n42266 = n79028 & n42265 ;
  assign n42267 = n41931 | n42266 ;
  assign n42268 = n65721 & n42267 ;
  assign n42269 = n41924 & n41932 ;
  assign n42270 = n9415 & n41746 ;
  assign n42271 = n78920 & n42270 ;
  assign n42272 = n9610 | n42271 ;
  assign n79119 = ~n42272 ;
  assign n42273 = n41935 & n79119 ;
  assign n42274 = n79028 & n42273 ;
  assign n42275 = n42269 | n42274 ;
  assign n42276 = n65686 & n42275 ;
  assign n79120 = ~n42274 ;
  assign n42291 = x66 & n79120 ;
  assign n79121 = ~n42269 ;
  assign n42292 = n79121 & n42291 ;
  assign n42293 = n42276 | n42292 ;
  assign n42277 = n79014 & n42016 ;
  assign n42278 = n41920 | n42277 ;
  assign n42279 = n79017 & n42278 ;
  assign n79122 = ~n42279 ;
  assign n42280 = n9950 & n79122 ;
  assign n79123 = ~n42280 ;
  assign n42281 = x30 & n79123 ;
  assign n42282 = n9956 & n79028 ;
  assign n42283 = n42281 | n42282 ;
  assign n42284 = x65 & n42283 ;
  assign n42285 = x65 | n42282 ;
  assign n42286 = n42281 | n42285 ;
  assign n79124 = ~n42284 ;
  assign n42287 = n79124 & n42286 ;
  assign n42289 = n9964 | n42287 ;
  assign n42290 = n65670 & n42283 ;
  assign n79125 = ~n42290 ;
  assign n42294 = n42289 & n79125 ;
  assign n42295 = n42293 | n42294 ;
  assign n79126 = ~n42276 ;
  assign n42296 = n79126 & n42295 ;
  assign n79127 = ~n42266 ;
  assign n42297 = x67 & n79127 ;
  assign n79128 = ~n41931 ;
  assign n42298 = n79128 & n42297 ;
  assign n42299 = n42268 | n42298 ;
  assign n42300 = n42296 | n42299 ;
  assign n79129 = ~n42268 ;
  assign n42304 = n79129 & n42300 ;
  assign n42305 = n42303 | n42304 ;
  assign n79130 = ~n42260 ;
  assign n42306 = n79130 & n42305 ;
  assign n79131 = ~n42251 ;
  assign n42307 = x69 & n79131 ;
  assign n79132 = ~n41925 ;
  assign n42308 = n79132 & n42307 ;
  assign n42309 = n42253 | n42308 ;
  assign n42310 = n42306 | n42309 ;
  assign n79133 = ~n42253 ;
  assign n42315 = n79133 & n42310 ;
  assign n42316 = n42313 | n42315 ;
  assign n79134 = ~n42245 ;
  assign n42317 = n79134 & n42316 ;
  assign n79135 = ~n42235 ;
  assign n42318 = x71 & n79135 ;
  assign n79136 = ~n41927 ;
  assign n42319 = n79136 & n42318 ;
  assign n42320 = n42237 | n42319 ;
  assign n42322 = n42317 | n42320 ;
  assign n79137 = ~n42237 ;
  assign n42327 = n79137 & n42322 ;
  assign n42328 = n42325 | n42327 ;
  assign n79138 = ~n42229 ;
  assign n42329 = n79138 & n42328 ;
  assign n79139 = ~n42219 ;
  assign n42330 = x73 & n79139 ;
  assign n79140 = ~n42214 ;
  assign n42331 = n79140 & n42330 ;
  assign n42332 = n42221 | n42331 ;
  assign n42334 = n42329 | n42332 ;
  assign n79141 = ~n42221 ;
  assign n42339 = n79141 & n42334 ;
  assign n42340 = n42337 | n42339 ;
  assign n79142 = ~n42213 ;
  assign n42341 = n79142 & n42340 ;
  assign n79143 = ~n42203 ;
  assign n42342 = x75 & n79143 ;
  assign n79144 = ~n42198 ;
  assign n42343 = n79144 & n42342 ;
  assign n42344 = n42205 | n42343 ;
  assign n42346 = n42341 | n42344 ;
  assign n79145 = ~n42205 ;
  assign n42351 = n79145 & n42346 ;
  assign n42352 = n42349 | n42351 ;
  assign n79146 = ~n42197 ;
  assign n42353 = n79146 & n42352 ;
  assign n79147 = ~n42187 ;
  assign n42354 = x77 & n79147 ;
  assign n79148 = ~n42182 ;
  assign n42355 = n79148 & n42354 ;
  assign n42356 = n42189 | n42355 ;
  assign n42358 = n42353 | n42356 ;
  assign n79149 = ~n42189 ;
  assign n42363 = n79149 & n42358 ;
  assign n42364 = n42361 | n42363 ;
  assign n79150 = ~n42181 ;
  assign n42365 = n79150 & n42364 ;
  assign n79151 = ~n42171 ;
  assign n42366 = x79 & n79151 ;
  assign n79152 = ~n42166 ;
  assign n42367 = n79152 & n42366 ;
  assign n42368 = n42173 | n42367 ;
  assign n42370 = n42365 | n42368 ;
  assign n79153 = ~n42173 ;
  assign n42375 = n79153 & n42370 ;
  assign n42376 = n42373 | n42375 ;
  assign n79154 = ~n42165 ;
  assign n42377 = n79154 & n42376 ;
  assign n79155 = ~n42155 ;
  assign n42378 = x81 & n79155 ;
  assign n79156 = ~n42150 ;
  assign n42379 = n79156 & n42378 ;
  assign n42380 = n42157 | n42379 ;
  assign n42382 = n42377 | n42380 ;
  assign n79157 = ~n42157 ;
  assign n42387 = n79157 & n42382 ;
  assign n42388 = n42385 | n42387 ;
  assign n79158 = ~n42149 ;
  assign n42389 = n79158 & n42388 ;
  assign n79159 = ~n42139 ;
  assign n42390 = x83 & n79159 ;
  assign n79160 = ~n42134 ;
  assign n42391 = n79160 & n42390 ;
  assign n42392 = n42141 | n42391 ;
  assign n42394 = n42389 | n42392 ;
  assign n79161 = ~n42141 ;
  assign n42399 = n79161 & n42394 ;
  assign n42400 = n42397 | n42399 ;
  assign n79162 = ~n42133 ;
  assign n42401 = n79162 & n42400 ;
  assign n79163 = ~n42123 ;
  assign n42402 = x85 & n79163 ;
  assign n79164 = ~n42118 ;
  assign n42403 = n79164 & n42402 ;
  assign n42404 = n42125 | n42403 ;
  assign n42406 = n42401 | n42404 ;
  assign n79165 = ~n42125 ;
  assign n42411 = n79165 & n42406 ;
  assign n42412 = n42409 | n42411 ;
  assign n79166 = ~n42117 ;
  assign n42413 = n79166 & n42412 ;
  assign n79167 = ~n42107 ;
  assign n42414 = x87 & n79167 ;
  assign n79168 = ~n42102 ;
  assign n42415 = n79168 & n42414 ;
  assign n42416 = n42109 | n42415 ;
  assign n42418 = n42413 | n42416 ;
  assign n79169 = ~n42109 ;
  assign n42423 = n79169 & n42418 ;
  assign n42424 = n42421 | n42423 ;
  assign n79170 = ~n42101 ;
  assign n42425 = n79170 & n42424 ;
  assign n79171 = ~n42091 ;
  assign n42426 = x89 & n79171 ;
  assign n79172 = ~n42086 ;
  assign n42427 = n79172 & n42426 ;
  assign n42428 = n42093 | n42427 ;
  assign n42430 = n42425 | n42428 ;
  assign n79173 = ~n42093 ;
  assign n42435 = n79173 & n42430 ;
  assign n42436 = n42433 | n42435 ;
  assign n79174 = ~n42085 ;
  assign n42437 = n79174 & n42436 ;
  assign n79175 = ~n42075 ;
  assign n42438 = x91 & n79175 ;
  assign n79176 = ~n42070 ;
  assign n42439 = n79176 & n42438 ;
  assign n42440 = n42077 | n42439 ;
  assign n42442 = n42437 | n42440 ;
  assign n79177 = ~n42077 ;
  assign n42447 = n79177 & n42442 ;
  assign n42448 = n42445 | n42447 ;
  assign n79178 = ~n42069 ;
  assign n42449 = n79178 & n42448 ;
  assign n79179 = ~n42059 ;
  assign n42450 = x93 & n79179 ;
  assign n79180 = ~n42054 ;
  assign n42451 = n79180 & n42450 ;
  assign n42452 = n42061 | n42451 ;
  assign n42454 = n42449 | n42452 ;
  assign n79181 = ~n42061 ;
  assign n42459 = n79181 & n42454 ;
  assign n42460 = n42457 | n42459 ;
  assign n79182 = ~n42053 ;
  assign n42461 = n79182 & n42460 ;
  assign n79183 = ~n42043 ;
  assign n42462 = x95 & n79183 ;
  assign n79184 = ~n42038 ;
  assign n42463 = n79184 & n42462 ;
  assign n42464 = n42045 | n42463 ;
  assign n42466 = n42461 | n42464 ;
  assign n79185 = ~n42045 ;
  assign n42471 = n79185 & n42466 ;
  assign n42472 = n42469 | n42471 ;
  assign n79186 = ~n42037 ;
  assign n42473 = n79186 & n42472 ;
  assign n79187 = ~n42021 ;
  assign n42474 = x97 & n79187 ;
  assign n79188 = ~n41930 ;
  assign n42475 = n79188 & n42474 ;
  assign n42476 = n42029 | n42475 ;
  assign n42478 = n42473 | n42476 ;
  assign n79189 = ~n42029 ;
  assign n42484 = n79189 & n42478 ;
  assign n42485 = n42483 | n42484 ;
  assign n79190 = ~n42028 ;
  assign n42486 = n79190 & n42485 ;
  assign n42487 = n10157 | n42486 ;
  assign n79191 = ~n42027 ;
  assign n42489 = n79191 & n42487 ;
  assign n79192 = ~n42484 ;
  assign n43022 = n42483 & n79192 ;
  assign n42491 = n9950 & n79028 ;
  assign n79193 = ~n42491 ;
  assign n42492 = x30 & n79193 ;
  assign n42493 = n42282 | n42492 ;
  assign n42494 = x65 & n42493 ;
  assign n79194 = ~n42494 ;
  assign n42495 = n42286 & n79194 ;
  assign n42496 = n9964 | n42495 ;
  assign n42497 = n79125 & n42496 ;
  assign n42498 = n42293 | n42497 ;
  assign n42499 = n79126 & n42498 ;
  assign n42500 = n42299 | n42499 ;
  assign n42501 = n79129 & n42500 ;
  assign n42502 = n42303 | n42501 ;
  assign n42503 = n79130 & n42502 ;
  assign n42504 = n42309 | n42503 ;
  assign n42505 = n79133 & n42504 ;
  assign n42506 = n42313 | n42505 ;
  assign n42507 = n79134 & n42506 ;
  assign n42508 = n42320 | n42507 ;
  assign n42509 = n79137 & n42508 ;
  assign n42510 = n42325 | n42509 ;
  assign n42511 = n79138 & n42510 ;
  assign n42512 = n42332 | n42511 ;
  assign n42513 = n79141 & n42512 ;
  assign n42514 = n42337 | n42513 ;
  assign n42515 = n79142 & n42514 ;
  assign n42516 = n42344 | n42515 ;
  assign n42517 = n79145 & n42516 ;
  assign n42518 = n42349 | n42517 ;
  assign n42519 = n79146 & n42518 ;
  assign n42520 = n42356 | n42519 ;
  assign n42521 = n79149 & n42520 ;
  assign n42522 = n42361 | n42521 ;
  assign n42523 = n79150 & n42522 ;
  assign n42524 = n42368 | n42523 ;
  assign n42525 = n79153 & n42524 ;
  assign n42526 = n42373 | n42525 ;
  assign n42527 = n79154 & n42526 ;
  assign n42528 = n42380 | n42527 ;
  assign n42529 = n79157 & n42528 ;
  assign n42530 = n42385 | n42529 ;
  assign n42531 = n79158 & n42530 ;
  assign n42532 = n42392 | n42531 ;
  assign n42533 = n79161 & n42532 ;
  assign n42534 = n42397 | n42533 ;
  assign n42535 = n79162 & n42534 ;
  assign n42536 = n42404 | n42535 ;
  assign n42537 = n79165 & n42536 ;
  assign n42538 = n42409 | n42537 ;
  assign n42539 = n79166 & n42538 ;
  assign n42540 = n42416 | n42539 ;
  assign n42541 = n79169 & n42540 ;
  assign n42542 = n42421 | n42541 ;
  assign n42543 = n79170 & n42542 ;
  assign n42544 = n42428 | n42543 ;
  assign n42545 = n79173 & n42544 ;
  assign n42546 = n42433 | n42545 ;
  assign n42547 = n79174 & n42546 ;
  assign n42548 = n42440 | n42547 ;
  assign n42549 = n79177 & n42548 ;
  assign n42550 = n42445 | n42549 ;
  assign n42551 = n79178 & n42550 ;
  assign n42552 = n42452 | n42551 ;
  assign n42553 = n79181 & n42552 ;
  assign n42554 = n42457 | n42553 ;
  assign n42555 = n79182 & n42554 ;
  assign n42556 = n42464 | n42555 ;
  assign n42557 = n79185 & n42556 ;
  assign n42558 = n42469 | n42557 ;
  assign n42560 = n79186 & n42558 ;
  assign n42826 = n42476 | n42560 ;
  assign n43023 = n42029 | n42483 ;
  assign n79195 = ~n43023 ;
  assign n43024 = n42826 & n79195 ;
  assign n43025 = n43022 | n43024 ;
  assign n43026 = n42487 | n43025 ;
  assign n79196 = ~n42489 ;
  assign n43027 = n79196 & n43026 ;
  assign n43035 = n68894 & n43027 ;
  assign n42490 = n42022 & n42487 ;
  assign n42477 = n42037 | n42476 ;
  assign n79197 = ~n42477 ;
  assign n42559 = n79197 & n42558 ;
  assign n79198 = ~n42560 ;
  assign n42561 = n42476 & n79198 ;
  assign n42562 = n42559 | n42561 ;
  assign n42563 = n68894 & n42562 ;
  assign n79199 = ~n42486 ;
  assign n42564 = n79199 & n42563 ;
  assign n42565 = n42490 | n42564 ;
  assign n42566 = n68716 & n42565 ;
  assign n42567 = n42036 & n42487 ;
  assign n42470 = n42045 | n42469 ;
  assign n79200 = ~n42470 ;
  assign n42568 = n42466 & n79200 ;
  assign n79201 = ~n42471 ;
  assign n42569 = n42469 & n79201 ;
  assign n42570 = n42568 | n42569 ;
  assign n42571 = n68894 & n42570 ;
  assign n42572 = n79199 & n42571 ;
  assign n42573 = n42567 | n42572 ;
  assign n42574 = n68545 & n42573 ;
  assign n42575 = n42044 & n42487 ;
  assign n42465 = n42053 | n42464 ;
  assign n79202 = ~n42465 ;
  assign n42576 = n79202 & n42554 ;
  assign n79203 = ~n42555 ;
  assign n42577 = n42464 & n79203 ;
  assign n42578 = n42576 | n42577 ;
  assign n42579 = n68894 & n42578 ;
  assign n42580 = n79199 & n42579 ;
  assign n42581 = n42575 | n42580 ;
  assign n42582 = n68438 & n42581 ;
  assign n42583 = n42052 & n42487 ;
  assign n42458 = n42061 | n42457 ;
  assign n79204 = ~n42458 ;
  assign n42584 = n42454 & n79204 ;
  assign n79205 = ~n42459 ;
  assign n42585 = n42457 & n79205 ;
  assign n42586 = n42584 | n42585 ;
  assign n42587 = n68894 & n42586 ;
  assign n42588 = n79199 & n42587 ;
  assign n42589 = n42583 | n42588 ;
  assign n42590 = n68214 & n42589 ;
  assign n42591 = n42060 & n42487 ;
  assign n42453 = n42069 | n42452 ;
  assign n79206 = ~n42453 ;
  assign n42592 = n79206 & n42550 ;
  assign n79207 = ~n42551 ;
  assign n42593 = n42452 & n79207 ;
  assign n42594 = n42592 | n42593 ;
  assign n42595 = n68894 & n42594 ;
  assign n42596 = n79199 & n42595 ;
  assign n42597 = n42591 | n42596 ;
  assign n42598 = n68058 & n42597 ;
  assign n42599 = n42068 & n42487 ;
  assign n42446 = n42077 | n42445 ;
  assign n79208 = ~n42446 ;
  assign n42600 = n42442 & n79208 ;
  assign n79209 = ~n42447 ;
  assign n42601 = n42445 & n79209 ;
  assign n42602 = n42600 | n42601 ;
  assign n42603 = n68894 & n42602 ;
  assign n42604 = n79199 & n42603 ;
  assign n42605 = n42599 | n42604 ;
  assign n42606 = n67986 & n42605 ;
  assign n42607 = n42076 & n42487 ;
  assign n42441 = n42085 | n42440 ;
  assign n79210 = ~n42441 ;
  assign n42608 = n79210 & n42546 ;
  assign n79211 = ~n42547 ;
  assign n42609 = n42440 & n79211 ;
  assign n42610 = n42608 | n42609 ;
  assign n42611 = n68894 & n42610 ;
  assign n42612 = n79199 & n42611 ;
  assign n42613 = n42607 | n42612 ;
  assign n42614 = n67763 & n42613 ;
  assign n42615 = n42084 & n42487 ;
  assign n42434 = n42093 | n42433 ;
  assign n79212 = ~n42434 ;
  assign n42616 = n42430 & n79212 ;
  assign n79213 = ~n42435 ;
  assign n42617 = n42433 & n79213 ;
  assign n42618 = n42616 | n42617 ;
  assign n42619 = n68894 & n42618 ;
  assign n42620 = n79199 & n42619 ;
  assign n42621 = n42615 | n42620 ;
  assign n42622 = n67622 & n42621 ;
  assign n42623 = n42092 & n42487 ;
  assign n42429 = n42101 | n42428 ;
  assign n79214 = ~n42429 ;
  assign n42624 = n79214 & n42542 ;
  assign n79215 = ~n42543 ;
  assign n42625 = n42428 & n79215 ;
  assign n42626 = n42624 | n42625 ;
  assign n42627 = n68894 & n42626 ;
  assign n42628 = n79199 & n42627 ;
  assign n42629 = n42623 | n42628 ;
  assign n42630 = n67531 & n42629 ;
  assign n42631 = n42100 & n42487 ;
  assign n42422 = n42109 | n42421 ;
  assign n79216 = ~n42422 ;
  assign n42632 = n42418 & n79216 ;
  assign n79217 = ~n42423 ;
  assign n42633 = n42421 & n79217 ;
  assign n42634 = n42632 | n42633 ;
  assign n42635 = n68894 & n42634 ;
  assign n42636 = n79199 & n42635 ;
  assign n42637 = n42631 | n42636 ;
  assign n42638 = n67348 & n42637 ;
  assign n42639 = n42108 & n42487 ;
  assign n42417 = n42117 | n42416 ;
  assign n79218 = ~n42417 ;
  assign n42640 = n79218 & n42538 ;
  assign n79219 = ~n42539 ;
  assign n42641 = n42416 & n79219 ;
  assign n42642 = n42640 | n42641 ;
  assign n42643 = n68894 & n42642 ;
  assign n42644 = n79199 & n42643 ;
  assign n42645 = n42639 | n42644 ;
  assign n42646 = n67222 & n42645 ;
  assign n42647 = n42116 & n42487 ;
  assign n42410 = n42125 | n42409 ;
  assign n79220 = ~n42410 ;
  assign n42648 = n42406 & n79220 ;
  assign n79221 = ~n42411 ;
  assign n42649 = n42409 & n79221 ;
  assign n42650 = n42648 | n42649 ;
  assign n42651 = n68894 & n42650 ;
  assign n42652 = n79199 & n42651 ;
  assign n42653 = n42647 | n42652 ;
  assign n42654 = n67164 & n42653 ;
  assign n42655 = n42124 & n42487 ;
  assign n42405 = n42133 | n42404 ;
  assign n79222 = ~n42405 ;
  assign n42656 = n79222 & n42534 ;
  assign n79223 = ~n42535 ;
  assign n42657 = n42404 & n79223 ;
  assign n42658 = n42656 | n42657 ;
  assign n42659 = n68894 & n42658 ;
  assign n42660 = n79199 & n42659 ;
  assign n42661 = n42655 | n42660 ;
  assign n42662 = n66979 & n42661 ;
  assign n42663 = n42132 & n42487 ;
  assign n42398 = n42141 | n42397 ;
  assign n79224 = ~n42398 ;
  assign n42664 = n42394 & n79224 ;
  assign n79225 = ~n42399 ;
  assign n42665 = n42397 & n79225 ;
  assign n42666 = n42664 | n42665 ;
  assign n42667 = n68894 & n42666 ;
  assign n42668 = n79199 & n42667 ;
  assign n42669 = n42663 | n42668 ;
  assign n42670 = n66868 & n42669 ;
  assign n42671 = n42140 & n42487 ;
  assign n42393 = n42149 | n42392 ;
  assign n79226 = ~n42393 ;
  assign n42672 = n79226 & n42530 ;
  assign n79227 = ~n42531 ;
  assign n42673 = n42392 & n79227 ;
  assign n42674 = n42672 | n42673 ;
  assign n42675 = n68894 & n42674 ;
  assign n42676 = n79199 & n42675 ;
  assign n42677 = n42671 | n42676 ;
  assign n42678 = n66797 & n42677 ;
  assign n42679 = n42148 & n42487 ;
  assign n42386 = n42157 | n42385 ;
  assign n79228 = ~n42386 ;
  assign n42680 = n42382 & n79228 ;
  assign n79229 = ~n42387 ;
  assign n42681 = n42385 & n79229 ;
  assign n42682 = n42680 | n42681 ;
  assign n42683 = n68894 & n42682 ;
  assign n42684 = n79199 & n42683 ;
  assign n42685 = n42679 | n42684 ;
  assign n42686 = n66654 & n42685 ;
  assign n42687 = n42156 & n42487 ;
  assign n42381 = n42165 | n42380 ;
  assign n79230 = ~n42381 ;
  assign n42688 = n79230 & n42526 ;
  assign n79231 = ~n42527 ;
  assign n42689 = n42380 & n79231 ;
  assign n42690 = n42688 | n42689 ;
  assign n42691 = n68894 & n42690 ;
  assign n42692 = n79199 & n42691 ;
  assign n42693 = n42687 | n42692 ;
  assign n42694 = n66560 & n42693 ;
  assign n42695 = n42164 & n42487 ;
  assign n42374 = n42173 | n42373 ;
  assign n79232 = ~n42374 ;
  assign n42696 = n42370 & n79232 ;
  assign n79233 = ~n42375 ;
  assign n42697 = n42373 & n79233 ;
  assign n42698 = n42696 | n42697 ;
  assign n42699 = n68894 & n42698 ;
  assign n42700 = n79199 & n42699 ;
  assign n42701 = n42695 | n42700 ;
  assign n42702 = n66505 & n42701 ;
  assign n42703 = n42172 & n42487 ;
  assign n42369 = n42181 | n42368 ;
  assign n79234 = ~n42369 ;
  assign n42704 = n79234 & n42522 ;
  assign n79235 = ~n42523 ;
  assign n42705 = n42368 & n79235 ;
  assign n42706 = n42704 | n42705 ;
  assign n42707 = n68894 & n42706 ;
  assign n42708 = n79199 & n42707 ;
  assign n42709 = n42703 | n42708 ;
  assign n42710 = n66379 & n42709 ;
  assign n42711 = n42180 & n42487 ;
  assign n42362 = n42189 | n42361 ;
  assign n79236 = ~n42362 ;
  assign n42712 = n42358 & n79236 ;
  assign n79237 = ~n42363 ;
  assign n42713 = n42361 & n79237 ;
  assign n42714 = n42712 | n42713 ;
  assign n42715 = n68894 & n42714 ;
  assign n42716 = n79199 & n42715 ;
  assign n42717 = n42711 | n42716 ;
  assign n42718 = n66299 & n42717 ;
  assign n42719 = n42188 & n42487 ;
  assign n42357 = n42197 | n42356 ;
  assign n79238 = ~n42357 ;
  assign n42720 = n79238 & n42518 ;
  assign n79239 = ~n42519 ;
  assign n42721 = n42356 & n79239 ;
  assign n42722 = n42720 | n42721 ;
  assign n42723 = n68894 & n42722 ;
  assign n42724 = n79199 & n42723 ;
  assign n42725 = n42719 | n42724 ;
  assign n42726 = n66244 & n42725 ;
  assign n42727 = n42196 & n42487 ;
  assign n42350 = n42205 | n42349 ;
  assign n79240 = ~n42350 ;
  assign n42728 = n42346 & n79240 ;
  assign n79241 = ~n42351 ;
  assign n42729 = n42349 & n79241 ;
  assign n42730 = n42728 | n42729 ;
  assign n42731 = n68894 & n42730 ;
  assign n42732 = n79199 & n42731 ;
  assign n42733 = n42727 | n42732 ;
  assign n42734 = n66145 & n42733 ;
  assign n42735 = n42204 & n42487 ;
  assign n42345 = n42213 | n42344 ;
  assign n79242 = ~n42345 ;
  assign n42736 = n79242 & n42514 ;
  assign n79243 = ~n42515 ;
  assign n42737 = n42344 & n79243 ;
  assign n42738 = n42736 | n42737 ;
  assign n42739 = n68894 & n42738 ;
  assign n42740 = n79199 & n42739 ;
  assign n42741 = n42735 | n42740 ;
  assign n42742 = n66081 & n42741 ;
  assign n42743 = n42212 & n42487 ;
  assign n42338 = n42221 | n42337 ;
  assign n79244 = ~n42338 ;
  assign n42744 = n42334 & n79244 ;
  assign n79245 = ~n42339 ;
  assign n42745 = n42337 & n79245 ;
  assign n42746 = n42744 | n42745 ;
  assign n42747 = n68894 & n42746 ;
  assign n42748 = n79199 & n42747 ;
  assign n42749 = n42743 | n42748 ;
  assign n42750 = n66043 & n42749 ;
  assign n42751 = n42220 & n42487 ;
  assign n42333 = n42229 | n42332 ;
  assign n79246 = ~n42333 ;
  assign n42752 = n79246 & n42510 ;
  assign n79247 = ~n42511 ;
  assign n42753 = n42332 & n79247 ;
  assign n42754 = n42752 | n42753 ;
  assign n42755 = n68894 & n42754 ;
  assign n42756 = n79199 & n42755 ;
  assign n42757 = n42751 | n42756 ;
  assign n42758 = n65960 & n42757 ;
  assign n42759 = n42228 & n42487 ;
  assign n42326 = n42237 | n42325 ;
  assign n79248 = ~n42326 ;
  assign n42760 = n42322 & n79248 ;
  assign n79249 = ~n42327 ;
  assign n42761 = n42325 & n79249 ;
  assign n42762 = n42760 | n42761 ;
  assign n42763 = n68894 & n42762 ;
  assign n42764 = n79199 & n42763 ;
  assign n42765 = n42759 | n42764 ;
  assign n42766 = n65909 & n42765 ;
  assign n42767 = n42236 & n42487 ;
  assign n42321 = n42245 | n42320 ;
  assign n79250 = ~n42321 ;
  assign n42768 = n79250 & n42506 ;
  assign n79251 = ~n42507 ;
  assign n42769 = n42320 & n79251 ;
  assign n42770 = n42768 | n42769 ;
  assign n42771 = n68894 & n42770 ;
  assign n42772 = n79199 & n42771 ;
  assign n42773 = n42767 | n42772 ;
  assign n42774 = n65877 & n42773 ;
  assign n42775 = n42244 & n42487 ;
  assign n42314 = n42253 | n42313 ;
  assign n79252 = ~n42314 ;
  assign n42776 = n79252 & n42504 ;
  assign n79253 = ~n42315 ;
  assign n42777 = n42313 & n79253 ;
  assign n42778 = n42776 | n42777 ;
  assign n42779 = n68894 & n42778 ;
  assign n42780 = n79199 & n42779 ;
  assign n42781 = n42775 | n42780 ;
  assign n42782 = n65820 & n42781 ;
  assign n42783 = n42252 & n42487 ;
  assign n42784 = n42260 | n42309 ;
  assign n79254 = ~n42784 ;
  assign n42785 = n42502 & n79254 ;
  assign n79255 = ~n42503 ;
  assign n42786 = n42309 & n79255 ;
  assign n42787 = n42785 | n42786 ;
  assign n42788 = n68894 & n42787 ;
  assign n42789 = n79199 & n42788 ;
  assign n42790 = n42783 | n42789 ;
  assign n42791 = n65791 & n42790 ;
  assign n42792 = n42259 & n42487 ;
  assign n42793 = n42268 | n42303 ;
  assign n79256 = ~n42793 ;
  assign n42794 = n42500 & n79256 ;
  assign n79257 = ~n42304 ;
  assign n42795 = n42303 & n79257 ;
  assign n42796 = n42794 | n42795 ;
  assign n42797 = n68894 & n42796 ;
  assign n42798 = n79199 & n42797 ;
  assign n42799 = n42792 | n42798 ;
  assign n42800 = n65772 & n42799 ;
  assign n42801 = n42267 & n42487 ;
  assign n42802 = n42276 | n42299 ;
  assign n79258 = ~n42802 ;
  assign n42803 = n42498 & n79258 ;
  assign n79259 = ~n42499 ;
  assign n42804 = n42299 & n79259 ;
  assign n42805 = n42803 | n42804 ;
  assign n42806 = n68894 & n42805 ;
  assign n42807 = n79199 & n42806 ;
  assign n42808 = n42801 | n42807 ;
  assign n42809 = n65746 & n42808 ;
  assign n42810 = n42275 & n42487 ;
  assign n79260 = ~n42497 ;
  assign n42811 = n42293 & n79260 ;
  assign n42812 = n42290 | n42293 ;
  assign n79261 = ~n42812 ;
  assign n42813 = n42496 & n79261 ;
  assign n42814 = n42811 | n42813 ;
  assign n42815 = n68894 & n42814 ;
  assign n42816 = n79199 & n42815 ;
  assign n42817 = n42810 | n42816 ;
  assign n42818 = n65721 & n42817 ;
  assign n42488 = n42283 & n42487 ;
  assign n42288 = n9964 & n42286 ;
  assign n42819 = n42288 & n79194 ;
  assign n42820 = n10157 | n42819 ;
  assign n79262 = ~n42820 ;
  assign n42821 = n42496 & n79262 ;
  assign n42822 = n79199 & n42821 ;
  assign n42823 = n42488 | n42822 ;
  assign n42824 = n65686 & n42823 ;
  assign n42825 = n10522 & n79199 ;
  assign n42827 = n79189 & n42826 ;
  assign n42828 = n42483 | n42827 ;
  assign n42829 = n79190 & n42828 ;
  assign n79263 = ~n42829 ;
  assign n42830 = n10516 & n79263 ;
  assign n79264 = ~n42830 ;
  assign n42831 = x29 & n79264 ;
  assign n42832 = n42825 | n42831 ;
  assign n42840 = n65670 & n42832 ;
  assign n42833 = n10516 & n79199 ;
  assign n79265 = ~n42833 ;
  assign n42834 = x29 & n79265 ;
  assign n42835 = n42825 | n42834 ;
  assign n42836 = x65 & n42835 ;
  assign n42837 = x65 | n42825 ;
  assign n42838 = n42834 | n42837 ;
  assign n79266 = ~n42836 ;
  assign n42839 = n79266 & n42838 ;
  assign n42841 = n10529 | n42839 ;
  assign n79267 = ~n42840 ;
  assign n42842 = n79267 & n42841 ;
  assign n79268 = ~n42822 ;
  assign n42843 = x66 & n79268 ;
  assign n79269 = ~n42488 ;
  assign n42844 = n79269 & n42843 ;
  assign n42845 = n42842 | n42844 ;
  assign n79270 = ~n42824 ;
  assign n42846 = n79270 & n42845 ;
  assign n79271 = ~n42816 ;
  assign n42847 = x67 & n79271 ;
  assign n79272 = ~n42810 ;
  assign n42848 = n79272 & n42847 ;
  assign n42849 = n42818 | n42848 ;
  assign n42850 = n42846 | n42849 ;
  assign n79273 = ~n42818 ;
  assign n42851 = n79273 & n42850 ;
  assign n79274 = ~n42807 ;
  assign n42852 = x68 & n79274 ;
  assign n79275 = ~n42801 ;
  assign n42853 = n79275 & n42852 ;
  assign n42854 = n42809 | n42853 ;
  assign n42855 = n42851 | n42854 ;
  assign n79276 = ~n42809 ;
  assign n42856 = n79276 & n42855 ;
  assign n79277 = ~n42798 ;
  assign n42857 = x69 & n79277 ;
  assign n79278 = ~n42792 ;
  assign n42858 = n79278 & n42857 ;
  assign n42859 = n42800 | n42858 ;
  assign n42860 = n42856 | n42859 ;
  assign n79279 = ~n42800 ;
  assign n42861 = n79279 & n42860 ;
  assign n79280 = ~n42789 ;
  assign n42862 = x70 & n79280 ;
  assign n79281 = ~n42783 ;
  assign n42863 = n79281 & n42862 ;
  assign n42864 = n42791 | n42863 ;
  assign n42866 = n42861 | n42864 ;
  assign n79282 = ~n42791 ;
  assign n42867 = n79282 & n42866 ;
  assign n79283 = ~n42780 ;
  assign n42868 = x71 & n79283 ;
  assign n79284 = ~n42775 ;
  assign n42869 = n79284 & n42868 ;
  assign n42870 = n42782 | n42869 ;
  assign n42871 = n42867 | n42870 ;
  assign n79285 = ~n42782 ;
  assign n42872 = n79285 & n42871 ;
  assign n79286 = ~n42772 ;
  assign n42873 = x72 & n79286 ;
  assign n79287 = ~n42767 ;
  assign n42874 = n79287 & n42873 ;
  assign n42875 = n42774 | n42874 ;
  assign n42877 = n42872 | n42875 ;
  assign n79288 = ~n42774 ;
  assign n42878 = n79288 & n42877 ;
  assign n79289 = ~n42764 ;
  assign n42879 = x73 & n79289 ;
  assign n79290 = ~n42759 ;
  assign n42880 = n79290 & n42879 ;
  assign n42881 = n42766 | n42880 ;
  assign n42882 = n42878 | n42881 ;
  assign n79291 = ~n42766 ;
  assign n42883 = n79291 & n42882 ;
  assign n79292 = ~n42756 ;
  assign n42884 = x74 & n79292 ;
  assign n79293 = ~n42751 ;
  assign n42885 = n79293 & n42884 ;
  assign n42886 = n42758 | n42885 ;
  assign n42888 = n42883 | n42886 ;
  assign n79294 = ~n42758 ;
  assign n42889 = n79294 & n42888 ;
  assign n79295 = ~n42748 ;
  assign n42890 = x75 & n79295 ;
  assign n79296 = ~n42743 ;
  assign n42891 = n79296 & n42890 ;
  assign n42892 = n42750 | n42891 ;
  assign n42893 = n42889 | n42892 ;
  assign n79297 = ~n42750 ;
  assign n42894 = n79297 & n42893 ;
  assign n79298 = ~n42740 ;
  assign n42895 = x76 & n79298 ;
  assign n79299 = ~n42735 ;
  assign n42896 = n79299 & n42895 ;
  assign n42897 = n42742 | n42896 ;
  assign n42899 = n42894 | n42897 ;
  assign n79300 = ~n42742 ;
  assign n42900 = n79300 & n42899 ;
  assign n79301 = ~n42732 ;
  assign n42901 = x77 & n79301 ;
  assign n79302 = ~n42727 ;
  assign n42902 = n79302 & n42901 ;
  assign n42903 = n42734 | n42902 ;
  assign n42904 = n42900 | n42903 ;
  assign n79303 = ~n42734 ;
  assign n42905 = n79303 & n42904 ;
  assign n79304 = ~n42724 ;
  assign n42906 = x78 & n79304 ;
  assign n79305 = ~n42719 ;
  assign n42907 = n79305 & n42906 ;
  assign n42908 = n42726 | n42907 ;
  assign n42910 = n42905 | n42908 ;
  assign n79306 = ~n42726 ;
  assign n42911 = n79306 & n42910 ;
  assign n79307 = ~n42716 ;
  assign n42912 = x79 & n79307 ;
  assign n79308 = ~n42711 ;
  assign n42913 = n79308 & n42912 ;
  assign n42914 = n42718 | n42913 ;
  assign n42915 = n42911 | n42914 ;
  assign n79309 = ~n42718 ;
  assign n42916 = n79309 & n42915 ;
  assign n79310 = ~n42708 ;
  assign n42917 = x80 & n79310 ;
  assign n79311 = ~n42703 ;
  assign n42918 = n79311 & n42917 ;
  assign n42919 = n42710 | n42918 ;
  assign n42921 = n42916 | n42919 ;
  assign n79312 = ~n42710 ;
  assign n42922 = n79312 & n42921 ;
  assign n79313 = ~n42700 ;
  assign n42923 = x81 & n79313 ;
  assign n79314 = ~n42695 ;
  assign n42924 = n79314 & n42923 ;
  assign n42925 = n42702 | n42924 ;
  assign n42926 = n42922 | n42925 ;
  assign n79315 = ~n42702 ;
  assign n42927 = n79315 & n42926 ;
  assign n79316 = ~n42692 ;
  assign n42928 = x82 & n79316 ;
  assign n79317 = ~n42687 ;
  assign n42929 = n79317 & n42928 ;
  assign n42930 = n42694 | n42929 ;
  assign n42932 = n42927 | n42930 ;
  assign n79318 = ~n42694 ;
  assign n42933 = n79318 & n42932 ;
  assign n79319 = ~n42684 ;
  assign n42934 = x83 & n79319 ;
  assign n79320 = ~n42679 ;
  assign n42935 = n79320 & n42934 ;
  assign n42936 = n42686 | n42935 ;
  assign n42937 = n42933 | n42936 ;
  assign n79321 = ~n42686 ;
  assign n42938 = n79321 & n42937 ;
  assign n79322 = ~n42676 ;
  assign n42939 = x84 & n79322 ;
  assign n79323 = ~n42671 ;
  assign n42940 = n79323 & n42939 ;
  assign n42941 = n42678 | n42940 ;
  assign n42943 = n42938 | n42941 ;
  assign n79324 = ~n42678 ;
  assign n42944 = n79324 & n42943 ;
  assign n79325 = ~n42668 ;
  assign n42945 = x85 & n79325 ;
  assign n79326 = ~n42663 ;
  assign n42946 = n79326 & n42945 ;
  assign n42947 = n42670 | n42946 ;
  assign n42948 = n42944 | n42947 ;
  assign n79327 = ~n42670 ;
  assign n42949 = n79327 & n42948 ;
  assign n79328 = ~n42660 ;
  assign n42950 = x86 & n79328 ;
  assign n79329 = ~n42655 ;
  assign n42951 = n79329 & n42950 ;
  assign n42952 = n42662 | n42951 ;
  assign n42954 = n42949 | n42952 ;
  assign n79330 = ~n42662 ;
  assign n42955 = n79330 & n42954 ;
  assign n79331 = ~n42652 ;
  assign n42956 = x87 & n79331 ;
  assign n79332 = ~n42647 ;
  assign n42957 = n79332 & n42956 ;
  assign n42958 = n42654 | n42957 ;
  assign n42959 = n42955 | n42958 ;
  assign n79333 = ~n42654 ;
  assign n42960 = n79333 & n42959 ;
  assign n79334 = ~n42644 ;
  assign n42961 = x88 & n79334 ;
  assign n79335 = ~n42639 ;
  assign n42962 = n79335 & n42961 ;
  assign n42963 = n42646 | n42962 ;
  assign n42965 = n42960 | n42963 ;
  assign n79336 = ~n42646 ;
  assign n42966 = n79336 & n42965 ;
  assign n79337 = ~n42636 ;
  assign n42967 = x89 & n79337 ;
  assign n79338 = ~n42631 ;
  assign n42968 = n79338 & n42967 ;
  assign n42969 = n42638 | n42968 ;
  assign n42970 = n42966 | n42969 ;
  assign n79339 = ~n42638 ;
  assign n42971 = n79339 & n42970 ;
  assign n79340 = ~n42628 ;
  assign n42972 = x90 & n79340 ;
  assign n79341 = ~n42623 ;
  assign n42973 = n79341 & n42972 ;
  assign n42974 = n42630 | n42973 ;
  assign n42976 = n42971 | n42974 ;
  assign n79342 = ~n42630 ;
  assign n42977 = n79342 & n42976 ;
  assign n79343 = ~n42620 ;
  assign n42978 = x91 & n79343 ;
  assign n79344 = ~n42615 ;
  assign n42979 = n79344 & n42978 ;
  assign n42980 = n42622 | n42979 ;
  assign n42981 = n42977 | n42980 ;
  assign n79345 = ~n42622 ;
  assign n42982 = n79345 & n42981 ;
  assign n79346 = ~n42612 ;
  assign n42983 = x92 & n79346 ;
  assign n79347 = ~n42607 ;
  assign n42984 = n79347 & n42983 ;
  assign n42985 = n42614 | n42984 ;
  assign n42987 = n42982 | n42985 ;
  assign n79348 = ~n42614 ;
  assign n42988 = n79348 & n42987 ;
  assign n79349 = ~n42604 ;
  assign n42989 = x93 & n79349 ;
  assign n79350 = ~n42599 ;
  assign n42990 = n79350 & n42989 ;
  assign n42991 = n42606 | n42990 ;
  assign n42992 = n42988 | n42991 ;
  assign n79351 = ~n42606 ;
  assign n42993 = n79351 & n42992 ;
  assign n79352 = ~n42596 ;
  assign n42994 = x94 & n79352 ;
  assign n79353 = ~n42591 ;
  assign n42995 = n79353 & n42994 ;
  assign n42996 = n42598 | n42995 ;
  assign n42998 = n42993 | n42996 ;
  assign n79354 = ~n42598 ;
  assign n42999 = n79354 & n42998 ;
  assign n79355 = ~n42588 ;
  assign n43000 = x95 & n79355 ;
  assign n79356 = ~n42583 ;
  assign n43001 = n79356 & n43000 ;
  assign n43002 = n42590 | n43001 ;
  assign n43003 = n42999 | n43002 ;
  assign n79357 = ~n42590 ;
  assign n43004 = n79357 & n43003 ;
  assign n79358 = ~n42580 ;
  assign n43005 = x96 & n79358 ;
  assign n79359 = ~n42575 ;
  assign n43006 = n79359 & n43005 ;
  assign n43007 = n42582 | n43006 ;
  assign n43009 = n43004 | n43007 ;
  assign n79360 = ~n42582 ;
  assign n43010 = n79360 & n43009 ;
  assign n79361 = ~n42572 ;
  assign n43011 = x97 & n79361 ;
  assign n79362 = ~n42567 ;
  assign n43012 = n79362 & n43011 ;
  assign n43013 = n42574 | n43012 ;
  assign n43014 = n43010 | n43013 ;
  assign n79363 = ~n42574 ;
  assign n43015 = n79363 & n43014 ;
  assign n79364 = ~n42564 ;
  assign n43016 = x98 & n79364 ;
  assign n79365 = ~n42490 ;
  assign n43017 = n79365 & n43016 ;
  assign n43018 = n42566 | n43017 ;
  assign n43020 = n43015 | n43018 ;
  assign n79366 = ~n42566 ;
  assign n43021 = n79366 & n43020 ;
  assign n43028 = n68993 & n43027 ;
  assign n79367 = ~n42487 ;
  assign n43029 = n79367 & n43025 ;
  assign n43030 = n42027 & n42487 ;
  assign n79368 = ~n43030 ;
  assign n43031 = x99 & n79368 ;
  assign n79369 = ~n43029 ;
  assign n43032 = n79369 & n43031 ;
  assign n43033 = n380 | n43032 ;
  assign n43034 = n43028 | n43033 ;
  assign n43036 = n43021 | n43034 ;
  assign n79370 = ~n43035 ;
  assign n43037 = n79370 & n43036 ;
  assign n79371 = ~n43015 ;
  assign n43019 = n79371 & n43018 ;
  assign n43040 = x65 & n42832 ;
  assign n79372 = ~n43040 ;
  assign n43041 = n42838 & n79372 ;
  assign n43042 = n10529 | n43041 ;
  assign n43043 = n79267 & n43042 ;
  assign n43044 = n42824 | n42844 ;
  assign n43046 = n43043 | n43044 ;
  assign n43047 = n79270 & n43046 ;
  assign n43048 = n42848 | n43047 ;
  assign n43050 = n79273 & n43048 ;
  assign n43052 = n42854 | n43050 ;
  assign n43053 = n79276 & n43052 ;
  assign n43055 = n42859 | n43053 ;
  assign n43056 = n79279 & n43055 ;
  assign n43057 = n42864 | n43056 ;
  assign n43058 = n79282 & n43057 ;
  assign n43059 = n42870 | n43058 ;
  assign n43061 = n79285 & n43059 ;
  assign n43062 = n42875 | n43061 ;
  assign n43063 = n79288 & n43062 ;
  assign n43064 = n42881 | n43063 ;
  assign n43066 = n79291 & n43064 ;
  assign n43067 = n42886 | n43066 ;
  assign n43068 = n79294 & n43067 ;
  assign n43069 = n42892 | n43068 ;
  assign n43071 = n79297 & n43069 ;
  assign n43072 = n42897 | n43071 ;
  assign n43073 = n79300 & n43072 ;
  assign n43074 = n42903 | n43073 ;
  assign n43076 = n79303 & n43074 ;
  assign n43077 = n42908 | n43076 ;
  assign n43078 = n79306 & n43077 ;
  assign n43079 = n42914 | n43078 ;
  assign n43081 = n79309 & n43079 ;
  assign n43082 = n42919 | n43081 ;
  assign n43083 = n79312 & n43082 ;
  assign n43084 = n42925 | n43083 ;
  assign n43086 = n79315 & n43084 ;
  assign n43087 = n42930 | n43086 ;
  assign n43088 = n79318 & n43087 ;
  assign n43089 = n42936 | n43088 ;
  assign n43091 = n79321 & n43089 ;
  assign n43092 = n42941 | n43091 ;
  assign n43093 = n79324 & n43092 ;
  assign n43094 = n42947 | n43093 ;
  assign n43096 = n79327 & n43094 ;
  assign n43097 = n42952 | n43096 ;
  assign n43098 = n79330 & n43097 ;
  assign n43099 = n42958 | n43098 ;
  assign n43101 = n79333 & n43099 ;
  assign n43102 = n42963 | n43101 ;
  assign n43103 = n79336 & n43102 ;
  assign n43104 = n42969 | n43103 ;
  assign n43106 = n79339 & n43104 ;
  assign n43107 = n42974 | n43106 ;
  assign n43108 = n79342 & n43107 ;
  assign n43109 = n42980 | n43108 ;
  assign n43111 = n79345 & n43109 ;
  assign n43112 = n42985 | n43111 ;
  assign n43113 = n79348 & n43112 ;
  assign n43114 = n42991 | n43113 ;
  assign n43116 = n79351 & n43114 ;
  assign n43117 = n42996 | n43116 ;
  assign n43118 = n79354 & n43117 ;
  assign n43119 = n43002 | n43118 ;
  assign n43121 = n79357 & n43119 ;
  assign n43122 = n43007 | n43121 ;
  assign n43123 = n79360 & n43122 ;
  assign n43124 = n43013 | n43123 ;
  assign n43126 = n42574 | n43018 ;
  assign n79373 = ~n43126 ;
  assign n43127 = n43124 & n79373 ;
  assign n43128 = n43019 | n43127 ;
  assign n79374 = ~n43037 ;
  assign n43129 = n79374 & n43128 ;
  assign n43130 = n79363 & n43124 ;
  assign n43131 = n43018 | n43130 ;
  assign n43132 = n79366 & n43131 ;
  assign n43133 = n43034 | n43132 ;
  assign n43134 = n42565 & n79370 ;
  assign n43135 = n43133 & n43134 ;
  assign n43136 = n43129 | n43135 ;
  assign n43137 = n42566 | n43032 ;
  assign n43138 = n43028 | n43137 ;
  assign n79375 = ~n43138 ;
  assign n43139 = n43020 & n79375 ;
  assign n43140 = n43028 | n43032 ;
  assign n79376 = ~n43132 ;
  assign n43141 = n79376 & n43140 ;
  assign n43142 = n43139 | n43141 ;
  assign n43143 = n79374 & n43142 ;
  assign n43144 = n10157 & n42027 ;
  assign n43145 = n43133 & n43144 ;
  assign n43146 = n43143 | n43145 ;
  assign n43147 = n69075 & n43146 ;
  assign n79377 = ~n43145 ;
  assign n43626 = x100 & n79377 ;
  assign n79378 = ~n43143 ;
  assign n43627 = n79378 & n43626 ;
  assign n43628 = n43147 | n43627 ;
  assign n43148 = n68993 & n43136 ;
  assign n79379 = ~n43123 ;
  assign n43125 = n43013 & n79379 ;
  assign n43149 = n42582 | n43013 ;
  assign n79380 = ~n43149 ;
  assign n43150 = n43009 & n79380 ;
  assign n43151 = n43125 | n43150 ;
  assign n43152 = n79374 & n43151 ;
  assign n43153 = n42573 & n79370 ;
  assign n43154 = n43133 & n43153 ;
  assign n43155 = n43152 | n43154 ;
  assign n43156 = n68716 & n43155 ;
  assign n79381 = ~n43154 ;
  assign n43614 = x98 & n79381 ;
  assign n79382 = ~n43152 ;
  assign n43615 = n79382 & n43614 ;
  assign n43616 = n43156 | n43615 ;
  assign n79383 = ~n43004 ;
  assign n43008 = n79383 & n43007 ;
  assign n43157 = n42590 | n43007 ;
  assign n79384 = ~n43157 ;
  assign n43158 = n43119 & n79384 ;
  assign n43159 = n43008 | n43158 ;
  assign n43160 = n79374 & n43159 ;
  assign n43161 = n42581 & n79370 ;
  assign n43162 = n43133 & n43161 ;
  assign n43163 = n43160 | n43162 ;
  assign n43164 = n68545 & n43163 ;
  assign n79385 = ~n43118 ;
  assign n43120 = n43002 & n79385 ;
  assign n43165 = n42598 | n43002 ;
  assign n79386 = ~n43165 ;
  assign n43166 = n42998 & n79386 ;
  assign n43167 = n43120 | n43166 ;
  assign n43168 = n79374 & n43167 ;
  assign n43169 = n42589 & n79370 ;
  assign n43170 = n43133 & n43169 ;
  assign n43171 = n43168 | n43170 ;
  assign n43172 = n68438 & n43171 ;
  assign n79387 = ~n43170 ;
  assign n43602 = x96 & n79387 ;
  assign n79388 = ~n43168 ;
  assign n43603 = n79388 & n43602 ;
  assign n43604 = n43172 | n43603 ;
  assign n79389 = ~n42993 ;
  assign n42997 = n79389 & n42996 ;
  assign n43173 = n42606 | n42996 ;
  assign n79390 = ~n43173 ;
  assign n43174 = n43114 & n79390 ;
  assign n43175 = n42997 | n43174 ;
  assign n43176 = n79374 & n43175 ;
  assign n43177 = n42597 & n79370 ;
  assign n43178 = n43133 & n43177 ;
  assign n43179 = n43176 | n43178 ;
  assign n43180 = n68214 & n43179 ;
  assign n79391 = ~n43113 ;
  assign n43115 = n42991 & n79391 ;
  assign n43181 = n42614 | n42991 ;
  assign n79392 = ~n43181 ;
  assign n43182 = n42987 & n79392 ;
  assign n43183 = n43115 | n43182 ;
  assign n43184 = n79374 & n43183 ;
  assign n43185 = n42605 & n79370 ;
  assign n43186 = n43133 & n43185 ;
  assign n43187 = n43184 | n43186 ;
  assign n43188 = n68058 & n43187 ;
  assign n79393 = ~n43186 ;
  assign n43590 = x94 & n79393 ;
  assign n79394 = ~n43184 ;
  assign n43591 = n79394 & n43590 ;
  assign n43592 = n43188 | n43591 ;
  assign n79395 = ~n42982 ;
  assign n42986 = n79395 & n42985 ;
  assign n43189 = n42622 | n42985 ;
  assign n79396 = ~n43189 ;
  assign n43190 = n43109 & n79396 ;
  assign n43191 = n42986 | n43190 ;
  assign n43192 = n79374 & n43191 ;
  assign n43193 = n42613 & n79370 ;
  assign n43194 = n43133 & n43193 ;
  assign n43195 = n43192 | n43194 ;
  assign n43196 = n67986 & n43195 ;
  assign n79397 = ~n43108 ;
  assign n43110 = n42980 & n79397 ;
  assign n43197 = n42630 | n42980 ;
  assign n79398 = ~n43197 ;
  assign n43198 = n42976 & n79398 ;
  assign n43199 = n43110 | n43198 ;
  assign n43200 = n79374 & n43199 ;
  assign n43201 = n42621 & n79370 ;
  assign n43202 = n43133 & n43201 ;
  assign n43203 = n43200 | n43202 ;
  assign n43204 = n67763 & n43203 ;
  assign n79399 = ~n43202 ;
  assign n43578 = x92 & n79399 ;
  assign n79400 = ~n43200 ;
  assign n43579 = n79400 & n43578 ;
  assign n43580 = n43204 | n43579 ;
  assign n79401 = ~n42971 ;
  assign n42975 = n79401 & n42974 ;
  assign n43205 = n42638 | n42974 ;
  assign n79402 = ~n43205 ;
  assign n43206 = n43104 & n79402 ;
  assign n43207 = n42975 | n43206 ;
  assign n43208 = n79374 & n43207 ;
  assign n43209 = n42629 & n79370 ;
  assign n43210 = n43133 & n43209 ;
  assign n43211 = n43208 | n43210 ;
  assign n43212 = n67622 & n43211 ;
  assign n79403 = ~n43103 ;
  assign n43105 = n42969 & n79403 ;
  assign n43213 = n42646 | n42969 ;
  assign n79404 = ~n43213 ;
  assign n43214 = n42965 & n79404 ;
  assign n43215 = n43105 | n43214 ;
  assign n43216 = n79374 & n43215 ;
  assign n43217 = n42637 & n79370 ;
  assign n43218 = n43133 & n43217 ;
  assign n43219 = n43216 | n43218 ;
  assign n43220 = n67531 & n43219 ;
  assign n79405 = ~n43218 ;
  assign n43566 = x90 & n79405 ;
  assign n79406 = ~n43216 ;
  assign n43567 = n79406 & n43566 ;
  assign n43568 = n43220 | n43567 ;
  assign n79407 = ~n42960 ;
  assign n42964 = n79407 & n42963 ;
  assign n43221 = n42654 | n42963 ;
  assign n79408 = ~n43221 ;
  assign n43222 = n43099 & n79408 ;
  assign n43223 = n42964 | n43222 ;
  assign n43224 = n79374 & n43223 ;
  assign n43225 = n42645 & n79370 ;
  assign n43226 = n43133 & n43225 ;
  assign n43227 = n43224 | n43226 ;
  assign n43228 = n67348 & n43227 ;
  assign n79409 = ~n43098 ;
  assign n43100 = n42958 & n79409 ;
  assign n43229 = n42662 | n42958 ;
  assign n79410 = ~n43229 ;
  assign n43230 = n42954 & n79410 ;
  assign n43231 = n43100 | n43230 ;
  assign n43232 = n79374 & n43231 ;
  assign n43233 = n42653 & n79370 ;
  assign n43234 = n43133 & n43233 ;
  assign n43235 = n43232 | n43234 ;
  assign n43236 = n67222 & n43235 ;
  assign n79411 = ~n43234 ;
  assign n43554 = x88 & n79411 ;
  assign n79412 = ~n43232 ;
  assign n43555 = n79412 & n43554 ;
  assign n43556 = n43236 | n43555 ;
  assign n79413 = ~n42949 ;
  assign n42953 = n79413 & n42952 ;
  assign n43237 = n42670 | n42952 ;
  assign n79414 = ~n43237 ;
  assign n43238 = n43094 & n79414 ;
  assign n43239 = n42953 | n43238 ;
  assign n43240 = n79374 & n43239 ;
  assign n43241 = n42661 & n79370 ;
  assign n43242 = n43133 & n43241 ;
  assign n43243 = n43240 | n43242 ;
  assign n43244 = n67164 & n43243 ;
  assign n79415 = ~n43093 ;
  assign n43095 = n42947 & n79415 ;
  assign n43245 = n42678 | n42947 ;
  assign n79416 = ~n43245 ;
  assign n43246 = n42943 & n79416 ;
  assign n43247 = n43095 | n43246 ;
  assign n43248 = n79374 & n43247 ;
  assign n43249 = n42669 & n79370 ;
  assign n43250 = n43133 & n43249 ;
  assign n43251 = n43248 | n43250 ;
  assign n43252 = n66979 & n43251 ;
  assign n79417 = ~n43250 ;
  assign n43542 = x86 & n79417 ;
  assign n79418 = ~n43248 ;
  assign n43543 = n79418 & n43542 ;
  assign n43544 = n43252 | n43543 ;
  assign n79419 = ~n42938 ;
  assign n42942 = n79419 & n42941 ;
  assign n43253 = n42686 | n42941 ;
  assign n79420 = ~n43253 ;
  assign n43254 = n43089 & n79420 ;
  assign n43255 = n42942 | n43254 ;
  assign n43256 = n79374 & n43255 ;
  assign n43257 = n42677 & n79370 ;
  assign n43258 = n43133 & n43257 ;
  assign n43259 = n43256 | n43258 ;
  assign n43260 = n66868 & n43259 ;
  assign n79421 = ~n43088 ;
  assign n43090 = n42936 & n79421 ;
  assign n43261 = n42694 | n42936 ;
  assign n79422 = ~n43261 ;
  assign n43262 = n42932 & n79422 ;
  assign n43263 = n43090 | n43262 ;
  assign n43264 = n79374 & n43263 ;
  assign n43265 = n42685 & n79370 ;
  assign n43266 = n43133 & n43265 ;
  assign n43267 = n43264 | n43266 ;
  assign n43268 = n66797 & n43267 ;
  assign n79423 = ~n43266 ;
  assign n43530 = x84 & n79423 ;
  assign n79424 = ~n43264 ;
  assign n43531 = n79424 & n43530 ;
  assign n43532 = n43268 | n43531 ;
  assign n79425 = ~n42927 ;
  assign n42931 = n79425 & n42930 ;
  assign n43269 = n42702 | n42930 ;
  assign n79426 = ~n43269 ;
  assign n43270 = n43084 & n79426 ;
  assign n43271 = n42931 | n43270 ;
  assign n43272 = n79374 & n43271 ;
  assign n43273 = n42693 & n79370 ;
  assign n43274 = n43133 & n43273 ;
  assign n43275 = n43272 | n43274 ;
  assign n43276 = n66654 & n43275 ;
  assign n79427 = ~n43083 ;
  assign n43085 = n42925 & n79427 ;
  assign n43277 = n42710 | n42925 ;
  assign n79428 = ~n43277 ;
  assign n43278 = n42921 & n79428 ;
  assign n43279 = n43085 | n43278 ;
  assign n43280 = n79374 & n43279 ;
  assign n43281 = n42701 & n79370 ;
  assign n43282 = n43133 & n43281 ;
  assign n43283 = n43280 | n43282 ;
  assign n43284 = n66560 & n43283 ;
  assign n79429 = ~n43282 ;
  assign n43518 = x82 & n79429 ;
  assign n79430 = ~n43280 ;
  assign n43519 = n79430 & n43518 ;
  assign n43520 = n43284 | n43519 ;
  assign n79431 = ~n42916 ;
  assign n42920 = n79431 & n42919 ;
  assign n43285 = n42718 | n42919 ;
  assign n79432 = ~n43285 ;
  assign n43286 = n43079 & n79432 ;
  assign n43287 = n42920 | n43286 ;
  assign n43288 = n79374 & n43287 ;
  assign n43289 = n42709 & n79370 ;
  assign n43290 = n43133 & n43289 ;
  assign n43291 = n43288 | n43290 ;
  assign n43292 = n66505 & n43291 ;
  assign n79433 = ~n43078 ;
  assign n43080 = n42914 & n79433 ;
  assign n43293 = n42726 | n42914 ;
  assign n79434 = ~n43293 ;
  assign n43294 = n42910 & n79434 ;
  assign n43295 = n43080 | n43294 ;
  assign n43296 = n79374 & n43295 ;
  assign n43297 = n42717 & n79370 ;
  assign n43298 = n43133 & n43297 ;
  assign n43299 = n43296 | n43298 ;
  assign n43300 = n66379 & n43299 ;
  assign n79435 = ~n43298 ;
  assign n43506 = x80 & n79435 ;
  assign n79436 = ~n43296 ;
  assign n43507 = n79436 & n43506 ;
  assign n43508 = n43300 | n43507 ;
  assign n79437 = ~n42905 ;
  assign n42909 = n79437 & n42908 ;
  assign n43301 = n42734 | n42908 ;
  assign n79438 = ~n43301 ;
  assign n43302 = n43074 & n79438 ;
  assign n43303 = n42909 | n43302 ;
  assign n43304 = n79374 & n43303 ;
  assign n43305 = n42725 & n79370 ;
  assign n43306 = n43133 & n43305 ;
  assign n43307 = n43304 | n43306 ;
  assign n43308 = n66299 & n43307 ;
  assign n79439 = ~n43073 ;
  assign n43075 = n42903 & n79439 ;
  assign n43309 = n42742 | n42903 ;
  assign n79440 = ~n43309 ;
  assign n43310 = n42899 & n79440 ;
  assign n43311 = n43075 | n43310 ;
  assign n43312 = n79374 & n43311 ;
  assign n43313 = n42733 & n79370 ;
  assign n43314 = n43133 & n43313 ;
  assign n43315 = n43312 | n43314 ;
  assign n43316 = n66244 & n43315 ;
  assign n79441 = ~n43314 ;
  assign n43494 = x78 & n79441 ;
  assign n79442 = ~n43312 ;
  assign n43495 = n79442 & n43494 ;
  assign n43496 = n43316 | n43495 ;
  assign n79443 = ~n42894 ;
  assign n42898 = n79443 & n42897 ;
  assign n43317 = n42750 | n42897 ;
  assign n79444 = ~n43317 ;
  assign n43318 = n43069 & n79444 ;
  assign n43319 = n42898 | n43318 ;
  assign n43320 = n79374 & n43319 ;
  assign n43321 = n42741 & n79370 ;
  assign n43322 = n43133 & n43321 ;
  assign n43323 = n43320 | n43322 ;
  assign n43324 = n66145 & n43323 ;
  assign n79445 = ~n43068 ;
  assign n43070 = n42892 & n79445 ;
  assign n43325 = n42758 | n42892 ;
  assign n79446 = ~n43325 ;
  assign n43326 = n42888 & n79446 ;
  assign n43327 = n43070 | n43326 ;
  assign n43328 = n79374 & n43327 ;
  assign n43329 = n42749 & n79370 ;
  assign n43330 = n43133 & n43329 ;
  assign n43331 = n43328 | n43330 ;
  assign n43332 = n66081 & n43331 ;
  assign n79447 = ~n43330 ;
  assign n43482 = x76 & n79447 ;
  assign n79448 = ~n43328 ;
  assign n43483 = n79448 & n43482 ;
  assign n43484 = n43332 | n43483 ;
  assign n79449 = ~n42883 ;
  assign n42887 = n79449 & n42886 ;
  assign n43333 = n42766 | n42886 ;
  assign n79450 = ~n43333 ;
  assign n43334 = n43064 & n79450 ;
  assign n43335 = n42887 | n43334 ;
  assign n43336 = n79374 & n43335 ;
  assign n43337 = n42757 & n79370 ;
  assign n43338 = n43133 & n43337 ;
  assign n43339 = n43336 | n43338 ;
  assign n43340 = n66043 & n43339 ;
  assign n79451 = ~n43063 ;
  assign n43065 = n42881 & n79451 ;
  assign n43341 = n42774 | n42881 ;
  assign n79452 = ~n43341 ;
  assign n43342 = n42877 & n79452 ;
  assign n43343 = n43065 | n43342 ;
  assign n43344 = n79374 & n43343 ;
  assign n43345 = n42765 & n79370 ;
  assign n43346 = n43133 & n43345 ;
  assign n43347 = n43344 | n43346 ;
  assign n43348 = n65960 & n43347 ;
  assign n79453 = ~n43346 ;
  assign n43470 = x74 & n79453 ;
  assign n79454 = ~n43344 ;
  assign n43471 = n79454 & n43470 ;
  assign n43472 = n43348 | n43471 ;
  assign n79455 = ~n42872 ;
  assign n42876 = n79455 & n42875 ;
  assign n43349 = n42782 | n42875 ;
  assign n79456 = ~n43349 ;
  assign n43350 = n43059 & n79456 ;
  assign n43351 = n42876 | n43350 ;
  assign n43352 = n79374 & n43351 ;
  assign n43353 = n42773 & n79370 ;
  assign n43354 = n43133 & n43353 ;
  assign n43355 = n43352 | n43354 ;
  assign n43356 = n65909 & n43355 ;
  assign n79457 = ~n43058 ;
  assign n43060 = n42870 & n79457 ;
  assign n43357 = n42791 | n42870 ;
  assign n79458 = ~n43357 ;
  assign n43358 = n42866 & n79458 ;
  assign n43359 = n43060 | n43358 ;
  assign n43360 = n79374 & n43359 ;
  assign n43361 = n42781 & n79370 ;
  assign n43362 = n43133 & n43361 ;
  assign n43363 = n43360 | n43362 ;
  assign n43364 = n65877 & n43363 ;
  assign n79459 = ~n43362 ;
  assign n43458 = x72 & n79459 ;
  assign n79460 = ~n43360 ;
  assign n43459 = n79460 & n43458 ;
  assign n43460 = n43364 | n43459 ;
  assign n79461 = ~n42861 ;
  assign n42865 = n79461 & n42864 ;
  assign n43365 = n42800 | n42864 ;
  assign n79462 = ~n43365 ;
  assign n43366 = n43055 & n79462 ;
  assign n43367 = n42865 | n43366 ;
  assign n43368 = n79374 & n43367 ;
  assign n43369 = n42790 & n79370 ;
  assign n43370 = n43133 & n43369 ;
  assign n43371 = n43368 | n43370 ;
  assign n43372 = n65820 & n43371 ;
  assign n79463 = ~n43053 ;
  assign n43054 = n42859 & n79463 ;
  assign n43373 = n42809 | n42859 ;
  assign n79464 = ~n43373 ;
  assign n43374 = n42855 & n79464 ;
  assign n43375 = n43054 | n43374 ;
  assign n43376 = n79374 & n43375 ;
  assign n43377 = n42799 & n79370 ;
  assign n43378 = n43133 & n43377 ;
  assign n43379 = n43376 | n43378 ;
  assign n43380 = n65791 & n43379 ;
  assign n79465 = ~n43378 ;
  assign n43446 = x70 & n79465 ;
  assign n79466 = ~n43376 ;
  assign n43447 = n79466 & n43446 ;
  assign n43448 = n43380 | n43447 ;
  assign n79467 = ~n42851 ;
  assign n43051 = n79467 & n42854 ;
  assign n43381 = n42849 | n43047 ;
  assign n43382 = n42818 | n42854 ;
  assign n79468 = ~n43382 ;
  assign n43383 = n43381 & n79468 ;
  assign n43384 = n43051 | n43383 ;
  assign n43385 = n79374 & n43384 ;
  assign n43386 = n42808 & n79370 ;
  assign n43387 = n43133 & n43386 ;
  assign n43388 = n43385 | n43387 ;
  assign n43389 = n65772 & n43388 ;
  assign n79469 = ~n43047 ;
  assign n43049 = n42849 & n79469 ;
  assign n43390 = n42824 | n42849 ;
  assign n79470 = ~n43390 ;
  assign n43391 = n43046 & n79470 ;
  assign n43392 = n43049 | n43391 ;
  assign n43393 = n79374 & n43392 ;
  assign n43394 = n42817 & n79370 ;
  assign n43395 = n43133 & n43394 ;
  assign n43396 = n43393 | n43395 ;
  assign n43397 = n65746 & n43396 ;
  assign n79471 = ~n43395 ;
  assign n43435 = x68 & n79471 ;
  assign n79472 = ~n43393 ;
  assign n43436 = n79472 & n43435 ;
  assign n43437 = n43397 | n43436 ;
  assign n79473 = ~n42842 ;
  assign n43045 = n79473 & n43044 ;
  assign n43398 = n42840 | n43044 ;
  assign n79474 = ~n43398 ;
  assign n43399 = n42841 & n79474 ;
  assign n43400 = n43045 | n43399 ;
  assign n43401 = n79374 & n43400 ;
  assign n43402 = n42823 & n79370 ;
  assign n43403 = n43133 & n43402 ;
  assign n43404 = n43401 | n43403 ;
  assign n43405 = n65721 & n43404 ;
  assign n43406 = n10529 & n42838 ;
  assign n43407 = n79372 & n43406 ;
  assign n79475 = ~n43407 ;
  assign n43408 = n42841 & n79475 ;
  assign n43409 = n79374 & n43408 ;
  assign n43410 = n42832 & n79370 ;
  assign n43411 = n43133 & n43410 ;
  assign n43412 = n43409 | n43411 ;
  assign n43413 = n65686 & n43412 ;
  assign n79476 = ~n43411 ;
  assign n43425 = x66 & n79476 ;
  assign n79477 = ~n43409 ;
  assign n43426 = n79477 & n43425 ;
  assign n43427 = n43413 | n43426 ;
  assign n43039 = n10529 & n79374 ;
  assign n43038 = x64 & n79374 ;
  assign n79478 = ~n43038 ;
  assign n43414 = x28 & n79478 ;
  assign n43415 = n43039 | n43414 ;
  assign n43416 = x65 & n43415 ;
  assign n43417 = n79370 & n43133 ;
  assign n79479 = ~n43417 ;
  assign n43418 = n10529 & n79479 ;
  assign n43419 = x65 | n43418 ;
  assign n43420 = n43414 | n43419 ;
  assign n79480 = ~n43416 ;
  assign n43421 = n79480 & n43420 ;
  assign n43423 = n11115 | n43421 ;
  assign n43424 = n65670 & n43415 ;
  assign n79481 = ~n43424 ;
  assign n43428 = n43423 & n79481 ;
  assign n43429 = n43427 | n43428 ;
  assign n79482 = ~n43413 ;
  assign n43430 = n79482 & n43429 ;
  assign n79483 = ~n43403 ;
  assign n43431 = x67 & n79483 ;
  assign n79484 = ~n43401 ;
  assign n43432 = n79484 & n43431 ;
  assign n43433 = n43405 | n43432 ;
  assign n43434 = n43430 | n43433 ;
  assign n79485 = ~n43405 ;
  assign n43438 = n79485 & n43434 ;
  assign n43439 = n43437 | n43438 ;
  assign n79486 = ~n43397 ;
  assign n43440 = n79486 & n43439 ;
  assign n79487 = ~n43387 ;
  assign n43441 = x69 & n79487 ;
  assign n79488 = ~n43385 ;
  assign n43442 = n79488 & n43441 ;
  assign n43443 = n43389 | n43442 ;
  assign n43445 = n43440 | n43443 ;
  assign n79489 = ~n43389 ;
  assign n43450 = n79489 & n43445 ;
  assign n43451 = n43448 | n43450 ;
  assign n79490 = ~n43380 ;
  assign n43452 = n79490 & n43451 ;
  assign n79491 = ~n43370 ;
  assign n43453 = x71 & n79491 ;
  assign n79492 = ~n43368 ;
  assign n43454 = n79492 & n43453 ;
  assign n43455 = n43372 | n43454 ;
  assign n43457 = n43452 | n43455 ;
  assign n79493 = ~n43372 ;
  assign n43462 = n79493 & n43457 ;
  assign n43463 = n43460 | n43462 ;
  assign n79494 = ~n43364 ;
  assign n43464 = n79494 & n43463 ;
  assign n79495 = ~n43354 ;
  assign n43465 = x73 & n79495 ;
  assign n79496 = ~n43352 ;
  assign n43466 = n79496 & n43465 ;
  assign n43467 = n43356 | n43466 ;
  assign n43469 = n43464 | n43467 ;
  assign n79497 = ~n43356 ;
  assign n43474 = n79497 & n43469 ;
  assign n43475 = n43472 | n43474 ;
  assign n79498 = ~n43348 ;
  assign n43476 = n79498 & n43475 ;
  assign n79499 = ~n43338 ;
  assign n43477 = x75 & n79499 ;
  assign n79500 = ~n43336 ;
  assign n43478 = n79500 & n43477 ;
  assign n43479 = n43340 | n43478 ;
  assign n43481 = n43476 | n43479 ;
  assign n79501 = ~n43340 ;
  assign n43486 = n79501 & n43481 ;
  assign n43487 = n43484 | n43486 ;
  assign n79502 = ~n43332 ;
  assign n43488 = n79502 & n43487 ;
  assign n79503 = ~n43322 ;
  assign n43489 = x77 & n79503 ;
  assign n79504 = ~n43320 ;
  assign n43490 = n79504 & n43489 ;
  assign n43491 = n43324 | n43490 ;
  assign n43493 = n43488 | n43491 ;
  assign n79505 = ~n43324 ;
  assign n43498 = n79505 & n43493 ;
  assign n43499 = n43496 | n43498 ;
  assign n79506 = ~n43316 ;
  assign n43500 = n79506 & n43499 ;
  assign n79507 = ~n43306 ;
  assign n43501 = x79 & n79507 ;
  assign n79508 = ~n43304 ;
  assign n43502 = n79508 & n43501 ;
  assign n43503 = n43308 | n43502 ;
  assign n43505 = n43500 | n43503 ;
  assign n79509 = ~n43308 ;
  assign n43510 = n79509 & n43505 ;
  assign n43511 = n43508 | n43510 ;
  assign n79510 = ~n43300 ;
  assign n43512 = n79510 & n43511 ;
  assign n79511 = ~n43290 ;
  assign n43513 = x81 & n79511 ;
  assign n79512 = ~n43288 ;
  assign n43514 = n79512 & n43513 ;
  assign n43515 = n43292 | n43514 ;
  assign n43517 = n43512 | n43515 ;
  assign n79513 = ~n43292 ;
  assign n43522 = n79513 & n43517 ;
  assign n43523 = n43520 | n43522 ;
  assign n79514 = ~n43284 ;
  assign n43524 = n79514 & n43523 ;
  assign n79515 = ~n43274 ;
  assign n43525 = x83 & n79515 ;
  assign n79516 = ~n43272 ;
  assign n43526 = n79516 & n43525 ;
  assign n43527 = n43276 | n43526 ;
  assign n43529 = n43524 | n43527 ;
  assign n79517 = ~n43276 ;
  assign n43534 = n79517 & n43529 ;
  assign n43535 = n43532 | n43534 ;
  assign n79518 = ~n43268 ;
  assign n43536 = n79518 & n43535 ;
  assign n79519 = ~n43258 ;
  assign n43537 = x85 & n79519 ;
  assign n79520 = ~n43256 ;
  assign n43538 = n79520 & n43537 ;
  assign n43539 = n43260 | n43538 ;
  assign n43541 = n43536 | n43539 ;
  assign n79521 = ~n43260 ;
  assign n43546 = n79521 & n43541 ;
  assign n43547 = n43544 | n43546 ;
  assign n79522 = ~n43252 ;
  assign n43548 = n79522 & n43547 ;
  assign n79523 = ~n43242 ;
  assign n43549 = x87 & n79523 ;
  assign n79524 = ~n43240 ;
  assign n43550 = n79524 & n43549 ;
  assign n43551 = n43244 | n43550 ;
  assign n43553 = n43548 | n43551 ;
  assign n79525 = ~n43244 ;
  assign n43558 = n79525 & n43553 ;
  assign n43559 = n43556 | n43558 ;
  assign n79526 = ~n43236 ;
  assign n43560 = n79526 & n43559 ;
  assign n79527 = ~n43226 ;
  assign n43561 = x89 & n79527 ;
  assign n79528 = ~n43224 ;
  assign n43562 = n79528 & n43561 ;
  assign n43563 = n43228 | n43562 ;
  assign n43565 = n43560 | n43563 ;
  assign n79529 = ~n43228 ;
  assign n43570 = n79529 & n43565 ;
  assign n43571 = n43568 | n43570 ;
  assign n79530 = ~n43220 ;
  assign n43572 = n79530 & n43571 ;
  assign n79531 = ~n43210 ;
  assign n43573 = x91 & n79531 ;
  assign n79532 = ~n43208 ;
  assign n43574 = n79532 & n43573 ;
  assign n43575 = n43212 | n43574 ;
  assign n43577 = n43572 | n43575 ;
  assign n79533 = ~n43212 ;
  assign n43582 = n79533 & n43577 ;
  assign n43583 = n43580 | n43582 ;
  assign n79534 = ~n43204 ;
  assign n43584 = n79534 & n43583 ;
  assign n79535 = ~n43194 ;
  assign n43585 = x93 & n79535 ;
  assign n79536 = ~n43192 ;
  assign n43586 = n79536 & n43585 ;
  assign n43587 = n43196 | n43586 ;
  assign n43589 = n43584 | n43587 ;
  assign n79537 = ~n43196 ;
  assign n43594 = n79537 & n43589 ;
  assign n43595 = n43592 | n43594 ;
  assign n79538 = ~n43188 ;
  assign n43596 = n79538 & n43595 ;
  assign n79539 = ~n43178 ;
  assign n43597 = x95 & n79539 ;
  assign n79540 = ~n43176 ;
  assign n43598 = n79540 & n43597 ;
  assign n43599 = n43180 | n43598 ;
  assign n43601 = n43596 | n43599 ;
  assign n79541 = ~n43180 ;
  assign n43606 = n79541 & n43601 ;
  assign n43607 = n43604 | n43606 ;
  assign n79542 = ~n43172 ;
  assign n43608 = n79542 & n43607 ;
  assign n79543 = ~n43162 ;
  assign n43609 = x97 & n79543 ;
  assign n79544 = ~n43160 ;
  assign n43610 = n79544 & n43609 ;
  assign n43611 = n43164 | n43610 ;
  assign n43613 = n43608 | n43611 ;
  assign n79545 = ~n43164 ;
  assign n43618 = n79545 & n43613 ;
  assign n43619 = n43616 | n43618 ;
  assign n79546 = ~n43156 ;
  assign n43620 = n79546 & n43619 ;
  assign n79547 = ~n43135 ;
  assign n43621 = x99 & n79547 ;
  assign n79548 = ~n43129 ;
  assign n43622 = n79548 & n43621 ;
  assign n43623 = n43148 | n43622 ;
  assign n43625 = n43620 | n43623 ;
  assign n79549 = ~n43148 ;
  assign n43629 = n79549 & n43625 ;
  assign n43630 = n43628 | n43629 ;
  assign n79550 = ~n43147 ;
  assign n43631 = n79550 & n43630 ;
  assign n43632 = n469 | n43631 ;
  assign n43635 = n43136 & n43632 ;
  assign n43624 = n43156 | n43623 ;
  assign n43636 = x64 & n79479 ;
  assign n79551 = ~n43636 ;
  assign n43637 = x28 & n79551 ;
  assign n43638 = n43039 | n43637 ;
  assign n43639 = x65 & n43638 ;
  assign n79552 = ~n43639 ;
  assign n43640 = n43420 & n79552 ;
  assign n43641 = n11115 | n43640 ;
  assign n43642 = n79481 & n43641 ;
  assign n43644 = n43427 | n43642 ;
  assign n43645 = n79482 & n43644 ;
  assign n43646 = n43433 | n43645 ;
  assign n43647 = n79485 & n43646 ;
  assign n43648 = n43437 | n43647 ;
  assign n43649 = n79486 & n43648 ;
  assign n43650 = n43443 | n43649 ;
  assign n43651 = n79489 & n43650 ;
  assign n43652 = n43448 | n43651 ;
  assign n43653 = n79490 & n43652 ;
  assign n43654 = n43455 | n43653 ;
  assign n43655 = n79493 & n43654 ;
  assign n43656 = n43460 | n43655 ;
  assign n43657 = n79494 & n43656 ;
  assign n43658 = n43467 | n43657 ;
  assign n43659 = n79497 & n43658 ;
  assign n43660 = n43472 | n43659 ;
  assign n43661 = n79498 & n43660 ;
  assign n43662 = n43479 | n43661 ;
  assign n43663 = n79501 & n43662 ;
  assign n43664 = n43484 | n43663 ;
  assign n43665 = n79502 & n43664 ;
  assign n43666 = n43491 | n43665 ;
  assign n43667 = n79505 & n43666 ;
  assign n43668 = n43496 | n43667 ;
  assign n43669 = n79506 & n43668 ;
  assign n43670 = n43503 | n43669 ;
  assign n43671 = n79509 & n43670 ;
  assign n43672 = n43508 | n43671 ;
  assign n43673 = n79510 & n43672 ;
  assign n43674 = n43515 | n43673 ;
  assign n43675 = n79513 & n43674 ;
  assign n43676 = n43520 | n43675 ;
  assign n43677 = n79514 & n43676 ;
  assign n43678 = n43527 | n43677 ;
  assign n43679 = n79517 & n43678 ;
  assign n43680 = n43532 | n43679 ;
  assign n43681 = n79518 & n43680 ;
  assign n43682 = n43539 | n43681 ;
  assign n43683 = n79521 & n43682 ;
  assign n43684 = n43544 | n43683 ;
  assign n43685 = n79522 & n43684 ;
  assign n43686 = n43551 | n43685 ;
  assign n43687 = n79525 & n43686 ;
  assign n43688 = n43556 | n43687 ;
  assign n43689 = n79526 & n43688 ;
  assign n43690 = n43563 | n43689 ;
  assign n43691 = n79529 & n43690 ;
  assign n43692 = n43568 | n43691 ;
  assign n43693 = n79530 & n43692 ;
  assign n43694 = n43575 | n43693 ;
  assign n43695 = n79533 & n43694 ;
  assign n43696 = n43580 | n43695 ;
  assign n43697 = n79534 & n43696 ;
  assign n43698 = n43587 | n43697 ;
  assign n43699 = n79537 & n43698 ;
  assign n43700 = n43592 | n43699 ;
  assign n43701 = n79538 & n43700 ;
  assign n43702 = n43599 | n43701 ;
  assign n43703 = n79541 & n43702 ;
  assign n43704 = n43604 | n43703 ;
  assign n43705 = n79542 & n43704 ;
  assign n43706 = n43611 | n43705 ;
  assign n43707 = n79545 & n43706 ;
  assign n43708 = n43616 | n43707 ;
  assign n79553 = ~n43624 ;
  assign n43709 = n79553 & n43708 ;
  assign n43710 = n79546 & n43708 ;
  assign n79554 = ~n43710 ;
  assign n43711 = n43623 & n79554 ;
  assign n43712 = n43709 | n43711 ;
  assign n43713 = n65845 & n43712 ;
  assign n79555 = ~n43631 ;
  assign n43714 = n79555 & n43713 ;
  assign n43715 = n43635 | n43714 ;
  assign n79556 = ~n43146 ;
  assign n43634 = n79556 & n43632 ;
  assign n79557 = ~n43629 ;
  assign n43718 = n43628 & n79557 ;
  assign n43716 = n43623 | n43710 ;
  assign n43719 = n43148 | n43628 ;
  assign n79558 = ~n43719 ;
  assign n43720 = n43716 & n79558 ;
  assign n43721 = n43718 | n43720 ;
  assign n43722 = n43632 | n43721 ;
  assign n79559 = ~n43634 ;
  assign n43723 = n79559 & n43722 ;
  assign n43724 = n69261 & n43723 ;
  assign n43725 = n69075 & n43715 ;
  assign n43726 = n43155 & n43632 ;
  assign n43617 = n43164 | n43616 ;
  assign n79560 = ~n43617 ;
  assign n43727 = n43613 & n79560 ;
  assign n79561 = ~n43618 ;
  assign n43728 = n43616 & n79561 ;
  assign n43729 = n43727 | n43728 ;
  assign n43730 = n65845 & n43729 ;
  assign n43731 = n79555 & n43730 ;
  assign n43732 = n43726 | n43731 ;
  assign n43733 = n68993 & n43732 ;
  assign n43734 = n43163 & n43632 ;
  assign n43612 = n43172 | n43611 ;
  assign n79562 = ~n43612 ;
  assign n43735 = n79562 & n43704 ;
  assign n79563 = ~n43705 ;
  assign n43736 = n43611 & n79563 ;
  assign n43737 = n43735 | n43736 ;
  assign n43738 = n65845 & n43737 ;
  assign n43739 = n79555 & n43738 ;
  assign n43740 = n43734 | n43739 ;
  assign n43741 = n68716 & n43740 ;
  assign n43742 = n43171 & n43632 ;
  assign n43605 = n43180 | n43604 ;
  assign n79564 = ~n43605 ;
  assign n43743 = n43601 & n79564 ;
  assign n79565 = ~n43606 ;
  assign n43744 = n43604 & n79565 ;
  assign n43745 = n43743 | n43744 ;
  assign n43746 = n65845 & n43745 ;
  assign n43747 = n79555 & n43746 ;
  assign n43748 = n43742 | n43747 ;
  assign n43749 = n68545 & n43748 ;
  assign n43750 = n43179 & n43632 ;
  assign n43600 = n43188 | n43599 ;
  assign n79566 = ~n43600 ;
  assign n43751 = n79566 & n43700 ;
  assign n79567 = ~n43701 ;
  assign n43752 = n43599 & n79567 ;
  assign n43753 = n43751 | n43752 ;
  assign n43754 = n65845 & n43753 ;
  assign n43755 = n79555 & n43754 ;
  assign n43756 = n43750 | n43755 ;
  assign n43757 = n68438 & n43756 ;
  assign n43758 = n43187 & n43632 ;
  assign n43593 = n43196 | n43592 ;
  assign n79568 = ~n43593 ;
  assign n43759 = n43589 & n79568 ;
  assign n79569 = ~n43594 ;
  assign n43760 = n43592 & n79569 ;
  assign n43761 = n43759 | n43760 ;
  assign n43762 = n65845 & n43761 ;
  assign n43763 = n79555 & n43762 ;
  assign n43764 = n43758 | n43763 ;
  assign n43765 = n68214 & n43764 ;
  assign n43766 = n43195 & n43632 ;
  assign n43588 = n43204 | n43587 ;
  assign n79570 = ~n43588 ;
  assign n43767 = n79570 & n43696 ;
  assign n79571 = ~n43697 ;
  assign n43768 = n43587 & n79571 ;
  assign n43769 = n43767 | n43768 ;
  assign n43770 = n65845 & n43769 ;
  assign n43771 = n79555 & n43770 ;
  assign n43772 = n43766 | n43771 ;
  assign n43773 = n68058 & n43772 ;
  assign n43774 = n43203 & n43632 ;
  assign n43581 = n43212 | n43580 ;
  assign n79572 = ~n43581 ;
  assign n43775 = n43577 & n79572 ;
  assign n79573 = ~n43582 ;
  assign n43776 = n43580 & n79573 ;
  assign n43777 = n43775 | n43776 ;
  assign n43778 = n65845 & n43777 ;
  assign n43779 = n79555 & n43778 ;
  assign n43780 = n43774 | n43779 ;
  assign n43781 = n67986 & n43780 ;
  assign n43782 = n43211 & n43632 ;
  assign n43576 = n43220 | n43575 ;
  assign n79574 = ~n43576 ;
  assign n43783 = n79574 & n43692 ;
  assign n79575 = ~n43693 ;
  assign n43784 = n43575 & n79575 ;
  assign n43785 = n43783 | n43784 ;
  assign n43786 = n65845 & n43785 ;
  assign n43787 = n79555 & n43786 ;
  assign n43788 = n43782 | n43787 ;
  assign n43789 = n67763 & n43788 ;
  assign n43790 = n43219 & n43632 ;
  assign n43569 = n43228 | n43568 ;
  assign n79576 = ~n43569 ;
  assign n43791 = n43565 & n79576 ;
  assign n79577 = ~n43570 ;
  assign n43792 = n43568 & n79577 ;
  assign n43793 = n43791 | n43792 ;
  assign n43794 = n65845 & n43793 ;
  assign n43795 = n79555 & n43794 ;
  assign n43796 = n43790 | n43795 ;
  assign n43797 = n67622 & n43796 ;
  assign n43798 = n43227 & n43632 ;
  assign n43564 = n43236 | n43563 ;
  assign n79578 = ~n43564 ;
  assign n43799 = n79578 & n43688 ;
  assign n79579 = ~n43689 ;
  assign n43800 = n43563 & n79579 ;
  assign n43801 = n43799 | n43800 ;
  assign n43802 = n65845 & n43801 ;
  assign n43803 = n79555 & n43802 ;
  assign n43804 = n43798 | n43803 ;
  assign n43805 = n67531 & n43804 ;
  assign n43806 = n43235 & n43632 ;
  assign n43557 = n43244 | n43556 ;
  assign n79580 = ~n43557 ;
  assign n43807 = n43553 & n79580 ;
  assign n79581 = ~n43558 ;
  assign n43808 = n43556 & n79581 ;
  assign n43809 = n43807 | n43808 ;
  assign n43810 = n65845 & n43809 ;
  assign n43811 = n79555 & n43810 ;
  assign n43812 = n43806 | n43811 ;
  assign n43813 = n67348 & n43812 ;
  assign n43814 = n43243 & n43632 ;
  assign n43552 = n43252 | n43551 ;
  assign n79582 = ~n43552 ;
  assign n43815 = n79582 & n43684 ;
  assign n79583 = ~n43685 ;
  assign n43816 = n43551 & n79583 ;
  assign n43817 = n43815 | n43816 ;
  assign n43818 = n65845 & n43817 ;
  assign n43819 = n79555 & n43818 ;
  assign n43820 = n43814 | n43819 ;
  assign n43821 = n67222 & n43820 ;
  assign n43822 = n43251 & n43632 ;
  assign n43545 = n43260 | n43544 ;
  assign n79584 = ~n43545 ;
  assign n43823 = n43541 & n79584 ;
  assign n79585 = ~n43546 ;
  assign n43824 = n43544 & n79585 ;
  assign n43825 = n43823 | n43824 ;
  assign n43826 = n65845 & n43825 ;
  assign n43827 = n79555 & n43826 ;
  assign n43828 = n43822 | n43827 ;
  assign n43829 = n67164 & n43828 ;
  assign n43830 = n43259 & n43632 ;
  assign n43540 = n43268 | n43539 ;
  assign n79586 = ~n43540 ;
  assign n43831 = n79586 & n43680 ;
  assign n79587 = ~n43681 ;
  assign n43832 = n43539 & n79587 ;
  assign n43833 = n43831 | n43832 ;
  assign n43834 = n65845 & n43833 ;
  assign n43835 = n79555 & n43834 ;
  assign n43836 = n43830 | n43835 ;
  assign n43837 = n66979 & n43836 ;
  assign n43838 = n43267 & n43632 ;
  assign n43533 = n43276 | n43532 ;
  assign n79588 = ~n43533 ;
  assign n43839 = n43529 & n79588 ;
  assign n79589 = ~n43534 ;
  assign n43840 = n43532 & n79589 ;
  assign n43841 = n43839 | n43840 ;
  assign n43842 = n65845 & n43841 ;
  assign n43843 = n79555 & n43842 ;
  assign n43844 = n43838 | n43843 ;
  assign n43845 = n66868 & n43844 ;
  assign n43846 = n43275 & n43632 ;
  assign n43528 = n43284 | n43527 ;
  assign n79590 = ~n43528 ;
  assign n43847 = n79590 & n43676 ;
  assign n79591 = ~n43677 ;
  assign n43848 = n43527 & n79591 ;
  assign n43849 = n43847 | n43848 ;
  assign n43850 = n65845 & n43849 ;
  assign n43851 = n79555 & n43850 ;
  assign n43852 = n43846 | n43851 ;
  assign n43853 = n66797 & n43852 ;
  assign n43854 = n43283 & n43632 ;
  assign n43521 = n43292 | n43520 ;
  assign n79592 = ~n43521 ;
  assign n43855 = n43517 & n79592 ;
  assign n79593 = ~n43522 ;
  assign n43856 = n43520 & n79593 ;
  assign n43857 = n43855 | n43856 ;
  assign n43858 = n65845 & n43857 ;
  assign n43859 = n79555 & n43858 ;
  assign n43860 = n43854 | n43859 ;
  assign n43861 = n66654 & n43860 ;
  assign n43862 = n43291 & n43632 ;
  assign n43516 = n43300 | n43515 ;
  assign n79594 = ~n43516 ;
  assign n43863 = n79594 & n43672 ;
  assign n79595 = ~n43673 ;
  assign n43864 = n43515 & n79595 ;
  assign n43865 = n43863 | n43864 ;
  assign n43866 = n65845 & n43865 ;
  assign n43867 = n79555 & n43866 ;
  assign n43868 = n43862 | n43867 ;
  assign n43869 = n66560 & n43868 ;
  assign n43870 = n43299 & n43632 ;
  assign n43509 = n43308 | n43508 ;
  assign n79596 = ~n43509 ;
  assign n43871 = n43505 & n79596 ;
  assign n79597 = ~n43510 ;
  assign n43872 = n43508 & n79597 ;
  assign n43873 = n43871 | n43872 ;
  assign n43874 = n65845 & n43873 ;
  assign n43875 = n79555 & n43874 ;
  assign n43876 = n43870 | n43875 ;
  assign n43877 = n66505 & n43876 ;
  assign n43878 = n43307 & n43632 ;
  assign n43504 = n43316 | n43503 ;
  assign n79598 = ~n43504 ;
  assign n43879 = n79598 & n43668 ;
  assign n79599 = ~n43669 ;
  assign n43880 = n43503 & n79599 ;
  assign n43881 = n43879 | n43880 ;
  assign n43882 = n65845 & n43881 ;
  assign n43883 = n79555 & n43882 ;
  assign n43884 = n43878 | n43883 ;
  assign n43885 = n66379 & n43884 ;
  assign n43886 = n43315 & n43632 ;
  assign n43497 = n43324 | n43496 ;
  assign n79600 = ~n43497 ;
  assign n43887 = n43493 & n79600 ;
  assign n79601 = ~n43498 ;
  assign n43888 = n43496 & n79601 ;
  assign n43889 = n43887 | n43888 ;
  assign n43890 = n65845 & n43889 ;
  assign n43891 = n79555 & n43890 ;
  assign n43892 = n43886 | n43891 ;
  assign n43893 = n66299 & n43892 ;
  assign n43894 = n43323 & n43632 ;
  assign n43492 = n43332 | n43491 ;
  assign n79602 = ~n43492 ;
  assign n43895 = n79602 & n43664 ;
  assign n79603 = ~n43665 ;
  assign n43896 = n43491 & n79603 ;
  assign n43897 = n43895 | n43896 ;
  assign n43898 = n65845 & n43897 ;
  assign n43899 = n79555 & n43898 ;
  assign n43900 = n43894 | n43899 ;
  assign n43901 = n66244 & n43900 ;
  assign n43902 = n43331 & n43632 ;
  assign n43485 = n43340 | n43484 ;
  assign n79604 = ~n43485 ;
  assign n43903 = n43481 & n79604 ;
  assign n79605 = ~n43486 ;
  assign n43904 = n43484 & n79605 ;
  assign n43905 = n43903 | n43904 ;
  assign n43906 = n65845 & n43905 ;
  assign n43907 = n79555 & n43906 ;
  assign n43908 = n43902 | n43907 ;
  assign n43909 = n66145 & n43908 ;
  assign n43910 = n43339 & n43632 ;
  assign n43480 = n43348 | n43479 ;
  assign n79606 = ~n43480 ;
  assign n43911 = n79606 & n43660 ;
  assign n79607 = ~n43661 ;
  assign n43912 = n43479 & n79607 ;
  assign n43913 = n43911 | n43912 ;
  assign n43914 = n65845 & n43913 ;
  assign n43915 = n79555 & n43914 ;
  assign n43916 = n43910 | n43915 ;
  assign n43917 = n66081 & n43916 ;
  assign n43918 = n43347 & n43632 ;
  assign n43473 = n43356 | n43472 ;
  assign n79608 = ~n43473 ;
  assign n43919 = n43469 & n79608 ;
  assign n79609 = ~n43474 ;
  assign n43920 = n43472 & n79609 ;
  assign n43921 = n43919 | n43920 ;
  assign n43922 = n65845 & n43921 ;
  assign n43923 = n79555 & n43922 ;
  assign n43924 = n43918 | n43923 ;
  assign n43925 = n66043 & n43924 ;
  assign n43926 = n43355 & n43632 ;
  assign n43468 = n43364 | n43467 ;
  assign n79610 = ~n43468 ;
  assign n43927 = n79610 & n43656 ;
  assign n79611 = ~n43657 ;
  assign n43928 = n43467 & n79611 ;
  assign n43929 = n43927 | n43928 ;
  assign n43930 = n65845 & n43929 ;
  assign n43931 = n79555 & n43930 ;
  assign n43932 = n43926 | n43931 ;
  assign n43933 = n65960 & n43932 ;
  assign n43934 = n43363 & n43632 ;
  assign n43461 = n43372 | n43460 ;
  assign n79612 = ~n43461 ;
  assign n43935 = n43457 & n79612 ;
  assign n79613 = ~n43462 ;
  assign n43936 = n43460 & n79613 ;
  assign n43937 = n43935 | n43936 ;
  assign n43938 = n65845 & n43937 ;
  assign n43939 = n79555 & n43938 ;
  assign n43940 = n43934 | n43939 ;
  assign n43941 = n65909 & n43940 ;
  assign n43942 = n43371 & n43632 ;
  assign n43456 = n43380 | n43455 ;
  assign n79614 = ~n43456 ;
  assign n43943 = n79614 & n43652 ;
  assign n79615 = ~n43653 ;
  assign n43944 = n43455 & n79615 ;
  assign n43945 = n43943 | n43944 ;
  assign n43946 = n65845 & n43945 ;
  assign n43947 = n79555 & n43946 ;
  assign n43948 = n43942 | n43947 ;
  assign n43949 = n65877 & n43948 ;
  assign n43950 = n43379 & n43632 ;
  assign n43449 = n43389 | n43448 ;
  assign n79616 = ~n43449 ;
  assign n43951 = n43445 & n79616 ;
  assign n79617 = ~n43450 ;
  assign n43952 = n43448 & n79617 ;
  assign n43953 = n43951 | n43952 ;
  assign n43954 = n65845 & n43953 ;
  assign n43955 = n79555 & n43954 ;
  assign n43956 = n43950 | n43955 ;
  assign n43957 = n65820 & n43956 ;
  assign n43958 = n43388 & n43632 ;
  assign n43444 = n43397 | n43443 ;
  assign n79618 = ~n43444 ;
  assign n43959 = n79618 & n43648 ;
  assign n79619 = ~n43649 ;
  assign n43960 = n43443 & n79619 ;
  assign n43961 = n43959 | n43960 ;
  assign n43962 = n65845 & n43961 ;
  assign n43963 = n79555 & n43962 ;
  assign n43964 = n43958 | n43963 ;
  assign n43965 = n65791 & n43964 ;
  assign n43966 = n43396 & n43632 ;
  assign n43967 = n43405 | n43437 ;
  assign n79620 = ~n43967 ;
  assign n43968 = n43434 & n79620 ;
  assign n79621 = ~n43438 ;
  assign n43969 = n43437 & n79621 ;
  assign n43970 = n43968 | n43969 ;
  assign n43971 = n65845 & n43970 ;
  assign n43972 = n79555 & n43971 ;
  assign n43973 = n43966 | n43972 ;
  assign n43974 = n65772 & n43973 ;
  assign n43975 = n43404 & n43632 ;
  assign n43976 = n43413 | n43433 ;
  assign n79622 = ~n43976 ;
  assign n43977 = n43429 & n79622 ;
  assign n79623 = ~n43645 ;
  assign n43978 = n43433 & n79623 ;
  assign n43979 = n43977 | n43978 ;
  assign n43980 = n65845 & n43979 ;
  assign n43981 = n79555 & n43980 ;
  assign n43982 = n43975 | n43981 ;
  assign n43983 = n65746 & n43982 ;
  assign n43984 = n43412 & n43632 ;
  assign n43643 = n43424 | n43427 ;
  assign n79624 = ~n43643 ;
  assign n43985 = n43641 & n79624 ;
  assign n79625 = ~n43428 ;
  assign n43986 = n43427 & n79625 ;
  assign n43987 = n43985 | n43986 ;
  assign n43988 = n65845 & n43987 ;
  assign n43989 = n79555 & n43988 ;
  assign n43990 = n43984 | n43989 ;
  assign n43991 = n65721 & n43990 ;
  assign n43633 = n43415 & n43632 ;
  assign n43422 = n11115 & n43420 ;
  assign n43993 = n43422 & n79552 ;
  assign n43994 = n469 | n43993 ;
  assign n79626 = ~n43994 ;
  assign n43995 = n43641 & n79626 ;
  assign n43996 = n79555 & n43995 ;
  assign n43997 = n43633 | n43996 ;
  assign n43998 = n65686 & n43997 ;
  assign n43992 = n11697 & n79555 ;
  assign n43999 = n11692 & n79555 ;
  assign n79627 = ~n43999 ;
  assign n44000 = x27 & n79627 ;
  assign n44001 = n43992 | n44000 ;
  assign n44002 = n65670 & n44001 ;
  assign n43717 = n79549 & n43716 ;
  assign n44004 = n43628 | n43717 ;
  assign n44005 = n79550 & n44004 ;
  assign n79628 = ~n44005 ;
  assign n44006 = n11692 & n79628 ;
  assign n79629 = ~n44006 ;
  assign n44007 = x27 & n79629 ;
  assign n44008 = n43992 | n44007 ;
  assign n44010 = x65 & n44008 ;
  assign n44009 = x65 | n43992 ;
  assign n44011 = n44000 | n44009 ;
  assign n79630 = ~n44010 ;
  assign n44012 = n79630 & n44011 ;
  assign n44013 = n11708 | n44012 ;
  assign n79631 = ~n44002 ;
  assign n44014 = n79631 & n44013 ;
  assign n79632 = ~n43996 ;
  assign n44015 = x66 & n79632 ;
  assign n79633 = ~n43633 ;
  assign n44016 = n79633 & n44015 ;
  assign n44017 = n43998 | n44016 ;
  assign n44018 = n44014 | n44017 ;
  assign n79634 = ~n43998 ;
  assign n44019 = n79634 & n44018 ;
  assign n79635 = ~n43989 ;
  assign n44020 = x67 & n79635 ;
  assign n79636 = ~n43984 ;
  assign n44021 = n79636 & n44020 ;
  assign n44022 = n44019 | n44021 ;
  assign n79637 = ~n43991 ;
  assign n44023 = n79637 & n44022 ;
  assign n79638 = ~n43981 ;
  assign n44024 = x68 & n79638 ;
  assign n79639 = ~n43975 ;
  assign n44025 = n79639 & n44024 ;
  assign n44026 = n43983 | n44025 ;
  assign n44027 = n44023 | n44026 ;
  assign n79640 = ~n43983 ;
  assign n44028 = n79640 & n44027 ;
  assign n79641 = ~n43972 ;
  assign n44029 = x69 & n79641 ;
  assign n79642 = ~n43966 ;
  assign n44030 = n79642 & n44029 ;
  assign n44031 = n43974 | n44030 ;
  assign n44032 = n44028 | n44031 ;
  assign n79643 = ~n43974 ;
  assign n44033 = n79643 & n44032 ;
  assign n79644 = ~n43963 ;
  assign n44034 = x70 & n79644 ;
  assign n79645 = ~n43958 ;
  assign n44035 = n79645 & n44034 ;
  assign n44036 = n43965 | n44035 ;
  assign n44037 = n44033 | n44036 ;
  assign n79646 = ~n43965 ;
  assign n44038 = n79646 & n44037 ;
  assign n79647 = ~n43955 ;
  assign n44039 = x71 & n79647 ;
  assign n79648 = ~n43950 ;
  assign n44040 = n79648 & n44039 ;
  assign n44041 = n43957 | n44040 ;
  assign n44043 = n44038 | n44041 ;
  assign n79649 = ~n43957 ;
  assign n44044 = n79649 & n44043 ;
  assign n79650 = ~n43947 ;
  assign n44045 = x72 & n79650 ;
  assign n79651 = ~n43942 ;
  assign n44046 = n79651 & n44045 ;
  assign n44047 = n43949 | n44046 ;
  assign n44048 = n44044 | n44047 ;
  assign n79652 = ~n43949 ;
  assign n44049 = n79652 & n44048 ;
  assign n79653 = ~n43939 ;
  assign n44050 = x73 & n79653 ;
  assign n79654 = ~n43934 ;
  assign n44051 = n79654 & n44050 ;
  assign n44052 = n43941 | n44051 ;
  assign n44054 = n44049 | n44052 ;
  assign n79655 = ~n43941 ;
  assign n44055 = n79655 & n44054 ;
  assign n79656 = ~n43931 ;
  assign n44056 = x74 & n79656 ;
  assign n79657 = ~n43926 ;
  assign n44057 = n79657 & n44056 ;
  assign n44058 = n43933 | n44057 ;
  assign n44059 = n44055 | n44058 ;
  assign n79658 = ~n43933 ;
  assign n44060 = n79658 & n44059 ;
  assign n79659 = ~n43923 ;
  assign n44061 = x75 & n79659 ;
  assign n79660 = ~n43918 ;
  assign n44062 = n79660 & n44061 ;
  assign n44063 = n43925 | n44062 ;
  assign n44065 = n44060 | n44063 ;
  assign n79661 = ~n43925 ;
  assign n44066 = n79661 & n44065 ;
  assign n79662 = ~n43915 ;
  assign n44067 = x76 & n79662 ;
  assign n79663 = ~n43910 ;
  assign n44068 = n79663 & n44067 ;
  assign n44069 = n43917 | n44068 ;
  assign n44070 = n44066 | n44069 ;
  assign n79664 = ~n43917 ;
  assign n44071 = n79664 & n44070 ;
  assign n79665 = ~n43907 ;
  assign n44072 = x77 & n79665 ;
  assign n79666 = ~n43902 ;
  assign n44073 = n79666 & n44072 ;
  assign n44074 = n43909 | n44073 ;
  assign n44076 = n44071 | n44074 ;
  assign n79667 = ~n43909 ;
  assign n44077 = n79667 & n44076 ;
  assign n79668 = ~n43899 ;
  assign n44078 = x78 & n79668 ;
  assign n79669 = ~n43894 ;
  assign n44079 = n79669 & n44078 ;
  assign n44080 = n43901 | n44079 ;
  assign n44081 = n44077 | n44080 ;
  assign n79670 = ~n43901 ;
  assign n44082 = n79670 & n44081 ;
  assign n79671 = ~n43891 ;
  assign n44083 = x79 & n79671 ;
  assign n79672 = ~n43886 ;
  assign n44084 = n79672 & n44083 ;
  assign n44085 = n43893 | n44084 ;
  assign n44087 = n44082 | n44085 ;
  assign n79673 = ~n43893 ;
  assign n44088 = n79673 & n44087 ;
  assign n79674 = ~n43883 ;
  assign n44089 = x80 & n79674 ;
  assign n79675 = ~n43878 ;
  assign n44090 = n79675 & n44089 ;
  assign n44091 = n43885 | n44090 ;
  assign n44092 = n44088 | n44091 ;
  assign n79676 = ~n43885 ;
  assign n44093 = n79676 & n44092 ;
  assign n79677 = ~n43875 ;
  assign n44094 = x81 & n79677 ;
  assign n79678 = ~n43870 ;
  assign n44095 = n79678 & n44094 ;
  assign n44096 = n43877 | n44095 ;
  assign n44098 = n44093 | n44096 ;
  assign n79679 = ~n43877 ;
  assign n44099 = n79679 & n44098 ;
  assign n79680 = ~n43867 ;
  assign n44100 = x82 & n79680 ;
  assign n79681 = ~n43862 ;
  assign n44101 = n79681 & n44100 ;
  assign n44102 = n43869 | n44101 ;
  assign n44103 = n44099 | n44102 ;
  assign n79682 = ~n43869 ;
  assign n44104 = n79682 & n44103 ;
  assign n79683 = ~n43859 ;
  assign n44105 = x83 & n79683 ;
  assign n79684 = ~n43854 ;
  assign n44106 = n79684 & n44105 ;
  assign n44107 = n43861 | n44106 ;
  assign n44109 = n44104 | n44107 ;
  assign n79685 = ~n43861 ;
  assign n44110 = n79685 & n44109 ;
  assign n79686 = ~n43851 ;
  assign n44111 = x84 & n79686 ;
  assign n79687 = ~n43846 ;
  assign n44112 = n79687 & n44111 ;
  assign n44113 = n43853 | n44112 ;
  assign n44114 = n44110 | n44113 ;
  assign n79688 = ~n43853 ;
  assign n44115 = n79688 & n44114 ;
  assign n79689 = ~n43843 ;
  assign n44116 = x85 & n79689 ;
  assign n79690 = ~n43838 ;
  assign n44117 = n79690 & n44116 ;
  assign n44118 = n43845 | n44117 ;
  assign n44120 = n44115 | n44118 ;
  assign n79691 = ~n43845 ;
  assign n44121 = n79691 & n44120 ;
  assign n79692 = ~n43835 ;
  assign n44122 = x86 & n79692 ;
  assign n79693 = ~n43830 ;
  assign n44123 = n79693 & n44122 ;
  assign n44124 = n43837 | n44123 ;
  assign n44125 = n44121 | n44124 ;
  assign n79694 = ~n43837 ;
  assign n44126 = n79694 & n44125 ;
  assign n79695 = ~n43827 ;
  assign n44127 = x87 & n79695 ;
  assign n79696 = ~n43822 ;
  assign n44128 = n79696 & n44127 ;
  assign n44129 = n43829 | n44128 ;
  assign n44131 = n44126 | n44129 ;
  assign n79697 = ~n43829 ;
  assign n44132 = n79697 & n44131 ;
  assign n79698 = ~n43819 ;
  assign n44133 = x88 & n79698 ;
  assign n79699 = ~n43814 ;
  assign n44134 = n79699 & n44133 ;
  assign n44135 = n43821 | n44134 ;
  assign n44136 = n44132 | n44135 ;
  assign n79700 = ~n43821 ;
  assign n44137 = n79700 & n44136 ;
  assign n79701 = ~n43811 ;
  assign n44138 = x89 & n79701 ;
  assign n79702 = ~n43806 ;
  assign n44139 = n79702 & n44138 ;
  assign n44140 = n43813 | n44139 ;
  assign n44142 = n44137 | n44140 ;
  assign n79703 = ~n43813 ;
  assign n44143 = n79703 & n44142 ;
  assign n79704 = ~n43803 ;
  assign n44144 = x90 & n79704 ;
  assign n79705 = ~n43798 ;
  assign n44145 = n79705 & n44144 ;
  assign n44146 = n43805 | n44145 ;
  assign n44147 = n44143 | n44146 ;
  assign n79706 = ~n43805 ;
  assign n44148 = n79706 & n44147 ;
  assign n79707 = ~n43795 ;
  assign n44149 = x91 & n79707 ;
  assign n79708 = ~n43790 ;
  assign n44150 = n79708 & n44149 ;
  assign n44151 = n43797 | n44150 ;
  assign n44153 = n44148 | n44151 ;
  assign n79709 = ~n43797 ;
  assign n44154 = n79709 & n44153 ;
  assign n79710 = ~n43787 ;
  assign n44155 = x92 & n79710 ;
  assign n79711 = ~n43782 ;
  assign n44156 = n79711 & n44155 ;
  assign n44157 = n43789 | n44156 ;
  assign n44158 = n44154 | n44157 ;
  assign n79712 = ~n43789 ;
  assign n44159 = n79712 & n44158 ;
  assign n79713 = ~n43779 ;
  assign n44160 = x93 & n79713 ;
  assign n79714 = ~n43774 ;
  assign n44161 = n79714 & n44160 ;
  assign n44162 = n43781 | n44161 ;
  assign n44164 = n44159 | n44162 ;
  assign n79715 = ~n43781 ;
  assign n44165 = n79715 & n44164 ;
  assign n79716 = ~n43771 ;
  assign n44166 = x94 & n79716 ;
  assign n79717 = ~n43766 ;
  assign n44167 = n79717 & n44166 ;
  assign n44168 = n43773 | n44167 ;
  assign n44169 = n44165 | n44168 ;
  assign n79718 = ~n43773 ;
  assign n44170 = n79718 & n44169 ;
  assign n79719 = ~n43763 ;
  assign n44171 = x95 & n79719 ;
  assign n79720 = ~n43758 ;
  assign n44172 = n79720 & n44171 ;
  assign n44173 = n43765 | n44172 ;
  assign n44175 = n44170 | n44173 ;
  assign n79721 = ~n43765 ;
  assign n44176 = n79721 & n44175 ;
  assign n79722 = ~n43755 ;
  assign n44177 = x96 & n79722 ;
  assign n79723 = ~n43750 ;
  assign n44178 = n79723 & n44177 ;
  assign n44179 = n43757 | n44178 ;
  assign n44180 = n44176 | n44179 ;
  assign n79724 = ~n43757 ;
  assign n44181 = n79724 & n44180 ;
  assign n79725 = ~n43747 ;
  assign n44182 = x97 & n79725 ;
  assign n79726 = ~n43742 ;
  assign n44183 = n79726 & n44182 ;
  assign n44184 = n43749 | n44183 ;
  assign n44186 = n44181 | n44184 ;
  assign n79727 = ~n43749 ;
  assign n44187 = n79727 & n44186 ;
  assign n79728 = ~n43739 ;
  assign n44188 = x98 & n79728 ;
  assign n79729 = ~n43734 ;
  assign n44189 = n79729 & n44188 ;
  assign n44190 = n43741 | n44189 ;
  assign n44191 = n44187 | n44190 ;
  assign n79730 = ~n43741 ;
  assign n44192 = n79730 & n44191 ;
  assign n79731 = ~n43731 ;
  assign n44193 = x99 & n79731 ;
  assign n79732 = ~n43726 ;
  assign n44194 = n79732 & n44193 ;
  assign n44195 = n43733 | n44194 ;
  assign n44197 = n44192 | n44195 ;
  assign n79733 = ~n43733 ;
  assign n44198 = n79733 & n44197 ;
  assign n79734 = ~n43714 ;
  assign n44199 = x100 & n79734 ;
  assign n79735 = ~n43635 ;
  assign n44200 = n79735 & n44199 ;
  assign n44201 = n43725 | n44200 ;
  assign n44202 = n44198 | n44201 ;
  assign n79736 = ~n43725 ;
  assign n44203 = n79736 & n44202 ;
  assign n79737 = ~n43632 ;
  assign n44204 = n79737 & n43721 ;
  assign n44205 = n43146 & n43632 ;
  assign n79738 = ~n44205 ;
  assign n44206 = x101 & n79738 ;
  assign n79739 = ~n44204 ;
  assign n44207 = n79739 & n44206 ;
  assign n44208 = n43724 | n44207 ;
  assign n44210 = n44203 | n44208 ;
  assign n79740 = ~n43724 ;
  assign n44211 = n79740 & n44210 ;
  assign n44212 = n11929 | n44211 ;
  assign n44213 = n43715 & n44212 ;
  assign n44215 = n65670 & n44008 ;
  assign n44003 = x65 & n44001 ;
  assign n79741 = ~n44003 ;
  assign n44214 = n79741 & n44011 ;
  assign n44216 = n11708 | n44214 ;
  assign n79742 = ~n44215 ;
  assign n44217 = n79742 & n44216 ;
  assign n44218 = n44017 | n44217 ;
  assign n44219 = n79634 & n44218 ;
  assign n44220 = n43991 | n44021 ;
  assign n44222 = n44219 | n44220 ;
  assign n44223 = n79637 & n44222 ;
  assign n44225 = n44026 | n44223 ;
  assign n44226 = n79640 & n44225 ;
  assign n44228 = n44031 | n44226 ;
  assign n44229 = n79643 & n44228 ;
  assign n44230 = n44036 | n44229 ;
  assign n44232 = n79646 & n44230 ;
  assign n44233 = n44041 | n44232 ;
  assign n44234 = n79649 & n44233 ;
  assign n44235 = n44047 | n44234 ;
  assign n44237 = n79652 & n44235 ;
  assign n44238 = n44052 | n44237 ;
  assign n44239 = n79655 & n44238 ;
  assign n44240 = n44058 | n44239 ;
  assign n44242 = n79658 & n44240 ;
  assign n44243 = n44063 | n44242 ;
  assign n44244 = n79661 & n44243 ;
  assign n44245 = n44069 | n44244 ;
  assign n44247 = n79664 & n44245 ;
  assign n44248 = n44074 | n44247 ;
  assign n44249 = n79667 & n44248 ;
  assign n44250 = n44080 | n44249 ;
  assign n44252 = n79670 & n44250 ;
  assign n44253 = n44085 | n44252 ;
  assign n44254 = n79673 & n44253 ;
  assign n44255 = n44091 | n44254 ;
  assign n44257 = n79676 & n44255 ;
  assign n44258 = n44096 | n44257 ;
  assign n44259 = n79679 & n44258 ;
  assign n44260 = n44102 | n44259 ;
  assign n44262 = n79682 & n44260 ;
  assign n44263 = n44107 | n44262 ;
  assign n44264 = n79685 & n44263 ;
  assign n44265 = n44113 | n44264 ;
  assign n44267 = n79688 & n44265 ;
  assign n44268 = n44118 | n44267 ;
  assign n44269 = n79691 & n44268 ;
  assign n44270 = n44124 | n44269 ;
  assign n44272 = n79694 & n44270 ;
  assign n44273 = n44129 | n44272 ;
  assign n44274 = n79697 & n44273 ;
  assign n44275 = n44135 | n44274 ;
  assign n44277 = n79700 & n44275 ;
  assign n44278 = n44140 | n44277 ;
  assign n44279 = n79703 & n44278 ;
  assign n44280 = n44146 | n44279 ;
  assign n44282 = n79706 & n44280 ;
  assign n44283 = n44151 | n44282 ;
  assign n44284 = n79709 & n44283 ;
  assign n44285 = n44157 | n44284 ;
  assign n44287 = n79712 & n44285 ;
  assign n44288 = n44162 | n44287 ;
  assign n44289 = n79715 & n44288 ;
  assign n44290 = n44168 | n44289 ;
  assign n44292 = n79718 & n44290 ;
  assign n44293 = n44173 | n44292 ;
  assign n44294 = n79721 & n44293 ;
  assign n44295 = n44179 | n44294 ;
  assign n44297 = n79724 & n44295 ;
  assign n44298 = n44184 | n44297 ;
  assign n44299 = n79727 & n44298 ;
  assign n44300 = n44190 | n44299 ;
  assign n44302 = n79730 & n44300 ;
  assign n44303 = n44195 | n44302 ;
  assign n44304 = n79733 & n44303 ;
  assign n79743 = ~n44304 ;
  assign n44305 = n44201 & n79743 ;
  assign n44307 = n43733 | n44201 ;
  assign n79744 = ~n44307 ;
  assign n44308 = n44197 & n79744 ;
  assign n44309 = n44305 | n44308 ;
  assign n44310 = n69455 & n44309 ;
  assign n79745 = ~n44211 ;
  assign n44311 = n79745 & n44310 ;
  assign n44312 = n44213 | n44311 ;
  assign n44313 = n69261 & n44312 ;
  assign n79746 = ~n44311 ;
  assign n44792 = x101 & n79746 ;
  assign n79747 = ~n44213 ;
  assign n44793 = n79747 & n44792 ;
  assign n44794 = n44313 | n44793 ;
  assign n44314 = n43732 & n44212 ;
  assign n79748 = ~n44192 ;
  assign n44196 = n79748 & n44195 ;
  assign n44315 = n43741 | n44195 ;
  assign n79749 = ~n44315 ;
  assign n44316 = n44300 & n79749 ;
  assign n44317 = n44196 | n44316 ;
  assign n44318 = n69455 & n44317 ;
  assign n44319 = n79745 & n44318 ;
  assign n44320 = n44314 | n44319 ;
  assign n44321 = n69075 & n44320 ;
  assign n44322 = n43740 & n44212 ;
  assign n79750 = ~n44299 ;
  assign n44301 = n44190 & n79750 ;
  assign n44323 = n43749 | n44190 ;
  assign n79751 = ~n44323 ;
  assign n44324 = n44186 & n79751 ;
  assign n44325 = n44301 | n44324 ;
  assign n44326 = n69455 & n44325 ;
  assign n44327 = n79745 & n44326 ;
  assign n44328 = n44322 | n44327 ;
  assign n44329 = n68993 & n44328 ;
  assign n79752 = ~n44327 ;
  assign n44781 = x99 & n79752 ;
  assign n79753 = ~n44322 ;
  assign n44782 = n79753 & n44781 ;
  assign n44783 = n44329 | n44782 ;
  assign n44330 = n43748 & n44212 ;
  assign n79754 = ~n44181 ;
  assign n44185 = n79754 & n44184 ;
  assign n44331 = n43757 | n44184 ;
  assign n79755 = ~n44331 ;
  assign n44332 = n44295 & n79755 ;
  assign n44333 = n44185 | n44332 ;
  assign n44334 = n69455 & n44333 ;
  assign n44335 = n79745 & n44334 ;
  assign n44336 = n44330 | n44335 ;
  assign n44337 = n68716 & n44336 ;
  assign n44338 = n43756 & n44212 ;
  assign n79756 = ~n44294 ;
  assign n44296 = n44179 & n79756 ;
  assign n44339 = n43765 | n44179 ;
  assign n79757 = ~n44339 ;
  assign n44340 = n44175 & n79757 ;
  assign n44341 = n44296 | n44340 ;
  assign n44342 = n69455 & n44341 ;
  assign n44343 = n79745 & n44342 ;
  assign n44344 = n44338 | n44343 ;
  assign n44345 = n68545 & n44344 ;
  assign n79758 = ~n44343 ;
  assign n44771 = x97 & n79758 ;
  assign n79759 = ~n44338 ;
  assign n44772 = n79759 & n44771 ;
  assign n44773 = n44345 | n44772 ;
  assign n44346 = n43764 & n44212 ;
  assign n79760 = ~n44170 ;
  assign n44174 = n79760 & n44173 ;
  assign n44347 = n43773 | n44173 ;
  assign n79761 = ~n44347 ;
  assign n44348 = n44290 & n79761 ;
  assign n44349 = n44174 | n44348 ;
  assign n44350 = n69455 & n44349 ;
  assign n44351 = n79745 & n44350 ;
  assign n44352 = n44346 | n44351 ;
  assign n44353 = n68438 & n44352 ;
  assign n44354 = n43772 & n44212 ;
  assign n79762 = ~n44289 ;
  assign n44291 = n44168 & n79762 ;
  assign n44355 = n43781 | n44168 ;
  assign n79763 = ~n44355 ;
  assign n44356 = n44164 & n79763 ;
  assign n44357 = n44291 | n44356 ;
  assign n44358 = n69455 & n44357 ;
  assign n44359 = n79745 & n44358 ;
  assign n44360 = n44354 | n44359 ;
  assign n44361 = n68214 & n44360 ;
  assign n79764 = ~n44359 ;
  assign n44761 = x95 & n79764 ;
  assign n79765 = ~n44354 ;
  assign n44762 = n79765 & n44761 ;
  assign n44763 = n44361 | n44762 ;
  assign n44362 = n43780 & n44212 ;
  assign n79766 = ~n44159 ;
  assign n44163 = n79766 & n44162 ;
  assign n44363 = n43789 | n44162 ;
  assign n79767 = ~n44363 ;
  assign n44364 = n44285 & n79767 ;
  assign n44365 = n44163 | n44364 ;
  assign n44366 = n69455 & n44365 ;
  assign n44367 = n79745 & n44366 ;
  assign n44368 = n44362 | n44367 ;
  assign n44369 = n68058 & n44368 ;
  assign n44370 = n43788 & n44212 ;
  assign n79768 = ~n44284 ;
  assign n44286 = n44157 & n79768 ;
  assign n44371 = n43797 | n44157 ;
  assign n79769 = ~n44371 ;
  assign n44372 = n44153 & n79769 ;
  assign n44373 = n44286 | n44372 ;
  assign n44374 = n69455 & n44373 ;
  assign n44375 = n79745 & n44374 ;
  assign n44376 = n44370 | n44375 ;
  assign n44377 = n67986 & n44376 ;
  assign n79770 = ~n44375 ;
  assign n44751 = x93 & n79770 ;
  assign n79771 = ~n44370 ;
  assign n44752 = n79771 & n44751 ;
  assign n44753 = n44377 | n44752 ;
  assign n44378 = n43796 & n44212 ;
  assign n79772 = ~n44148 ;
  assign n44152 = n79772 & n44151 ;
  assign n44379 = n43805 | n44151 ;
  assign n79773 = ~n44379 ;
  assign n44380 = n44280 & n79773 ;
  assign n44381 = n44152 | n44380 ;
  assign n44382 = n69455 & n44381 ;
  assign n44383 = n79745 & n44382 ;
  assign n44384 = n44378 | n44383 ;
  assign n44385 = n67763 & n44384 ;
  assign n44386 = n43804 & n44212 ;
  assign n79774 = ~n44279 ;
  assign n44281 = n44146 & n79774 ;
  assign n44387 = n43813 | n44146 ;
  assign n79775 = ~n44387 ;
  assign n44388 = n44142 & n79775 ;
  assign n44389 = n44281 | n44388 ;
  assign n44390 = n69455 & n44389 ;
  assign n44391 = n79745 & n44390 ;
  assign n44392 = n44386 | n44391 ;
  assign n44393 = n67622 & n44392 ;
  assign n79776 = ~n44391 ;
  assign n44740 = x91 & n79776 ;
  assign n79777 = ~n44386 ;
  assign n44741 = n79777 & n44740 ;
  assign n44742 = n44393 | n44741 ;
  assign n44394 = n43812 & n44212 ;
  assign n79778 = ~n44137 ;
  assign n44141 = n79778 & n44140 ;
  assign n44395 = n43821 | n44140 ;
  assign n79779 = ~n44395 ;
  assign n44396 = n44275 & n79779 ;
  assign n44397 = n44141 | n44396 ;
  assign n44398 = n69455 & n44397 ;
  assign n44399 = n79745 & n44398 ;
  assign n44400 = n44394 | n44399 ;
  assign n44401 = n67531 & n44400 ;
  assign n44402 = n43820 & n44212 ;
  assign n79780 = ~n44274 ;
  assign n44276 = n44135 & n79780 ;
  assign n44403 = n43829 | n44135 ;
  assign n79781 = ~n44403 ;
  assign n44404 = n44131 & n79781 ;
  assign n44405 = n44276 | n44404 ;
  assign n44406 = n69455 & n44405 ;
  assign n44407 = n79745 & n44406 ;
  assign n44408 = n44402 | n44407 ;
  assign n44409 = n67348 & n44408 ;
  assign n79782 = ~n44407 ;
  assign n44729 = x89 & n79782 ;
  assign n79783 = ~n44402 ;
  assign n44730 = n79783 & n44729 ;
  assign n44731 = n44409 | n44730 ;
  assign n44410 = n43828 & n44212 ;
  assign n79784 = ~n44126 ;
  assign n44130 = n79784 & n44129 ;
  assign n44411 = n43837 | n44129 ;
  assign n79785 = ~n44411 ;
  assign n44412 = n44270 & n79785 ;
  assign n44413 = n44130 | n44412 ;
  assign n44414 = n69455 & n44413 ;
  assign n44415 = n79745 & n44414 ;
  assign n44416 = n44410 | n44415 ;
  assign n44417 = n67222 & n44416 ;
  assign n44418 = n43836 & n44212 ;
  assign n79786 = ~n44269 ;
  assign n44271 = n44124 & n79786 ;
  assign n44419 = n43845 | n44124 ;
  assign n79787 = ~n44419 ;
  assign n44420 = n44120 & n79787 ;
  assign n44421 = n44271 | n44420 ;
  assign n44422 = n69455 & n44421 ;
  assign n44423 = n79745 & n44422 ;
  assign n44424 = n44418 | n44423 ;
  assign n44425 = n67164 & n44424 ;
  assign n79788 = ~n44423 ;
  assign n44718 = x87 & n79788 ;
  assign n79789 = ~n44418 ;
  assign n44719 = n79789 & n44718 ;
  assign n44720 = n44425 | n44719 ;
  assign n44426 = n43844 & n44212 ;
  assign n79790 = ~n44115 ;
  assign n44119 = n79790 & n44118 ;
  assign n44427 = n43853 | n44118 ;
  assign n79791 = ~n44427 ;
  assign n44428 = n44265 & n79791 ;
  assign n44429 = n44119 | n44428 ;
  assign n44430 = n69455 & n44429 ;
  assign n44431 = n79745 & n44430 ;
  assign n44432 = n44426 | n44431 ;
  assign n44433 = n66979 & n44432 ;
  assign n44434 = n43852 & n44212 ;
  assign n79792 = ~n44264 ;
  assign n44266 = n44113 & n79792 ;
  assign n44435 = n43861 | n44113 ;
  assign n79793 = ~n44435 ;
  assign n44436 = n44109 & n79793 ;
  assign n44437 = n44266 | n44436 ;
  assign n44438 = n69455 & n44437 ;
  assign n44439 = n79745 & n44438 ;
  assign n44440 = n44434 | n44439 ;
  assign n44441 = n66868 & n44440 ;
  assign n79794 = ~n44439 ;
  assign n44708 = x85 & n79794 ;
  assign n79795 = ~n44434 ;
  assign n44709 = n79795 & n44708 ;
  assign n44710 = n44441 | n44709 ;
  assign n44442 = n43860 & n44212 ;
  assign n79796 = ~n44104 ;
  assign n44108 = n79796 & n44107 ;
  assign n44443 = n43869 | n44107 ;
  assign n79797 = ~n44443 ;
  assign n44444 = n44260 & n79797 ;
  assign n44445 = n44108 | n44444 ;
  assign n44446 = n69455 & n44445 ;
  assign n44447 = n79745 & n44446 ;
  assign n44448 = n44442 | n44447 ;
  assign n44449 = n66797 & n44448 ;
  assign n44450 = n43868 & n44212 ;
  assign n79798 = ~n44259 ;
  assign n44261 = n44102 & n79798 ;
  assign n44451 = n43877 | n44102 ;
  assign n79799 = ~n44451 ;
  assign n44452 = n44098 & n79799 ;
  assign n44453 = n44261 | n44452 ;
  assign n44454 = n69455 & n44453 ;
  assign n44455 = n79745 & n44454 ;
  assign n44456 = n44450 | n44455 ;
  assign n44457 = n66654 & n44456 ;
  assign n79800 = ~n44455 ;
  assign n44698 = x83 & n79800 ;
  assign n79801 = ~n44450 ;
  assign n44699 = n79801 & n44698 ;
  assign n44700 = n44457 | n44699 ;
  assign n44458 = n43876 & n44212 ;
  assign n79802 = ~n44093 ;
  assign n44097 = n79802 & n44096 ;
  assign n44459 = n43885 | n44096 ;
  assign n79803 = ~n44459 ;
  assign n44460 = n44255 & n79803 ;
  assign n44461 = n44097 | n44460 ;
  assign n44462 = n69455 & n44461 ;
  assign n44463 = n79745 & n44462 ;
  assign n44464 = n44458 | n44463 ;
  assign n44465 = n66560 & n44464 ;
  assign n44466 = n43884 & n44212 ;
  assign n79804 = ~n44254 ;
  assign n44256 = n44091 & n79804 ;
  assign n44467 = n43893 | n44091 ;
  assign n79805 = ~n44467 ;
  assign n44468 = n44087 & n79805 ;
  assign n44469 = n44256 | n44468 ;
  assign n44470 = n69455 & n44469 ;
  assign n44471 = n79745 & n44470 ;
  assign n44472 = n44466 | n44471 ;
  assign n44473 = n66505 & n44472 ;
  assign n79806 = ~n44471 ;
  assign n44688 = x81 & n79806 ;
  assign n79807 = ~n44466 ;
  assign n44689 = n79807 & n44688 ;
  assign n44690 = n44473 | n44689 ;
  assign n44474 = n43892 & n44212 ;
  assign n79808 = ~n44082 ;
  assign n44086 = n79808 & n44085 ;
  assign n44475 = n43901 | n44085 ;
  assign n79809 = ~n44475 ;
  assign n44476 = n44250 & n79809 ;
  assign n44477 = n44086 | n44476 ;
  assign n44478 = n69455 & n44477 ;
  assign n44479 = n79745 & n44478 ;
  assign n44480 = n44474 | n44479 ;
  assign n44481 = n66379 & n44480 ;
  assign n44482 = n43900 & n44212 ;
  assign n79810 = ~n44249 ;
  assign n44251 = n44080 & n79810 ;
  assign n44483 = n43909 | n44080 ;
  assign n79811 = ~n44483 ;
  assign n44484 = n44076 & n79811 ;
  assign n44485 = n44251 | n44484 ;
  assign n44486 = n69455 & n44485 ;
  assign n44487 = n79745 & n44486 ;
  assign n44488 = n44482 | n44487 ;
  assign n44489 = n66299 & n44488 ;
  assign n79812 = ~n44487 ;
  assign n44678 = x79 & n79812 ;
  assign n79813 = ~n44482 ;
  assign n44679 = n79813 & n44678 ;
  assign n44680 = n44489 | n44679 ;
  assign n44490 = n43908 & n44212 ;
  assign n79814 = ~n44071 ;
  assign n44075 = n79814 & n44074 ;
  assign n44491 = n43917 | n44074 ;
  assign n79815 = ~n44491 ;
  assign n44492 = n44245 & n79815 ;
  assign n44493 = n44075 | n44492 ;
  assign n44494 = n69455 & n44493 ;
  assign n44495 = n79745 & n44494 ;
  assign n44496 = n44490 | n44495 ;
  assign n44497 = n66244 & n44496 ;
  assign n44498 = n43916 & n44212 ;
  assign n79816 = ~n44244 ;
  assign n44246 = n44069 & n79816 ;
  assign n44499 = n43925 | n44069 ;
  assign n79817 = ~n44499 ;
  assign n44500 = n44065 & n79817 ;
  assign n44501 = n44246 | n44500 ;
  assign n44502 = n69455 & n44501 ;
  assign n44503 = n79745 & n44502 ;
  assign n44504 = n44498 | n44503 ;
  assign n44505 = n66145 & n44504 ;
  assign n79818 = ~n44503 ;
  assign n44667 = x77 & n79818 ;
  assign n79819 = ~n44498 ;
  assign n44668 = n79819 & n44667 ;
  assign n44669 = n44505 | n44668 ;
  assign n44506 = n43924 & n44212 ;
  assign n79820 = ~n44060 ;
  assign n44064 = n79820 & n44063 ;
  assign n44507 = n43933 | n44063 ;
  assign n79821 = ~n44507 ;
  assign n44508 = n44240 & n79821 ;
  assign n44509 = n44064 | n44508 ;
  assign n44510 = n69455 & n44509 ;
  assign n44511 = n79745 & n44510 ;
  assign n44512 = n44506 | n44511 ;
  assign n44513 = n66081 & n44512 ;
  assign n44514 = n43932 & n44212 ;
  assign n79822 = ~n44239 ;
  assign n44241 = n44058 & n79822 ;
  assign n44515 = n43941 | n44058 ;
  assign n79823 = ~n44515 ;
  assign n44516 = n44054 & n79823 ;
  assign n44517 = n44241 | n44516 ;
  assign n44518 = n69455 & n44517 ;
  assign n44519 = n79745 & n44518 ;
  assign n44520 = n44514 | n44519 ;
  assign n44521 = n66043 & n44520 ;
  assign n79824 = ~n44519 ;
  assign n44657 = x75 & n79824 ;
  assign n79825 = ~n44514 ;
  assign n44658 = n79825 & n44657 ;
  assign n44659 = n44521 | n44658 ;
  assign n44522 = n43940 & n44212 ;
  assign n79826 = ~n44049 ;
  assign n44053 = n79826 & n44052 ;
  assign n44523 = n43949 | n44052 ;
  assign n79827 = ~n44523 ;
  assign n44524 = n44235 & n79827 ;
  assign n44525 = n44053 | n44524 ;
  assign n44526 = n69455 & n44525 ;
  assign n44527 = n79745 & n44526 ;
  assign n44528 = n44522 | n44527 ;
  assign n44529 = n65960 & n44528 ;
  assign n44530 = n43948 & n44212 ;
  assign n79828 = ~n44234 ;
  assign n44236 = n44047 & n79828 ;
  assign n44531 = n43957 | n44047 ;
  assign n79829 = ~n44531 ;
  assign n44532 = n44043 & n79829 ;
  assign n44533 = n44236 | n44532 ;
  assign n44534 = n69455 & n44533 ;
  assign n44535 = n79745 & n44534 ;
  assign n44536 = n44530 | n44535 ;
  assign n44537 = n65909 & n44536 ;
  assign n79830 = ~n44535 ;
  assign n44647 = x73 & n79830 ;
  assign n79831 = ~n44530 ;
  assign n44648 = n79831 & n44647 ;
  assign n44649 = n44537 | n44648 ;
  assign n44538 = n43956 & n44212 ;
  assign n79832 = ~n44038 ;
  assign n44042 = n79832 & n44041 ;
  assign n44539 = n43965 | n44041 ;
  assign n79833 = ~n44539 ;
  assign n44540 = n44230 & n79833 ;
  assign n44541 = n44042 | n44540 ;
  assign n44542 = n69455 & n44541 ;
  assign n44543 = n79745 & n44542 ;
  assign n44544 = n44538 | n44543 ;
  assign n44545 = n65877 & n44544 ;
  assign n44546 = n43964 & n44212 ;
  assign n79834 = ~n44229 ;
  assign n44231 = n44036 & n79834 ;
  assign n44547 = n43974 | n44036 ;
  assign n79835 = ~n44547 ;
  assign n44548 = n44032 & n79835 ;
  assign n44549 = n44231 | n44548 ;
  assign n44550 = n69455 & n44549 ;
  assign n44551 = n79745 & n44550 ;
  assign n44552 = n44546 | n44551 ;
  assign n44553 = n65820 & n44552 ;
  assign n79836 = ~n44551 ;
  assign n44637 = x71 & n79836 ;
  assign n79837 = ~n44546 ;
  assign n44638 = n79837 & n44637 ;
  assign n44639 = n44553 | n44638 ;
  assign n44554 = n43973 & n44212 ;
  assign n79838 = ~n44028 ;
  assign n44227 = n79838 & n44031 ;
  assign n44555 = n43983 | n44031 ;
  assign n79839 = ~n44555 ;
  assign n44556 = n44027 & n79839 ;
  assign n44557 = n44227 | n44556 ;
  assign n44558 = n69455 & n44557 ;
  assign n44559 = n79745 & n44558 ;
  assign n44560 = n44554 | n44559 ;
  assign n44561 = n65791 & n44560 ;
  assign n44562 = n43982 & n44212 ;
  assign n79840 = ~n44223 ;
  assign n44224 = n44026 & n79840 ;
  assign n44563 = n44019 | n44220 ;
  assign n44564 = n43991 | n44026 ;
  assign n79841 = ~n44564 ;
  assign n44565 = n44563 & n79841 ;
  assign n44566 = n44224 | n44565 ;
  assign n44567 = n69455 & n44566 ;
  assign n44568 = n79745 & n44567 ;
  assign n44569 = n44562 | n44568 ;
  assign n44570 = n65772 & n44569 ;
  assign n79842 = ~n44568 ;
  assign n44627 = x69 & n79842 ;
  assign n79843 = ~n44562 ;
  assign n44628 = n79843 & n44627 ;
  assign n44629 = n44570 | n44628 ;
  assign n44571 = n43990 & n44212 ;
  assign n79844 = ~n44019 ;
  assign n44221 = n79844 & n44220 ;
  assign n44572 = n43998 | n44220 ;
  assign n79845 = ~n44572 ;
  assign n44573 = n44018 & n79845 ;
  assign n44574 = n44221 | n44573 ;
  assign n44575 = n69455 & n44574 ;
  assign n44576 = n79745 & n44575 ;
  assign n44577 = n44571 | n44576 ;
  assign n44578 = n65746 & n44577 ;
  assign n44579 = n43997 & n44212 ;
  assign n44580 = n44017 | n44215 ;
  assign n79846 = ~n44580 ;
  assign n44581 = n44216 & n79846 ;
  assign n79847 = ~n44217 ;
  assign n44582 = n44017 & n79847 ;
  assign n44583 = n44581 | n44582 ;
  assign n44584 = n69455 & n44583 ;
  assign n44585 = n79745 & n44584 ;
  assign n44586 = n44579 | n44585 ;
  assign n44588 = n65721 & n44586 ;
  assign n79848 = ~n44585 ;
  assign n44587 = x67 & n79848 ;
  assign n79849 = ~n44579 ;
  assign n44618 = n79849 & n44587 ;
  assign n44619 = n44588 | n44618 ;
  assign n44589 = n44001 & n44212 ;
  assign n44590 = n11708 & n44011 ;
  assign n44591 = n79630 & n44590 ;
  assign n44592 = n11929 | n44591 ;
  assign n79850 = ~n44592 ;
  assign n44593 = n44216 & n79850 ;
  assign n44594 = n79745 & n44593 ;
  assign n44595 = n44589 | n44594 ;
  assign n44596 = n65686 & n44595 ;
  assign n44597 = n12300 & n79745 ;
  assign n79851 = ~n44597 ;
  assign n44598 = x26 & n79851 ;
  assign n44599 = n12312 & n79745 ;
  assign n44600 = n44598 | n44599 ;
  assign n44601 = x65 & n44600 ;
  assign n44306 = n44201 | n44304 ;
  assign n44602 = n79736 & n44306 ;
  assign n44603 = n44208 | n44602 ;
  assign n44604 = n79740 & n44603 ;
  assign n79852 = ~n44604 ;
  assign n44605 = n12300 & n79852 ;
  assign n79853 = ~n44605 ;
  assign n44606 = x26 & n79853 ;
  assign n44607 = x65 | n44599 ;
  assign n44608 = n44606 | n44607 ;
  assign n79854 = ~n44601 ;
  assign n44609 = n79854 & n44608 ;
  assign n44610 = n12319 | n44609 ;
  assign n44611 = n44599 | n44606 ;
  assign n44612 = n65670 & n44611 ;
  assign n79855 = ~n44612 ;
  assign n44613 = n44610 & n79855 ;
  assign n79856 = ~n44594 ;
  assign n44614 = x66 & n79856 ;
  assign n79857 = ~n44589 ;
  assign n44615 = n79857 & n44614 ;
  assign n44616 = n44596 | n44615 ;
  assign n44617 = n44613 | n44616 ;
  assign n79858 = ~n44596 ;
  assign n44620 = n79858 & n44617 ;
  assign n44621 = n44619 | n44620 ;
  assign n79859 = ~n44588 ;
  assign n44622 = n79859 & n44621 ;
  assign n79860 = ~n44576 ;
  assign n44623 = x68 & n79860 ;
  assign n79861 = ~n44571 ;
  assign n44624 = n79861 & n44623 ;
  assign n44625 = n44578 | n44624 ;
  assign n44626 = n44622 | n44625 ;
  assign n79862 = ~n44578 ;
  assign n44630 = n79862 & n44626 ;
  assign n44631 = n44629 | n44630 ;
  assign n79863 = ~n44570 ;
  assign n44632 = n79863 & n44631 ;
  assign n79864 = ~n44559 ;
  assign n44633 = x70 & n79864 ;
  assign n79865 = ~n44554 ;
  assign n44634 = n79865 & n44633 ;
  assign n44635 = n44561 | n44634 ;
  assign n44636 = n44632 | n44635 ;
  assign n79866 = ~n44561 ;
  assign n44640 = n79866 & n44636 ;
  assign n44641 = n44639 | n44640 ;
  assign n79867 = ~n44553 ;
  assign n44642 = n79867 & n44641 ;
  assign n79868 = ~n44543 ;
  assign n44643 = x72 & n79868 ;
  assign n79869 = ~n44538 ;
  assign n44644 = n79869 & n44643 ;
  assign n44645 = n44545 | n44644 ;
  assign n44646 = n44642 | n44645 ;
  assign n79870 = ~n44545 ;
  assign n44650 = n79870 & n44646 ;
  assign n44651 = n44649 | n44650 ;
  assign n79871 = ~n44537 ;
  assign n44652 = n79871 & n44651 ;
  assign n79872 = ~n44527 ;
  assign n44653 = x74 & n79872 ;
  assign n79873 = ~n44522 ;
  assign n44654 = n79873 & n44653 ;
  assign n44655 = n44529 | n44654 ;
  assign n44656 = n44652 | n44655 ;
  assign n79874 = ~n44529 ;
  assign n44660 = n79874 & n44656 ;
  assign n44661 = n44659 | n44660 ;
  assign n79875 = ~n44521 ;
  assign n44662 = n79875 & n44661 ;
  assign n79876 = ~n44511 ;
  assign n44663 = x76 & n79876 ;
  assign n79877 = ~n44506 ;
  assign n44664 = n79877 & n44663 ;
  assign n44665 = n44513 | n44664 ;
  assign n44666 = n44662 | n44665 ;
  assign n79878 = ~n44513 ;
  assign n44671 = n79878 & n44666 ;
  assign n44672 = n44669 | n44671 ;
  assign n79879 = ~n44505 ;
  assign n44673 = n79879 & n44672 ;
  assign n79880 = ~n44495 ;
  assign n44674 = x78 & n79880 ;
  assign n79881 = ~n44490 ;
  assign n44675 = n79881 & n44674 ;
  assign n44676 = n44497 | n44675 ;
  assign n44677 = n44673 | n44676 ;
  assign n79882 = ~n44497 ;
  assign n44681 = n79882 & n44677 ;
  assign n44682 = n44680 | n44681 ;
  assign n79883 = ~n44489 ;
  assign n44683 = n79883 & n44682 ;
  assign n79884 = ~n44479 ;
  assign n44684 = x80 & n79884 ;
  assign n79885 = ~n44474 ;
  assign n44685 = n79885 & n44684 ;
  assign n44686 = n44481 | n44685 ;
  assign n44687 = n44683 | n44686 ;
  assign n79886 = ~n44481 ;
  assign n44691 = n79886 & n44687 ;
  assign n44692 = n44690 | n44691 ;
  assign n79887 = ~n44473 ;
  assign n44693 = n79887 & n44692 ;
  assign n79888 = ~n44463 ;
  assign n44694 = x82 & n79888 ;
  assign n79889 = ~n44458 ;
  assign n44695 = n79889 & n44694 ;
  assign n44696 = n44465 | n44695 ;
  assign n44697 = n44693 | n44696 ;
  assign n79890 = ~n44465 ;
  assign n44701 = n79890 & n44697 ;
  assign n44702 = n44700 | n44701 ;
  assign n79891 = ~n44457 ;
  assign n44703 = n79891 & n44702 ;
  assign n79892 = ~n44447 ;
  assign n44704 = x84 & n79892 ;
  assign n79893 = ~n44442 ;
  assign n44705 = n79893 & n44704 ;
  assign n44706 = n44449 | n44705 ;
  assign n44707 = n44703 | n44706 ;
  assign n79894 = ~n44449 ;
  assign n44711 = n79894 & n44707 ;
  assign n44712 = n44710 | n44711 ;
  assign n79895 = ~n44441 ;
  assign n44713 = n79895 & n44712 ;
  assign n79896 = ~n44431 ;
  assign n44714 = x86 & n79896 ;
  assign n79897 = ~n44426 ;
  assign n44715 = n79897 & n44714 ;
  assign n44716 = n44433 | n44715 ;
  assign n44717 = n44713 | n44716 ;
  assign n79898 = ~n44433 ;
  assign n44721 = n79898 & n44717 ;
  assign n44722 = n44720 | n44721 ;
  assign n79899 = ~n44425 ;
  assign n44723 = n79899 & n44722 ;
  assign n79900 = ~n44415 ;
  assign n44724 = x88 & n79900 ;
  assign n79901 = ~n44410 ;
  assign n44725 = n79901 & n44724 ;
  assign n44726 = n44417 | n44725 ;
  assign n44728 = n44723 | n44726 ;
  assign n79902 = ~n44417 ;
  assign n44733 = n79902 & n44728 ;
  assign n44734 = n44731 | n44733 ;
  assign n79903 = ~n44409 ;
  assign n44735 = n79903 & n44734 ;
  assign n79904 = ~n44399 ;
  assign n44736 = x90 & n79904 ;
  assign n79905 = ~n44394 ;
  assign n44737 = n79905 & n44736 ;
  assign n44738 = n44401 | n44737 ;
  assign n44739 = n44735 | n44738 ;
  assign n79906 = ~n44401 ;
  assign n44744 = n79906 & n44739 ;
  assign n44745 = n44742 | n44744 ;
  assign n79907 = ~n44393 ;
  assign n44746 = n79907 & n44745 ;
  assign n79908 = ~n44383 ;
  assign n44747 = x92 & n79908 ;
  assign n79909 = ~n44378 ;
  assign n44748 = n79909 & n44747 ;
  assign n44749 = n44385 | n44748 ;
  assign n44750 = n44746 | n44749 ;
  assign n79910 = ~n44385 ;
  assign n44754 = n79910 & n44750 ;
  assign n44755 = n44753 | n44754 ;
  assign n79911 = ~n44377 ;
  assign n44756 = n79911 & n44755 ;
  assign n79912 = ~n44367 ;
  assign n44757 = x94 & n79912 ;
  assign n79913 = ~n44362 ;
  assign n44758 = n79913 & n44757 ;
  assign n44759 = n44369 | n44758 ;
  assign n44760 = n44756 | n44759 ;
  assign n79914 = ~n44369 ;
  assign n44764 = n79914 & n44760 ;
  assign n44765 = n44763 | n44764 ;
  assign n79915 = ~n44361 ;
  assign n44766 = n79915 & n44765 ;
  assign n79916 = ~n44351 ;
  assign n44767 = x96 & n79916 ;
  assign n79917 = ~n44346 ;
  assign n44768 = n79917 & n44767 ;
  assign n44769 = n44353 | n44768 ;
  assign n44770 = n44766 | n44769 ;
  assign n79918 = ~n44353 ;
  assign n44774 = n79918 & n44770 ;
  assign n44775 = n44773 | n44774 ;
  assign n79919 = ~n44345 ;
  assign n44776 = n79919 & n44775 ;
  assign n79920 = ~n44335 ;
  assign n44777 = x98 & n79920 ;
  assign n79921 = ~n44330 ;
  assign n44778 = n79921 & n44777 ;
  assign n44779 = n44337 | n44778 ;
  assign n44780 = n44776 | n44779 ;
  assign n79922 = ~n44337 ;
  assign n44784 = n79922 & n44780 ;
  assign n44785 = n44783 | n44784 ;
  assign n79923 = ~n44329 ;
  assign n44786 = n79923 & n44785 ;
  assign n79924 = ~n44319 ;
  assign n44787 = x100 & n79924 ;
  assign n79925 = ~n44314 ;
  assign n44788 = n79925 & n44787 ;
  assign n44789 = n44321 | n44788 ;
  assign n44791 = n44786 | n44789 ;
  assign n79926 = ~n44321 ;
  assign n44795 = n79926 & n44791 ;
  assign n44796 = n44794 | n44795 ;
  assign n79927 = ~n44313 ;
  assign n44797 = n79927 & n44796 ;
  assign n79928 = ~n44203 ;
  assign n44209 = n79928 & n44208 ;
  assign n44798 = n43725 | n44208 ;
  assign n79929 = ~n44798 ;
  assign n44799 = n44306 & n79929 ;
  assign n44800 = n44209 | n44799 ;
  assign n44801 = n44212 | n44800 ;
  assign n79930 = ~n43723 ;
  assign n44802 = n79930 & n44212 ;
  assign n79931 = ~n44802 ;
  assign n44803 = n44801 & n79931 ;
  assign n44804 = n69528 & n44803 ;
  assign n79932 = ~n44212 ;
  assign n44805 = n79932 & n44800 ;
  assign n44806 = n43723 & n44212 ;
  assign n79933 = ~n44806 ;
  assign n44807 = x102 & n79933 ;
  assign n79934 = ~n44805 ;
  assign n44808 = n79934 & n44807 ;
  assign n44809 = n12531 | n44808 ;
  assign n44810 = n44804 | n44809 ;
  assign n44811 = n44797 | n44810 ;
  assign n44812 = n69455 & n44803 ;
  assign n79935 = ~n44812 ;
  assign n44813 = n44811 & n79935 ;
  assign n44897 = n44313 | n44808 ;
  assign n44898 = n44804 | n44897 ;
  assign n79936 = ~n44898 ;
  assign n44899 = n44796 & n79936 ;
  assign n44900 = n44804 | n44808 ;
  assign n79937 = ~n44797 ;
  assign n44901 = n79937 & n44900 ;
  assign n44902 = n44899 | n44901 ;
  assign n79938 = ~n44813 ;
  assign n44903 = n79938 & n44902 ;
  assign n44904 = n11929 & n43723 ;
  assign n44905 = n44811 & n44904 ;
  assign n44906 = n44903 | n44905 ;
  assign n44907 = n69656 & n44906 ;
  assign n79939 = ~n44795 ;
  assign n44889 = n44794 & n79939 ;
  assign n44815 = x65 & n44611 ;
  assign n79940 = ~n44815 ;
  assign n44816 = n44608 & n79940 ;
  assign n44817 = n12319 | n44816 ;
  assign n44818 = n79855 & n44817 ;
  assign n44819 = n44616 | n44818 ;
  assign n44820 = n79858 & n44819 ;
  assign n44821 = n44619 | n44820 ;
  assign n44822 = n79859 & n44821 ;
  assign n44823 = n44625 | n44822 ;
  assign n44824 = n79862 & n44823 ;
  assign n44825 = n44629 | n44824 ;
  assign n44826 = n79863 & n44825 ;
  assign n44827 = n44635 | n44826 ;
  assign n44828 = n79866 & n44827 ;
  assign n44829 = n44639 | n44828 ;
  assign n44830 = n79867 & n44829 ;
  assign n44831 = n44645 | n44830 ;
  assign n44832 = n79870 & n44831 ;
  assign n44833 = n44649 | n44832 ;
  assign n44834 = n79871 & n44833 ;
  assign n44835 = n44655 | n44834 ;
  assign n44836 = n79874 & n44835 ;
  assign n44837 = n44659 | n44836 ;
  assign n44838 = n79875 & n44837 ;
  assign n44839 = n44665 | n44838 ;
  assign n44840 = n79878 & n44839 ;
  assign n44841 = n44669 | n44840 ;
  assign n44842 = n79879 & n44841 ;
  assign n44843 = n44676 | n44842 ;
  assign n44844 = n79882 & n44843 ;
  assign n44845 = n44680 | n44844 ;
  assign n44846 = n79883 & n44845 ;
  assign n44847 = n44686 | n44846 ;
  assign n44848 = n79886 & n44847 ;
  assign n44849 = n44690 | n44848 ;
  assign n44850 = n79887 & n44849 ;
  assign n44851 = n44696 | n44850 ;
  assign n44852 = n79890 & n44851 ;
  assign n44853 = n44700 | n44852 ;
  assign n44854 = n79891 & n44853 ;
  assign n44855 = n44706 | n44854 ;
  assign n44856 = n79894 & n44855 ;
  assign n44857 = n44710 | n44856 ;
  assign n44858 = n79895 & n44857 ;
  assign n44859 = n44716 | n44858 ;
  assign n44860 = n79898 & n44859 ;
  assign n44861 = n44720 | n44860 ;
  assign n44862 = n79899 & n44861 ;
  assign n44863 = n44726 | n44862 ;
  assign n44864 = n79902 & n44863 ;
  assign n44865 = n44731 | n44864 ;
  assign n44866 = n79903 & n44865 ;
  assign n44867 = n44738 | n44866 ;
  assign n44868 = n79906 & n44867 ;
  assign n44869 = n44742 | n44868 ;
  assign n44870 = n79907 & n44869 ;
  assign n44871 = n44749 | n44870 ;
  assign n44872 = n79910 & n44871 ;
  assign n44873 = n44753 | n44872 ;
  assign n44874 = n79911 & n44873 ;
  assign n44875 = n44759 | n44874 ;
  assign n44876 = n79914 & n44875 ;
  assign n44877 = n44763 | n44876 ;
  assign n44878 = n79915 & n44877 ;
  assign n44879 = n44769 | n44878 ;
  assign n44880 = n79918 & n44879 ;
  assign n44881 = n44773 | n44880 ;
  assign n44882 = n79919 & n44881 ;
  assign n44883 = n44779 | n44882 ;
  assign n44884 = n79922 & n44883 ;
  assign n44885 = n44783 | n44884 ;
  assign n44886 = n79923 & n44885 ;
  assign n44887 = n44789 | n44886 ;
  assign n44890 = n44321 | n44794 ;
  assign n79941 = ~n44890 ;
  assign n44891 = n44887 & n79941 ;
  assign n44892 = n44889 | n44891 ;
  assign n44893 = n79938 & n44892 ;
  assign n44894 = n44312 & n79935 ;
  assign n44895 = n44811 & n44894 ;
  assign n44896 = n44893 | n44895 ;
  assign n44908 = n69528 & n44896 ;
  assign n79942 = ~n44886 ;
  assign n44909 = n44789 & n79942 ;
  assign n44790 = n44329 | n44789 ;
  assign n79943 = ~n44790 ;
  assign n44910 = n79943 & n44885 ;
  assign n44911 = n44909 | n44910 ;
  assign n44912 = n79938 & n44911 ;
  assign n44913 = n44320 & n79935 ;
  assign n44914 = n44811 & n44913 ;
  assign n44915 = n44912 | n44914 ;
  assign n44916 = n69261 & n44915 ;
  assign n79944 = ~n44784 ;
  assign n44917 = n44783 & n79944 ;
  assign n44918 = n44337 | n44783 ;
  assign n79945 = ~n44918 ;
  assign n44919 = n44883 & n79945 ;
  assign n44920 = n44917 | n44919 ;
  assign n44921 = n79938 & n44920 ;
  assign n44922 = n44328 & n79935 ;
  assign n44923 = n44811 & n44922 ;
  assign n44924 = n44921 | n44923 ;
  assign n44925 = n69075 & n44924 ;
  assign n79946 = ~n44882 ;
  assign n44926 = n44779 & n79946 ;
  assign n44927 = n44345 | n44779 ;
  assign n79947 = ~n44927 ;
  assign n44928 = n44775 & n79947 ;
  assign n44929 = n44926 | n44928 ;
  assign n44930 = n79938 & n44929 ;
  assign n44931 = n44336 & n79935 ;
  assign n44932 = n44811 & n44931 ;
  assign n44933 = n44930 | n44932 ;
  assign n44934 = n68993 & n44933 ;
  assign n79948 = ~n44774 ;
  assign n44935 = n44773 & n79948 ;
  assign n44936 = n44353 | n44773 ;
  assign n79949 = ~n44936 ;
  assign n44937 = n44879 & n79949 ;
  assign n44938 = n44935 | n44937 ;
  assign n44939 = n79938 & n44938 ;
  assign n44940 = n44344 & n79935 ;
  assign n44941 = n44811 & n44940 ;
  assign n44942 = n44939 | n44941 ;
  assign n44943 = n68716 & n44942 ;
  assign n79950 = ~n44878 ;
  assign n44944 = n44769 & n79950 ;
  assign n44945 = n44361 | n44769 ;
  assign n79951 = ~n44945 ;
  assign n44946 = n44765 & n79951 ;
  assign n44947 = n44944 | n44946 ;
  assign n44948 = n79938 & n44947 ;
  assign n44949 = n44352 & n79935 ;
  assign n44950 = n44811 & n44949 ;
  assign n44951 = n44948 | n44950 ;
  assign n44952 = n68545 & n44951 ;
  assign n79952 = ~n44764 ;
  assign n44953 = n44763 & n79952 ;
  assign n44954 = n44369 | n44763 ;
  assign n79953 = ~n44954 ;
  assign n44955 = n44875 & n79953 ;
  assign n44956 = n44953 | n44955 ;
  assign n44957 = n79938 & n44956 ;
  assign n44958 = n44360 & n79935 ;
  assign n44959 = n44811 & n44958 ;
  assign n44960 = n44957 | n44959 ;
  assign n44961 = n68438 & n44960 ;
  assign n79954 = ~n44874 ;
  assign n44962 = n44759 & n79954 ;
  assign n44963 = n44377 | n44759 ;
  assign n79955 = ~n44963 ;
  assign n44964 = n44755 & n79955 ;
  assign n44965 = n44962 | n44964 ;
  assign n44966 = n79938 & n44965 ;
  assign n44967 = n44368 & n79935 ;
  assign n44968 = n44811 & n44967 ;
  assign n44969 = n44966 | n44968 ;
  assign n44970 = n68214 & n44969 ;
  assign n79956 = ~n44754 ;
  assign n44971 = n44753 & n79956 ;
  assign n44972 = n44385 | n44753 ;
  assign n79957 = ~n44972 ;
  assign n44973 = n44871 & n79957 ;
  assign n44974 = n44971 | n44973 ;
  assign n44975 = n79938 & n44974 ;
  assign n44976 = n44376 & n79935 ;
  assign n44977 = n44811 & n44976 ;
  assign n44978 = n44975 | n44977 ;
  assign n44979 = n68058 & n44978 ;
  assign n79958 = ~n44870 ;
  assign n44980 = n44749 & n79958 ;
  assign n44981 = n44393 | n44749 ;
  assign n79959 = ~n44981 ;
  assign n44982 = n44745 & n79959 ;
  assign n44983 = n44980 | n44982 ;
  assign n44984 = n79938 & n44983 ;
  assign n44985 = n44384 & n79935 ;
  assign n44986 = n44811 & n44985 ;
  assign n44987 = n44984 | n44986 ;
  assign n44988 = n67986 & n44987 ;
  assign n79960 = ~n44744 ;
  assign n44989 = n44742 & n79960 ;
  assign n44743 = n44401 | n44742 ;
  assign n79961 = ~n44743 ;
  assign n44990 = n44739 & n79961 ;
  assign n44991 = n44989 | n44990 ;
  assign n44992 = n79938 & n44991 ;
  assign n44993 = n44392 & n79935 ;
  assign n44994 = n44811 & n44993 ;
  assign n44995 = n44992 | n44994 ;
  assign n44996 = n67763 & n44995 ;
  assign n79962 = ~n44866 ;
  assign n44997 = n44738 & n79962 ;
  assign n44998 = n44409 | n44738 ;
  assign n79963 = ~n44998 ;
  assign n44999 = n44734 & n79963 ;
  assign n45000 = n44997 | n44999 ;
  assign n45001 = n79938 & n45000 ;
  assign n45002 = n44400 & n79935 ;
  assign n45003 = n44811 & n45002 ;
  assign n45004 = n45001 | n45003 ;
  assign n45005 = n67622 & n45004 ;
  assign n79964 = ~n44733 ;
  assign n45006 = n44731 & n79964 ;
  assign n44732 = n44417 | n44731 ;
  assign n79965 = ~n44732 ;
  assign n45007 = n44728 & n79965 ;
  assign n45008 = n45006 | n45007 ;
  assign n45009 = n79938 & n45008 ;
  assign n45010 = n44408 & n79935 ;
  assign n45011 = n44811 & n45010 ;
  assign n45012 = n45009 | n45011 ;
  assign n45013 = n67531 & n45012 ;
  assign n79966 = ~n44862 ;
  assign n45014 = n44726 & n79966 ;
  assign n44727 = n44425 | n44726 ;
  assign n79967 = ~n44727 ;
  assign n45015 = n79967 & n44861 ;
  assign n45016 = n45014 | n45015 ;
  assign n45017 = n79938 & n45016 ;
  assign n45018 = n44416 & n79935 ;
  assign n45019 = n44811 & n45018 ;
  assign n45020 = n45017 | n45019 ;
  assign n45021 = n67348 & n45020 ;
  assign n79968 = ~n44721 ;
  assign n45022 = n44720 & n79968 ;
  assign n45023 = n44433 | n44720 ;
  assign n79969 = ~n45023 ;
  assign n45024 = n44859 & n79969 ;
  assign n45025 = n45022 | n45024 ;
  assign n45026 = n79938 & n45025 ;
  assign n45027 = n44424 & n79935 ;
  assign n45028 = n44811 & n45027 ;
  assign n45029 = n45026 | n45028 ;
  assign n45030 = n67222 & n45029 ;
  assign n79970 = ~n44858 ;
  assign n45031 = n44716 & n79970 ;
  assign n45032 = n44441 | n44716 ;
  assign n79971 = ~n45032 ;
  assign n45033 = n44712 & n79971 ;
  assign n45034 = n45031 | n45033 ;
  assign n45035 = n79938 & n45034 ;
  assign n45036 = n44432 & n79935 ;
  assign n45037 = n44811 & n45036 ;
  assign n45038 = n45035 | n45037 ;
  assign n45039 = n67164 & n45038 ;
  assign n79972 = ~n44711 ;
  assign n45040 = n44710 & n79972 ;
  assign n45041 = n44449 | n44710 ;
  assign n79973 = ~n45041 ;
  assign n45042 = n44855 & n79973 ;
  assign n45043 = n45040 | n45042 ;
  assign n45044 = n79938 & n45043 ;
  assign n45045 = n44440 & n79935 ;
  assign n45046 = n44811 & n45045 ;
  assign n45047 = n45044 | n45046 ;
  assign n45048 = n66979 & n45047 ;
  assign n79974 = ~n44854 ;
  assign n45049 = n44706 & n79974 ;
  assign n45050 = n44457 | n44706 ;
  assign n79975 = ~n45050 ;
  assign n45051 = n44702 & n79975 ;
  assign n45052 = n45049 | n45051 ;
  assign n45053 = n79938 & n45052 ;
  assign n45054 = n44448 & n79935 ;
  assign n45055 = n44811 & n45054 ;
  assign n45056 = n45053 | n45055 ;
  assign n45057 = n66868 & n45056 ;
  assign n79976 = ~n44701 ;
  assign n45058 = n44700 & n79976 ;
  assign n45059 = n44465 | n44700 ;
  assign n79977 = ~n45059 ;
  assign n45060 = n44851 & n79977 ;
  assign n45061 = n45058 | n45060 ;
  assign n45062 = n79938 & n45061 ;
  assign n45063 = n44456 & n79935 ;
  assign n45064 = n44811 & n45063 ;
  assign n45065 = n45062 | n45064 ;
  assign n45066 = n66797 & n45065 ;
  assign n79978 = ~n44850 ;
  assign n45067 = n44696 & n79978 ;
  assign n45068 = n44473 | n44696 ;
  assign n79979 = ~n45068 ;
  assign n45069 = n44692 & n79979 ;
  assign n45070 = n45067 | n45069 ;
  assign n45071 = n79938 & n45070 ;
  assign n45072 = n44464 & n79935 ;
  assign n45073 = n44811 & n45072 ;
  assign n45074 = n45071 | n45073 ;
  assign n45075 = n66654 & n45074 ;
  assign n79980 = ~n44691 ;
  assign n45076 = n44690 & n79980 ;
  assign n45077 = n44481 | n44690 ;
  assign n79981 = ~n45077 ;
  assign n45078 = n44847 & n79981 ;
  assign n45079 = n45076 | n45078 ;
  assign n45080 = n79938 & n45079 ;
  assign n45081 = n44472 & n79935 ;
  assign n45082 = n44811 & n45081 ;
  assign n45083 = n45080 | n45082 ;
  assign n45084 = n66560 & n45083 ;
  assign n79982 = ~n44846 ;
  assign n45085 = n44686 & n79982 ;
  assign n45086 = n44489 | n44686 ;
  assign n79983 = ~n45086 ;
  assign n45087 = n44682 & n79983 ;
  assign n45088 = n45085 | n45087 ;
  assign n45089 = n79938 & n45088 ;
  assign n45090 = n44480 & n79935 ;
  assign n45091 = n44811 & n45090 ;
  assign n45092 = n45089 | n45091 ;
  assign n45093 = n66505 & n45092 ;
  assign n79984 = ~n44681 ;
  assign n45094 = n44680 & n79984 ;
  assign n45095 = n44497 | n44680 ;
  assign n79985 = ~n45095 ;
  assign n45096 = n44843 & n79985 ;
  assign n45097 = n45094 | n45096 ;
  assign n45098 = n79938 & n45097 ;
  assign n45099 = n44488 & n79935 ;
  assign n45100 = n44811 & n45099 ;
  assign n45101 = n45098 | n45100 ;
  assign n45102 = n66379 & n45101 ;
  assign n79986 = ~n44842 ;
  assign n45103 = n44676 & n79986 ;
  assign n45104 = n44505 | n44676 ;
  assign n79987 = ~n45104 ;
  assign n45105 = n44672 & n79987 ;
  assign n45106 = n45103 | n45105 ;
  assign n45107 = n79938 & n45106 ;
  assign n45108 = n44496 & n79935 ;
  assign n45109 = n44811 & n45108 ;
  assign n45110 = n45107 | n45109 ;
  assign n45111 = n66299 & n45110 ;
  assign n79988 = ~n44671 ;
  assign n45112 = n44669 & n79988 ;
  assign n44670 = n44513 | n44669 ;
  assign n79989 = ~n44670 ;
  assign n45113 = n44666 & n79989 ;
  assign n45114 = n45112 | n45113 ;
  assign n45115 = n79938 & n45114 ;
  assign n45116 = n44504 & n79935 ;
  assign n45117 = n44811 & n45116 ;
  assign n45118 = n45115 | n45117 ;
  assign n45119 = n66244 & n45118 ;
  assign n79990 = ~n44838 ;
  assign n45120 = n44665 & n79990 ;
  assign n45121 = n44521 | n44665 ;
  assign n79991 = ~n45121 ;
  assign n45122 = n44661 & n79991 ;
  assign n45123 = n45120 | n45122 ;
  assign n45124 = n79938 & n45123 ;
  assign n45125 = n44512 & n79935 ;
  assign n45126 = n44811 & n45125 ;
  assign n45127 = n45124 | n45126 ;
  assign n45128 = n66145 & n45127 ;
  assign n79992 = ~n44660 ;
  assign n45129 = n44659 & n79992 ;
  assign n45130 = n44529 | n44659 ;
  assign n79993 = ~n45130 ;
  assign n45131 = n44835 & n79993 ;
  assign n45132 = n45129 | n45131 ;
  assign n45133 = n79938 & n45132 ;
  assign n45134 = n44520 & n79935 ;
  assign n45135 = n44811 & n45134 ;
  assign n45136 = n45133 | n45135 ;
  assign n45137 = n66081 & n45136 ;
  assign n79994 = ~n44834 ;
  assign n45138 = n44655 & n79994 ;
  assign n45139 = n44537 | n44655 ;
  assign n79995 = ~n45139 ;
  assign n45140 = n44651 & n79995 ;
  assign n45141 = n45138 | n45140 ;
  assign n45142 = n79938 & n45141 ;
  assign n45143 = n44528 & n79935 ;
  assign n45144 = n44811 & n45143 ;
  assign n45145 = n45142 | n45144 ;
  assign n45146 = n66043 & n45145 ;
  assign n79996 = ~n44650 ;
  assign n45147 = n44649 & n79996 ;
  assign n45148 = n44545 | n44649 ;
  assign n79997 = ~n45148 ;
  assign n45149 = n44831 & n79997 ;
  assign n45150 = n45147 | n45149 ;
  assign n45151 = n79938 & n45150 ;
  assign n45152 = n44536 & n79935 ;
  assign n45153 = n44811 & n45152 ;
  assign n45154 = n45151 | n45153 ;
  assign n45155 = n65960 & n45154 ;
  assign n79998 = ~n44830 ;
  assign n45156 = n44645 & n79998 ;
  assign n45157 = n44553 | n44645 ;
  assign n79999 = ~n45157 ;
  assign n45158 = n44641 & n79999 ;
  assign n45159 = n45156 | n45158 ;
  assign n45160 = n79938 & n45159 ;
  assign n45161 = n44544 & n79935 ;
  assign n45162 = n44811 & n45161 ;
  assign n45163 = n45160 | n45162 ;
  assign n45164 = n65909 & n45163 ;
  assign n80000 = ~n44640 ;
  assign n45165 = n44639 & n80000 ;
  assign n45166 = n44561 | n44639 ;
  assign n80001 = ~n45166 ;
  assign n45167 = n44827 & n80001 ;
  assign n45168 = n45165 | n45167 ;
  assign n45169 = n79938 & n45168 ;
  assign n45170 = n44552 & n79935 ;
  assign n45171 = n44811 & n45170 ;
  assign n45172 = n45169 | n45171 ;
  assign n45173 = n65877 & n45172 ;
  assign n80002 = ~n44826 ;
  assign n45174 = n44635 & n80002 ;
  assign n45175 = n44570 | n44635 ;
  assign n80003 = ~n45175 ;
  assign n45176 = n44631 & n80003 ;
  assign n45177 = n45174 | n45176 ;
  assign n45178 = n79938 & n45177 ;
  assign n45179 = n44560 & n79935 ;
  assign n45180 = n44811 & n45179 ;
  assign n45181 = n45178 | n45180 ;
  assign n45182 = n65820 & n45181 ;
  assign n80004 = ~n44630 ;
  assign n45183 = n44629 & n80004 ;
  assign n45184 = n44578 | n44629 ;
  assign n80005 = ~n45184 ;
  assign n45185 = n44823 & n80005 ;
  assign n45186 = n45183 | n45185 ;
  assign n45187 = n79938 & n45186 ;
  assign n45188 = n44569 & n79935 ;
  assign n45189 = n44811 & n45188 ;
  assign n45190 = n45187 | n45189 ;
  assign n45191 = n65791 & n45190 ;
  assign n80006 = ~n44822 ;
  assign n45193 = n44625 & n80006 ;
  assign n45192 = n44588 | n44625 ;
  assign n80007 = ~n45192 ;
  assign n45194 = n44821 & n80007 ;
  assign n45195 = n45193 | n45194 ;
  assign n45196 = n79938 & n45195 ;
  assign n45197 = n44577 & n79935 ;
  assign n45198 = n44811 & n45197 ;
  assign n45199 = n45196 | n45198 ;
  assign n45200 = n65772 & n45199 ;
  assign n80008 = ~n44620 ;
  assign n45202 = n44619 & n80008 ;
  assign n45201 = n44596 | n44619 ;
  assign n80009 = ~n45201 ;
  assign n45203 = n44617 & n80009 ;
  assign n45204 = n45202 | n45203 ;
  assign n45205 = n79938 & n45204 ;
  assign n45206 = n44586 & n79935 ;
  assign n45207 = n44811 & n45206 ;
  assign n45208 = n45205 | n45207 ;
  assign n45209 = n65746 & n45208 ;
  assign n80010 = ~n44818 ;
  assign n45211 = n44616 & n80010 ;
  assign n45210 = n44612 | n44616 ;
  assign n80011 = ~n45210 ;
  assign n45212 = n44817 & n80011 ;
  assign n45213 = n45211 | n45212 ;
  assign n45214 = n79938 & n45213 ;
  assign n45215 = n44595 & n79935 ;
  assign n45216 = n44811 & n45215 ;
  assign n45217 = n45214 | n45216 ;
  assign n45218 = n65721 & n45217 ;
  assign n45219 = n12319 & n44608 ;
  assign n45220 = n79940 & n45219 ;
  assign n80012 = ~n45220 ;
  assign n45221 = n44817 & n80012 ;
  assign n45222 = n79938 & n45221 ;
  assign n45223 = n44611 & n79935 ;
  assign n45224 = n44811 & n45223 ;
  assign n45225 = n45222 | n45224 ;
  assign n45226 = n65686 & n45225 ;
  assign n44814 = n12319 & n79938 ;
  assign n45233 = x64 & n79938 ;
  assign n80013 = ~n45233 ;
  assign n45234 = x25 & n80013 ;
  assign n45235 = n44814 | n45234 ;
  assign n45237 = x65 & n45235 ;
  assign n44888 = n79926 & n44887 ;
  assign n45227 = n44794 | n44888 ;
  assign n45228 = n79927 & n45227 ;
  assign n45229 = n44810 | n45228 ;
  assign n45230 = n79935 & n45229 ;
  assign n80014 = ~n45230 ;
  assign n45231 = x64 & n80014 ;
  assign n80015 = ~n45231 ;
  assign n45232 = x25 & n80015 ;
  assign n45236 = x65 | n44814 ;
  assign n45238 = n45232 | n45236 ;
  assign n80016 = ~n45237 ;
  assign n45239 = n80016 & n45238 ;
  assign n45240 = n12955 | n45239 ;
  assign n45241 = n65670 & n45235 ;
  assign n80017 = ~n45241 ;
  assign n45242 = n45240 & n80017 ;
  assign n80018 = ~n45224 ;
  assign n45243 = x66 & n80018 ;
  assign n80019 = ~n45222 ;
  assign n45244 = n80019 & n45243 ;
  assign n45245 = n45226 | n45244 ;
  assign n45246 = n45242 | n45245 ;
  assign n80020 = ~n45226 ;
  assign n45247 = n80020 & n45246 ;
  assign n80021 = ~n45216 ;
  assign n45248 = x67 & n80021 ;
  assign n80022 = ~n45214 ;
  assign n45249 = n80022 & n45248 ;
  assign n45250 = n45247 | n45249 ;
  assign n80023 = ~n45218 ;
  assign n45251 = n80023 & n45250 ;
  assign n80024 = ~n45207 ;
  assign n45252 = x68 & n80024 ;
  assign n80025 = ~n45205 ;
  assign n45253 = n80025 & n45252 ;
  assign n45254 = n45209 | n45253 ;
  assign n45255 = n45251 | n45254 ;
  assign n80026 = ~n45209 ;
  assign n45256 = n80026 & n45255 ;
  assign n80027 = ~n45198 ;
  assign n45257 = x69 & n80027 ;
  assign n80028 = ~n45196 ;
  assign n45258 = n80028 & n45257 ;
  assign n45259 = n45256 | n45258 ;
  assign n80029 = ~n45200 ;
  assign n45260 = n80029 & n45259 ;
  assign n80030 = ~n45189 ;
  assign n45261 = x70 & n80030 ;
  assign n80031 = ~n45187 ;
  assign n45262 = n80031 & n45261 ;
  assign n45263 = n45191 | n45262 ;
  assign n45264 = n45260 | n45263 ;
  assign n80032 = ~n45191 ;
  assign n45265 = n80032 & n45264 ;
  assign n80033 = ~n45180 ;
  assign n45266 = x71 & n80033 ;
  assign n80034 = ~n45178 ;
  assign n45267 = n80034 & n45266 ;
  assign n45268 = n45182 | n45267 ;
  assign n45271 = n45265 | n45268 ;
  assign n80035 = ~n45182 ;
  assign n45272 = n80035 & n45271 ;
  assign n80036 = ~n45171 ;
  assign n45273 = x72 & n80036 ;
  assign n80037 = ~n45169 ;
  assign n45274 = n80037 & n45273 ;
  assign n45275 = n45173 | n45274 ;
  assign n45276 = n45272 | n45275 ;
  assign n80038 = ~n45173 ;
  assign n45277 = n80038 & n45276 ;
  assign n80039 = ~n45162 ;
  assign n45278 = x73 & n80039 ;
  assign n80040 = ~n45160 ;
  assign n45279 = n80040 & n45278 ;
  assign n45280 = n45164 | n45279 ;
  assign n45282 = n45277 | n45280 ;
  assign n80041 = ~n45164 ;
  assign n45283 = n80041 & n45282 ;
  assign n80042 = ~n45153 ;
  assign n45284 = x74 & n80042 ;
  assign n80043 = ~n45151 ;
  assign n45285 = n80043 & n45284 ;
  assign n45286 = n45155 | n45285 ;
  assign n45287 = n45283 | n45286 ;
  assign n80044 = ~n45155 ;
  assign n45288 = n80044 & n45287 ;
  assign n80045 = ~n45144 ;
  assign n45289 = x75 & n80045 ;
  assign n80046 = ~n45142 ;
  assign n45290 = n80046 & n45289 ;
  assign n45291 = n45146 | n45290 ;
  assign n45293 = n45288 | n45291 ;
  assign n80047 = ~n45146 ;
  assign n45294 = n80047 & n45293 ;
  assign n80048 = ~n45135 ;
  assign n45295 = x76 & n80048 ;
  assign n80049 = ~n45133 ;
  assign n45296 = n80049 & n45295 ;
  assign n45297 = n45137 | n45296 ;
  assign n45298 = n45294 | n45297 ;
  assign n80050 = ~n45137 ;
  assign n45299 = n80050 & n45298 ;
  assign n80051 = ~n45126 ;
  assign n45300 = x77 & n80051 ;
  assign n80052 = ~n45124 ;
  assign n45301 = n80052 & n45300 ;
  assign n45302 = n45128 | n45301 ;
  assign n45304 = n45299 | n45302 ;
  assign n80053 = ~n45128 ;
  assign n45305 = n80053 & n45304 ;
  assign n80054 = ~n45117 ;
  assign n45306 = x78 & n80054 ;
  assign n80055 = ~n45115 ;
  assign n45307 = n80055 & n45306 ;
  assign n45308 = n45119 | n45307 ;
  assign n45309 = n45305 | n45308 ;
  assign n80056 = ~n45119 ;
  assign n45310 = n80056 & n45309 ;
  assign n80057 = ~n45109 ;
  assign n45311 = x79 & n80057 ;
  assign n80058 = ~n45107 ;
  assign n45312 = n80058 & n45311 ;
  assign n45313 = n45111 | n45312 ;
  assign n45315 = n45310 | n45313 ;
  assign n80059 = ~n45111 ;
  assign n45316 = n80059 & n45315 ;
  assign n80060 = ~n45100 ;
  assign n45317 = x80 & n80060 ;
  assign n80061 = ~n45098 ;
  assign n45318 = n80061 & n45317 ;
  assign n45319 = n45102 | n45318 ;
  assign n45320 = n45316 | n45319 ;
  assign n80062 = ~n45102 ;
  assign n45321 = n80062 & n45320 ;
  assign n80063 = ~n45091 ;
  assign n45322 = x81 & n80063 ;
  assign n80064 = ~n45089 ;
  assign n45323 = n80064 & n45322 ;
  assign n45324 = n45093 | n45323 ;
  assign n45326 = n45321 | n45324 ;
  assign n80065 = ~n45093 ;
  assign n45327 = n80065 & n45326 ;
  assign n80066 = ~n45082 ;
  assign n45328 = x82 & n80066 ;
  assign n80067 = ~n45080 ;
  assign n45329 = n80067 & n45328 ;
  assign n45330 = n45084 | n45329 ;
  assign n45331 = n45327 | n45330 ;
  assign n80068 = ~n45084 ;
  assign n45332 = n80068 & n45331 ;
  assign n80069 = ~n45073 ;
  assign n45333 = x83 & n80069 ;
  assign n80070 = ~n45071 ;
  assign n45334 = n80070 & n45333 ;
  assign n45335 = n45075 | n45334 ;
  assign n45337 = n45332 | n45335 ;
  assign n80071 = ~n45075 ;
  assign n45338 = n80071 & n45337 ;
  assign n80072 = ~n45064 ;
  assign n45339 = x84 & n80072 ;
  assign n80073 = ~n45062 ;
  assign n45340 = n80073 & n45339 ;
  assign n45341 = n45066 | n45340 ;
  assign n45342 = n45338 | n45341 ;
  assign n80074 = ~n45066 ;
  assign n45343 = n80074 & n45342 ;
  assign n80075 = ~n45055 ;
  assign n45344 = x85 & n80075 ;
  assign n80076 = ~n45053 ;
  assign n45345 = n80076 & n45344 ;
  assign n45346 = n45057 | n45345 ;
  assign n45348 = n45343 | n45346 ;
  assign n80077 = ~n45057 ;
  assign n45349 = n80077 & n45348 ;
  assign n80078 = ~n45046 ;
  assign n45350 = x86 & n80078 ;
  assign n80079 = ~n45044 ;
  assign n45351 = n80079 & n45350 ;
  assign n45352 = n45048 | n45351 ;
  assign n45353 = n45349 | n45352 ;
  assign n80080 = ~n45048 ;
  assign n45354 = n80080 & n45353 ;
  assign n80081 = ~n45037 ;
  assign n45355 = x87 & n80081 ;
  assign n80082 = ~n45035 ;
  assign n45356 = n80082 & n45355 ;
  assign n45357 = n45039 | n45356 ;
  assign n45359 = n45354 | n45357 ;
  assign n80083 = ~n45039 ;
  assign n45360 = n80083 & n45359 ;
  assign n80084 = ~n45028 ;
  assign n45361 = x88 & n80084 ;
  assign n80085 = ~n45026 ;
  assign n45362 = n80085 & n45361 ;
  assign n45363 = n45030 | n45362 ;
  assign n45364 = n45360 | n45363 ;
  assign n80086 = ~n45030 ;
  assign n45365 = n80086 & n45364 ;
  assign n80087 = ~n45019 ;
  assign n45366 = x89 & n80087 ;
  assign n80088 = ~n45017 ;
  assign n45367 = n80088 & n45366 ;
  assign n45368 = n45021 | n45367 ;
  assign n45370 = n45365 | n45368 ;
  assign n80089 = ~n45021 ;
  assign n45371 = n80089 & n45370 ;
  assign n80090 = ~n45011 ;
  assign n45372 = x90 & n80090 ;
  assign n80091 = ~n45009 ;
  assign n45373 = n80091 & n45372 ;
  assign n45374 = n45013 | n45373 ;
  assign n45375 = n45371 | n45374 ;
  assign n80092 = ~n45013 ;
  assign n45376 = n80092 & n45375 ;
  assign n80093 = ~n45003 ;
  assign n45377 = x91 & n80093 ;
  assign n80094 = ~n45001 ;
  assign n45378 = n80094 & n45377 ;
  assign n45379 = n45005 | n45378 ;
  assign n45381 = n45376 | n45379 ;
  assign n80095 = ~n45005 ;
  assign n45382 = n80095 & n45381 ;
  assign n80096 = ~n44994 ;
  assign n45383 = x92 & n80096 ;
  assign n80097 = ~n44992 ;
  assign n45384 = n80097 & n45383 ;
  assign n45385 = n44996 | n45384 ;
  assign n45386 = n45382 | n45385 ;
  assign n80098 = ~n44996 ;
  assign n45387 = n80098 & n45386 ;
  assign n80099 = ~n44986 ;
  assign n45388 = x93 & n80099 ;
  assign n80100 = ~n44984 ;
  assign n45389 = n80100 & n45388 ;
  assign n45390 = n44988 | n45389 ;
  assign n45392 = n45387 | n45390 ;
  assign n80101 = ~n44988 ;
  assign n45393 = n80101 & n45392 ;
  assign n80102 = ~n44977 ;
  assign n45394 = x94 & n80102 ;
  assign n80103 = ~n44975 ;
  assign n45395 = n80103 & n45394 ;
  assign n45396 = n44979 | n45395 ;
  assign n45397 = n45393 | n45396 ;
  assign n80104 = ~n44979 ;
  assign n45398 = n80104 & n45397 ;
  assign n80105 = ~n44968 ;
  assign n45399 = x95 & n80105 ;
  assign n80106 = ~n44966 ;
  assign n45400 = n80106 & n45399 ;
  assign n45401 = n44970 | n45400 ;
  assign n45403 = n45398 | n45401 ;
  assign n80107 = ~n44970 ;
  assign n45404 = n80107 & n45403 ;
  assign n80108 = ~n44959 ;
  assign n45405 = x96 & n80108 ;
  assign n80109 = ~n44957 ;
  assign n45406 = n80109 & n45405 ;
  assign n45407 = n44961 | n45406 ;
  assign n45408 = n45404 | n45407 ;
  assign n80110 = ~n44961 ;
  assign n45409 = n80110 & n45408 ;
  assign n80111 = ~n44950 ;
  assign n45410 = x97 & n80111 ;
  assign n80112 = ~n44948 ;
  assign n45411 = n80112 & n45410 ;
  assign n45412 = n44952 | n45411 ;
  assign n45414 = n45409 | n45412 ;
  assign n80113 = ~n44952 ;
  assign n45415 = n80113 & n45414 ;
  assign n80114 = ~n44941 ;
  assign n45416 = x98 & n80114 ;
  assign n80115 = ~n44939 ;
  assign n45417 = n80115 & n45416 ;
  assign n45418 = n44943 | n45417 ;
  assign n45419 = n45415 | n45418 ;
  assign n80116 = ~n44943 ;
  assign n45420 = n80116 & n45419 ;
  assign n80117 = ~n44932 ;
  assign n45421 = x99 & n80117 ;
  assign n80118 = ~n44930 ;
  assign n45422 = n80118 & n45421 ;
  assign n45423 = n44934 | n45422 ;
  assign n45425 = n45420 | n45423 ;
  assign n80119 = ~n44934 ;
  assign n45426 = n80119 & n45425 ;
  assign n80120 = ~n44923 ;
  assign n45427 = x100 & n80120 ;
  assign n80121 = ~n44921 ;
  assign n45428 = n80121 & n45427 ;
  assign n45429 = n44925 | n45428 ;
  assign n45430 = n45426 | n45429 ;
  assign n80122 = ~n44925 ;
  assign n45431 = n80122 & n45430 ;
  assign n80123 = ~n44914 ;
  assign n45432 = x101 & n80123 ;
  assign n80124 = ~n44912 ;
  assign n45433 = n80124 & n45432 ;
  assign n45434 = n44916 | n45433 ;
  assign n45436 = n45431 | n45434 ;
  assign n80125 = ~n44916 ;
  assign n45437 = n80125 & n45436 ;
  assign n80126 = ~n44895 ;
  assign n45438 = x102 & n80126 ;
  assign n80127 = ~n44893 ;
  assign n45439 = n80127 & n45438 ;
  assign n45440 = n44908 | n45439 ;
  assign n45441 = n45437 | n45440 ;
  assign n80128 = ~n44908 ;
  assign n45442 = n80128 & n45441 ;
  assign n80129 = ~n44905 ;
  assign n45443 = x103 & n80129 ;
  assign n80130 = ~n44903 ;
  assign n45444 = n80130 & n45443 ;
  assign n45445 = n44907 | n45444 ;
  assign n45447 = n45442 | n45445 ;
  assign n80131 = ~n44907 ;
  assign n45448 = n80131 & n45447 ;
  assign n45449 = n13184 | n45448 ;
  assign n80132 = ~n44906 ;
  assign n45450 = n80132 & n45449 ;
  assign n80133 = ~n45442 ;
  assign n45446 = n80133 & n45445 ;
  assign n45457 = n44814 | n45232 ;
  assign n45458 = x65 & n45457 ;
  assign n80134 = ~n45458 ;
  assign n45459 = n45238 & n80134 ;
  assign n45460 = n12955 | n45459 ;
  assign n45461 = n80017 & n45460 ;
  assign n45462 = n45245 | n45461 ;
  assign n45463 = n80020 & n45462 ;
  assign n45464 = n45218 | n45249 ;
  assign n45466 = n45463 | n45464 ;
  assign n45467 = n80023 & n45466 ;
  assign n45468 = n45253 | n45467 ;
  assign n45470 = n80026 & n45468 ;
  assign n45471 = n45200 | n45258 ;
  assign n45473 = n45470 | n45471 ;
  assign n45474 = n80029 & n45473 ;
  assign n45475 = n45262 | n45474 ;
  assign n45477 = n80032 & n45475 ;
  assign n45478 = n45268 | n45477 ;
  assign n45479 = n80035 & n45478 ;
  assign n45480 = n45275 | n45479 ;
  assign n45482 = n80038 & n45480 ;
  assign n45483 = n45280 | n45482 ;
  assign n45484 = n80041 & n45483 ;
  assign n45485 = n45286 | n45484 ;
  assign n45487 = n80044 & n45485 ;
  assign n45488 = n45291 | n45487 ;
  assign n45489 = n80047 & n45488 ;
  assign n45490 = n45297 | n45489 ;
  assign n45492 = n80050 & n45490 ;
  assign n45493 = n45302 | n45492 ;
  assign n45494 = n80053 & n45493 ;
  assign n45495 = n45308 | n45494 ;
  assign n45497 = n80056 & n45495 ;
  assign n45498 = n45313 | n45497 ;
  assign n45499 = n80059 & n45498 ;
  assign n45500 = n45319 | n45499 ;
  assign n45502 = n80062 & n45500 ;
  assign n45503 = n45324 | n45502 ;
  assign n45504 = n80065 & n45503 ;
  assign n45505 = n45330 | n45504 ;
  assign n45507 = n80068 & n45505 ;
  assign n45508 = n45335 | n45507 ;
  assign n45509 = n80071 & n45508 ;
  assign n45510 = n45341 | n45509 ;
  assign n45512 = n80074 & n45510 ;
  assign n45513 = n45346 | n45512 ;
  assign n45514 = n80077 & n45513 ;
  assign n45515 = n45352 | n45514 ;
  assign n45517 = n80080 & n45515 ;
  assign n45518 = n45357 | n45517 ;
  assign n45519 = n80083 & n45518 ;
  assign n45520 = n45363 | n45519 ;
  assign n45522 = n80086 & n45520 ;
  assign n45523 = n45368 | n45522 ;
  assign n45524 = n80089 & n45523 ;
  assign n45525 = n45374 | n45524 ;
  assign n45527 = n80092 & n45525 ;
  assign n45528 = n45379 | n45527 ;
  assign n45529 = n80095 & n45528 ;
  assign n45530 = n45385 | n45529 ;
  assign n45532 = n80098 & n45530 ;
  assign n45533 = n45390 | n45532 ;
  assign n45534 = n80101 & n45533 ;
  assign n45535 = n45396 | n45534 ;
  assign n45537 = n80104 & n45535 ;
  assign n45538 = n45401 | n45537 ;
  assign n45539 = n80107 & n45538 ;
  assign n45540 = n45407 | n45539 ;
  assign n45542 = n80110 & n45540 ;
  assign n45543 = n45412 | n45542 ;
  assign n45544 = n80113 & n45543 ;
  assign n45545 = n45418 | n45544 ;
  assign n45547 = n80116 & n45545 ;
  assign n45548 = n45423 | n45547 ;
  assign n45549 = n80119 & n45548 ;
  assign n45550 = n45429 | n45549 ;
  assign n45552 = n80122 & n45550 ;
  assign n45553 = n45434 | n45552 ;
  assign n45554 = n80125 & n45553 ;
  assign n45556 = n45440 | n45554 ;
  assign n45563 = n44908 | n45445 ;
  assign n80135 = ~n45563 ;
  assign n45564 = n45556 & n80135 ;
  assign n45565 = n45446 | n45564 ;
  assign n45566 = n45449 | n45565 ;
  assign n80136 = ~n45450 ;
  assign n45567 = n80136 & n45566 ;
  assign n45568 = n69857 & n45567 ;
  assign n80137 = ~n45449 ;
  assign n46102 = n80137 & n45565 ;
  assign n46103 = n44906 & n45449 ;
  assign n80138 = ~n46103 ;
  assign n46104 = x104 & n80138 ;
  assign n80139 = ~n46102 ;
  assign n46105 = n80139 & n46104 ;
  assign n46106 = n45568 | n46105 ;
  assign n45455 = n44896 & n45449 ;
  assign n80140 = ~n45554 ;
  assign n45555 = n45440 & n80140 ;
  assign n45557 = n44916 | n45440 ;
  assign n80141 = ~n45557 ;
  assign n45558 = n45436 & n80141 ;
  assign n45559 = n45555 | n45558 ;
  assign n45560 = n69851 & n45559 ;
  assign n80142 = ~n45448 ;
  assign n45561 = n80142 & n45560 ;
  assign n45562 = n45455 | n45561 ;
  assign n45569 = n69656 & n45562 ;
  assign n45570 = n44915 & n45449 ;
  assign n80143 = ~n45431 ;
  assign n45435 = n80143 & n45434 ;
  assign n45571 = n44925 | n45434 ;
  assign n80144 = ~n45571 ;
  assign n45572 = n45550 & n80144 ;
  assign n45573 = n45435 | n45572 ;
  assign n45574 = n69851 & n45573 ;
  assign n45575 = n80142 & n45574 ;
  assign n45576 = n45570 | n45575 ;
  assign n45577 = n69528 & n45576 ;
  assign n80145 = ~n45575 ;
  assign n46090 = x102 & n80145 ;
  assign n80146 = ~n45570 ;
  assign n46091 = n80146 & n46090 ;
  assign n46092 = n45577 | n46091 ;
  assign n45578 = n44924 & n45449 ;
  assign n80147 = ~n45549 ;
  assign n45551 = n45429 & n80147 ;
  assign n45579 = n44934 | n45429 ;
  assign n80148 = ~n45579 ;
  assign n45580 = n45425 & n80148 ;
  assign n45581 = n45551 | n45580 ;
  assign n45582 = n69851 & n45581 ;
  assign n45583 = n80142 & n45582 ;
  assign n45584 = n45578 | n45583 ;
  assign n45585 = n69261 & n45584 ;
  assign n45586 = n44933 & n45449 ;
  assign n80149 = ~n45420 ;
  assign n45424 = n80149 & n45423 ;
  assign n45587 = n44943 | n45423 ;
  assign n80150 = ~n45587 ;
  assign n45588 = n45545 & n80150 ;
  assign n45589 = n45424 | n45588 ;
  assign n45590 = n69851 & n45589 ;
  assign n45591 = n80142 & n45590 ;
  assign n45592 = n45586 | n45591 ;
  assign n45593 = n69075 & n45592 ;
  assign n80151 = ~n45591 ;
  assign n46078 = x100 & n80151 ;
  assign n80152 = ~n45586 ;
  assign n46079 = n80152 & n46078 ;
  assign n46080 = n45593 | n46079 ;
  assign n45594 = n44942 & n45449 ;
  assign n80153 = ~n45544 ;
  assign n45546 = n45418 & n80153 ;
  assign n45595 = n44952 | n45418 ;
  assign n80154 = ~n45595 ;
  assign n45596 = n45414 & n80154 ;
  assign n45597 = n45546 | n45596 ;
  assign n45598 = n69851 & n45597 ;
  assign n45599 = n80142 & n45598 ;
  assign n45600 = n45594 | n45599 ;
  assign n45601 = n68993 & n45600 ;
  assign n45602 = n44951 & n45449 ;
  assign n80155 = ~n45409 ;
  assign n45413 = n80155 & n45412 ;
  assign n45603 = n44961 | n45412 ;
  assign n80156 = ~n45603 ;
  assign n45604 = n45540 & n80156 ;
  assign n45605 = n45413 | n45604 ;
  assign n45606 = n69851 & n45605 ;
  assign n45607 = n80142 & n45606 ;
  assign n45608 = n45602 | n45607 ;
  assign n45609 = n68716 & n45608 ;
  assign n80157 = ~n45607 ;
  assign n46066 = x98 & n80157 ;
  assign n80158 = ~n45602 ;
  assign n46067 = n80158 & n46066 ;
  assign n46068 = n45609 | n46067 ;
  assign n45610 = n44960 & n45449 ;
  assign n80159 = ~n45539 ;
  assign n45541 = n45407 & n80159 ;
  assign n45611 = n44970 | n45407 ;
  assign n80160 = ~n45611 ;
  assign n45612 = n45403 & n80160 ;
  assign n45613 = n45541 | n45612 ;
  assign n45614 = n69851 & n45613 ;
  assign n45615 = n80142 & n45614 ;
  assign n45616 = n45610 | n45615 ;
  assign n45617 = n68545 & n45616 ;
  assign n45618 = n44969 & n45449 ;
  assign n80161 = ~n45398 ;
  assign n45402 = n80161 & n45401 ;
  assign n45619 = n44979 | n45401 ;
  assign n80162 = ~n45619 ;
  assign n45620 = n45535 & n80162 ;
  assign n45621 = n45402 | n45620 ;
  assign n45622 = n69851 & n45621 ;
  assign n45623 = n80142 & n45622 ;
  assign n45624 = n45618 | n45623 ;
  assign n45625 = n68438 & n45624 ;
  assign n80163 = ~n45623 ;
  assign n46054 = x96 & n80163 ;
  assign n80164 = ~n45618 ;
  assign n46055 = n80164 & n46054 ;
  assign n46056 = n45625 | n46055 ;
  assign n45626 = n44978 & n45449 ;
  assign n80165 = ~n45534 ;
  assign n45536 = n45396 & n80165 ;
  assign n45627 = n44988 | n45396 ;
  assign n80166 = ~n45627 ;
  assign n45628 = n45392 & n80166 ;
  assign n45629 = n45536 | n45628 ;
  assign n45630 = n69851 & n45629 ;
  assign n45631 = n80142 & n45630 ;
  assign n45632 = n45626 | n45631 ;
  assign n45633 = n68214 & n45632 ;
  assign n45634 = n44987 & n45449 ;
  assign n80167 = ~n45387 ;
  assign n45391 = n80167 & n45390 ;
  assign n45635 = n44996 | n45390 ;
  assign n80168 = ~n45635 ;
  assign n45636 = n45530 & n80168 ;
  assign n45637 = n45391 | n45636 ;
  assign n45638 = n69851 & n45637 ;
  assign n45639 = n80142 & n45638 ;
  assign n45640 = n45634 | n45639 ;
  assign n45641 = n68058 & n45640 ;
  assign n80169 = ~n45639 ;
  assign n46042 = x94 & n80169 ;
  assign n80170 = ~n45634 ;
  assign n46043 = n80170 & n46042 ;
  assign n46044 = n45641 | n46043 ;
  assign n45642 = n44995 & n45449 ;
  assign n80171 = ~n45529 ;
  assign n45531 = n45385 & n80171 ;
  assign n45643 = n45005 | n45385 ;
  assign n80172 = ~n45643 ;
  assign n45644 = n45381 & n80172 ;
  assign n45645 = n45531 | n45644 ;
  assign n45646 = n69851 & n45645 ;
  assign n45647 = n80142 & n45646 ;
  assign n45648 = n45642 | n45647 ;
  assign n45649 = n67986 & n45648 ;
  assign n45650 = n45004 & n45449 ;
  assign n80173 = ~n45376 ;
  assign n45380 = n80173 & n45379 ;
  assign n45651 = n45013 | n45379 ;
  assign n80174 = ~n45651 ;
  assign n45652 = n45525 & n80174 ;
  assign n45653 = n45380 | n45652 ;
  assign n45654 = n69851 & n45653 ;
  assign n45655 = n80142 & n45654 ;
  assign n45656 = n45650 | n45655 ;
  assign n45657 = n67763 & n45656 ;
  assign n80175 = ~n45655 ;
  assign n46030 = x92 & n80175 ;
  assign n80176 = ~n45650 ;
  assign n46031 = n80176 & n46030 ;
  assign n46032 = n45657 | n46031 ;
  assign n45658 = n45012 & n45449 ;
  assign n80177 = ~n45524 ;
  assign n45526 = n45374 & n80177 ;
  assign n45659 = n45021 | n45374 ;
  assign n80178 = ~n45659 ;
  assign n45660 = n45370 & n80178 ;
  assign n45661 = n45526 | n45660 ;
  assign n45662 = n69851 & n45661 ;
  assign n45663 = n80142 & n45662 ;
  assign n45664 = n45658 | n45663 ;
  assign n45665 = n67622 & n45664 ;
  assign n45666 = n45020 & n45449 ;
  assign n80179 = ~n45365 ;
  assign n45369 = n80179 & n45368 ;
  assign n45667 = n45030 | n45368 ;
  assign n80180 = ~n45667 ;
  assign n45668 = n45520 & n80180 ;
  assign n45669 = n45369 | n45668 ;
  assign n45670 = n69851 & n45669 ;
  assign n45671 = n80142 & n45670 ;
  assign n45672 = n45666 | n45671 ;
  assign n45673 = n67531 & n45672 ;
  assign n80181 = ~n45671 ;
  assign n46018 = x90 & n80181 ;
  assign n80182 = ~n45666 ;
  assign n46019 = n80182 & n46018 ;
  assign n46020 = n45673 | n46019 ;
  assign n45674 = n45029 & n45449 ;
  assign n80183 = ~n45519 ;
  assign n45521 = n45363 & n80183 ;
  assign n45675 = n45039 | n45363 ;
  assign n80184 = ~n45675 ;
  assign n45676 = n45359 & n80184 ;
  assign n45677 = n45521 | n45676 ;
  assign n45678 = n69851 & n45677 ;
  assign n45679 = n80142 & n45678 ;
  assign n45680 = n45674 | n45679 ;
  assign n45681 = n67348 & n45680 ;
  assign n45682 = n45038 & n45449 ;
  assign n80185 = ~n45354 ;
  assign n45358 = n80185 & n45357 ;
  assign n45683 = n45048 | n45357 ;
  assign n80186 = ~n45683 ;
  assign n45684 = n45515 & n80186 ;
  assign n45685 = n45358 | n45684 ;
  assign n45686 = n69851 & n45685 ;
  assign n45687 = n80142 & n45686 ;
  assign n45688 = n45682 | n45687 ;
  assign n45689 = n67222 & n45688 ;
  assign n80187 = ~n45687 ;
  assign n46006 = x88 & n80187 ;
  assign n80188 = ~n45682 ;
  assign n46007 = n80188 & n46006 ;
  assign n46008 = n45689 | n46007 ;
  assign n45690 = n45047 & n45449 ;
  assign n80189 = ~n45514 ;
  assign n45516 = n45352 & n80189 ;
  assign n45691 = n45057 | n45352 ;
  assign n80190 = ~n45691 ;
  assign n45692 = n45348 & n80190 ;
  assign n45693 = n45516 | n45692 ;
  assign n45694 = n69851 & n45693 ;
  assign n45695 = n80142 & n45694 ;
  assign n45696 = n45690 | n45695 ;
  assign n45697 = n67164 & n45696 ;
  assign n45698 = n45056 & n45449 ;
  assign n80191 = ~n45343 ;
  assign n45347 = n80191 & n45346 ;
  assign n45699 = n45066 | n45346 ;
  assign n80192 = ~n45699 ;
  assign n45700 = n45510 & n80192 ;
  assign n45701 = n45347 | n45700 ;
  assign n45702 = n69851 & n45701 ;
  assign n45703 = n80142 & n45702 ;
  assign n45704 = n45698 | n45703 ;
  assign n45705 = n66979 & n45704 ;
  assign n80193 = ~n45703 ;
  assign n45994 = x86 & n80193 ;
  assign n80194 = ~n45698 ;
  assign n45995 = n80194 & n45994 ;
  assign n45996 = n45705 | n45995 ;
  assign n45706 = n45065 & n45449 ;
  assign n80195 = ~n45509 ;
  assign n45511 = n45341 & n80195 ;
  assign n45707 = n45075 | n45341 ;
  assign n80196 = ~n45707 ;
  assign n45708 = n45337 & n80196 ;
  assign n45709 = n45511 | n45708 ;
  assign n45710 = n69851 & n45709 ;
  assign n45711 = n80142 & n45710 ;
  assign n45712 = n45706 | n45711 ;
  assign n45713 = n66868 & n45712 ;
  assign n45714 = n45074 & n45449 ;
  assign n80197 = ~n45332 ;
  assign n45336 = n80197 & n45335 ;
  assign n45715 = n45084 | n45335 ;
  assign n80198 = ~n45715 ;
  assign n45716 = n45505 & n80198 ;
  assign n45717 = n45336 | n45716 ;
  assign n45718 = n69851 & n45717 ;
  assign n45719 = n80142 & n45718 ;
  assign n45720 = n45714 | n45719 ;
  assign n45721 = n66797 & n45720 ;
  assign n80199 = ~n45719 ;
  assign n45982 = x84 & n80199 ;
  assign n80200 = ~n45714 ;
  assign n45983 = n80200 & n45982 ;
  assign n45984 = n45721 | n45983 ;
  assign n45722 = n45083 & n45449 ;
  assign n80201 = ~n45504 ;
  assign n45506 = n45330 & n80201 ;
  assign n45723 = n45093 | n45330 ;
  assign n80202 = ~n45723 ;
  assign n45724 = n45326 & n80202 ;
  assign n45725 = n45506 | n45724 ;
  assign n45726 = n69851 & n45725 ;
  assign n45727 = n80142 & n45726 ;
  assign n45728 = n45722 | n45727 ;
  assign n45729 = n66654 & n45728 ;
  assign n45730 = n45092 & n45449 ;
  assign n80203 = ~n45321 ;
  assign n45325 = n80203 & n45324 ;
  assign n45731 = n45102 | n45324 ;
  assign n80204 = ~n45731 ;
  assign n45732 = n45500 & n80204 ;
  assign n45733 = n45325 | n45732 ;
  assign n45734 = n69851 & n45733 ;
  assign n45735 = n80142 & n45734 ;
  assign n45736 = n45730 | n45735 ;
  assign n45737 = n66560 & n45736 ;
  assign n80205 = ~n45735 ;
  assign n45970 = x82 & n80205 ;
  assign n80206 = ~n45730 ;
  assign n45971 = n80206 & n45970 ;
  assign n45972 = n45737 | n45971 ;
  assign n45738 = n45101 & n45449 ;
  assign n80207 = ~n45499 ;
  assign n45501 = n45319 & n80207 ;
  assign n45739 = n45111 | n45319 ;
  assign n80208 = ~n45739 ;
  assign n45740 = n45315 & n80208 ;
  assign n45741 = n45501 | n45740 ;
  assign n45742 = n69851 & n45741 ;
  assign n45743 = n80142 & n45742 ;
  assign n45744 = n45738 | n45743 ;
  assign n45745 = n66505 & n45744 ;
  assign n45746 = n45110 & n45449 ;
  assign n80209 = ~n45310 ;
  assign n45314 = n80209 & n45313 ;
  assign n45747 = n45119 | n45313 ;
  assign n80210 = ~n45747 ;
  assign n45748 = n45495 & n80210 ;
  assign n45749 = n45314 | n45748 ;
  assign n45750 = n69851 & n45749 ;
  assign n45751 = n80142 & n45750 ;
  assign n45752 = n45746 | n45751 ;
  assign n45753 = n66379 & n45752 ;
  assign n80211 = ~n45751 ;
  assign n45958 = x80 & n80211 ;
  assign n80212 = ~n45746 ;
  assign n45959 = n80212 & n45958 ;
  assign n45960 = n45753 | n45959 ;
  assign n45754 = n45118 & n45449 ;
  assign n80213 = ~n45494 ;
  assign n45496 = n45308 & n80213 ;
  assign n45755 = n45128 | n45308 ;
  assign n80214 = ~n45755 ;
  assign n45756 = n45304 & n80214 ;
  assign n45757 = n45496 | n45756 ;
  assign n45758 = n69851 & n45757 ;
  assign n45759 = n80142 & n45758 ;
  assign n45760 = n45754 | n45759 ;
  assign n45761 = n66299 & n45760 ;
  assign n45762 = n45127 & n45449 ;
  assign n80215 = ~n45299 ;
  assign n45303 = n80215 & n45302 ;
  assign n45763 = n45137 | n45302 ;
  assign n80216 = ~n45763 ;
  assign n45764 = n45490 & n80216 ;
  assign n45765 = n45303 | n45764 ;
  assign n45766 = n69851 & n45765 ;
  assign n45767 = n80142 & n45766 ;
  assign n45768 = n45762 | n45767 ;
  assign n45769 = n66244 & n45768 ;
  assign n80217 = ~n45767 ;
  assign n45946 = x78 & n80217 ;
  assign n80218 = ~n45762 ;
  assign n45947 = n80218 & n45946 ;
  assign n45948 = n45769 | n45947 ;
  assign n45770 = n45136 & n45449 ;
  assign n80219 = ~n45489 ;
  assign n45491 = n45297 & n80219 ;
  assign n45771 = n45146 | n45297 ;
  assign n80220 = ~n45771 ;
  assign n45772 = n45293 & n80220 ;
  assign n45773 = n45491 | n45772 ;
  assign n45774 = n69851 & n45773 ;
  assign n45775 = n80142 & n45774 ;
  assign n45776 = n45770 | n45775 ;
  assign n45777 = n66145 & n45776 ;
  assign n45778 = n45145 & n45449 ;
  assign n80221 = ~n45288 ;
  assign n45292 = n80221 & n45291 ;
  assign n45779 = n45155 | n45291 ;
  assign n80222 = ~n45779 ;
  assign n45780 = n45485 & n80222 ;
  assign n45781 = n45292 | n45780 ;
  assign n45782 = n69851 & n45781 ;
  assign n45783 = n80142 & n45782 ;
  assign n45784 = n45778 | n45783 ;
  assign n45785 = n66081 & n45784 ;
  assign n80223 = ~n45783 ;
  assign n45934 = x76 & n80223 ;
  assign n80224 = ~n45778 ;
  assign n45935 = n80224 & n45934 ;
  assign n45936 = n45785 | n45935 ;
  assign n45786 = n45154 & n45449 ;
  assign n80225 = ~n45484 ;
  assign n45486 = n45286 & n80225 ;
  assign n45787 = n45164 | n45286 ;
  assign n80226 = ~n45787 ;
  assign n45788 = n45282 & n80226 ;
  assign n45789 = n45486 | n45788 ;
  assign n45790 = n69851 & n45789 ;
  assign n45791 = n80142 & n45790 ;
  assign n45792 = n45786 | n45791 ;
  assign n45793 = n66043 & n45792 ;
  assign n45794 = n45163 & n45449 ;
  assign n80227 = ~n45277 ;
  assign n45281 = n80227 & n45280 ;
  assign n45795 = n45173 | n45280 ;
  assign n80228 = ~n45795 ;
  assign n45796 = n45480 & n80228 ;
  assign n45797 = n45281 | n45796 ;
  assign n45798 = n69851 & n45797 ;
  assign n45799 = n80142 & n45798 ;
  assign n45800 = n45794 | n45799 ;
  assign n45801 = n65960 & n45800 ;
  assign n80229 = ~n45799 ;
  assign n45922 = x74 & n80229 ;
  assign n80230 = ~n45794 ;
  assign n45923 = n80230 & n45922 ;
  assign n45924 = n45801 | n45923 ;
  assign n45802 = n45172 & n45449 ;
  assign n80231 = ~n45479 ;
  assign n45481 = n45275 & n80231 ;
  assign n45803 = n45182 | n45275 ;
  assign n80232 = ~n45803 ;
  assign n45804 = n45271 & n80232 ;
  assign n45805 = n45481 | n45804 ;
  assign n45806 = n69851 & n45805 ;
  assign n45807 = n80142 & n45806 ;
  assign n45808 = n45802 | n45807 ;
  assign n45809 = n65909 & n45808 ;
  assign n45810 = n45181 & n45449 ;
  assign n80233 = ~n45265 ;
  assign n45269 = n80233 & n45268 ;
  assign n45270 = n45191 | n45268 ;
  assign n45811 = n45263 | n45474 ;
  assign n80234 = ~n45270 ;
  assign n45812 = n80234 & n45811 ;
  assign n45813 = n45269 | n45812 ;
  assign n45814 = n69851 & n45813 ;
  assign n45815 = n80142 & n45814 ;
  assign n45816 = n45810 | n45815 ;
  assign n45817 = n65877 & n45816 ;
  assign n80235 = ~n45815 ;
  assign n45910 = x72 & n80235 ;
  assign n80236 = ~n45810 ;
  assign n45911 = n80236 & n45910 ;
  assign n45912 = n45817 | n45911 ;
  assign n45451 = n45190 & n45449 ;
  assign n80237 = ~n45474 ;
  assign n45476 = n45263 & n80237 ;
  assign n45818 = n45256 | n45471 ;
  assign n45819 = n45200 | n45263 ;
  assign n80238 = ~n45819 ;
  assign n45820 = n45818 & n80238 ;
  assign n45821 = n45476 | n45820 ;
  assign n45822 = n69851 & n45821 ;
  assign n45823 = n80142 & n45822 ;
  assign n45824 = n45451 | n45823 ;
  assign n45825 = n65820 & n45824 ;
  assign n45452 = n45199 & n45449 ;
  assign n80239 = ~n45256 ;
  assign n45472 = n80239 & n45471 ;
  assign n45826 = n45254 | n45467 ;
  assign n45827 = n45209 | n45471 ;
  assign n80240 = ~n45827 ;
  assign n45828 = n45826 & n80240 ;
  assign n45829 = n45472 | n45828 ;
  assign n45830 = n69851 & n45829 ;
  assign n45831 = n80142 & n45830 ;
  assign n45832 = n45452 | n45831 ;
  assign n45833 = n65791 & n45832 ;
  assign n80241 = ~n45831 ;
  assign n45899 = x70 & n80241 ;
  assign n80242 = ~n45452 ;
  assign n45900 = n80242 & n45899 ;
  assign n45901 = n45833 | n45900 ;
  assign n45453 = n45208 & n45449 ;
  assign n80243 = ~n45467 ;
  assign n45469 = n45254 & n80243 ;
  assign n45834 = n45247 | n45464 ;
  assign n45835 = n45218 | n45254 ;
  assign n80244 = ~n45835 ;
  assign n45836 = n45834 & n80244 ;
  assign n45837 = n45469 | n45836 ;
  assign n45838 = n69851 & n45837 ;
  assign n45839 = n80142 & n45838 ;
  assign n45840 = n45453 | n45839 ;
  assign n45841 = n65772 & n45840 ;
  assign n45454 = n45217 & n45449 ;
  assign n80245 = ~n45247 ;
  assign n45465 = n80245 & n45464 ;
  assign n45842 = n45226 | n45464 ;
  assign n80246 = ~n45842 ;
  assign n45843 = n45246 & n80246 ;
  assign n45844 = n45465 | n45843 ;
  assign n45845 = n69851 & n45844 ;
  assign n45846 = n80142 & n45845 ;
  assign n45847 = n45454 | n45846 ;
  assign n45848 = n65746 & n45847 ;
  assign n80247 = ~n45846 ;
  assign n45889 = x68 & n80247 ;
  assign n80248 = ~n45454 ;
  assign n45890 = n80248 & n45889 ;
  assign n45891 = n45848 | n45890 ;
  assign n45456 = n45225 & n45449 ;
  assign n45849 = n45241 | n45245 ;
  assign n80249 = ~n45849 ;
  assign n45850 = n45460 & n80249 ;
  assign n80250 = ~n45461 ;
  assign n45851 = n45245 & n80250 ;
  assign n45852 = n45850 | n45851 ;
  assign n45853 = n69851 & n45852 ;
  assign n45854 = n80142 & n45853 ;
  assign n45855 = n45456 | n45854 ;
  assign n45856 = n65721 & n45855 ;
  assign n45857 = n45449 & n45457 ;
  assign n45858 = n12955 & n45238 ;
  assign n45859 = n80016 & n45858 ;
  assign n45860 = n13184 | n45859 ;
  assign n80251 = ~n45860 ;
  assign n45861 = n45460 & n80251 ;
  assign n45862 = n80142 & n45861 ;
  assign n45863 = n45857 | n45862 ;
  assign n45864 = n65686 & n45863 ;
  assign n80252 = ~n45862 ;
  assign n45879 = x66 & n80252 ;
  assign n80253 = ~n45857 ;
  assign n45880 = n80253 & n45879 ;
  assign n45881 = n45864 | n45880 ;
  assign n45865 = n80128 & n45556 ;
  assign n45866 = n45445 | n45865 ;
  assign n45867 = n80131 & n45866 ;
  assign n80254 = ~n45867 ;
  assign n45868 = n13583 & n80254 ;
  assign n80255 = ~n45868 ;
  assign n45869 = x24 & n80255 ;
  assign n45870 = n13588 & n80142 ;
  assign n45871 = n45869 | n45870 ;
  assign n45872 = x65 & n45871 ;
  assign n45873 = x65 | n45870 ;
  assign n45874 = n45869 | n45873 ;
  assign n80256 = ~n45872 ;
  assign n45875 = n80256 & n45874 ;
  assign n45877 = n13596 | n45875 ;
  assign n45878 = n65670 & n45871 ;
  assign n80257 = ~n45878 ;
  assign n45882 = n45877 & n80257 ;
  assign n45883 = n45881 | n45882 ;
  assign n80258 = ~n45864 ;
  assign n45884 = n80258 & n45883 ;
  assign n80259 = ~n45854 ;
  assign n45885 = x67 & n80259 ;
  assign n80260 = ~n45456 ;
  assign n45886 = n80260 & n45885 ;
  assign n45887 = n45856 | n45886 ;
  assign n45888 = n45884 | n45887 ;
  assign n80261 = ~n45856 ;
  assign n45892 = n80261 & n45888 ;
  assign n45893 = n45891 | n45892 ;
  assign n80262 = ~n45848 ;
  assign n45894 = n80262 & n45893 ;
  assign n80263 = ~n45839 ;
  assign n45895 = x69 & n80263 ;
  assign n80264 = ~n45453 ;
  assign n45896 = n80264 & n45895 ;
  assign n45897 = n45841 | n45896 ;
  assign n45898 = n45894 | n45897 ;
  assign n80265 = ~n45841 ;
  assign n45902 = n80265 & n45898 ;
  assign n45903 = n45901 | n45902 ;
  assign n80266 = ~n45833 ;
  assign n45904 = n80266 & n45903 ;
  assign n80267 = ~n45823 ;
  assign n45905 = x71 & n80267 ;
  assign n80268 = ~n45451 ;
  assign n45906 = n80268 & n45905 ;
  assign n45907 = n45825 | n45906 ;
  assign n45909 = n45904 | n45907 ;
  assign n80269 = ~n45825 ;
  assign n45914 = n80269 & n45909 ;
  assign n45915 = n45912 | n45914 ;
  assign n80270 = ~n45817 ;
  assign n45916 = n80270 & n45915 ;
  assign n80271 = ~n45807 ;
  assign n45917 = x73 & n80271 ;
  assign n80272 = ~n45802 ;
  assign n45918 = n80272 & n45917 ;
  assign n45919 = n45809 | n45918 ;
  assign n45921 = n45916 | n45919 ;
  assign n80273 = ~n45809 ;
  assign n45926 = n80273 & n45921 ;
  assign n45927 = n45924 | n45926 ;
  assign n80274 = ~n45801 ;
  assign n45928 = n80274 & n45927 ;
  assign n80275 = ~n45791 ;
  assign n45929 = x75 & n80275 ;
  assign n80276 = ~n45786 ;
  assign n45930 = n80276 & n45929 ;
  assign n45931 = n45793 | n45930 ;
  assign n45933 = n45928 | n45931 ;
  assign n80277 = ~n45793 ;
  assign n45938 = n80277 & n45933 ;
  assign n45939 = n45936 | n45938 ;
  assign n80278 = ~n45785 ;
  assign n45940 = n80278 & n45939 ;
  assign n80279 = ~n45775 ;
  assign n45941 = x77 & n80279 ;
  assign n80280 = ~n45770 ;
  assign n45942 = n80280 & n45941 ;
  assign n45943 = n45777 | n45942 ;
  assign n45945 = n45940 | n45943 ;
  assign n80281 = ~n45777 ;
  assign n45950 = n80281 & n45945 ;
  assign n45951 = n45948 | n45950 ;
  assign n80282 = ~n45769 ;
  assign n45952 = n80282 & n45951 ;
  assign n80283 = ~n45759 ;
  assign n45953 = x79 & n80283 ;
  assign n80284 = ~n45754 ;
  assign n45954 = n80284 & n45953 ;
  assign n45955 = n45761 | n45954 ;
  assign n45957 = n45952 | n45955 ;
  assign n80285 = ~n45761 ;
  assign n45962 = n80285 & n45957 ;
  assign n45963 = n45960 | n45962 ;
  assign n80286 = ~n45753 ;
  assign n45964 = n80286 & n45963 ;
  assign n80287 = ~n45743 ;
  assign n45965 = x81 & n80287 ;
  assign n80288 = ~n45738 ;
  assign n45966 = n80288 & n45965 ;
  assign n45967 = n45745 | n45966 ;
  assign n45969 = n45964 | n45967 ;
  assign n80289 = ~n45745 ;
  assign n45974 = n80289 & n45969 ;
  assign n45975 = n45972 | n45974 ;
  assign n80290 = ~n45737 ;
  assign n45976 = n80290 & n45975 ;
  assign n80291 = ~n45727 ;
  assign n45977 = x83 & n80291 ;
  assign n80292 = ~n45722 ;
  assign n45978 = n80292 & n45977 ;
  assign n45979 = n45729 | n45978 ;
  assign n45981 = n45976 | n45979 ;
  assign n80293 = ~n45729 ;
  assign n45986 = n80293 & n45981 ;
  assign n45987 = n45984 | n45986 ;
  assign n80294 = ~n45721 ;
  assign n45988 = n80294 & n45987 ;
  assign n80295 = ~n45711 ;
  assign n45989 = x85 & n80295 ;
  assign n80296 = ~n45706 ;
  assign n45990 = n80296 & n45989 ;
  assign n45991 = n45713 | n45990 ;
  assign n45993 = n45988 | n45991 ;
  assign n80297 = ~n45713 ;
  assign n45998 = n80297 & n45993 ;
  assign n45999 = n45996 | n45998 ;
  assign n80298 = ~n45705 ;
  assign n46000 = n80298 & n45999 ;
  assign n80299 = ~n45695 ;
  assign n46001 = x87 & n80299 ;
  assign n80300 = ~n45690 ;
  assign n46002 = n80300 & n46001 ;
  assign n46003 = n45697 | n46002 ;
  assign n46005 = n46000 | n46003 ;
  assign n80301 = ~n45697 ;
  assign n46010 = n80301 & n46005 ;
  assign n46011 = n46008 | n46010 ;
  assign n80302 = ~n45689 ;
  assign n46012 = n80302 & n46011 ;
  assign n80303 = ~n45679 ;
  assign n46013 = x89 & n80303 ;
  assign n80304 = ~n45674 ;
  assign n46014 = n80304 & n46013 ;
  assign n46015 = n45681 | n46014 ;
  assign n46017 = n46012 | n46015 ;
  assign n80305 = ~n45681 ;
  assign n46022 = n80305 & n46017 ;
  assign n46023 = n46020 | n46022 ;
  assign n80306 = ~n45673 ;
  assign n46024 = n80306 & n46023 ;
  assign n80307 = ~n45663 ;
  assign n46025 = x91 & n80307 ;
  assign n80308 = ~n45658 ;
  assign n46026 = n80308 & n46025 ;
  assign n46027 = n45665 | n46026 ;
  assign n46029 = n46024 | n46027 ;
  assign n80309 = ~n45665 ;
  assign n46034 = n80309 & n46029 ;
  assign n46035 = n46032 | n46034 ;
  assign n80310 = ~n45657 ;
  assign n46036 = n80310 & n46035 ;
  assign n80311 = ~n45647 ;
  assign n46037 = x93 & n80311 ;
  assign n80312 = ~n45642 ;
  assign n46038 = n80312 & n46037 ;
  assign n46039 = n45649 | n46038 ;
  assign n46041 = n46036 | n46039 ;
  assign n80313 = ~n45649 ;
  assign n46046 = n80313 & n46041 ;
  assign n46047 = n46044 | n46046 ;
  assign n80314 = ~n45641 ;
  assign n46048 = n80314 & n46047 ;
  assign n80315 = ~n45631 ;
  assign n46049 = x95 & n80315 ;
  assign n80316 = ~n45626 ;
  assign n46050 = n80316 & n46049 ;
  assign n46051 = n45633 | n46050 ;
  assign n46053 = n46048 | n46051 ;
  assign n80317 = ~n45633 ;
  assign n46058 = n80317 & n46053 ;
  assign n46059 = n46056 | n46058 ;
  assign n80318 = ~n45625 ;
  assign n46060 = n80318 & n46059 ;
  assign n80319 = ~n45615 ;
  assign n46061 = x97 & n80319 ;
  assign n80320 = ~n45610 ;
  assign n46062 = n80320 & n46061 ;
  assign n46063 = n45617 | n46062 ;
  assign n46065 = n46060 | n46063 ;
  assign n80321 = ~n45617 ;
  assign n46070 = n80321 & n46065 ;
  assign n46071 = n46068 | n46070 ;
  assign n80322 = ~n45609 ;
  assign n46072 = n80322 & n46071 ;
  assign n80323 = ~n45599 ;
  assign n46073 = x99 & n80323 ;
  assign n80324 = ~n45594 ;
  assign n46074 = n80324 & n46073 ;
  assign n46075 = n45601 | n46074 ;
  assign n46077 = n46072 | n46075 ;
  assign n80325 = ~n45601 ;
  assign n46082 = n80325 & n46077 ;
  assign n46083 = n46080 | n46082 ;
  assign n80326 = ~n45593 ;
  assign n46084 = n80326 & n46083 ;
  assign n80327 = ~n45583 ;
  assign n46085 = x101 & n80327 ;
  assign n80328 = ~n45578 ;
  assign n46086 = n80328 & n46085 ;
  assign n46087 = n45585 | n46086 ;
  assign n46089 = n46084 | n46087 ;
  assign n80329 = ~n45585 ;
  assign n46094 = n80329 & n46089 ;
  assign n46095 = n46092 | n46094 ;
  assign n80330 = ~n45577 ;
  assign n46096 = n80330 & n46095 ;
  assign n80331 = ~n45561 ;
  assign n46097 = x103 & n80331 ;
  assign n80332 = ~n45455 ;
  assign n46098 = n80332 & n46097 ;
  assign n46099 = n45569 | n46098 ;
  assign n46101 = n46096 | n46099 ;
  assign n80333 = ~n45569 ;
  assign n46107 = n80333 & n46101 ;
  assign n46108 = n46106 | n46107 ;
  assign n80334 = ~n45568 ;
  assign n46109 = n80334 & n46108 ;
  assign n46110 = n13820 | n46109 ;
  assign n80335 = ~n45567 ;
  assign n46112 = n80335 & n46110 ;
  assign n80336 = ~n46107 ;
  assign n46739 = n46106 & n80336 ;
  assign n46115 = n13583 & n80142 ;
  assign n80337 = ~n46115 ;
  assign n46116 = x24 & n80337 ;
  assign n46117 = n45870 | n46116 ;
  assign n46118 = x65 & n46117 ;
  assign n80338 = ~n46118 ;
  assign n46119 = n45874 & n80338 ;
  assign n46120 = n13596 | n46119 ;
  assign n46121 = n80257 & n46120 ;
  assign n46122 = n45881 | n46121 ;
  assign n46123 = n80258 & n46122 ;
  assign n46124 = n45887 | n46123 ;
  assign n46125 = n80261 & n46124 ;
  assign n46126 = n45891 | n46125 ;
  assign n46127 = n80262 & n46126 ;
  assign n46128 = n45897 | n46127 ;
  assign n46129 = n80265 & n46128 ;
  assign n46130 = n45901 | n46129 ;
  assign n46131 = n80266 & n46130 ;
  assign n46132 = n45907 | n46131 ;
  assign n46133 = n80269 & n46132 ;
  assign n46134 = n45912 | n46133 ;
  assign n46135 = n80270 & n46134 ;
  assign n46136 = n45919 | n46135 ;
  assign n46137 = n80273 & n46136 ;
  assign n46138 = n45924 | n46137 ;
  assign n46139 = n80274 & n46138 ;
  assign n46140 = n45931 | n46139 ;
  assign n46141 = n80277 & n46140 ;
  assign n46142 = n45936 | n46141 ;
  assign n46143 = n80278 & n46142 ;
  assign n46144 = n45943 | n46143 ;
  assign n46145 = n80281 & n46144 ;
  assign n46146 = n45948 | n46145 ;
  assign n46147 = n80282 & n46146 ;
  assign n46148 = n45955 | n46147 ;
  assign n46149 = n80285 & n46148 ;
  assign n46150 = n45960 | n46149 ;
  assign n46151 = n80286 & n46150 ;
  assign n46152 = n45967 | n46151 ;
  assign n46153 = n80289 & n46152 ;
  assign n46154 = n45972 | n46153 ;
  assign n46155 = n80290 & n46154 ;
  assign n46156 = n45979 | n46155 ;
  assign n46157 = n80293 & n46156 ;
  assign n46158 = n45984 | n46157 ;
  assign n46159 = n80294 & n46158 ;
  assign n46160 = n45991 | n46159 ;
  assign n46161 = n80297 & n46160 ;
  assign n46162 = n45996 | n46161 ;
  assign n46163 = n80298 & n46162 ;
  assign n46164 = n46003 | n46163 ;
  assign n46165 = n80301 & n46164 ;
  assign n46166 = n46008 | n46165 ;
  assign n46167 = n80302 & n46166 ;
  assign n46168 = n46015 | n46167 ;
  assign n46169 = n80305 & n46168 ;
  assign n46170 = n46020 | n46169 ;
  assign n46171 = n80306 & n46170 ;
  assign n46172 = n46027 | n46171 ;
  assign n46173 = n80309 & n46172 ;
  assign n46174 = n46032 | n46173 ;
  assign n46175 = n80310 & n46174 ;
  assign n46176 = n46039 | n46175 ;
  assign n46177 = n80313 & n46176 ;
  assign n46178 = n46044 | n46177 ;
  assign n46179 = n80314 & n46178 ;
  assign n46180 = n46051 | n46179 ;
  assign n46181 = n80317 & n46180 ;
  assign n46182 = n46056 | n46181 ;
  assign n46183 = n80318 & n46182 ;
  assign n46184 = n46063 | n46183 ;
  assign n46185 = n80321 & n46184 ;
  assign n46186 = n46068 | n46185 ;
  assign n46187 = n80322 & n46186 ;
  assign n46188 = n46075 | n46187 ;
  assign n46189 = n80325 & n46188 ;
  assign n46190 = n46080 | n46189 ;
  assign n46191 = n80326 & n46190 ;
  assign n46192 = n46087 | n46191 ;
  assign n46193 = n80329 & n46192 ;
  assign n46194 = n46092 | n46193 ;
  assign n46196 = n80330 & n46194 ;
  assign n46510 = n46099 | n46196 ;
  assign n46740 = n45569 | n46106 ;
  assign n80339 = ~n46740 ;
  assign n46741 = n46510 & n80339 ;
  assign n46742 = n46739 | n46741 ;
  assign n46743 = n46110 | n46742 ;
  assign n80340 = ~n46112 ;
  assign n46744 = n80340 & n46743 ;
  assign n46752 = n70059 & n46744 ;
  assign n46113 = n45562 & n46110 ;
  assign n46100 = n45577 | n46099 ;
  assign n80341 = ~n46100 ;
  assign n46195 = n80341 & n46194 ;
  assign n80342 = ~n46196 ;
  assign n46197 = n46099 & n80342 ;
  assign n46198 = n46195 | n46197 ;
  assign n46199 = n70059 & n46198 ;
  assign n80343 = ~n46109 ;
  assign n46200 = n80343 & n46199 ;
  assign n46201 = n46113 | n46200 ;
  assign n46202 = n69857 & n46201 ;
  assign n46203 = n45576 & n46110 ;
  assign n46093 = n45585 | n46092 ;
  assign n80344 = ~n46093 ;
  assign n46204 = n46089 & n80344 ;
  assign n80345 = ~n46094 ;
  assign n46205 = n46092 & n80345 ;
  assign n46206 = n46204 | n46205 ;
  assign n46207 = n70059 & n46206 ;
  assign n46208 = n80343 & n46207 ;
  assign n46209 = n46203 | n46208 ;
  assign n46210 = n69656 & n46209 ;
  assign n46211 = n45584 & n46110 ;
  assign n46088 = n45593 | n46087 ;
  assign n80346 = ~n46088 ;
  assign n46212 = n80346 & n46190 ;
  assign n80347 = ~n46191 ;
  assign n46213 = n46087 & n80347 ;
  assign n46214 = n46212 | n46213 ;
  assign n46215 = n70059 & n46214 ;
  assign n46216 = n80343 & n46215 ;
  assign n46217 = n46211 | n46216 ;
  assign n46218 = n69528 & n46217 ;
  assign n46219 = n45592 & n46110 ;
  assign n46081 = n45601 | n46080 ;
  assign n80348 = ~n46081 ;
  assign n46220 = n46077 & n80348 ;
  assign n80349 = ~n46082 ;
  assign n46221 = n46080 & n80349 ;
  assign n46222 = n46220 | n46221 ;
  assign n46223 = n70059 & n46222 ;
  assign n46224 = n80343 & n46223 ;
  assign n46225 = n46219 | n46224 ;
  assign n46226 = n69261 & n46225 ;
  assign n46227 = n45600 & n46110 ;
  assign n46076 = n45609 | n46075 ;
  assign n80350 = ~n46076 ;
  assign n46228 = n80350 & n46186 ;
  assign n80351 = ~n46187 ;
  assign n46229 = n46075 & n80351 ;
  assign n46230 = n46228 | n46229 ;
  assign n46231 = n70059 & n46230 ;
  assign n46232 = n80343 & n46231 ;
  assign n46233 = n46227 | n46232 ;
  assign n46234 = n69075 & n46233 ;
  assign n46235 = n45608 & n46110 ;
  assign n46069 = n45617 | n46068 ;
  assign n80352 = ~n46069 ;
  assign n46236 = n46065 & n80352 ;
  assign n80353 = ~n46070 ;
  assign n46237 = n46068 & n80353 ;
  assign n46238 = n46236 | n46237 ;
  assign n46239 = n70059 & n46238 ;
  assign n46240 = n80343 & n46239 ;
  assign n46241 = n46235 | n46240 ;
  assign n46242 = n68993 & n46241 ;
  assign n46243 = n45616 & n46110 ;
  assign n46064 = n45625 | n46063 ;
  assign n80354 = ~n46064 ;
  assign n46244 = n80354 & n46182 ;
  assign n80355 = ~n46183 ;
  assign n46245 = n46063 & n80355 ;
  assign n46246 = n46244 | n46245 ;
  assign n46247 = n70059 & n46246 ;
  assign n46248 = n80343 & n46247 ;
  assign n46249 = n46243 | n46248 ;
  assign n46250 = n68716 & n46249 ;
  assign n46251 = n45624 & n46110 ;
  assign n46057 = n45633 | n46056 ;
  assign n80356 = ~n46057 ;
  assign n46252 = n46053 & n80356 ;
  assign n80357 = ~n46058 ;
  assign n46253 = n46056 & n80357 ;
  assign n46254 = n46252 | n46253 ;
  assign n46255 = n70059 & n46254 ;
  assign n46256 = n80343 & n46255 ;
  assign n46257 = n46251 | n46256 ;
  assign n46258 = n68545 & n46257 ;
  assign n46259 = n45632 & n46110 ;
  assign n46052 = n45641 | n46051 ;
  assign n80358 = ~n46052 ;
  assign n46260 = n80358 & n46178 ;
  assign n80359 = ~n46179 ;
  assign n46261 = n46051 & n80359 ;
  assign n46262 = n46260 | n46261 ;
  assign n46263 = n70059 & n46262 ;
  assign n46264 = n80343 & n46263 ;
  assign n46265 = n46259 | n46264 ;
  assign n46266 = n68438 & n46265 ;
  assign n46267 = n45640 & n46110 ;
  assign n46045 = n45649 | n46044 ;
  assign n80360 = ~n46045 ;
  assign n46268 = n46041 & n80360 ;
  assign n80361 = ~n46046 ;
  assign n46269 = n46044 & n80361 ;
  assign n46270 = n46268 | n46269 ;
  assign n46271 = n70059 & n46270 ;
  assign n46272 = n80343 & n46271 ;
  assign n46273 = n46267 | n46272 ;
  assign n46274 = n68214 & n46273 ;
  assign n46275 = n45648 & n46110 ;
  assign n46040 = n45657 | n46039 ;
  assign n80362 = ~n46040 ;
  assign n46276 = n80362 & n46174 ;
  assign n80363 = ~n46175 ;
  assign n46277 = n46039 & n80363 ;
  assign n46278 = n46276 | n46277 ;
  assign n46279 = n70059 & n46278 ;
  assign n46280 = n80343 & n46279 ;
  assign n46281 = n46275 | n46280 ;
  assign n46282 = n68058 & n46281 ;
  assign n46283 = n45656 & n46110 ;
  assign n46033 = n45665 | n46032 ;
  assign n80364 = ~n46033 ;
  assign n46284 = n46029 & n80364 ;
  assign n80365 = ~n46034 ;
  assign n46285 = n46032 & n80365 ;
  assign n46286 = n46284 | n46285 ;
  assign n46287 = n70059 & n46286 ;
  assign n46288 = n80343 & n46287 ;
  assign n46289 = n46283 | n46288 ;
  assign n46290 = n67986 & n46289 ;
  assign n46291 = n45664 & n46110 ;
  assign n46028 = n45673 | n46027 ;
  assign n80366 = ~n46028 ;
  assign n46292 = n80366 & n46170 ;
  assign n80367 = ~n46171 ;
  assign n46293 = n46027 & n80367 ;
  assign n46294 = n46292 | n46293 ;
  assign n46295 = n70059 & n46294 ;
  assign n46296 = n80343 & n46295 ;
  assign n46297 = n46291 | n46296 ;
  assign n46298 = n67763 & n46297 ;
  assign n46299 = n45672 & n46110 ;
  assign n46021 = n45681 | n46020 ;
  assign n80368 = ~n46021 ;
  assign n46300 = n46017 & n80368 ;
  assign n80369 = ~n46022 ;
  assign n46301 = n46020 & n80369 ;
  assign n46302 = n46300 | n46301 ;
  assign n46303 = n70059 & n46302 ;
  assign n46304 = n80343 & n46303 ;
  assign n46305 = n46299 | n46304 ;
  assign n46306 = n67622 & n46305 ;
  assign n46307 = n45680 & n46110 ;
  assign n46016 = n45689 | n46015 ;
  assign n80370 = ~n46016 ;
  assign n46308 = n80370 & n46166 ;
  assign n80371 = ~n46167 ;
  assign n46309 = n46015 & n80371 ;
  assign n46310 = n46308 | n46309 ;
  assign n46311 = n70059 & n46310 ;
  assign n46312 = n80343 & n46311 ;
  assign n46313 = n46307 | n46312 ;
  assign n46314 = n67531 & n46313 ;
  assign n46315 = n45688 & n46110 ;
  assign n46009 = n45697 | n46008 ;
  assign n80372 = ~n46009 ;
  assign n46316 = n46005 & n80372 ;
  assign n80373 = ~n46010 ;
  assign n46317 = n46008 & n80373 ;
  assign n46318 = n46316 | n46317 ;
  assign n46319 = n70059 & n46318 ;
  assign n46320 = n80343 & n46319 ;
  assign n46321 = n46315 | n46320 ;
  assign n46322 = n67348 & n46321 ;
  assign n46323 = n45696 & n46110 ;
  assign n46004 = n45705 | n46003 ;
  assign n80374 = ~n46004 ;
  assign n46324 = n80374 & n46162 ;
  assign n80375 = ~n46163 ;
  assign n46325 = n46003 & n80375 ;
  assign n46326 = n46324 | n46325 ;
  assign n46327 = n70059 & n46326 ;
  assign n46328 = n80343 & n46327 ;
  assign n46329 = n46323 | n46328 ;
  assign n46330 = n67222 & n46329 ;
  assign n46331 = n45704 & n46110 ;
  assign n45997 = n45713 | n45996 ;
  assign n80376 = ~n45997 ;
  assign n46332 = n45993 & n80376 ;
  assign n80377 = ~n45998 ;
  assign n46333 = n45996 & n80377 ;
  assign n46334 = n46332 | n46333 ;
  assign n46335 = n70059 & n46334 ;
  assign n46336 = n80343 & n46335 ;
  assign n46337 = n46331 | n46336 ;
  assign n46338 = n67164 & n46337 ;
  assign n46339 = n45712 & n46110 ;
  assign n45992 = n45721 | n45991 ;
  assign n80378 = ~n45992 ;
  assign n46340 = n80378 & n46158 ;
  assign n80379 = ~n46159 ;
  assign n46341 = n45991 & n80379 ;
  assign n46342 = n46340 | n46341 ;
  assign n46343 = n70059 & n46342 ;
  assign n46344 = n80343 & n46343 ;
  assign n46345 = n46339 | n46344 ;
  assign n46346 = n66979 & n46345 ;
  assign n46347 = n45720 & n46110 ;
  assign n45985 = n45729 | n45984 ;
  assign n80380 = ~n45985 ;
  assign n46348 = n45981 & n80380 ;
  assign n80381 = ~n45986 ;
  assign n46349 = n45984 & n80381 ;
  assign n46350 = n46348 | n46349 ;
  assign n46351 = n70059 & n46350 ;
  assign n46352 = n80343 & n46351 ;
  assign n46353 = n46347 | n46352 ;
  assign n46354 = n66868 & n46353 ;
  assign n46355 = n45728 & n46110 ;
  assign n45980 = n45737 | n45979 ;
  assign n80382 = ~n45980 ;
  assign n46356 = n80382 & n46154 ;
  assign n80383 = ~n46155 ;
  assign n46357 = n45979 & n80383 ;
  assign n46358 = n46356 | n46357 ;
  assign n46359 = n70059 & n46358 ;
  assign n46360 = n80343 & n46359 ;
  assign n46361 = n46355 | n46360 ;
  assign n46362 = n66797 & n46361 ;
  assign n46363 = n45736 & n46110 ;
  assign n45973 = n45745 | n45972 ;
  assign n80384 = ~n45973 ;
  assign n46364 = n45969 & n80384 ;
  assign n80385 = ~n45974 ;
  assign n46365 = n45972 & n80385 ;
  assign n46366 = n46364 | n46365 ;
  assign n46367 = n70059 & n46366 ;
  assign n46368 = n80343 & n46367 ;
  assign n46369 = n46363 | n46368 ;
  assign n46370 = n66654 & n46369 ;
  assign n46371 = n45744 & n46110 ;
  assign n45968 = n45753 | n45967 ;
  assign n80386 = ~n45968 ;
  assign n46372 = n80386 & n46150 ;
  assign n80387 = ~n46151 ;
  assign n46373 = n45967 & n80387 ;
  assign n46374 = n46372 | n46373 ;
  assign n46375 = n70059 & n46374 ;
  assign n46376 = n80343 & n46375 ;
  assign n46377 = n46371 | n46376 ;
  assign n46378 = n66560 & n46377 ;
  assign n46379 = n45752 & n46110 ;
  assign n45961 = n45761 | n45960 ;
  assign n80388 = ~n45961 ;
  assign n46380 = n45957 & n80388 ;
  assign n80389 = ~n45962 ;
  assign n46381 = n45960 & n80389 ;
  assign n46382 = n46380 | n46381 ;
  assign n46383 = n70059 & n46382 ;
  assign n46384 = n80343 & n46383 ;
  assign n46385 = n46379 | n46384 ;
  assign n46386 = n66505 & n46385 ;
  assign n46387 = n45760 & n46110 ;
  assign n45956 = n45769 | n45955 ;
  assign n80390 = ~n45956 ;
  assign n46388 = n80390 & n46146 ;
  assign n80391 = ~n46147 ;
  assign n46389 = n45955 & n80391 ;
  assign n46390 = n46388 | n46389 ;
  assign n46391 = n70059 & n46390 ;
  assign n46392 = n80343 & n46391 ;
  assign n46393 = n46387 | n46392 ;
  assign n46394 = n66379 & n46393 ;
  assign n46395 = n45768 & n46110 ;
  assign n45949 = n45777 | n45948 ;
  assign n80392 = ~n45949 ;
  assign n46396 = n45945 & n80392 ;
  assign n80393 = ~n45950 ;
  assign n46397 = n45948 & n80393 ;
  assign n46398 = n46396 | n46397 ;
  assign n46399 = n70059 & n46398 ;
  assign n46400 = n80343 & n46399 ;
  assign n46401 = n46395 | n46400 ;
  assign n46402 = n66299 & n46401 ;
  assign n46403 = n45776 & n46110 ;
  assign n45944 = n45785 | n45943 ;
  assign n80394 = ~n45944 ;
  assign n46404 = n80394 & n46142 ;
  assign n80395 = ~n46143 ;
  assign n46405 = n45943 & n80395 ;
  assign n46406 = n46404 | n46405 ;
  assign n46407 = n70059 & n46406 ;
  assign n46408 = n80343 & n46407 ;
  assign n46409 = n46403 | n46408 ;
  assign n46410 = n66244 & n46409 ;
  assign n46411 = n45784 & n46110 ;
  assign n45937 = n45793 | n45936 ;
  assign n80396 = ~n45937 ;
  assign n46412 = n45933 & n80396 ;
  assign n80397 = ~n45938 ;
  assign n46413 = n45936 & n80397 ;
  assign n46414 = n46412 | n46413 ;
  assign n46415 = n70059 & n46414 ;
  assign n46416 = n80343 & n46415 ;
  assign n46417 = n46411 | n46416 ;
  assign n46418 = n66145 & n46417 ;
  assign n46419 = n45792 & n46110 ;
  assign n45932 = n45801 | n45931 ;
  assign n80398 = ~n45932 ;
  assign n46420 = n80398 & n46138 ;
  assign n80399 = ~n46139 ;
  assign n46421 = n45931 & n80399 ;
  assign n46422 = n46420 | n46421 ;
  assign n46423 = n70059 & n46422 ;
  assign n46424 = n80343 & n46423 ;
  assign n46425 = n46419 | n46424 ;
  assign n46426 = n66081 & n46425 ;
  assign n46427 = n45800 & n46110 ;
  assign n45925 = n45809 | n45924 ;
  assign n80400 = ~n45925 ;
  assign n46428 = n45921 & n80400 ;
  assign n80401 = ~n45926 ;
  assign n46429 = n45924 & n80401 ;
  assign n46430 = n46428 | n46429 ;
  assign n46431 = n70059 & n46430 ;
  assign n46432 = n80343 & n46431 ;
  assign n46433 = n46427 | n46432 ;
  assign n46434 = n66043 & n46433 ;
  assign n46435 = n45808 & n46110 ;
  assign n45920 = n45817 | n45919 ;
  assign n80402 = ~n45920 ;
  assign n46436 = n80402 & n46134 ;
  assign n80403 = ~n46135 ;
  assign n46437 = n45919 & n80403 ;
  assign n46438 = n46436 | n46437 ;
  assign n46439 = n70059 & n46438 ;
  assign n46440 = n80343 & n46439 ;
  assign n46441 = n46435 | n46440 ;
  assign n46442 = n65960 & n46441 ;
  assign n46443 = n45816 & n46110 ;
  assign n45913 = n45825 | n45912 ;
  assign n80404 = ~n45913 ;
  assign n46444 = n45909 & n80404 ;
  assign n80405 = ~n45914 ;
  assign n46445 = n45912 & n80405 ;
  assign n46446 = n46444 | n46445 ;
  assign n46447 = n70059 & n46446 ;
  assign n46448 = n80343 & n46447 ;
  assign n46449 = n46443 | n46448 ;
  assign n46450 = n65909 & n46449 ;
  assign n46451 = n45824 & n46110 ;
  assign n45908 = n45833 | n45907 ;
  assign n80406 = ~n45908 ;
  assign n46452 = n80406 & n46130 ;
  assign n80407 = ~n46131 ;
  assign n46453 = n45907 & n80407 ;
  assign n46454 = n46452 | n46453 ;
  assign n46455 = n70059 & n46454 ;
  assign n46456 = n80343 & n46455 ;
  assign n46457 = n46451 | n46456 ;
  assign n46458 = n65877 & n46457 ;
  assign n46459 = n45832 & n46110 ;
  assign n46114 = n45841 | n45901 ;
  assign n80408 = ~n46114 ;
  assign n46460 = n80408 & n46128 ;
  assign n80409 = ~n45902 ;
  assign n46461 = n45901 & n80409 ;
  assign n46462 = n46460 | n46461 ;
  assign n46463 = n70059 & n46462 ;
  assign n46464 = n80343 & n46463 ;
  assign n46465 = n46459 | n46464 ;
  assign n46466 = n65820 & n46465 ;
  assign n46467 = n45840 & n46110 ;
  assign n46468 = n45848 | n45897 ;
  assign n80410 = ~n46468 ;
  assign n46469 = n46126 & n80410 ;
  assign n80411 = ~n46127 ;
  assign n46470 = n45897 & n80411 ;
  assign n46471 = n46469 | n46470 ;
  assign n46472 = n70059 & n46471 ;
  assign n46473 = n80343 & n46472 ;
  assign n46474 = n46467 | n46473 ;
  assign n46475 = n65791 & n46474 ;
  assign n46476 = n45847 & n46110 ;
  assign n46477 = n45856 | n45891 ;
  assign n80412 = ~n46477 ;
  assign n46478 = n46124 & n80412 ;
  assign n80413 = ~n45892 ;
  assign n46479 = n45891 & n80413 ;
  assign n46480 = n46478 | n46479 ;
  assign n46481 = n70059 & n46480 ;
  assign n46482 = n80343 & n46481 ;
  assign n46483 = n46476 | n46482 ;
  assign n46484 = n65772 & n46483 ;
  assign n46485 = n45855 & n46110 ;
  assign n46486 = n45864 | n45887 ;
  assign n80414 = ~n46486 ;
  assign n46487 = n46122 & n80414 ;
  assign n80415 = ~n46123 ;
  assign n46488 = n45887 & n80415 ;
  assign n46489 = n46487 | n46488 ;
  assign n46490 = n70059 & n46489 ;
  assign n46491 = n80343 & n46490 ;
  assign n46492 = n46485 | n46491 ;
  assign n46493 = n65746 & n46492 ;
  assign n46494 = n45863 & n46110 ;
  assign n80416 = ~n46121 ;
  assign n46495 = n45881 & n80416 ;
  assign n46496 = n45878 | n45881 ;
  assign n80417 = ~n46496 ;
  assign n46497 = n46120 & n80417 ;
  assign n46498 = n46495 | n46497 ;
  assign n46499 = n70059 & n46498 ;
  assign n46500 = n80343 & n46499 ;
  assign n46501 = n46494 | n46500 ;
  assign n46502 = n65721 & n46501 ;
  assign n46111 = n45871 & n46110 ;
  assign n45876 = n13596 & n45874 ;
  assign n46503 = n45876 & n80338 ;
  assign n46504 = n13820 | n46503 ;
  assign n80418 = ~n46504 ;
  assign n46505 = n46120 & n80418 ;
  assign n46506 = n80343 & n46505 ;
  assign n46507 = n46111 | n46506 ;
  assign n46508 = n65686 & n46507 ;
  assign n46509 = n14248 & n80343 ;
  assign n46511 = n80333 & n46510 ;
  assign n46512 = n46106 | n46511 ;
  assign n46513 = n80334 & n46512 ;
  assign n80419 = ~n46513 ;
  assign n46514 = n14243 & n80419 ;
  assign n80420 = ~n46514 ;
  assign n46515 = x23 & n80420 ;
  assign n46516 = n46509 | n46515 ;
  assign n46524 = n65670 & n46516 ;
  assign n46517 = n14243 & n80343 ;
  assign n80421 = ~n46517 ;
  assign n46518 = x23 & n80421 ;
  assign n46519 = n46509 | n46518 ;
  assign n46520 = x65 & n46519 ;
  assign n46521 = x65 | n46509 ;
  assign n46522 = n46518 | n46521 ;
  assign n80422 = ~n46520 ;
  assign n46523 = n80422 & n46522 ;
  assign n46525 = n14255 | n46523 ;
  assign n80423 = ~n46524 ;
  assign n46526 = n80423 & n46525 ;
  assign n80424 = ~n46506 ;
  assign n46527 = x66 & n80424 ;
  assign n80425 = ~n46111 ;
  assign n46528 = n80425 & n46527 ;
  assign n46529 = n46526 | n46528 ;
  assign n80426 = ~n46508 ;
  assign n46530 = n80426 & n46529 ;
  assign n80427 = ~n46500 ;
  assign n46531 = x67 & n80427 ;
  assign n80428 = ~n46494 ;
  assign n46532 = n80428 & n46531 ;
  assign n46533 = n46502 | n46532 ;
  assign n46534 = n46530 | n46533 ;
  assign n80429 = ~n46502 ;
  assign n46535 = n80429 & n46534 ;
  assign n80430 = ~n46491 ;
  assign n46536 = x68 & n80430 ;
  assign n80431 = ~n46485 ;
  assign n46537 = n80431 & n46536 ;
  assign n46538 = n46493 | n46537 ;
  assign n46539 = n46535 | n46538 ;
  assign n80432 = ~n46493 ;
  assign n46540 = n80432 & n46539 ;
  assign n80433 = ~n46482 ;
  assign n46541 = x69 & n80433 ;
  assign n80434 = ~n46476 ;
  assign n46542 = n80434 & n46541 ;
  assign n46543 = n46484 | n46542 ;
  assign n46544 = n46540 | n46543 ;
  assign n80435 = ~n46484 ;
  assign n46545 = n80435 & n46544 ;
  assign n80436 = ~n46473 ;
  assign n46546 = x70 & n80436 ;
  assign n80437 = ~n46467 ;
  assign n46547 = n80437 & n46546 ;
  assign n46548 = n46475 | n46547 ;
  assign n46550 = n46545 | n46548 ;
  assign n80438 = ~n46475 ;
  assign n46551 = n80438 & n46550 ;
  assign n80439 = ~n46464 ;
  assign n46552 = x71 & n80439 ;
  assign n80440 = ~n46459 ;
  assign n46553 = n80440 & n46552 ;
  assign n46554 = n46466 | n46553 ;
  assign n46555 = n46551 | n46554 ;
  assign n80441 = ~n46466 ;
  assign n46556 = n80441 & n46555 ;
  assign n80442 = ~n46456 ;
  assign n46557 = x72 & n80442 ;
  assign n80443 = ~n46451 ;
  assign n46558 = n80443 & n46557 ;
  assign n46559 = n46458 | n46558 ;
  assign n46561 = n46556 | n46559 ;
  assign n80444 = ~n46458 ;
  assign n46562 = n80444 & n46561 ;
  assign n80445 = ~n46448 ;
  assign n46563 = x73 & n80445 ;
  assign n80446 = ~n46443 ;
  assign n46564 = n80446 & n46563 ;
  assign n46565 = n46450 | n46564 ;
  assign n46566 = n46562 | n46565 ;
  assign n80447 = ~n46450 ;
  assign n46567 = n80447 & n46566 ;
  assign n80448 = ~n46440 ;
  assign n46568 = x74 & n80448 ;
  assign n80449 = ~n46435 ;
  assign n46569 = n80449 & n46568 ;
  assign n46570 = n46442 | n46569 ;
  assign n46572 = n46567 | n46570 ;
  assign n80450 = ~n46442 ;
  assign n46573 = n80450 & n46572 ;
  assign n80451 = ~n46432 ;
  assign n46574 = x75 & n80451 ;
  assign n80452 = ~n46427 ;
  assign n46575 = n80452 & n46574 ;
  assign n46576 = n46434 | n46575 ;
  assign n46577 = n46573 | n46576 ;
  assign n80453 = ~n46434 ;
  assign n46578 = n80453 & n46577 ;
  assign n80454 = ~n46424 ;
  assign n46579 = x76 & n80454 ;
  assign n80455 = ~n46419 ;
  assign n46580 = n80455 & n46579 ;
  assign n46581 = n46426 | n46580 ;
  assign n46583 = n46578 | n46581 ;
  assign n80456 = ~n46426 ;
  assign n46584 = n80456 & n46583 ;
  assign n80457 = ~n46416 ;
  assign n46585 = x77 & n80457 ;
  assign n80458 = ~n46411 ;
  assign n46586 = n80458 & n46585 ;
  assign n46587 = n46418 | n46586 ;
  assign n46588 = n46584 | n46587 ;
  assign n80459 = ~n46418 ;
  assign n46589 = n80459 & n46588 ;
  assign n80460 = ~n46408 ;
  assign n46590 = x78 & n80460 ;
  assign n80461 = ~n46403 ;
  assign n46591 = n80461 & n46590 ;
  assign n46592 = n46410 | n46591 ;
  assign n46594 = n46589 | n46592 ;
  assign n80462 = ~n46410 ;
  assign n46595 = n80462 & n46594 ;
  assign n80463 = ~n46400 ;
  assign n46596 = x79 & n80463 ;
  assign n80464 = ~n46395 ;
  assign n46597 = n80464 & n46596 ;
  assign n46598 = n46402 | n46597 ;
  assign n46599 = n46595 | n46598 ;
  assign n80465 = ~n46402 ;
  assign n46600 = n80465 & n46599 ;
  assign n80466 = ~n46392 ;
  assign n46601 = x80 & n80466 ;
  assign n80467 = ~n46387 ;
  assign n46602 = n80467 & n46601 ;
  assign n46603 = n46394 | n46602 ;
  assign n46605 = n46600 | n46603 ;
  assign n80468 = ~n46394 ;
  assign n46606 = n80468 & n46605 ;
  assign n80469 = ~n46384 ;
  assign n46607 = x81 & n80469 ;
  assign n80470 = ~n46379 ;
  assign n46608 = n80470 & n46607 ;
  assign n46609 = n46386 | n46608 ;
  assign n46610 = n46606 | n46609 ;
  assign n80471 = ~n46386 ;
  assign n46611 = n80471 & n46610 ;
  assign n80472 = ~n46376 ;
  assign n46612 = x82 & n80472 ;
  assign n80473 = ~n46371 ;
  assign n46613 = n80473 & n46612 ;
  assign n46614 = n46378 | n46613 ;
  assign n46616 = n46611 | n46614 ;
  assign n80474 = ~n46378 ;
  assign n46617 = n80474 & n46616 ;
  assign n80475 = ~n46368 ;
  assign n46618 = x83 & n80475 ;
  assign n80476 = ~n46363 ;
  assign n46619 = n80476 & n46618 ;
  assign n46620 = n46370 | n46619 ;
  assign n46621 = n46617 | n46620 ;
  assign n80477 = ~n46370 ;
  assign n46622 = n80477 & n46621 ;
  assign n80478 = ~n46360 ;
  assign n46623 = x84 & n80478 ;
  assign n80479 = ~n46355 ;
  assign n46624 = n80479 & n46623 ;
  assign n46625 = n46362 | n46624 ;
  assign n46627 = n46622 | n46625 ;
  assign n80480 = ~n46362 ;
  assign n46628 = n80480 & n46627 ;
  assign n80481 = ~n46352 ;
  assign n46629 = x85 & n80481 ;
  assign n80482 = ~n46347 ;
  assign n46630 = n80482 & n46629 ;
  assign n46631 = n46354 | n46630 ;
  assign n46632 = n46628 | n46631 ;
  assign n80483 = ~n46354 ;
  assign n46633 = n80483 & n46632 ;
  assign n80484 = ~n46344 ;
  assign n46634 = x86 & n80484 ;
  assign n80485 = ~n46339 ;
  assign n46635 = n80485 & n46634 ;
  assign n46636 = n46346 | n46635 ;
  assign n46638 = n46633 | n46636 ;
  assign n80486 = ~n46346 ;
  assign n46639 = n80486 & n46638 ;
  assign n80487 = ~n46336 ;
  assign n46640 = x87 & n80487 ;
  assign n80488 = ~n46331 ;
  assign n46641 = n80488 & n46640 ;
  assign n46642 = n46338 | n46641 ;
  assign n46643 = n46639 | n46642 ;
  assign n80489 = ~n46338 ;
  assign n46644 = n80489 & n46643 ;
  assign n80490 = ~n46328 ;
  assign n46645 = x88 & n80490 ;
  assign n80491 = ~n46323 ;
  assign n46646 = n80491 & n46645 ;
  assign n46647 = n46330 | n46646 ;
  assign n46649 = n46644 | n46647 ;
  assign n80492 = ~n46330 ;
  assign n46650 = n80492 & n46649 ;
  assign n80493 = ~n46320 ;
  assign n46651 = x89 & n80493 ;
  assign n80494 = ~n46315 ;
  assign n46652 = n80494 & n46651 ;
  assign n46653 = n46322 | n46652 ;
  assign n46654 = n46650 | n46653 ;
  assign n80495 = ~n46322 ;
  assign n46655 = n80495 & n46654 ;
  assign n80496 = ~n46312 ;
  assign n46656 = x90 & n80496 ;
  assign n80497 = ~n46307 ;
  assign n46657 = n80497 & n46656 ;
  assign n46658 = n46314 | n46657 ;
  assign n46660 = n46655 | n46658 ;
  assign n80498 = ~n46314 ;
  assign n46661 = n80498 & n46660 ;
  assign n80499 = ~n46304 ;
  assign n46662 = x91 & n80499 ;
  assign n80500 = ~n46299 ;
  assign n46663 = n80500 & n46662 ;
  assign n46664 = n46306 | n46663 ;
  assign n46665 = n46661 | n46664 ;
  assign n80501 = ~n46306 ;
  assign n46666 = n80501 & n46665 ;
  assign n80502 = ~n46296 ;
  assign n46667 = x92 & n80502 ;
  assign n80503 = ~n46291 ;
  assign n46668 = n80503 & n46667 ;
  assign n46669 = n46298 | n46668 ;
  assign n46671 = n46666 | n46669 ;
  assign n80504 = ~n46298 ;
  assign n46672 = n80504 & n46671 ;
  assign n80505 = ~n46288 ;
  assign n46673 = x93 & n80505 ;
  assign n80506 = ~n46283 ;
  assign n46674 = n80506 & n46673 ;
  assign n46675 = n46290 | n46674 ;
  assign n46676 = n46672 | n46675 ;
  assign n80507 = ~n46290 ;
  assign n46677 = n80507 & n46676 ;
  assign n80508 = ~n46280 ;
  assign n46678 = x94 & n80508 ;
  assign n80509 = ~n46275 ;
  assign n46679 = n80509 & n46678 ;
  assign n46680 = n46282 | n46679 ;
  assign n46682 = n46677 | n46680 ;
  assign n80510 = ~n46282 ;
  assign n46683 = n80510 & n46682 ;
  assign n80511 = ~n46272 ;
  assign n46684 = x95 & n80511 ;
  assign n80512 = ~n46267 ;
  assign n46685 = n80512 & n46684 ;
  assign n46686 = n46274 | n46685 ;
  assign n46687 = n46683 | n46686 ;
  assign n80513 = ~n46274 ;
  assign n46688 = n80513 & n46687 ;
  assign n80514 = ~n46264 ;
  assign n46689 = x96 & n80514 ;
  assign n80515 = ~n46259 ;
  assign n46690 = n80515 & n46689 ;
  assign n46691 = n46266 | n46690 ;
  assign n46693 = n46688 | n46691 ;
  assign n80516 = ~n46266 ;
  assign n46694 = n80516 & n46693 ;
  assign n80517 = ~n46256 ;
  assign n46695 = x97 & n80517 ;
  assign n80518 = ~n46251 ;
  assign n46696 = n80518 & n46695 ;
  assign n46697 = n46258 | n46696 ;
  assign n46698 = n46694 | n46697 ;
  assign n80519 = ~n46258 ;
  assign n46699 = n80519 & n46698 ;
  assign n80520 = ~n46248 ;
  assign n46700 = x98 & n80520 ;
  assign n80521 = ~n46243 ;
  assign n46701 = n80521 & n46700 ;
  assign n46702 = n46250 | n46701 ;
  assign n46704 = n46699 | n46702 ;
  assign n80522 = ~n46250 ;
  assign n46705 = n80522 & n46704 ;
  assign n80523 = ~n46240 ;
  assign n46706 = x99 & n80523 ;
  assign n80524 = ~n46235 ;
  assign n46707 = n80524 & n46706 ;
  assign n46708 = n46242 | n46707 ;
  assign n46709 = n46705 | n46708 ;
  assign n80525 = ~n46242 ;
  assign n46710 = n80525 & n46709 ;
  assign n80526 = ~n46232 ;
  assign n46711 = x100 & n80526 ;
  assign n80527 = ~n46227 ;
  assign n46712 = n80527 & n46711 ;
  assign n46713 = n46234 | n46712 ;
  assign n46715 = n46710 | n46713 ;
  assign n80528 = ~n46234 ;
  assign n46716 = n80528 & n46715 ;
  assign n80529 = ~n46224 ;
  assign n46717 = x101 & n80529 ;
  assign n80530 = ~n46219 ;
  assign n46718 = n80530 & n46717 ;
  assign n46719 = n46226 | n46718 ;
  assign n46720 = n46716 | n46719 ;
  assign n80531 = ~n46226 ;
  assign n46721 = n80531 & n46720 ;
  assign n80532 = ~n46216 ;
  assign n46722 = x102 & n80532 ;
  assign n80533 = ~n46211 ;
  assign n46723 = n80533 & n46722 ;
  assign n46724 = n46218 | n46723 ;
  assign n46726 = n46721 | n46724 ;
  assign n80534 = ~n46218 ;
  assign n46727 = n80534 & n46726 ;
  assign n80535 = ~n46208 ;
  assign n46728 = x103 & n80535 ;
  assign n80536 = ~n46203 ;
  assign n46729 = n80536 & n46728 ;
  assign n46730 = n46210 | n46729 ;
  assign n46731 = n46727 | n46730 ;
  assign n80537 = ~n46210 ;
  assign n46732 = n80537 & n46731 ;
  assign n80538 = ~n46200 ;
  assign n46733 = x104 & n80538 ;
  assign n80539 = ~n46113 ;
  assign n46734 = n80539 & n46733 ;
  assign n46735 = n46202 | n46734 ;
  assign n46737 = n46732 | n46735 ;
  assign n80540 = ~n46202 ;
  assign n46738 = n80540 & n46737 ;
  assign n46745 = n70176 & n46744 ;
  assign n80541 = ~n46110 ;
  assign n46746 = n80541 & n46742 ;
  assign n46747 = n45567 & n46110 ;
  assign n80542 = ~n46747 ;
  assign n46748 = x105 & n80542 ;
  assign n80543 = ~n46746 ;
  assign n46749 = n80543 & n46748 ;
  assign n46750 = n14472 | n46749 ;
  assign n46751 = n46745 | n46750 ;
  assign n46753 = n46738 | n46751 ;
  assign n80544 = ~n46752 ;
  assign n46754 = n80544 & n46753 ;
  assign n46869 = n46202 | n46749 ;
  assign n46870 = n46745 | n46869 ;
  assign n80545 = ~n46870 ;
  assign n46871 = n46737 & n80545 ;
  assign n46757 = x65 & n46516 ;
  assign n80546 = ~n46757 ;
  assign n46758 = n46522 & n80546 ;
  assign n46759 = n14255 | n46758 ;
  assign n46760 = n80423 & n46759 ;
  assign n46761 = n46508 | n46528 ;
  assign n46763 = n46760 | n46761 ;
  assign n46764 = n80426 & n46763 ;
  assign n46765 = n46532 | n46764 ;
  assign n46767 = n80429 & n46765 ;
  assign n46769 = n46538 | n46767 ;
  assign n46770 = n80432 & n46769 ;
  assign n46772 = n46543 | n46770 ;
  assign n46773 = n80435 & n46772 ;
  assign n46774 = n46548 | n46773 ;
  assign n46775 = n80438 & n46774 ;
  assign n46776 = n46554 | n46775 ;
  assign n46778 = n80441 & n46776 ;
  assign n46779 = n46559 | n46778 ;
  assign n46780 = n80444 & n46779 ;
  assign n46781 = n46565 | n46780 ;
  assign n46783 = n80447 & n46781 ;
  assign n46784 = n46570 | n46783 ;
  assign n46785 = n80450 & n46784 ;
  assign n46786 = n46576 | n46785 ;
  assign n46788 = n80453 & n46786 ;
  assign n46789 = n46581 | n46788 ;
  assign n46790 = n80456 & n46789 ;
  assign n46791 = n46587 | n46790 ;
  assign n46793 = n80459 & n46791 ;
  assign n46794 = n46592 | n46793 ;
  assign n46795 = n80462 & n46794 ;
  assign n46796 = n46598 | n46795 ;
  assign n46798 = n80465 & n46796 ;
  assign n46799 = n46603 | n46798 ;
  assign n46800 = n80468 & n46799 ;
  assign n46801 = n46609 | n46800 ;
  assign n46803 = n80471 & n46801 ;
  assign n46804 = n46614 | n46803 ;
  assign n46805 = n80474 & n46804 ;
  assign n46806 = n46620 | n46805 ;
  assign n46808 = n80477 & n46806 ;
  assign n46809 = n46625 | n46808 ;
  assign n46810 = n80480 & n46809 ;
  assign n46811 = n46631 | n46810 ;
  assign n46813 = n80483 & n46811 ;
  assign n46814 = n46636 | n46813 ;
  assign n46815 = n80486 & n46814 ;
  assign n46816 = n46642 | n46815 ;
  assign n46818 = n80489 & n46816 ;
  assign n46819 = n46647 | n46818 ;
  assign n46820 = n80492 & n46819 ;
  assign n46821 = n46653 | n46820 ;
  assign n46823 = n80495 & n46821 ;
  assign n46824 = n46658 | n46823 ;
  assign n46825 = n80498 & n46824 ;
  assign n46826 = n46664 | n46825 ;
  assign n46828 = n80501 & n46826 ;
  assign n46829 = n46669 | n46828 ;
  assign n46830 = n80504 & n46829 ;
  assign n46831 = n46675 | n46830 ;
  assign n46833 = n80507 & n46831 ;
  assign n46834 = n46680 | n46833 ;
  assign n46835 = n80510 & n46834 ;
  assign n46836 = n46686 | n46835 ;
  assign n46838 = n80513 & n46836 ;
  assign n46839 = n46691 | n46838 ;
  assign n46840 = n80516 & n46839 ;
  assign n46841 = n46697 | n46840 ;
  assign n46843 = n80519 & n46841 ;
  assign n46844 = n46702 | n46843 ;
  assign n46845 = n80522 & n46844 ;
  assign n46846 = n46708 | n46845 ;
  assign n46848 = n80525 & n46846 ;
  assign n46849 = n46713 | n46848 ;
  assign n46850 = n80528 & n46849 ;
  assign n46851 = n46719 | n46850 ;
  assign n46853 = n80531 & n46851 ;
  assign n46854 = n46724 | n46853 ;
  assign n46855 = n80534 & n46854 ;
  assign n46856 = n46730 | n46855 ;
  assign n46862 = n80537 & n46856 ;
  assign n46863 = n46735 | n46862 ;
  assign n46864 = n80540 & n46863 ;
  assign n46872 = n46745 | n46749 ;
  assign n80547 = ~n46864 ;
  assign n46873 = n80547 & n46872 ;
  assign n46874 = n46871 | n46873 ;
  assign n80548 = ~n46754 ;
  assign n46875 = n80548 & n46874 ;
  assign n46865 = n46751 | n46864 ;
  assign n46876 = n13820 & n45567 ;
  assign n46877 = n46865 & n46876 ;
  assign n46878 = n46875 | n46877 ;
  assign n46879 = n70276 & n46878 ;
  assign n80549 = ~n46877 ;
  assign n47442 = x106 & n80549 ;
  assign n80550 = ~n46875 ;
  assign n47443 = n80550 & n47442 ;
  assign n47444 = n46879 | n47443 ;
  assign n80551 = ~n46732 ;
  assign n46736 = n80551 & n46735 ;
  assign n46858 = n46210 | n46735 ;
  assign n80552 = ~n46858 ;
  assign n46859 = n46856 & n80552 ;
  assign n46860 = n46736 | n46859 ;
  assign n46861 = n80548 & n46860 ;
  assign n46866 = n46201 & n80544 ;
  assign n46867 = n46865 & n46866 ;
  assign n46868 = n46861 | n46867 ;
  assign n46880 = n70176 & n46868 ;
  assign n80553 = ~n46855 ;
  assign n46857 = n46730 & n80553 ;
  assign n46881 = n46218 | n46730 ;
  assign n80554 = ~n46881 ;
  assign n46882 = n46726 & n80554 ;
  assign n46883 = n46857 | n46882 ;
  assign n46884 = n80548 & n46883 ;
  assign n46885 = n46209 & n80544 ;
  assign n46886 = n46865 & n46885 ;
  assign n46887 = n46884 | n46886 ;
  assign n46888 = n69857 & n46887 ;
  assign n80555 = ~n46886 ;
  assign n47430 = x104 & n80555 ;
  assign n80556 = ~n46884 ;
  assign n47431 = n80556 & n47430 ;
  assign n47432 = n46888 | n47431 ;
  assign n80557 = ~n46721 ;
  assign n46725 = n80557 & n46724 ;
  assign n46889 = n46226 | n46724 ;
  assign n80558 = ~n46889 ;
  assign n46890 = n46851 & n80558 ;
  assign n46891 = n46725 | n46890 ;
  assign n46892 = n80548 & n46891 ;
  assign n46893 = n46217 & n80544 ;
  assign n46894 = n46865 & n46893 ;
  assign n46895 = n46892 | n46894 ;
  assign n46896 = n69656 & n46895 ;
  assign n80559 = ~n46850 ;
  assign n46852 = n46719 & n80559 ;
  assign n46897 = n46234 | n46719 ;
  assign n80560 = ~n46897 ;
  assign n46898 = n46715 & n80560 ;
  assign n46899 = n46852 | n46898 ;
  assign n46900 = n80548 & n46899 ;
  assign n46901 = n46225 & n80544 ;
  assign n46902 = n46865 & n46901 ;
  assign n46903 = n46900 | n46902 ;
  assign n46904 = n69528 & n46903 ;
  assign n80561 = ~n46902 ;
  assign n47418 = x102 & n80561 ;
  assign n80562 = ~n46900 ;
  assign n47419 = n80562 & n47418 ;
  assign n47420 = n46904 | n47419 ;
  assign n80563 = ~n46710 ;
  assign n46714 = n80563 & n46713 ;
  assign n46905 = n46242 | n46713 ;
  assign n80564 = ~n46905 ;
  assign n46906 = n46846 & n80564 ;
  assign n46907 = n46714 | n46906 ;
  assign n46908 = n80548 & n46907 ;
  assign n46909 = n46233 & n80544 ;
  assign n46910 = n46865 & n46909 ;
  assign n46911 = n46908 | n46910 ;
  assign n46912 = n69261 & n46911 ;
  assign n80565 = ~n46845 ;
  assign n46847 = n46708 & n80565 ;
  assign n46913 = n46250 | n46708 ;
  assign n80566 = ~n46913 ;
  assign n46914 = n46704 & n80566 ;
  assign n46915 = n46847 | n46914 ;
  assign n46916 = n80548 & n46915 ;
  assign n46917 = n46241 & n80544 ;
  assign n46918 = n46865 & n46917 ;
  assign n46919 = n46916 | n46918 ;
  assign n46920 = n69075 & n46919 ;
  assign n80567 = ~n46918 ;
  assign n47406 = x100 & n80567 ;
  assign n80568 = ~n46916 ;
  assign n47407 = n80568 & n47406 ;
  assign n47408 = n46920 | n47407 ;
  assign n80569 = ~n46699 ;
  assign n46703 = n80569 & n46702 ;
  assign n46921 = n46258 | n46702 ;
  assign n80570 = ~n46921 ;
  assign n46922 = n46841 & n80570 ;
  assign n46923 = n46703 | n46922 ;
  assign n46924 = n80548 & n46923 ;
  assign n46925 = n46249 & n80544 ;
  assign n46926 = n46865 & n46925 ;
  assign n46927 = n46924 | n46926 ;
  assign n46928 = n68993 & n46927 ;
  assign n80571 = ~n46840 ;
  assign n46842 = n46697 & n80571 ;
  assign n46929 = n46266 | n46697 ;
  assign n80572 = ~n46929 ;
  assign n46930 = n46693 & n80572 ;
  assign n46931 = n46842 | n46930 ;
  assign n46932 = n80548 & n46931 ;
  assign n46933 = n46257 & n80544 ;
  assign n46934 = n46865 & n46933 ;
  assign n46935 = n46932 | n46934 ;
  assign n46936 = n68716 & n46935 ;
  assign n80573 = ~n46934 ;
  assign n47394 = x98 & n80573 ;
  assign n80574 = ~n46932 ;
  assign n47395 = n80574 & n47394 ;
  assign n47396 = n46936 | n47395 ;
  assign n80575 = ~n46688 ;
  assign n46692 = n80575 & n46691 ;
  assign n46937 = n46274 | n46691 ;
  assign n80576 = ~n46937 ;
  assign n46938 = n46836 & n80576 ;
  assign n46939 = n46692 | n46938 ;
  assign n46940 = n80548 & n46939 ;
  assign n46941 = n46265 & n80544 ;
  assign n46942 = n46865 & n46941 ;
  assign n46943 = n46940 | n46942 ;
  assign n46944 = n68545 & n46943 ;
  assign n80577 = ~n46835 ;
  assign n46837 = n46686 & n80577 ;
  assign n46945 = n46282 | n46686 ;
  assign n80578 = ~n46945 ;
  assign n46946 = n46682 & n80578 ;
  assign n46947 = n46837 | n46946 ;
  assign n46948 = n80548 & n46947 ;
  assign n46949 = n46273 & n80544 ;
  assign n46950 = n46865 & n46949 ;
  assign n46951 = n46948 | n46950 ;
  assign n46952 = n68438 & n46951 ;
  assign n80579 = ~n46950 ;
  assign n47382 = x96 & n80579 ;
  assign n80580 = ~n46948 ;
  assign n47383 = n80580 & n47382 ;
  assign n47384 = n46952 | n47383 ;
  assign n80581 = ~n46677 ;
  assign n46681 = n80581 & n46680 ;
  assign n46953 = n46290 | n46680 ;
  assign n80582 = ~n46953 ;
  assign n46954 = n46831 & n80582 ;
  assign n46955 = n46681 | n46954 ;
  assign n46956 = n80548 & n46955 ;
  assign n46957 = n46281 & n80544 ;
  assign n46958 = n46865 & n46957 ;
  assign n46959 = n46956 | n46958 ;
  assign n46960 = n68214 & n46959 ;
  assign n80583 = ~n46830 ;
  assign n46832 = n46675 & n80583 ;
  assign n46961 = n46298 | n46675 ;
  assign n80584 = ~n46961 ;
  assign n46962 = n46671 & n80584 ;
  assign n46963 = n46832 | n46962 ;
  assign n46964 = n80548 & n46963 ;
  assign n46965 = n46289 & n80544 ;
  assign n46966 = n46865 & n46965 ;
  assign n46967 = n46964 | n46966 ;
  assign n46968 = n68058 & n46967 ;
  assign n80585 = ~n46966 ;
  assign n47370 = x94 & n80585 ;
  assign n80586 = ~n46964 ;
  assign n47371 = n80586 & n47370 ;
  assign n47372 = n46968 | n47371 ;
  assign n80587 = ~n46666 ;
  assign n46670 = n80587 & n46669 ;
  assign n46969 = n46306 | n46669 ;
  assign n80588 = ~n46969 ;
  assign n46970 = n46826 & n80588 ;
  assign n46971 = n46670 | n46970 ;
  assign n46972 = n80548 & n46971 ;
  assign n46973 = n46297 & n80544 ;
  assign n46974 = n46865 & n46973 ;
  assign n46975 = n46972 | n46974 ;
  assign n46976 = n67986 & n46975 ;
  assign n80589 = ~n46825 ;
  assign n46827 = n46664 & n80589 ;
  assign n46977 = n46314 | n46664 ;
  assign n80590 = ~n46977 ;
  assign n46978 = n46660 & n80590 ;
  assign n46979 = n46827 | n46978 ;
  assign n46980 = n80548 & n46979 ;
  assign n46981 = n46305 & n80544 ;
  assign n46982 = n46865 & n46981 ;
  assign n46983 = n46980 | n46982 ;
  assign n46984 = n67763 & n46983 ;
  assign n80591 = ~n46982 ;
  assign n47358 = x92 & n80591 ;
  assign n80592 = ~n46980 ;
  assign n47359 = n80592 & n47358 ;
  assign n47360 = n46984 | n47359 ;
  assign n80593 = ~n46655 ;
  assign n46659 = n80593 & n46658 ;
  assign n46985 = n46322 | n46658 ;
  assign n80594 = ~n46985 ;
  assign n46986 = n46821 & n80594 ;
  assign n46987 = n46659 | n46986 ;
  assign n46988 = n80548 & n46987 ;
  assign n46989 = n46313 & n80544 ;
  assign n46990 = n46865 & n46989 ;
  assign n46991 = n46988 | n46990 ;
  assign n46992 = n67622 & n46991 ;
  assign n80595 = ~n46820 ;
  assign n46822 = n46653 & n80595 ;
  assign n46993 = n46330 | n46653 ;
  assign n80596 = ~n46993 ;
  assign n46994 = n46649 & n80596 ;
  assign n46995 = n46822 | n46994 ;
  assign n46996 = n80548 & n46995 ;
  assign n46997 = n46321 & n80544 ;
  assign n46998 = n46865 & n46997 ;
  assign n46999 = n46996 | n46998 ;
  assign n47000 = n67531 & n46999 ;
  assign n80597 = ~n46998 ;
  assign n47346 = x90 & n80597 ;
  assign n80598 = ~n46996 ;
  assign n47347 = n80598 & n47346 ;
  assign n47348 = n47000 | n47347 ;
  assign n80599 = ~n46644 ;
  assign n46648 = n80599 & n46647 ;
  assign n47001 = n46338 | n46647 ;
  assign n80600 = ~n47001 ;
  assign n47002 = n46816 & n80600 ;
  assign n47003 = n46648 | n47002 ;
  assign n47004 = n80548 & n47003 ;
  assign n47005 = n46329 & n80544 ;
  assign n47006 = n46865 & n47005 ;
  assign n47007 = n47004 | n47006 ;
  assign n47008 = n67348 & n47007 ;
  assign n80601 = ~n46815 ;
  assign n46817 = n46642 & n80601 ;
  assign n47009 = n46346 | n46642 ;
  assign n80602 = ~n47009 ;
  assign n47010 = n46638 & n80602 ;
  assign n47011 = n46817 | n47010 ;
  assign n47012 = n80548 & n47011 ;
  assign n47013 = n46337 & n80544 ;
  assign n47014 = n46865 & n47013 ;
  assign n47015 = n47012 | n47014 ;
  assign n47016 = n67222 & n47015 ;
  assign n80603 = ~n47014 ;
  assign n47334 = x88 & n80603 ;
  assign n80604 = ~n47012 ;
  assign n47335 = n80604 & n47334 ;
  assign n47336 = n47016 | n47335 ;
  assign n80605 = ~n46633 ;
  assign n46637 = n80605 & n46636 ;
  assign n47017 = n46354 | n46636 ;
  assign n80606 = ~n47017 ;
  assign n47018 = n46811 & n80606 ;
  assign n47019 = n46637 | n47018 ;
  assign n47020 = n80548 & n47019 ;
  assign n47021 = n46345 & n80544 ;
  assign n47022 = n46865 & n47021 ;
  assign n47023 = n47020 | n47022 ;
  assign n47024 = n67164 & n47023 ;
  assign n80607 = ~n46810 ;
  assign n46812 = n46631 & n80607 ;
  assign n47025 = n46362 | n46631 ;
  assign n80608 = ~n47025 ;
  assign n47026 = n46627 & n80608 ;
  assign n47027 = n46812 | n47026 ;
  assign n47028 = n80548 & n47027 ;
  assign n47029 = n46353 & n80544 ;
  assign n47030 = n46865 & n47029 ;
  assign n47031 = n47028 | n47030 ;
  assign n47032 = n66979 & n47031 ;
  assign n80609 = ~n47030 ;
  assign n47322 = x86 & n80609 ;
  assign n80610 = ~n47028 ;
  assign n47323 = n80610 & n47322 ;
  assign n47324 = n47032 | n47323 ;
  assign n80611 = ~n46622 ;
  assign n46626 = n80611 & n46625 ;
  assign n47033 = n46370 | n46625 ;
  assign n80612 = ~n47033 ;
  assign n47034 = n46806 & n80612 ;
  assign n47035 = n46626 | n47034 ;
  assign n47036 = n80548 & n47035 ;
  assign n47037 = n46361 & n80544 ;
  assign n47038 = n46865 & n47037 ;
  assign n47039 = n47036 | n47038 ;
  assign n47040 = n66868 & n47039 ;
  assign n80613 = ~n46805 ;
  assign n46807 = n46620 & n80613 ;
  assign n47041 = n46378 | n46620 ;
  assign n80614 = ~n47041 ;
  assign n47042 = n46616 & n80614 ;
  assign n47043 = n46807 | n47042 ;
  assign n47044 = n80548 & n47043 ;
  assign n47045 = n46369 & n80544 ;
  assign n47046 = n46865 & n47045 ;
  assign n47047 = n47044 | n47046 ;
  assign n47048 = n66797 & n47047 ;
  assign n80615 = ~n47046 ;
  assign n47310 = x84 & n80615 ;
  assign n80616 = ~n47044 ;
  assign n47311 = n80616 & n47310 ;
  assign n47312 = n47048 | n47311 ;
  assign n80617 = ~n46611 ;
  assign n46615 = n80617 & n46614 ;
  assign n47049 = n46386 | n46614 ;
  assign n80618 = ~n47049 ;
  assign n47050 = n46801 & n80618 ;
  assign n47051 = n46615 | n47050 ;
  assign n47052 = n80548 & n47051 ;
  assign n47053 = n46377 & n80544 ;
  assign n47054 = n46865 & n47053 ;
  assign n47055 = n47052 | n47054 ;
  assign n47056 = n66654 & n47055 ;
  assign n80619 = ~n46800 ;
  assign n46802 = n46609 & n80619 ;
  assign n47057 = n46394 | n46609 ;
  assign n80620 = ~n47057 ;
  assign n47058 = n46605 & n80620 ;
  assign n47059 = n46802 | n47058 ;
  assign n47060 = n80548 & n47059 ;
  assign n47061 = n46385 & n80544 ;
  assign n47062 = n46865 & n47061 ;
  assign n47063 = n47060 | n47062 ;
  assign n47064 = n66560 & n47063 ;
  assign n80621 = ~n47062 ;
  assign n47298 = x82 & n80621 ;
  assign n80622 = ~n47060 ;
  assign n47299 = n80622 & n47298 ;
  assign n47300 = n47064 | n47299 ;
  assign n80623 = ~n46600 ;
  assign n46604 = n80623 & n46603 ;
  assign n47065 = n46402 | n46603 ;
  assign n80624 = ~n47065 ;
  assign n47066 = n46796 & n80624 ;
  assign n47067 = n46604 | n47066 ;
  assign n47068 = n80548 & n47067 ;
  assign n47069 = n46393 & n80544 ;
  assign n47070 = n46865 & n47069 ;
  assign n47071 = n47068 | n47070 ;
  assign n47072 = n66505 & n47071 ;
  assign n80625 = ~n46795 ;
  assign n46797 = n46598 & n80625 ;
  assign n47073 = n46410 | n46598 ;
  assign n80626 = ~n47073 ;
  assign n47074 = n46594 & n80626 ;
  assign n47075 = n46797 | n47074 ;
  assign n47076 = n80548 & n47075 ;
  assign n47077 = n46401 & n80544 ;
  assign n47078 = n46865 & n47077 ;
  assign n47079 = n47076 | n47078 ;
  assign n47080 = n66379 & n47079 ;
  assign n80627 = ~n47078 ;
  assign n47286 = x80 & n80627 ;
  assign n80628 = ~n47076 ;
  assign n47287 = n80628 & n47286 ;
  assign n47288 = n47080 | n47287 ;
  assign n80629 = ~n46589 ;
  assign n46593 = n80629 & n46592 ;
  assign n47081 = n46418 | n46592 ;
  assign n80630 = ~n47081 ;
  assign n47082 = n46791 & n80630 ;
  assign n47083 = n46593 | n47082 ;
  assign n47084 = n80548 & n47083 ;
  assign n47085 = n46409 & n80544 ;
  assign n47086 = n46865 & n47085 ;
  assign n47087 = n47084 | n47086 ;
  assign n47088 = n66299 & n47087 ;
  assign n80631 = ~n46790 ;
  assign n46792 = n46587 & n80631 ;
  assign n47089 = n46426 | n46587 ;
  assign n80632 = ~n47089 ;
  assign n47090 = n46583 & n80632 ;
  assign n47091 = n46792 | n47090 ;
  assign n47092 = n80548 & n47091 ;
  assign n47093 = n46417 & n80544 ;
  assign n47094 = n46865 & n47093 ;
  assign n47095 = n47092 | n47094 ;
  assign n47096 = n66244 & n47095 ;
  assign n80633 = ~n47094 ;
  assign n47274 = x78 & n80633 ;
  assign n80634 = ~n47092 ;
  assign n47275 = n80634 & n47274 ;
  assign n47276 = n47096 | n47275 ;
  assign n80635 = ~n46578 ;
  assign n46582 = n80635 & n46581 ;
  assign n47097 = n46434 | n46581 ;
  assign n80636 = ~n47097 ;
  assign n47098 = n46786 & n80636 ;
  assign n47099 = n46582 | n47098 ;
  assign n47100 = n80548 & n47099 ;
  assign n47101 = n46425 & n80544 ;
  assign n47102 = n46865 & n47101 ;
  assign n47103 = n47100 | n47102 ;
  assign n47104 = n66145 & n47103 ;
  assign n80637 = ~n46785 ;
  assign n46787 = n46576 & n80637 ;
  assign n47105 = n46442 | n46576 ;
  assign n80638 = ~n47105 ;
  assign n47106 = n46572 & n80638 ;
  assign n47107 = n46787 | n47106 ;
  assign n47108 = n80548 & n47107 ;
  assign n47109 = n46433 & n80544 ;
  assign n47110 = n46865 & n47109 ;
  assign n47111 = n47108 | n47110 ;
  assign n47112 = n66081 & n47111 ;
  assign n80639 = ~n47110 ;
  assign n47262 = x76 & n80639 ;
  assign n80640 = ~n47108 ;
  assign n47263 = n80640 & n47262 ;
  assign n47264 = n47112 | n47263 ;
  assign n80641 = ~n46567 ;
  assign n46571 = n80641 & n46570 ;
  assign n47113 = n46450 | n46570 ;
  assign n80642 = ~n47113 ;
  assign n47114 = n46781 & n80642 ;
  assign n47115 = n46571 | n47114 ;
  assign n47116 = n80548 & n47115 ;
  assign n47117 = n46441 & n80544 ;
  assign n47118 = n46865 & n47117 ;
  assign n47119 = n47116 | n47118 ;
  assign n47120 = n66043 & n47119 ;
  assign n80643 = ~n46780 ;
  assign n46782 = n46565 & n80643 ;
  assign n47121 = n46458 | n46565 ;
  assign n80644 = ~n47121 ;
  assign n47122 = n46561 & n80644 ;
  assign n47123 = n46782 | n47122 ;
  assign n47124 = n80548 & n47123 ;
  assign n47125 = n46449 & n80544 ;
  assign n47126 = n46865 & n47125 ;
  assign n47127 = n47124 | n47126 ;
  assign n47128 = n65960 & n47127 ;
  assign n80645 = ~n47126 ;
  assign n47250 = x74 & n80645 ;
  assign n80646 = ~n47124 ;
  assign n47251 = n80646 & n47250 ;
  assign n47252 = n47128 | n47251 ;
  assign n80647 = ~n46556 ;
  assign n46560 = n80647 & n46559 ;
  assign n47129 = n46466 | n46559 ;
  assign n80648 = ~n47129 ;
  assign n47130 = n46776 & n80648 ;
  assign n47131 = n46560 | n47130 ;
  assign n47132 = n80548 & n47131 ;
  assign n47133 = n46457 & n80544 ;
  assign n47134 = n46865 & n47133 ;
  assign n47135 = n47132 | n47134 ;
  assign n47136 = n65909 & n47135 ;
  assign n80649 = ~n46775 ;
  assign n46777 = n46554 & n80649 ;
  assign n47137 = n46475 | n46554 ;
  assign n80650 = ~n47137 ;
  assign n47138 = n46550 & n80650 ;
  assign n47139 = n46777 | n47138 ;
  assign n47140 = n80548 & n47139 ;
  assign n47141 = n46465 & n80544 ;
  assign n47142 = n46865 & n47141 ;
  assign n47143 = n47140 | n47142 ;
  assign n47144 = n65877 & n47143 ;
  assign n80651 = ~n47142 ;
  assign n47238 = x72 & n80651 ;
  assign n80652 = ~n47140 ;
  assign n47239 = n80652 & n47238 ;
  assign n47240 = n47144 | n47239 ;
  assign n80653 = ~n46545 ;
  assign n46549 = n80653 & n46548 ;
  assign n47145 = n46484 | n46548 ;
  assign n80654 = ~n47145 ;
  assign n47146 = n46772 & n80654 ;
  assign n47147 = n46549 | n47146 ;
  assign n47148 = n80548 & n47147 ;
  assign n47149 = n46474 & n80544 ;
  assign n47150 = n46865 & n47149 ;
  assign n47151 = n47148 | n47150 ;
  assign n47152 = n65820 & n47151 ;
  assign n80655 = ~n46770 ;
  assign n46771 = n46543 & n80655 ;
  assign n47153 = n46493 | n46543 ;
  assign n80656 = ~n47153 ;
  assign n47154 = n46539 & n80656 ;
  assign n47155 = n46771 | n47154 ;
  assign n47156 = n80548 & n47155 ;
  assign n47157 = n46483 & n80544 ;
  assign n47158 = n46865 & n47157 ;
  assign n47159 = n47156 | n47158 ;
  assign n47160 = n65791 & n47159 ;
  assign n80657 = ~n47158 ;
  assign n47226 = x70 & n80657 ;
  assign n80658 = ~n47156 ;
  assign n47227 = n80658 & n47226 ;
  assign n47228 = n47160 | n47227 ;
  assign n80659 = ~n46535 ;
  assign n46768 = n80659 & n46538 ;
  assign n47161 = n46533 | n46764 ;
  assign n47162 = n46502 | n46538 ;
  assign n80660 = ~n47162 ;
  assign n47163 = n47161 & n80660 ;
  assign n47164 = n46768 | n47163 ;
  assign n47165 = n80548 & n47164 ;
  assign n47166 = n46492 & n80544 ;
  assign n47167 = n46865 & n47166 ;
  assign n47168 = n47165 | n47167 ;
  assign n47169 = n65772 & n47168 ;
  assign n80661 = ~n46764 ;
  assign n46766 = n46533 & n80661 ;
  assign n47170 = n46508 | n46533 ;
  assign n80662 = ~n47170 ;
  assign n47171 = n46763 & n80662 ;
  assign n47172 = n46766 | n47171 ;
  assign n47173 = n80548 & n47172 ;
  assign n47174 = n46501 & n80544 ;
  assign n47175 = n46865 & n47174 ;
  assign n47176 = n47173 | n47175 ;
  assign n47177 = n65746 & n47176 ;
  assign n80663 = ~n47175 ;
  assign n47215 = x68 & n80663 ;
  assign n80664 = ~n47173 ;
  assign n47216 = n80664 & n47215 ;
  assign n47217 = n47177 | n47216 ;
  assign n80665 = ~n46526 ;
  assign n46762 = n80665 & n46761 ;
  assign n47178 = n46524 | n46761 ;
  assign n80666 = ~n47178 ;
  assign n47179 = n46525 & n80666 ;
  assign n47180 = n46762 | n47179 ;
  assign n47181 = n80548 & n47180 ;
  assign n47182 = n46507 & n80544 ;
  assign n47183 = n46865 & n47182 ;
  assign n47184 = n47181 | n47183 ;
  assign n47185 = n65721 & n47184 ;
  assign n47186 = n14255 & n46522 ;
  assign n47187 = n80546 & n47186 ;
  assign n80667 = ~n47187 ;
  assign n47188 = n46525 & n80667 ;
  assign n47189 = n80548 & n47188 ;
  assign n47190 = n46516 & n80544 ;
  assign n47191 = n46865 & n47190 ;
  assign n47192 = n47189 | n47191 ;
  assign n47193 = n65686 & n47192 ;
  assign n80668 = ~n47191 ;
  assign n47205 = x66 & n80668 ;
  assign n80669 = ~n47189 ;
  assign n47206 = n80669 & n47205 ;
  assign n47207 = n47193 | n47206 ;
  assign n46756 = n14255 & n80548 ;
  assign n46755 = x64 & n80548 ;
  assign n80670 = ~n46755 ;
  assign n47194 = x22 & n80670 ;
  assign n47195 = n46756 | n47194 ;
  assign n47196 = x65 & n47195 ;
  assign n47197 = n80544 & n46865 ;
  assign n80671 = ~n47197 ;
  assign n47198 = n14255 & n80671 ;
  assign n47199 = x65 | n47198 ;
  assign n47200 = n47194 | n47199 ;
  assign n80672 = ~n47196 ;
  assign n47201 = n80672 & n47200 ;
  assign n47203 = n14940 | n47201 ;
  assign n47204 = n65670 & n47195 ;
  assign n80673 = ~n47204 ;
  assign n47208 = n47203 & n80673 ;
  assign n47209 = n47207 | n47208 ;
  assign n80674 = ~n47193 ;
  assign n47210 = n80674 & n47209 ;
  assign n80675 = ~n47183 ;
  assign n47211 = x67 & n80675 ;
  assign n80676 = ~n47181 ;
  assign n47212 = n80676 & n47211 ;
  assign n47213 = n47185 | n47212 ;
  assign n47214 = n47210 | n47213 ;
  assign n80677 = ~n47185 ;
  assign n47218 = n80677 & n47214 ;
  assign n47219 = n47217 | n47218 ;
  assign n80678 = ~n47177 ;
  assign n47220 = n80678 & n47219 ;
  assign n80679 = ~n47167 ;
  assign n47221 = x69 & n80679 ;
  assign n80680 = ~n47165 ;
  assign n47222 = n80680 & n47221 ;
  assign n47223 = n47169 | n47222 ;
  assign n47225 = n47220 | n47223 ;
  assign n80681 = ~n47169 ;
  assign n47230 = n80681 & n47225 ;
  assign n47231 = n47228 | n47230 ;
  assign n80682 = ~n47160 ;
  assign n47232 = n80682 & n47231 ;
  assign n80683 = ~n47150 ;
  assign n47233 = x71 & n80683 ;
  assign n80684 = ~n47148 ;
  assign n47234 = n80684 & n47233 ;
  assign n47235 = n47152 | n47234 ;
  assign n47237 = n47232 | n47235 ;
  assign n80685 = ~n47152 ;
  assign n47242 = n80685 & n47237 ;
  assign n47243 = n47240 | n47242 ;
  assign n80686 = ~n47144 ;
  assign n47244 = n80686 & n47243 ;
  assign n80687 = ~n47134 ;
  assign n47245 = x73 & n80687 ;
  assign n80688 = ~n47132 ;
  assign n47246 = n80688 & n47245 ;
  assign n47247 = n47136 | n47246 ;
  assign n47249 = n47244 | n47247 ;
  assign n80689 = ~n47136 ;
  assign n47254 = n80689 & n47249 ;
  assign n47255 = n47252 | n47254 ;
  assign n80690 = ~n47128 ;
  assign n47256 = n80690 & n47255 ;
  assign n80691 = ~n47118 ;
  assign n47257 = x75 & n80691 ;
  assign n80692 = ~n47116 ;
  assign n47258 = n80692 & n47257 ;
  assign n47259 = n47120 | n47258 ;
  assign n47261 = n47256 | n47259 ;
  assign n80693 = ~n47120 ;
  assign n47266 = n80693 & n47261 ;
  assign n47267 = n47264 | n47266 ;
  assign n80694 = ~n47112 ;
  assign n47268 = n80694 & n47267 ;
  assign n80695 = ~n47102 ;
  assign n47269 = x77 & n80695 ;
  assign n80696 = ~n47100 ;
  assign n47270 = n80696 & n47269 ;
  assign n47271 = n47104 | n47270 ;
  assign n47273 = n47268 | n47271 ;
  assign n80697 = ~n47104 ;
  assign n47278 = n80697 & n47273 ;
  assign n47279 = n47276 | n47278 ;
  assign n80698 = ~n47096 ;
  assign n47280 = n80698 & n47279 ;
  assign n80699 = ~n47086 ;
  assign n47281 = x79 & n80699 ;
  assign n80700 = ~n47084 ;
  assign n47282 = n80700 & n47281 ;
  assign n47283 = n47088 | n47282 ;
  assign n47285 = n47280 | n47283 ;
  assign n80701 = ~n47088 ;
  assign n47290 = n80701 & n47285 ;
  assign n47291 = n47288 | n47290 ;
  assign n80702 = ~n47080 ;
  assign n47292 = n80702 & n47291 ;
  assign n80703 = ~n47070 ;
  assign n47293 = x81 & n80703 ;
  assign n80704 = ~n47068 ;
  assign n47294 = n80704 & n47293 ;
  assign n47295 = n47072 | n47294 ;
  assign n47297 = n47292 | n47295 ;
  assign n80705 = ~n47072 ;
  assign n47302 = n80705 & n47297 ;
  assign n47303 = n47300 | n47302 ;
  assign n80706 = ~n47064 ;
  assign n47304 = n80706 & n47303 ;
  assign n80707 = ~n47054 ;
  assign n47305 = x83 & n80707 ;
  assign n80708 = ~n47052 ;
  assign n47306 = n80708 & n47305 ;
  assign n47307 = n47056 | n47306 ;
  assign n47309 = n47304 | n47307 ;
  assign n80709 = ~n47056 ;
  assign n47314 = n80709 & n47309 ;
  assign n47315 = n47312 | n47314 ;
  assign n80710 = ~n47048 ;
  assign n47316 = n80710 & n47315 ;
  assign n80711 = ~n47038 ;
  assign n47317 = x85 & n80711 ;
  assign n80712 = ~n47036 ;
  assign n47318 = n80712 & n47317 ;
  assign n47319 = n47040 | n47318 ;
  assign n47321 = n47316 | n47319 ;
  assign n80713 = ~n47040 ;
  assign n47326 = n80713 & n47321 ;
  assign n47327 = n47324 | n47326 ;
  assign n80714 = ~n47032 ;
  assign n47328 = n80714 & n47327 ;
  assign n80715 = ~n47022 ;
  assign n47329 = x87 & n80715 ;
  assign n80716 = ~n47020 ;
  assign n47330 = n80716 & n47329 ;
  assign n47331 = n47024 | n47330 ;
  assign n47333 = n47328 | n47331 ;
  assign n80717 = ~n47024 ;
  assign n47338 = n80717 & n47333 ;
  assign n47339 = n47336 | n47338 ;
  assign n80718 = ~n47016 ;
  assign n47340 = n80718 & n47339 ;
  assign n80719 = ~n47006 ;
  assign n47341 = x89 & n80719 ;
  assign n80720 = ~n47004 ;
  assign n47342 = n80720 & n47341 ;
  assign n47343 = n47008 | n47342 ;
  assign n47345 = n47340 | n47343 ;
  assign n80721 = ~n47008 ;
  assign n47350 = n80721 & n47345 ;
  assign n47351 = n47348 | n47350 ;
  assign n80722 = ~n47000 ;
  assign n47352 = n80722 & n47351 ;
  assign n80723 = ~n46990 ;
  assign n47353 = x91 & n80723 ;
  assign n80724 = ~n46988 ;
  assign n47354 = n80724 & n47353 ;
  assign n47355 = n46992 | n47354 ;
  assign n47357 = n47352 | n47355 ;
  assign n80725 = ~n46992 ;
  assign n47362 = n80725 & n47357 ;
  assign n47363 = n47360 | n47362 ;
  assign n80726 = ~n46984 ;
  assign n47364 = n80726 & n47363 ;
  assign n80727 = ~n46974 ;
  assign n47365 = x93 & n80727 ;
  assign n80728 = ~n46972 ;
  assign n47366 = n80728 & n47365 ;
  assign n47367 = n46976 | n47366 ;
  assign n47369 = n47364 | n47367 ;
  assign n80729 = ~n46976 ;
  assign n47374 = n80729 & n47369 ;
  assign n47375 = n47372 | n47374 ;
  assign n80730 = ~n46968 ;
  assign n47376 = n80730 & n47375 ;
  assign n80731 = ~n46958 ;
  assign n47377 = x95 & n80731 ;
  assign n80732 = ~n46956 ;
  assign n47378 = n80732 & n47377 ;
  assign n47379 = n46960 | n47378 ;
  assign n47381 = n47376 | n47379 ;
  assign n80733 = ~n46960 ;
  assign n47386 = n80733 & n47381 ;
  assign n47387 = n47384 | n47386 ;
  assign n80734 = ~n46952 ;
  assign n47388 = n80734 & n47387 ;
  assign n80735 = ~n46942 ;
  assign n47389 = x97 & n80735 ;
  assign n80736 = ~n46940 ;
  assign n47390 = n80736 & n47389 ;
  assign n47391 = n46944 | n47390 ;
  assign n47393 = n47388 | n47391 ;
  assign n80737 = ~n46944 ;
  assign n47398 = n80737 & n47393 ;
  assign n47399 = n47396 | n47398 ;
  assign n80738 = ~n46936 ;
  assign n47400 = n80738 & n47399 ;
  assign n80739 = ~n46926 ;
  assign n47401 = x99 & n80739 ;
  assign n80740 = ~n46924 ;
  assign n47402 = n80740 & n47401 ;
  assign n47403 = n46928 | n47402 ;
  assign n47405 = n47400 | n47403 ;
  assign n80741 = ~n46928 ;
  assign n47410 = n80741 & n47405 ;
  assign n47411 = n47408 | n47410 ;
  assign n80742 = ~n46920 ;
  assign n47412 = n80742 & n47411 ;
  assign n80743 = ~n46910 ;
  assign n47413 = x101 & n80743 ;
  assign n80744 = ~n46908 ;
  assign n47414 = n80744 & n47413 ;
  assign n47415 = n46912 | n47414 ;
  assign n47417 = n47412 | n47415 ;
  assign n80745 = ~n46912 ;
  assign n47422 = n80745 & n47417 ;
  assign n47423 = n47420 | n47422 ;
  assign n80746 = ~n46904 ;
  assign n47424 = n80746 & n47423 ;
  assign n80747 = ~n46894 ;
  assign n47425 = x103 & n80747 ;
  assign n80748 = ~n46892 ;
  assign n47426 = n80748 & n47425 ;
  assign n47427 = n46896 | n47426 ;
  assign n47429 = n47424 | n47427 ;
  assign n80749 = ~n46896 ;
  assign n47434 = n80749 & n47429 ;
  assign n47435 = n47432 | n47434 ;
  assign n80750 = ~n46888 ;
  assign n47436 = n80750 & n47435 ;
  assign n80751 = ~n46867 ;
  assign n47437 = x105 & n80751 ;
  assign n80752 = ~n46861 ;
  assign n47438 = n80752 & n47437 ;
  assign n47439 = n46880 | n47438 ;
  assign n47441 = n47436 | n47439 ;
  assign n80753 = ~n46880 ;
  assign n47445 = n80753 & n47441 ;
  assign n47446 = n47444 | n47445 ;
  assign n80754 = ~n46879 ;
  assign n47447 = n80754 & n47446 ;
  assign n47448 = n15167 | n47447 ;
  assign n80755 = ~n46878 ;
  assign n47450 = n80755 & n47448 ;
  assign n80756 = ~n47445 ;
  assign n48106 = n47444 & n80756 ;
  assign n47452 = x64 & n80671 ;
  assign n80757 = ~n47452 ;
  assign n47453 = x22 & n80757 ;
  assign n47454 = n46756 | n47453 ;
  assign n47455 = x65 & n47454 ;
  assign n80758 = ~n47455 ;
  assign n47456 = n47200 & n80758 ;
  assign n47457 = n14940 | n47456 ;
  assign n47458 = n80673 & n47457 ;
  assign n47460 = n47207 | n47458 ;
  assign n47461 = n80674 & n47460 ;
  assign n47462 = n47213 | n47461 ;
  assign n47463 = n80677 & n47462 ;
  assign n47464 = n47217 | n47463 ;
  assign n47465 = n80678 & n47464 ;
  assign n47466 = n47223 | n47465 ;
  assign n47467 = n80681 & n47466 ;
  assign n47468 = n47228 | n47467 ;
  assign n47469 = n80682 & n47468 ;
  assign n47470 = n47235 | n47469 ;
  assign n47471 = n80685 & n47470 ;
  assign n47472 = n47240 | n47471 ;
  assign n47473 = n80686 & n47472 ;
  assign n47474 = n47247 | n47473 ;
  assign n47475 = n80689 & n47474 ;
  assign n47476 = n47252 | n47475 ;
  assign n47477 = n80690 & n47476 ;
  assign n47478 = n47259 | n47477 ;
  assign n47479 = n80693 & n47478 ;
  assign n47480 = n47264 | n47479 ;
  assign n47481 = n80694 & n47480 ;
  assign n47482 = n47271 | n47481 ;
  assign n47483 = n80697 & n47482 ;
  assign n47484 = n47276 | n47483 ;
  assign n47485 = n80698 & n47484 ;
  assign n47486 = n47283 | n47485 ;
  assign n47487 = n80701 & n47486 ;
  assign n47488 = n47288 | n47487 ;
  assign n47489 = n80702 & n47488 ;
  assign n47490 = n47295 | n47489 ;
  assign n47491 = n80705 & n47490 ;
  assign n47492 = n47300 | n47491 ;
  assign n47493 = n80706 & n47492 ;
  assign n47494 = n47307 | n47493 ;
  assign n47495 = n80709 & n47494 ;
  assign n47496 = n47312 | n47495 ;
  assign n47497 = n80710 & n47496 ;
  assign n47498 = n47319 | n47497 ;
  assign n47499 = n80713 & n47498 ;
  assign n47500 = n47324 | n47499 ;
  assign n47501 = n80714 & n47500 ;
  assign n47502 = n47331 | n47501 ;
  assign n47503 = n80717 & n47502 ;
  assign n47504 = n47336 | n47503 ;
  assign n47505 = n80718 & n47504 ;
  assign n47506 = n47343 | n47505 ;
  assign n47507 = n80721 & n47506 ;
  assign n47508 = n47348 | n47507 ;
  assign n47509 = n80722 & n47508 ;
  assign n47510 = n47355 | n47509 ;
  assign n47511 = n80725 & n47510 ;
  assign n47512 = n47360 | n47511 ;
  assign n47513 = n80726 & n47512 ;
  assign n47514 = n47367 | n47513 ;
  assign n47515 = n80729 & n47514 ;
  assign n47516 = n47372 | n47515 ;
  assign n47517 = n80730 & n47516 ;
  assign n47518 = n47379 | n47517 ;
  assign n47519 = n80733 & n47518 ;
  assign n47520 = n47384 | n47519 ;
  assign n47521 = n80734 & n47520 ;
  assign n47522 = n47391 | n47521 ;
  assign n47523 = n80737 & n47522 ;
  assign n47524 = n47396 | n47523 ;
  assign n47525 = n80738 & n47524 ;
  assign n47526 = n47403 | n47525 ;
  assign n47527 = n80741 & n47526 ;
  assign n47528 = n47408 | n47527 ;
  assign n47529 = n80742 & n47528 ;
  assign n47530 = n47415 | n47529 ;
  assign n47531 = n80745 & n47530 ;
  assign n47532 = n47420 | n47531 ;
  assign n47533 = n80746 & n47532 ;
  assign n47534 = n47427 | n47533 ;
  assign n47535 = n80749 & n47534 ;
  assign n47536 = n47432 | n47535 ;
  assign n47538 = n80750 & n47536 ;
  assign n47866 = n47439 | n47538 ;
  assign n48107 = n46880 | n47444 ;
  assign n80759 = ~n48107 ;
  assign n48108 = n47866 & n80759 ;
  assign n48109 = n48106 | n48108 ;
  assign n48110 = n47448 | n48109 ;
  assign n80760 = ~n47450 ;
  assign n48111 = n80760 & n48110 ;
  assign n48119 = n70486 & n48111 ;
  assign n47451 = n46868 & n47448 ;
  assign n47440 = n46888 | n47439 ;
  assign n80761 = ~n47440 ;
  assign n47537 = n80761 & n47536 ;
  assign n80762 = ~n47538 ;
  assign n47539 = n47439 & n80762 ;
  assign n47540 = n47537 | n47539 ;
  assign n47541 = n70486 & n47540 ;
  assign n80763 = ~n47447 ;
  assign n47542 = n80763 & n47541 ;
  assign n47543 = n47451 | n47542 ;
  assign n47544 = n70276 & n47543 ;
  assign n47545 = n46887 & n47448 ;
  assign n47433 = n46896 | n47432 ;
  assign n80764 = ~n47433 ;
  assign n47546 = n47429 & n80764 ;
  assign n80765 = ~n47434 ;
  assign n47547 = n47432 & n80765 ;
  assign n47548 = n47546 | n47547 ;
  assign n47549 = n70486 & n47548 ;
  assign n47550 = n80763 & n47549 ;
  assign n47551 = n47545 | n47550 ;
  assign n47552 = n70176 & n47551 ;
  assign n47553 = n46895 & n47448 ;
  assign n47428 = n46904 | n47427 ;
  assign n80766 = ~n47428 ;
  assign n47554 = n80766 & n47532 ;
  assign n80767 = ~n47533 ;
  assign n47555 = n47427 & n80767 ;
  assign n47556 = n47554 | n47555 ;
  assign n47557 = n70486 & n47556 ;
  assign n47558 = n80763 & n47557 ;
  assign n47559 = n47553 | n47558 ;
  assign n47560 = n69857 & n47559 ;
  assign n47561 = n46903 & n47448 ;
  assign n47421 = n46912 | n47420 ;
  assign n80768 = ~n47421 ;
  assign n47562 = n47417 & n80768 ;
  assign n80769 = ~n47422 ;
  assign n47563 = n47420 & n80769 ;
  assign n47564 = n47562 | n47563 ;
  assign n47565 = n70486 & n47564 ;
  assign n47566 = n80763 & n47565 ;
  assign n47567 = n47561 | n47566 ;
  assign n47568 = n69656 & n47567 ;
  assign n47569 = n46911 & n47448 ;
  assign n47416 = n46920 | n47415 ;
  assign n80770 = ~n47416 ;
  assign n47570 = n80770 & n47528 ;
  assign n80771 = ~n47529 ;
  assign n47571 = n47415 & n80771 ;
  assign n47572 = n47570 | n47571 ;
  assign n47573 = n70486 & n47572 ;
  assign n47574 = n80763 & n47573 ;
  assign n47575 = n47569 | n47574 ;
  assign n47576 = n69528 & n47575 ;
  assign n47577 = n46919 & n47448 ;
  assign n47409 = n46928 | n47408 ;
  assign n80772 = ~n47409 ;
  assign n47578 = n47405 & n80772 ;
  assign n80773 = ~n47410 ;
  assign n47579 = n47408 & n80773 ;
  assign n47580 = n47578 | n47579 ;
  assign n47581 = n70486 & n47580 ;
  assign n47582 = n80763 & n47581 ;
  assign n47583 = n47577 | n47582 ;
  assign n47584 = n69261 & n47583 ;
  assign n47585 = n46927 & n47448 ;
  assign n47404 = n46936 | n47403 ;
  assign n80774 = ~n47404 ;
  assign n47586 = n80774 & n47524 ;
  assign n80775 = ~n47525 ;
  assign n47587 = n47403 & n80775 ;
  assign n47588 = n47586 | n47587 ;
  assign n47589 = n70486 & n47588 ;
  assign n47590 = n80763 & n47589 ;
  assign n47591 = n47585 | n47590 ;
  assign n47592 = n69075 & n47591 ;
  assign n47593 = n46935 & n47448 ;
  assign n47397 = n46944 | n47396 ;
  assign n80776 = ~n47397 ;
  assign n47594 = n47393 & n80776 ;
  assign n80777 = ~n47398 ;
  assign n47595 = n47396 & n80777 ;
  assign n47596 = n47594 | n47595 ;
  assign n47597 = n70486 & n47596 ;
  assign n47598 = n80763 & n47597 ;
  assign n47599 = n47593 | n47598 ;
  assign n47600 = n68993 & n47599 ;
  assign n47601 = n46943 & n47448 ;
  assign n47392 = n46952 | n47391 ;
  assign n80778 = ~n47392 ;
  assign n47602 = n80778 & n47520 ;
  assign n80779 = ~n47521 ;
  assign n47603 = n47391 & n80779 ;
  assign n47604 = n47602 | n47603 ;
  assign n47605 = n70486 & n47604 ;
  assign n47606 = n80763 & n47605 ;
  assign n47607 = n47601 | n47606 ;
  assign n47608 = n68716 & n47607 ;
  assign n47609 = n46951 & n47448 ;
  assign n47385 = n46960 | n47384 ;
  assign n80780 = ~n47385 ;
  assign n47610 = n47381 & n80780 ;
  assign n80781 = ~n47386 ;
  assign n47611 = n47384 & n80781 ;
  assign n47612 = n47610 | n47611 ;
  assign n47613 = n70486 & n47612 ;
  assign n47614 = n80763 & n47613 ;
  assign n47615 = n47609 | n47614 ;
  assign n47616 = n68545 & n47615 ;
  assign n47617 = n46959 & n47448 ;
  assign n47380 = n46968 | n47379 ;
  assign n80782 = ~n47380 ;
  assign n47618 = n80782 & n47516 ;
  assign n80783 = ~n47517 ;
  assign n47619 = n47379 & n80783 ;
  assign n47620 = n47618 | n47619 ;
  assign n47621 = n70486 & n47620 ;
  assign n47622 = n80763 & n47621 ;
  assign n47623 = n47617 | n47622 ;
  assign n47624 = n68438 & n47623 ;
  assign n47625 = n46967 & n47448 ;
  assign n47373 = n46976 | n47372 ;
  assign n80784 = ~n47373 ;
  assign n47626 = n47369 & n80784 ;
  assign n80785 = ~n47374 ;
  assign n47627 = n47372 & n80785 ;
  assign n47628 = n47626 | n47627 ;
  assign n47629 = n70486 & n47628 ;
  assign n47630 = n80763 & n47629 ;
  assign n47631 = n47625 | n47630 ;
  assign n47632 = n68214 & n47631 ;
  assign n47633 = n46975 & n47448 ;
  assign n47368 = n46984 | n47367 ;
  assign n80786 = ~n47368 ;
  assign n47634 = n80786 & n47512 ;
  assign n80787 = ~n47513 ;
  assign n47635 = n47367 & n80787 ;
  assign n47636 = n47634 | n47635 ;
  assign n47637 = n70486 & n47636 ;
  assign n47638 = n80763 & n47637 ;
  assign n47639 = n47633 | n47638 ;
  assign n47640 = n68058 & n47639 ;
  assign n47641 = n46983 & n47448 ;
  assign n47361 = n46992 | n47360 ;
  assign n80788 = ~n47361 ;
  assign n47642 = n47357 & n80788 ;
  assign n80789 = ~n47362 ;
  assign n47643 = n47360 & n80789 ;
  assign n47644 = n47642 | n47643 ;
  assign n47645 = n70486 & n47644 ;
  assign n47646 = n80763 & n47645 ;
  assign n47647 = n47641 | n47646 ;
  assign n47648 = n67986 & n47647 ;
  assign n47649 = n46991 & n47448 ;
  assign n47356 = n47000 | n47355 ;
  assign n80790 = ~n47356 ;
  assign n47650 = n80790 & n47508 ;
  assign n80791 = ~n47509 ;
  assign n47651 = n47355 & n80791 ;
  assign n47652 = n47650 | n47651 ;
  assign n47653 = n70486 & n47652 ;
  assign n47654 = n80763 & n47653 ;
  assign n47655 = n47649 | n47654 ;
  assign n47656 = n67763 & n47655 ;
  assign n47657 = n46999 & n47448 ;
  assign n47349 = n47008 | n47348 ;
  assign n80792 = ~n47349 ;
  assign n47658 = n47345 & n80792 ;
  assign n80793 = ~n47350 ;
  assign n47659 = n47348 & n80793 ;
  assign n47660 = n47658 | n47659 ;
  assign n47661 = n70486 & n47660 ;
  assign n47662 = n80763 & n47661 ;
  assign n47663 = n47657 | n47662 ;
  assign n47664 = n67622 & n47663 ;
  assign n47665 = n47007 & n47448 ;
  assign n47344 = n47016 | n47343 ;
  assign n80794 = ~n47344 ;
  assign n47666 = n80794 & n47504 ;
  assign n80795 = ~n47505 ;
  assign n47667 = n47343 & n80795 ;
  assign n47668 = n47666 | n47667 ;
  assign n47669 = n70486 & n47668 ;
  assign n47670 = n80763 & n47669 ;
  assign n47671 = n47665 | n47670 ;
  assign n47672 = n67531 & n47671 ;
  assign n47673 = n47015 & n47448 ;
  assign n47337 = n47024 | n47336 ;
  assign n80796 = ~n47337 ;
  assign n47674 = n47333 & n80796 ;
  assign n80797 = ~n47338 ;
  assign n47675 = n47336 & n80797 ;
  assign n47676 = n47674 | n47675 ;
  assign n47677 = n70486 & n47676 ;
  assign n47678 = n80763 & n47677 ;
  assign n47679 = n47673 | n47678 ;
  assign n47680 = n67348 & n47679 ;
  assign n47681 = n47023 & n47448 ;
  assign n47332 = n47032 | n47331 ;
  assign n80798 = ~n47332 ;
  assign n47682 = n80798 & n47500 ;
  assign n80799 = ~n47501 ;
  assign n47683 = n47331 & n80799 ;
  assign n47684 = n47682 | n47683 ;
  assign n47685 = n70486 & n47684 ;
  assign n47686 = n80763 & n47685 ;
  assign n47687 = n47681 | n47686 ;
  assign n47688 = n67222 & n47687 ;
  assign n47689 = n47031 & n47448 ;
  assign n47325 = n47040 | n47324 ;
  assign n80800 = ~n47325 ;
  assign n47690 = n47321 & n80800 ;
  assign n80801 = ~n47326 ;
  assign n47691 = n47324 & n80801 ;
  assign n47692 = n47690 | n47691 ;
  assign n47693 = n70486 & n47692 ;
  assign n47694 = n80763 & n47693 ;
  assign n47695 = n47689 | n47694 ;
  assign n47696 = n67164 & n47695 ;
  assign n47697 = n47039 & n47448 ;
  assign n47320 = n47048 | n47319 ;
  assign n80802 = ~n47320 ;
  assign n47698 = n80802 & n47496 ;
  assign n80803 = ~n47497 ;
  assign n47699 = n47319 & n80803 ;
  assign n47700 = n47698 | n47699 ;
  assign n47701 = n70486 & n47700 ;
  assign n47702 = n80763 & n47701 ;
  assign n47703 = n47697 | n47702 ;
  assign n47704 = n66979 & n47703 ;
  assign n47705 = n47047 & n47448 ;
  assign n47313 = n47056 | n47312 ;
  assign n80804 = ~n47313 ;
  assign n47706 = n47309 & n80804 ;
  assign n80805 = ~n47314 ;
  assign n47707 = n47312 & n80805 ;
  assign n47708 = n47706 | n47707 ;
  assign n47709 = n70486 & n47708 ;
  assign n47710 = n80763 & n47709 ;
  assign n47711 = n47705 | n47710 ;
  assign n47712 = n66868 & n47711 ;
  assign n47713 = n47055 & n47448 ;
  assign n47308 = n47064 | n47307 ;
  assign n80806 = ~n47308 ;
  assign n47714 = n80806 & n47492 ;
  assign n80807 = ~n47493 ;
  assign n47715 = n47307 & n80807 ;
  assign n47716 = n47714 | n47715 ;
  assign n47717 = n70486 & n47716 ;
  assign n47718 = n80763 & n47717 ;
  assign n47719 = n47713 | n47718 ;
  assign n47720 = n66797 & n47719 ;
  assign n47721 = n47063 & n47448 ;
  assign n47301 = n47072 | n47300 ;
  assign n80808 = ~n47301 ;
  assign n47722 = n47297 & n80808 ;
  assign n80809 = ~n47302 ;
  assign n47723 = n47300 & n80809 ;
  assign n47724 = n47722 | n47723 ;
  assign n47725 = n70486 & n47724 ;
  assign n47726 = n80763 & n47725 ;
  assign n47727 = n47721 | n47726 ;
  assign n47728 = n66654 & n47727 ;
  assign n47729 = n47071 & n47448 ;
  assign n47296 = n47080 | n47295 ;
  assign n80810 = ~n47296 ;
  assign n47730 = n80810 & n47488 ;
  assign n80811 = ~n47489 ;
  assign n47731 = n47295 & n80811 ;
  assign n47732 = n47730 | n47731 ;
  assign n47733 = n70486 & n47732 ;
  assign n47734 = n80763 & n47733 ;
  assign n47735 = n47729 | n47734 ;
  assign n47736 = n66560 & n47735 ;
  assign n47737 = n47079 & n47448 ;
  assign n47289 = n47088 | n47288 ;
  assign n80812 = ~n47289 ;
  assign n47738 = n47285 & n80812 ;
  assign n80813 = ~n47290 ;
  assign n47739 = n47288 & n80813 ;
  assign n47740 = n47738 | n47739 ;
  assign n47741 = n70486 & n47740 ;
  assign n47742 = n80763 & n47741 ;
  assign n47743 = n47737 | n47742 ;
  assign n47744 = n66505 & n47743 ;
  assign n47745 = n47087 & n47448 ;
  assign n47284 = n47096 | n47283 ;
  assign n80814 = ~n47284 ;
  assign n47746 = n80814 & n47484 ;
  assign n80815 = ~n47485 ;
  assign n47747 = n47283 & n80815 ;
  assign n47748 = n47746 | n47747 ;
  assign n47749 = n70486 & n47748 ;
  assign n47750 = n80763 & n47749 ;
  assign n47751 = n47745 | n47750 ;
  assign n47752 = n66379 & n47751 ;
  assign n47753 = n47095 & n47448 ;
  assign n47277 = n47104 | n47276 ;
  assign n80816 = ~n47277 ;
  assign n47754 = n47273 & n80816 ;
  assign n80817 = ~n47278 ;
  assign n47755 = n47276 & n80817 ;
  assign n47756 = n47754 | n47755 ;
  assign n47757 = n70486 & n47756 ;
  assign n47758 = n80763 & n47757 ;
  assign n47759 = n47753 | n47758 ;
  assign n47760 = n66299 & n47759 ;
  assign n47761 = n47103 & n47448 ;
  assign n47272 = n47112 | n47271 ;
  assign n80818 = ~n47272 ;
  assign n47762 = n80818 & n47480 ;
  assign n80819 = ~n47481 ;
  assign n47763 = n47271 & n80819 ;
  assign n47764 = n47762 | n47763 ;
  assign n47765 = n70486 & n47764 ;
  assign n47766 = n80763 & n47765 ;
  assign n47767 = n47761 | n47766 ;
  assign n47768 = n66244 & n47767 ;
  assign n47769 = n47111 & n47448 ;
  assign n47265 = n47120 | n47264 ;
  assign n80820 = ~n47265 ;
  assign n47770 = n47261 & n80820 ;
  assign n80821 = ~n47266 ;
  assign n47771 = n47264 & n80821 ;
  assign n47772 = n47770 | n47771 ;
  assign n47773 = n70486 & n47772 ;
  assign n47774 = n80763 & n47773 ;
  assign n47775 = n47769 | n47774 ;
  assign n47776 = n66145 & n47775 ;
  assign n47777 = n47119 & n47448 ;
  assign n47260 = n47128 | n47259 ;
  assign n80822 = ~n47260 ;
  assign n47778 = n80822 & n47476 ;
  assign n80823 = ~n47477 ;
  assign n47779 = n47259 & n80823 ;
  assign n47780 = n47778 | n47779 ;
  assign n47781 = n70486 & n47780 ;
  assign n47782 = n80763 & n47781 ;
  assign n47783 = n47777 | n47782 ;
  assign n47784 = n66081 & n47783 ;
  assign n47785 = n47127 & n47448 ;
  assign n47253 = n47136 | n47252 ;
  assign n80824 = ~n47253 ;
  assign n47786 = n47249 & n80824 ;
  assign n80825 = ~n47254 ;
  assign n47787 = n47252 & n80825 ;
  assign n47788 = n47786 | n47787 ;
  assign n47789 = n70486 & n47788 ;
  assign n47790 = n80763 & n47789 ;
  assign n47791 = n47785 | n47790 ;
  assign n47792 = n66043 & n47791 ;
  assign n47793 = n47135 & n47448 ;
  assign n47248 = n47144 | n47247 ;
  assign n80826 = ~n47248 ;
  assign n47794 = n80826 & n47472 ;
  assign n80827 = ~n47473 ;
  assign n47795 = n47247 & n80827 ;
  assign n47796 = n47794 | n47795 ;
  assign n47797 = n70486 & n47796 ;
  assign n47798 = n80763 & n47797 ;
  assign n47799 = n47793 | n47798 ;
  assign n47800 = n65960 & n47799 ;
  assign n47801 = n47143 & n47448 ;
  assign n47241 = n47152 | n47240 ;
  assign n80828 = ~n47241 ;
  assign n47802 = n47237 & n80828 ;
  assign n80829 = ~n47242 ;
  assign n47803 = n47240 & n80829 ;
  assign n47804 = n47802 | n47803 ;
  assign n47805 = n70486 & n47804 ;
  assign n47806 = n80763 & n47805 ;
  assign n47807 = n47801 | n47806 ;
  assign n47808 = n65909 & n47807 ;
  assign n47809 = n47151 & n47448 ;
  assign n47236 = n47160 | n47235 ;
  assign n80830 = ~n47236 ;
  assign n47810 = n80830 & n47468 ;
  assign n80831 = ~n47469 ;
  assign n47811 = n47235 & n80831 ;
  assign n47812 = n47810 | n47811 ;
  assign n47813 = n70486 & n47812 ;
  assign n47814 = n80763 & n47813 ;
  assign n47815 = n47809 | n47814 ;
  assign n47816 = n65877 & n47815 ;
  assign n47817 = n47159 & n47448 ;
  assign n47229 = n47169 | n47228 ;
  assign n80832 = ~n47229 ;
  assign n47818 = n47225 & n80832 ;
  assign n80833 = ~n47230 ;
  assign n47819 = n47228 & n80833 ;
  assign n47820 = n47818 | n47819 ;
  assign n47821 = n70486 & n47820 ;
  assign n47822 = n80763 & n47821 ;
  assign n47823 = n47817 | n47822 ;
  assign n47824 = n65820 & n47823 ;
  assign n47825 = n47168 & n47448 ;
  assign n47224 = n47177 | n47223 ;
  assign n80834 = ~n47224 ;
  assign n47826 = n80834 & n47464 ;
  assign n80835 = ~n47465 ;
  assign n47827 = n47223 & n80835 ;
  assign n47828 = n47826 | n47827 ;
  assign n47829 = n70486 & n47828 ;
  assign n47830 = n80763 & n47829 ;
  assign n47831 = n47825 | n47830 ;
  assign n47832 = n65791 & n47831 ;
  assign n47833 = n47176 & n47448 ;
  assign n47834 = n47185 | n47217 ;
  assign n80836 = ~n47834 ;
  assign n47835 = n47214 & n80836 ;
  assign n80837 = ~n47218 ;
  assign n47836 = n47217 & n80837 ;
  assign n47837 = n47835 | n47836 ;
  assign n47838 = n70486 & n47837 ;
  assign n47839 = n80763 & n47838 ;
  assign n47840 = n47833 | n47839 ;
  assign n47841 = n65772 & n47840 ;
  assign n47842 = n47184 & n47448 ;
  assign n47843 = n47193 | n47213 ;
  assign n80838 = ~n47843 ;
  assign n47844 = n47209 & n80838 ;
  assign n80839 = ~n47461 ;
  assign n47845 = n47213 & n80839 ;
  assign n47846 = n47844 | n47845 ;
  assign n47847 = n70486 & n47846 ;
  assign n47848 = n80763 & n47847 ;
  assign n47849 = n47842 | n47848 ;
  assign n47850 = n65746 & n47849 ;
  assign n47851 = n47192 & n47448 ;
  assign n47459 = n47204 | n47207 ;
  assign n80840 = ~n47459 ;
  assign n47852 = n47457 & n80840 ;
  assign n80841 = ~n47208 ;
  assign n47853 = n47207 & n80841 ;
  assign n47854 = n47852 | n47853 ;
  assign n47855 = n70486 & n47854 ;
  assign n47856 = n80763 & n47855 ;
  assign n47857 = n47851 | n47856 ;
  assign n47858 = n65721 & n47857 ;
  assign n47449 = n47195 & n47448 ;
  assign n47202 = n14940 & n47200 ;
  assign n47859 = n47202 & n80758 ;
  assign n47860 = n15167 | n47859 ;
  assign n80842 = ~n47860 ;
  assign n47861 = n47457 & n80842 ;
  assign n47862 = n80763 & n47861 ;
  assign n47863 = n47449 | n47862 ;
  assign n47864 = n65686 & n47863 ;
  assign n47865 = n15616 & n80763 ;
  assign n47867 = n80753 & n47866 ;
  assign n47868 = n47444 | n47867 ;
  assign n47869 = n80754 & n47868 ;
  assign n80843 = ~n47869 ;
  assign n47870 = n15611 & n80843 ;
  assign n80844 = ~n47870 ;
  assign n47871 = x21 & n80844 ;
  assign n47872 = n47865 | n47871 ;
  assign n47880 = n65670 & n47872 ;
  assign n47873 = n15611 & n80763 ;
  assign n80845 = ~n47873 ;
  assign n47874 = x21 & n80845 ;
  assign n47875 = n47865 | n47874 ;
  assign n47876 = x65 & n47875 ;
  assign n47877 = x65 | n47865 ;
  assign n47878 = n47874 | n47877 ;
  assign n80846 = ~n47876 ;
  assign n47879 = n80846 & n47878 ;
  assign n47881 = n15623 | n47879 ;
  assign n80847 = ~n47880 ;
  assign n47882 = n80847 & n47881 ;
  assign n80848 = ~n47862 ;
  assign n47883 = x66 & n80848 ;
  assign n80849 = ~n47449 ;
  assign n47884 = n80849 & n47883 ;
  assign n47885 = n47882 | n47884 ;
  assign n80850 = ~n47864 ;
  assign n47886 = n80850 & n47885 ;
  assign n80851 = ~n47856 ;
  assign n47887 = x67 & n80851 ;
  assign n80852 = ~n47851 ;
  assign n47888 = n80852 & n47887 ;
  assign n47889 = n47858 | n47888 ;
  assign n47890 = n47886 | n47889 ;
  assign n80853 = ~n47858 ;
  assign n47891 = n80853 & n47890 ;
  assign n80854 = ~n47848 ;
  assign n47892 = x68 & n80854 ;
  assign n80855 = ~n47842 ;
  assign n47893 = n80855 & n47892 ;
  assign n47894 = n47850 | n47893 ;
  assign n47895 = n47891 | n47894 ;
  assign n80856 = ~n47850 ;
  assign n47896 = n80856 & n47895 ;
  assign n80857 = ~n47839 ;
  assign n47897 = x69 & n80857 ;
  assign n80858 = ~n47833 ;
  assign n47898 = n80858 & n47897 ;
  assign n47899 = n47841 | n47898 ;
  assign n47900 = n47896 | n47899 ;
  assign n80859 = ~n47841 ;
  assign n47901 = n80859 & n47900 ;
  assign n80860 = ~n47830 ;
  assign n47902 = x70 & n80860 ;
  assign n80861 = ~n47825 ;
  assign n47903 = n80861 & n47902 ;
  assign n47904 = n47832 | n47903 ;
  assign n47906 = n47901 | n47904 ;
  assign n80862 = ~n47832 ;
  assign n47907 = n80862 & n47906 ;
  assign n80863 = ~n47822 ;
  assign n47908 = x71 & n80863 ;
  assign n80864 = ~n47817 ;
  assign n47909 = n80864 & n47908 ;
  assign n47910 = n47824 | n47909 ;
  assign n47911 = n47907 | n47910 ;
  assign n80865 = ~n47824 ;
  assign n47912 = n80865 & n47911 ;
  assign n80866 = ~n47814 ;
  assign n47913 = x72 & n80866 ;
  assign n80867 = ~n47809 ;
  assign n47914 = n80867 & n47913 ;
  assign n47915 = n47816 | n47914 ;
  assign n47917 = n47912 | n47915 ;
  assign n80868 = ~n47816 ;
  assign n47918 = n80868 & n47917 ;
  assign n80869 = ~n47806 ;
  assign n47919 = x73 & n80869 ;
  assign n80870 = ~n47801 ;
  assign n47920 = n80870 & n47919 ;
  assign n47921 = n47808 | n47920 ;
  assign n47922 = n47918 | n47921 ;
  assign n80871 = ~n47808 ;
  assign n47923 = n80871 & n47922 ;
  assign n80872 = ~n47798 ;
  assign n47924 = x74 & n80872 ;
  assign n80873 = ~n47793 ;
  assign n47925 = n80873 & n47924 ;
  assign n47926 = n47800 | n47925 ;
  assign n47928 = n47923 | n47926 ;
  assign n80874 = ~n47800 ;
  assign n47929 = n80874 & n47928 ;
  assign n80875 = ~n47790 ;
  assign n47930 = x75 & n80875 ;
  assign n80876 = ~n47785 ;
  assign n47931 = n80876 & n47930 ;
  assign n47932 = n47792 | n47931 ;
  assign n47933 = n47929 | n47932 ;
  assign n80877 = ~n47792 ;
  assign n47934 = n80877 & n47933 ;
  assign n80878 = ~n47782 ;
  assign n47935 = x76 & n80878 ;
  assign n80879 = ~n47777 ;
  assign n47936 = n80879 & n47935 ;
  assign n47937 = n47784 | n47936 ;
  assign n47939 = n47934 | n47937 ;
  assign n80880 = ~n47784 ;
  assign n47940 = n80880 & n47939 ;
  assign n80881 = ~n47774 ;
  assign n47941 = x77 & n80881 ;
  assign n80882 = ~n47769 ;
  assign n47942 = n80882 & n47941 ;
  assign n47943 = n47776 | n47942 ;
  assign n47944 = n47940 | n47943 ;
  assign n80883 = ~n47776 ;
  assign n47945 = n80883 & n47944 ;
  assign n80884 = ~n47766 ;
  assign n47946 = x78 & n80884 ;
  assign n80885 = ~n47761 ;
  assign n47947 = n80885 & n47946 ;
  assign n47948 = n47768 | n47947 ;
  assign n47950 = n47945 | n47948 ;
  assign n80886 = ~n47768 ;
  assign n47951 = n80886 & n47950 ;
  assign n80887 = ~n47758 ;
  assign n47952 = x79 & n80887 ;
  assign n80888 = ~n47753 ;
  assign n47953 = n80888 & n47952 ;
  assign n47954 = n47760 | n47953 ;
  assign n47955 = n47951 | n47954 ;
  assign n80889 = ~n47760 ;
  assign n47956 = n80889 & n47955 ;
  assign n80890 = ~n47750 ;
  assign n47957 = x80 & n80890 ;
  assign n80891 = ~n47745 ;
  assign n47958 = n80891 & n47957 ;
  assign n47959 = n47752 | n47958 ;
  assign n47961 = n47956 | n47959 ;
  assign n80892 = ~n47752 ;
  assign n47962 = n80892 & n47961 ;
  assign n80893 = ~n47742 ;
  assign n47963 = x81 & n80893 ;
  assign n80894 = ~n47737 ;
  assign n47964 = n80894 & n47963 ;
  assign n47965 = n47744 | n47964 ;
  assign n47966 = n47962 | n47965 ;
  assign n80895 = ~n47744 ;
  assign n47967 = n80895 & n47966 ;
  assign n80896 = ~n47734 ;
  assign n47968 = x82 & n80896 ;
  assign n80897 = ~n47729 ;
  assign n47969 = n80897 & n47968 ;
  assign n47970 = n47736 | n47969 ;
  assign n47972 = n47967 | n47970 ;
  assign n80898 = ~n47736 ;
  assign n47973 = n80898 & n47972 ;
  assign n80899 = ~n47726 ;
  assign n47974 = x83 & n80899 ;
  assign n80900 = ~n47721 ;
  assign n47975 = n80900 & n47974 ;
  assign n47976 = n47728 | n47975 ;
  assign n47977 = n47973 | n47976 ;
  assign n80901 = ~n47728 ;
  assign n47978 = n80901 & n47977 ;
  assign n80902 = ~n47718 ;
  assign n47979 = x84 & n80902 ;
  assign n80903 = ~n47713 ;
  assign n47980 = n80903 & n47979 ;
  assign n47981 = n47720 | n47980 ;
  assign n47983 = n47978 | n47981 ;
  assign n80904 = ~n47720 ;
  assign n47984 = n80904 & n47983 ;
  assign n80905 = ~n47710 ;
  assign n47985 = x85 & n80905 ;
  assign n80906 = ~n47705 ;
  assign n47986 = n80906 & n47985 ;
  assign n47987 = n47712 | n47986 ;
  assign n47988 = n47984 | n47987 ;
  assign n80907 = ~n47712 ;
  assign n47989 = n80907 & n47988 ;
  assign n80908 = ~n47702 ;
  assign n47990 = x86 & n80908 ;
  assign n80909 = ~n47697 ;
  assign n47991 = n80909 & n47990 ;
  assign n47992 = n47704 | n47991 ;
  assign n47994 = n47989 | n47992 ;
  assign n80910 = ~n47704 ;
  assign n47995 = n80910 & n47994 ;
  assign n80911 = ~n47694 ;
  assign n47996 = x87 & n80911 ;
  assign n80912 = ~n47689 ;
  assign n47997 = n80912 & n47996 ;
  assign n47998 = n47696 | n47997 ;
  assign n47999 = n47995 | n47998 ;
  assign n80913 = ~n47696 ;
  assign n48000 = n80913 & n47999 ;
  assign n80914 = ~n47686 ;
  assign n48001 = x88 & n80914 ;
  assign n80915 = ~n47681 ;
  assign n48002 = n80915 & n48001 ;
  assign n48003 = n47688 | n48002 ;
  assign n48005 = n48000 | n48003 ;
  assign n80916 = ~n47688 ;
  assign n48006 = n80916 & n48005 ;
  assign n80917 = ~n47678 ;
  assign n48007 = x89 & n80917 ;
  assign n80918 = ~n47673 ;
  assign n48008 = n80918 & n48007 ;
  assign n48009 = n47680 | n48008 ;
  assign n48010 = n48006 | n48009 ;
  assign n80919 = ~n47680 ;
  assign n48011 = n80919 & n48010 ;
  assign n80920 = ~n47670 ;
  assign n48012 = x90 & n80920 ;
  assign n80921 = ~n47665 ;
  assign n48013 = n80921 & n48012 ;
  assign n48014 = n47672 | n48013 ;
  assign n48016 = n48011 | n48014 ;
  assign n80922 = ~n47672 ;
  assign n48017 = n80922 & n48016 ;
  assign n80923 = ~n47662 ;
  assign n48018 = x91 & n80923 ;
  assign n80924 = ~n47657 ;
  assign n48019 = n80924 & n48018 ;
  assign n48020 = n47664 | n48019 ;
  assign n48021 = n48017 | n48020 ;
  assign n80925 = ~n47664 ;
  assign n48022 = n80925 & n48021 ;
  assign n80926 = ~n47654 ;
  assign n48023 = x92 & n80926 ;
  assign n80927 = ~n47649 ;
  assign n48024 = n80927 & n48023 ;
  assign n48025 = n47656 | n48024 ;
  assign n48027 = n48022 | n48025 ;
  assign n80928 = ~n47656 ;
  assign n48028 = n80928 & n48027 ;
  assign n80929 = ~n47646 ;
  assign n48029 = x93 & n80929 ;
  assign n80930 = ~n47641 ;
  assign n48030 = n80930 & n48029 ;
  assign n48031 = n47648 | n48030 ;
  assign n48032 = n48028 | n48031 ;
  assign n80931 = ~n47648 ;
  assign n48033 = n80931 & n48032 ;
  assign n80932 = ~n47638 ;
  assign n48034 = x94 & n80932 ;
  assign n80933 = ~n47633 ;
  assign n48035 = n80933 & n48034 ;
  assign n48036 = n47640 | n48035 ;
  assign n48038 = n48033 | n48036 ;
  assign n80934 = ~n47640 ;
  assign n48039 = n80934 & n48038 ;
  assign n80935 = ~n47630 ;
  assign n48040 = x95 & n80935 ;
  assign n80936 = ~n47625 ;
  assign n48041 = n80936 & n48040 ;
  assign n48042 = n47632 | n48041 ;
  assign n48043 = n48039 | n48042 ;
  assign n80937 = ~n47632 ;
  assign n48044 = n80937 & n48043 ;
  assign n80938 = ~n47622 ;
  assign n48045 = x96 & n80938 ;
  assign n80939 = ~n47617 ;
  assign n48046 = n80939 & n48045 ;
  assign n48047 = n47624 | n48046 ;
  assign n48049 = n48044 | n48047 ;
  assign n80940 = ~n47624 ;
  assign n48050 = n80940 & n48049 ;
  assign n80941 = ~n47614 ;
  assign n48051 = x97 & n80941 ;
  assign n80942 = ~n47609 ;
  assign n48052 = n80942 & n48051 ;
  assign n48053 = n47616 | n48052 ;
  assign n48054 = n48050 | n48053 ;
  assign n80943 = ~n47616 ;
  assign n48055 = n80943 & n48054 ;
  assign n80944 = ~n47606 ;
  assign n48056 = x98 & n80944 ;
  assign n80945 = ~n47601 ;
  assign n48057 = n80945 & n48056 ;
  assign n48058 = n47608 | n48057 ;
  assign n48060 = n48055 | n48058 ;
  assign n80946 = ~n47608 ;
  assign n48061 = n80946 & n48060 ;
  assign n80947 = ~n47598 ;
  assign n48062 = x99 & n80947 ;
  assign n80948 = ~n47593 ;
  assign n48063 = n80948 & n48062 ;
  assign n48064 = n47600 | n48063 ;
  assign n48065 = n48061 | n48064 ;
  assign n80949 = ~n47600 ;
  assign n48066 = n80949 & n48065 ;
  assign n80950 = ~n47590 ;
  assign n48067 = x100 & n80950 ;
  assign n80951 = ~n47585 ;
  assign n48068 = n80951 & n48067 ;
  assign n48069 = n47592 | n48068 ;
  assign n48071 = n48066 | n48069 ;
  assign n80952 = ~n47592 ;
  assign n48072 = n80952 & n48071 ;
  assign n80953 = ~n47582 ;
  assign n48073 = x101 & n80953 ;
  assign n80954 = ~n47577 ;
  assign n48074 = n80954 & n48073 ;
  assign n48075 = n47584 | n48074 ;
  assign n48076 = n48072 | n48075 ;
  assign n80955 = ~n47584 ;
  assign n48077 = n80955 & n48076 ;
  assign n80956 = ~n47574 ;
  assign n48078 = x102 & n80956 ;
  assign n80957 = ~n47569 ;
  assign n48079 = n80957 & n48078 ;
  assign n48080 = n47576 | n48079 ;
  assign n48082 = n48077 | n48080 ;
  assign n80958 = ~n47576 ;
  assign n48083 = n80958 & n48082 ;
  assign n80959 = ~n47566 ;
  assign n48084 = x103 & n80959 ;
  assign n80960 = ~n47561 ;
  assign n48085 = n80960 & n48084 ;
  assign n48086 = n47568 | n48085 ;
  assign n48087 = n48083 | n48086 ;
  assign n80961 = ~n47568 ;
  assign n48088 = n80961 & n48087 ;
  assign n80962 = ~n47558 ;
  assign n48089 = x104 & n80962 ;
  assign n80963 = ~n47553 ;
  assign n48090 = n80963 & n48089 ;
  assign n48091 = n47560 | n48090 ;
  assign n48093 = n48088 | n48091 ;
  assign n80964 = ~n47560 ;
  assign n48094 = n80964 & n48093 ;
  assign n80965 = ~n47550 ;
  assign n48095 = x105 & n80965 ;
  assign n80966 = ~n47545 ;
  assign n48096 = n80966 & n48095 ;
  assign n48097 = n47552 | n48096 ;
  assign n48098 = n48094 | n48097 ;
  assign n80967 = ~n47552 ;
  assign n48099 = n80967 & n48098 ;
  assign n80968 = ~n47542 ;
  assign n48100 = x106 & n80968 ;
  assign n80969 = ~n47451 ;
  assign n48101 = n80969 & n48100 ;
  assign n48102 = n47544 | n48101 ;
  assign n48104 = n48099 | n48102 ;
  assign n80970 = ~n47544 ;
  assign n48105 = n80970 & n48104 ;
  assign n48112 = n70609 & n48111 ;
  assign n80971 = ~n47448 ;
  assign n48113 = n80971 & n48109 ;
  assign n48114 = n46878 & n47448 ;
  assign n80972 = ~n48114 ;
  assign n48115 = x107 & n80972 ;
  assign n80973 = ~n48113 ;
  assign n48116 = n80973 & n48115 ;
  assign n48117 = n15856 | n48116 ;
  assign n48118 = n48112 | n48117 ;
  assign n48120 = n48105 | n48118 ;
  assign n80974 = ~n48119 ;
  assign n48121 = n80974 & n48120 ;
  assign n80975 = ~n48099 ;
  assign n48103 = n80975 & n48102 ;
  assign n48124 = x65 & n47872 ;
  assign n80976 = ~n48124 ;
  assign n48125 = n47878 & n80976 ;
  assign n48126 = n15623 | n48125 ;
  assign n48127 = n80847 & n48126 ;
  assign n48128 = n47864 | n47884 ;
  assign n48130 = n48127 | n48128 ;
  assign n48131 = n80850 & n48130 ;
  assign n48132 = n47888 | n48131 ;
  assign n48134 = n80853 & n48132 ;
  assign n48136 = n47894 | n48134 ;
  assign n48137 = n80856 & n48136 ;
  assign n48139 = n47899 | n48137 ;
  assign n48140 = n80859 & n48139 ;
  assign n48141 = n47904 | n48140 ;
  assign n48142 = n80862 & n48141 ;
  assign n48143 = n47910 | n48142 ;
  assign n48145 = n80865 & n48143 ;
  assign n48146 = n47915 | n48145 ;
  assign n48147 = n80868 & n48146 ;
  assign n48148 = n47921 | n48147 ;
  assign n48150 = n80871 & n48148 ;
  assign n48151 = n47926 | n48150 ;
  assign n48152 = n80874 & n48151 ;
  assign n48153 = n47932 | n48152 ;
  assign n48155 = n80877 & n48153 ;
  assign n48156 = n47937 | n48155 ;
  assign n48157 = n80880 & n48156 ;
  assign n48158 = n47943 | n48157 ;
  assign n48160 = n80883 & n48158 ;
  assign n48161 = n47948 | n48160 ;
  assign n48162 = n80886 & n48161 ;
  assign n48163 = n47954 | n48162 ;
  assign n48165 = n80889 & n48163 ;
  assign n48166 = n47959 | n48165 ;
  assign n48167 = n80892 & n48166 ;
  assign n48168 = n47965 | n48167 ;
  assign n48170 = n80895 & n48168 ;
  assign n48171 = n47970 | n48170 ;
  assign n48172 = n80898 & n48171 ;
  assign n48173 = n47976 | n48172 ;
  assign n48175 = n80901 & n48173 ;
  assign n48176 = n47981 | n48175 ;
  assign n48177 = n80904 & n48176 ;
  assign n48178 = n47987 | n48177 ;
  assign n48180 = n80907 & n48178 ;
  assign n48181 = n47992 | n48180 ;
  assign n48182 = n80910 & n48181 ;
  assign n48183 = n47998 | n48182 ;
  assign n48185 = n80913 & n48183 ;
  assign n48186 = n48003 | n48185 ;
  assign n48187 = n80916 & n48186 ;
  assign n48188 = n48009 | n48187 ;
  assign n48190 = n80919 & n48188 ;
  assign n48191 = n48014 | n48190 ;
  assign n48192 = n80922 & n48191 ;
  assign n48193 = n48020 | n48192 ;
  assign n48195 = n80925 & n48193 ;
  assign n48196 = n48025 | n48195 ;
  assign n48197 = n80928 & n48196 ;
  assign n48198 = n48031 | n48197 ;
  assign n48200 = n80931 & n48198 ;
  assign n48201 = n48036 | n48200 ;
  assign n48202 = n80934 & n48201 ;
  assign n48203 = n48042 | n48202 ;
  assign n48205 = n80937 & n48203 ;
  assign n48206 = n48047 | n48205 ;
  assign n48207 = n80940 & n48206 ;
  assign n48208 = n48053 | n48207 ;
  assign n48210 = n80943 & n48208 ;
  assign n48211 = n48058 | n48210 ;
  assign n48212 = n80946 & n48211 ;
  assign n48213 = n48064 | n48212 ;
  assign n48215 = n80949 & n48213 ;
  assign n48216 = n48069 | n48215 ;
  assign n48217 = n80952 & n48216 ;
  assign n48218 = n48075 | n48217 ;
  assign n48220 = n80955 & n48218 ;
  assign n48221 = n48080 | n48220 ;
  assign n48222 = n80958 & n48221 ;
  assign n48223 = n48086 | n48222 ;
  assign n48225 = n80961 & n48223 ;
  assign n48226 = n48091 | n48225 ;
  assign n48227 = n80964 & n48226 ;
  assign n48228 = n48097 | n48227 ;
  assign n48230 = n47552 | n48102 ;
  assign n80977 = ~n48230 ;
  assign n48231 = n48228 & n80977 ;
  assign n48232 = n48103 | n48231 ;
  assign n80978 = ~n48121 ;
  assign n48233 = n80978 & n48232 ;
  assign n48234 = n80967 & n48228 ;
  assign n48235 = n48102 | n48234 ;
  assign n48236 = n80970 & n48235 ;
  assign n48237 = n48118 | n48236 ;
  assign n48238 = n47543 & n80974 ;
  assign n48239 = n48237 & n48238 ;
  assign n48240 = n48233 | n48239 ;
  assign n48241 = n70609 & n48240 ;
  assign n80979 = ~n48239 ;
  assign n48794 = x107 & n80979 ;
  assign n80980 = ~n48233 ;
  assign n48795 = n80980 & n48794 ;
  assign n48796 = n48241 | n48795 ;
  assign n80981 = ~n48227 ;
  assign n48229 = n48097 & n80981 ;
  assign n48242 = n47560 | n48097 ;
  assign n80982 = ~n48242 ;
  assign n48243 = n48093 & n80982 ;
  assign n48244 = n48229 | n48243 ;
  assign n48245 = n80978 & n48244 ;
  assign n48246 = n47551 & n80974 ;
  assign n48247 = n48237 & n48246 ;
  assign n48248 = n48245 | n48247 ;
  assign n48249 = n70276 & n48248 ;
  assign n80983 = ~n48088 ;
  assign n48092 = n80983 & n48091 ;
  assign n48250 = n47568 | n48091 ;
  assign n80984 = ~n48250 ;
  assign n48251 = n48223 & n80984 ;
  assign n48252 = n48092 | n48251 ;
  assign n48253 = n80978 & n48252 ;
  assign n48254 = n47559 & n80974 ;
  assign n48255 = n48237 & n48254 ;
  assign n48256 = n48253 | n48255 ;
  assign n48257 = n70176 & n48256 ;
  assign n80985 = ~n48255 ;
  assign n48784 = x105 & n80985 ;
  assign n80986 = ~n48253 ;
  assign n48785 = n80986 & n48784 ;
  assign n48786 = n48257 | n48785 ;
  assign n80987 = ~n48222 ;
  assign n48224 = n48086 & n80987 ;
  assign n48258 = n47576 | n48086 ;
  assign n80988 = ~n48258 ;
  assign n48259 = n48082 & n80988 ;
  assign n48260 = n48224 | n48259 ;
  assign n48261 = n80978 & n48260 ;
  assign n48262 = n47567 & n80974 ;
  assign n48263 = n48237 & n48262 ;
  assign n48264 = n48261 | n48263 ;
  assign n48265 = n69857 & n48264 ;
  assign n80989 = ~n48077 ;
  assign n48081 = n80989 & n48080 ;
  assign n48266 = n47584 | n48080 ;
  assign n80990 = ~n48266 ;
  assign n48267 = n48218 & n80990 ;
  assign n48268 = n48081 | n48267 ;
  assign n48269 = n80978 & n48268 ;
  assign n48270 = n47575 & n80974 ;
  assign n48271 = n48237 & n48270 ;
  assign n48272 = n48269 | n48271 ;
  assign n48273 = n69656 & n48272 ;
  assign n80991 = ~n48271 ;
  assign n48773 = x103 & n80991 ;
  assign n80992 = ~n48269 ;
  assign n48774 = n80992 & n48773 ;
  assign n48775 = n48273 | n48774 ;
  assign n80993 = ~n48217 ;
  assign n48219 = n48075 & n80993 ;
  assign n48274 = n47592 | n48075 ;
  assign n80994 = ~n48274 ;
  assign n48275 = n48071 & n80994 ;
  assign n48276 = n48219 | n48275 ;
  assign n48277 = n80978 & n48276 ;
  assign n48278 = n47583 & n80974 ;
  assign n48279 = n48237 & n48278 ;
  assign n48280 = n48277 | n48279 ;
  assign n48281 = n69528 & n48280 ;
  assign n80995 = ~n48066 ;
  assign n48070 = n80995 & n48069 ;
  assign n48282 = n47600 | n48069 ;
  assign n80996 = ~n48282 ;
  assign n48283 = n48213 & n80996 ;
  assign n48284 = n48070 | n48283 ;
  assign n48285 = n80978 & n48284 ;
  assign n48286 = n47591 & n80974 ;
  assign n48287 = n48237 & n48286 ;
  assign n48288 = n48285 | n48287 ;
  assign n48289 = n69261 & n48288 ;
  assign n80997 = ~n48287 ;
  assign n48763 = x101 & n80997 ;
  assign n80998 = ~n48285 ;
  assign n48764 = n80998 & n48763 ;
  assign n48765 = n48289 | n48764 ;
  assign n80999 = ~n48212 ;
  assign n48214 = n48064 & n80999 ;
  assign n48290 = n47608 | n48064 ;
  assign n81000 = ~n48290 ;
  assign n48291 = n48060 & n81000 ;
  assign n48292 = n48214 | n48291 ;
  assign n48293 = n80978 & n48292 ;
  assign n48294 = n47599 & n80974 ;
  assign n48295 = n48237 & n48294 ;
  assign n48296 = n48293 | n48295 ;
  assign n48297 = n69075 & n48296 ;
  assign n81001 = ~n48055 ;
  assign n48059 = n81001 & n48058 ;
  assign n48298 = n47616 | n48058 ;
  assign n81002 = ~n48298 ;
  assign n48299 = n48208 & n81002 ;
  assign n48300 = n48059 | n48299 ;
  assign n48301 = n80978 & n48300 ;
  assign n48302 = n47607 & n80974 ;
  assign n48303 = n48237 & n48302 ;
  assign n48304 = n48301 | n48303 ;
  assign n48305 = n68993 & n48304 ;
  assign n81003 = ~n48303 ;
  assign n48753 = x99 & n81003 ;
  assign n81004 = ~n48301 ;
  assign n48754 = n81004 & n48753 ;
  assign n48755 = n48305 | n48754 ;
  assign n81005 = ~n48207 ;
  assign n48209 = n48053 & n81005 ;
  assign n48306 = n47624 | n48053 ;
  assign n81006 = ~n48306 ;
  assign n48307 = n48049 & n81006 ;
  assign n48308 = n48209 | n48307 ;
  assign n48309 = n80978 & n48308 ;
  assign n48310 = n47615 & n80974 ;
  assign n48311 = n48237 & n48310 ;
  assign n48312 = n48309 | n48311 ;
  assign n48313 = n68716 & n48312 ;
  assign n81007 = ~n48044 ;
  assign n48048 = n81007 & n48047 ;
  assign n48314 = n47632 | n48047 ;
  assign n81008 = ~n48314 ;
  assign n48315 = n48203 & n81008 ;
  assign n48316 = n48048 | n48315 ;
  assign n48317 = n80978 & n48316 ;
  assign n48318 = n47623 & n80974 ;
  assign n48319 = n48237 & n48318 ;
  assign n48320 = n48317 | n48319 ;
  assign n48321 = n68545 & n48320 ;
  assign n81009 = ~n48319 ;
  assign n48743 = x97 & n81009 ;
  assign n81010 = ~n48317 ;
  assign n48744 = n81010 & n48743 ;
  assign n48745 = n48321 | n48744 ;
  assign n81011 = ~n48202 ;
  assign n48204 = n48042 & n81011 ;
  assign n48322 = n47640 | n48042 ;
  assign n81012 = ~n48322 ;
  assign n48323 = n48038 & n81012 ;
  assign n48324 = n48204 | n48323 ;
  assign n48325 = n80978 & n48324 ;
  assign n48326 = n47631 & n80974 ;
  assign n48327 = n48237 & n48326 ;
  assign n48328 = n48325 | n48327 ;
  assign n48329 = n68438 & n48328 ;
  assign n81013 = ~n48033 ;
  assign n48037 = n81013 & n48036 ;
  assign n48330 = n47648 | n48036 ;
  assign n81014 = ~n48330 ;
  assign n48331 = n48198 & n81014 ;
  assign n48332 = n48037 | n48331 ;
  assign n48333 = n80978 & n48332 ;
  assign n48334 = n47639 & n80974 ;
  assign n48335 = n48237 & n48334 ;
  assign n48336 = n48333 | n48335 ;
  assign n48337 = n68214 & n48336 ;
  assign n81015 = ~n48335 ;
  assign n48733 = x95 & n81015 ;
  assign n81016 = ~n48333 ;
  assign n48734 = n81016 & n48733 ;
  assign n48735 = n48337 | n48734 ;
  assign n81017 = ~n48197 ;
  assign n48199 = n48031 & n81017 ;
  assign n48338 = n47656 | n48031 ;
  assign n81018 = ~n48338 ;
  assign n48339 = n48027 & n81018 ;
  assign n48340 = n48199 | n48339 ;
  assign n48341 = n80978 & n48340 ;
  assign n48342 = n47647 & n80974 ;
  assign n48343 = n48237 & n48342 ;
  assign n48344 = n48341 | n48343 ;
  assign n48345 = n68058 & n48344 ;
  assign n81019 = ~n48022 ;
  assign n48026 = n81019 & n48025 ;
  assign n48346 = n47664 | n48025 ;
  assign n81020 = ~n48346 ;
  assign n48347 = n48193 & n81020 ;
  assign n48348 = n48026 | n48347 ;
  assign n48349 = n80978 & n48348 ;
  assign n48350 = n47655 & n80974 ;
  assign n48351 = n48237 & n48350 ;
  assign n48352 = n48349 | n48351 ;
  assign n48353 = n67986 & n48352 ;
  assign n81021 = ~n48351 ;
  assign n48722 = x93 & n81021 ;
  assign n81022 = ~n48349 ;
  assign n48723 = n81022 & n48722 ;
  assign n48724 = n48353 | n48723 ;
  assign n81023 = ~n48192 ;
  assign n48194 = n48020 & n81023 ;
  assign n48354 = n47672 | n48020 ;
  assign n81024 = ~n48354 ;
  assign n48355 = n48016 & n81024 ;
  assign n48356 = n48194 | n48355 ;
  assign n48357 = n80978 & n48356 ;
  assign n48358 = n47663 & n80974 ;
  assign n48359 = n48237 & n48358 ;
  assign n48360 = n48357 | n48359 ;
  assign n48361 = n67763 & n48360 ;
  assign n81025 = ~n48011 ;
  assign n48015 = n81025 & n48014 ;
  assign n48362 = n47680 | n48014 ;
  assign n81026 = ~n48362 ;
  assign n48363 = n48188 & n81026 ;
  assign n48364 = n48015 | n48363 ;
  assign n48365 = n80978 & n48364 ;
  assign n48366 = n47671 & n80974 ;
  assign n48367 = n48237 & n48366 ;
  assign n48368 = n48365 | n48367 ;
  assign n48369 = n67622 & n48368 ;
  assign n81027 = ~n48367 ;
  assign n48712 = x91 & n81027 ;
  assign n81028 = ~n48365 ;
  assign n48713 = n81028 & n48712 ;
  assign n48714 = n48369 | n48713 ;
  assign n81029 = ~n48187 ;
  assign n48189 = n48009 & n81029 ;
  assign n48370 = n47688 | n48009 ;
  assign n81030 = ~n48370 ;
  assign n48371 = n48005 & n81030 ;
  assign n48372 = n48189 | n48371 ;
  assign n48373 = n80978 & n48372 ;
  assign n48374 = n47679 & n80974 ;
  assign n48375 = n48237 & n48374 ;
  assign n48376 = n48373 | n48375 ;
  assign n48377 = n67531 & n48376 ;
  assign n81031 = ~n48000 ;
  assign n48004 = n81031 & n48003 ;
  assign n48378 = n47696 | n48003 ;
  assign n81032 = ~n48378 ;
  assign n48379 = n48183 & n81032 ;
  assign n48380 = n48004 | n48379 ;
  assign n48381 = n80978 & n48380 ;
  assign n48382 = n47687 & n80974 ;
  assign n48383 = n48237 & n48382 ;
  assign n48384 = n48381 | n48383 ;
  assign n48385 = n67348 & n48384 ;
  assign n81033 = ~n48383 ;
  assign n48702 = x89 & n81033 ;
  assign n81034 = ~n48381 ;
  assign n48703 = n81034 & n48702 ;
  assign n48704 = n48385 | n48703 ;
  assign n81035 = ~n48182 ;
  assign n48184 = n47998 & n81035 ;
  assign n48386 = n47704 | n47998 ;
  assign n81036 = ~n48386 ;
  assign n48387 = n47994 & n81036 ;
  assign n48388 = n48184 | n48387 ;
  assign n48389 = n80978 & n48388 ;
  assign n48390 = n47695 & n80974 ;
  assign n48391 = n48237 & n48390 ;
  assign n48392 = n48389 | n48391 ;
  assign n48393 = n67222 & n48392 ;
  assign n81037 = ~n47989 ;
  assign n47993 = n81037 & n47992 ;
  assign n48394 = n47712 | n47992 ;
  assign n81038 = ~n48394 ;
  assign n48395 = n48178 & n81038 ;
  assign n48396 = n47993 | n48395 ;
  assign n48397 = n80978 & n48396 ;
  assign n48398 = n47703 & n80974 ;
  assign n48399 = n48237 & n48398 ;
  assign n48400 = n48397 | n48399 ;
  assign n48401 = n67164 & n48400 ;
  assign n81039 = ~n48399 ;
  assign n48692 = x87 & n81039 ;
  assign n81040 = ~n48397 ;
  assign n48693 = n81040 & n48692 ;
  assign n48694 = n48401 | n48693 ;
  assign n81041 = ~n48177 ;
  assign n48179 = n47987 & n81041 ;
  assign n48402 = n47720 | n47987 ;
  assign n81042 = ~n48402 ;
  assign n48403 = n47983 & n81042 ;
  assign n48404 = n48179 | n48403 ;
  assign n48405 = n80978 & n48404 ;
  assign n48406 = n47711 & n80974 ;
  assign n48407 = n48237 & n48406 ;
  assign n48408 = n48405 | n48407 ;
  assign n48409 = n66979 & n48408 ;
  assign n81043 = ~n47978 ;
  assign n47982 = n81043 & n47981 ;
  assign n48410 = n47728 | n47981 ;
  assign n81044 = ~n48410 ;
  assign n48411 = n48173 & n81044 ;
  assign n48412 = n47982 | n48411 ;
  assign n48413 = n80978 & n48412 ;
  assign n48414 = n47719 & n80974 ;
  assign n48415 = n48237 & n48414 ;
  assign n48416 = n48413 | n48415 ;
  assign n48417 = n66868 & n48416 ;
  assign n81045 = ~n48415 ;
  assign n48682 = x85 & n81045 ;
  assign n81046 = ~n48413 ;
  assign n48683 = n81046 & n48682 ;
  assign n48684 = n48417 | n48683 ;
  assign n81047 = ~n48172 ;
  assign n48174 = n47976 & n81047 ;
  assign n48418 = n47736 | n47976 ;
  assign n81048 = ~n48418 ;
  assign n48419 = n47972 & n81048 ;
  assign n48420 = n48174 | n48419 ;
  assign n48421 = n80978 & n48420 ;
  assign n48422 = n47727 & n80974 ;
  assign n48423 = n48237 & n48422 ;
  assign n48424 = n48421 | n48423 ;
  assign n48425 = n66797 & n48424 ;
  assign n81049 = ~n47967 ;
  assign n47971 = n81049 & n47970 ;
  assign n48426 = n47744 | n47970 ;
  assign n81050 = ~n48426 ;
  assign n48427 = n48168 & n81050 ;
  assign n48428 = n47971 | n48427 ;
  assign n48429 = n80978 & n48428 ;
  assign n48430 = n47735 & n80974 ;
  assign n48431 = n48237 & n48430 ;
  assign n48432 = n48429 | n48431 ;
  assign n48433 = n66654 & n48432 ;
  assign n81051 = ~n48431 ;
  assign n48672 = x83 & n81051 ;
  assign n81052 = ~n48429 ;
  assign n48673 = n81052 & n48672 ;
  assign n48674 = n48433 | n48673 ;
  assign n81053 = ~n48167 ;
  assign n48169 = n47965 & n81053 ;
  assign n48434 = n47752 | n47965 ;
  assign n81054 = ~n48434 ;
  assign n48435 = n47961 & n81054 ;
  assign n48436 = n48169 | n48435 ;
  assign n48437 = n80978 & n48436 ;
  assign n48438 = n47743 & n80974 ;
  assign n48439 = n48237 & n48438 ;
  assign n48440 = n48437 | n48439 ;
  assign n48441 = n66560 & n48440 ;
  assign n81055 = ~n47956 ;
  assign n47960 = n81055 & n47959 ;
  assign n48442 = n47760 | n47959 ;
  assign n81056 = ~n48442 ;
  assign n48443 = n48163 & n81056 ;
  assign n48444 = n47960 | n48443 ;
  assign n48445 = n80978 & n48444 ;
  assign n48446 = n47751 & n80974 ;
  assign n48447 = n48237 & n48446 ;
  assign n48448 = n48445 | n48447 ;
  assign n48449 = n66505 & n48448 ;
  assign n81057 = ~n48447 ;
  assign n48662 = x81 & n81057 ;
  assign n81058 = ~n48445 ;
  assign n48663 = n81058 & n48662 ;
  assign n48664 = n48449 | n48663 ;
  assign n81059 = ~n48162 ;
  assign n48164 = n47954 & n81059 ;
  assign n48450 = n47768 | n47954 ;
  assign n81060 = ~n48450 ;
  assign n48451 = n47950 & n81060 ;
  assign n48452 = n48164 | n48451 ;
  assign n48453 = n80978 & n48452 ;
  assign n48454 = n47759 & n80974 ;
  assign n48455 = n48237 & n48454 ;
  assign n48456 = n48453 | n48455 ;
  assign n48457 = n66379 & n48456 ;
  assign n81061 = ~n47945 ;
  assign n47949 = n81061 & n47948 ;
  assign n48458 = n47776 | n47948 ;
  assign n81062 = ~n48458 ;
  assign n48459 = n48158 & n81062 ;
  assign n48460 = n47949 | n48459 ;
  assign n48461 = n80978 & n48460 ;
  assign n48462 = n47767 & n80974 ;
  assign n48463 = n48237 & n48462 ;
  assign n48464 = n48461 | n48463 ;
  assign n48465 = n66299 & n48464 ;
  assign n81063 = ~n48463 ;
  assign n48652 = x79 & n81063 ;
  assign n81064 = ~n48461 ;
  assign n48653 = n81064 & n48652 ;
  assign n48654 = n48465 | n48653 ;
  assign n81065 = ~n48157 ;
  assign n48159 = n47943 & n81065 ;
  assign n48466 = n47784 | n47943 ;
  assign n81066 = ~n48466 ;
  assign n48467 = n47939 & n81066 ;
  assign n48468 = n48159 | n48467 ;
  assign n48469 = n80978 & n48468 ;
  assign n48470 = n47775 & n80974 ;
  assign n48471 = n48237 & n48470 ;
  assign n48472 = n48469 | n48471 ;
  assign n48473 = n66244 & n48472 ;
  assign n81067 = ~n47934 ;
  assign n47938 = n81067 & n47937 ;
  assign n48474 = n47792 | n47937 ;
  assign n81068 = ~n48474 ;
  assign n48475 = n48153 & n81068 ;
  assign n48476 = n47938 | n48475 ;
  assign n48477 = n80978 & n48476 ;
  assign n48478 = n47783 & n80974 ;
  assign n48479 = n48237 & n48478 ;
  assign n48480 = n48477 | n48479 ;
  assign n48481 = n66145 & n48480 ;
  assign n81069 = ~n48479 ;
  assign n48641 = x77 & n81069 ;
  assign n81070 = ~n48477 ;
  assign n48642 = n81070 & n48641 ;
  assign n48643 = n48481 | n48642 ;
  assign n81071 = ~n48152 ;
  assign n48154 = n47932 & n81071 ;
  assign n48482 = n47800 | n47932 ;
  assign n81072 = ~n48482 ;
  assign n48483 = n47928 & n81072 ;
  assign n48484 = n48154 | n48483 ;
  assign n48485 = n80978 & n48484 ;
  assign n48486 = n47791 & n80974 ;
  assign n48487 = n48237 & n48486 ;
  assign n48488 = n48485 | n48487 ;
  assign n48489 = n66081 & n48488 ;
  assign n81073 = ~n47923 ;
  assign n47927 = n81073 & n47926 ;
  assign n48490 = n47808 | n47926 ;
  assign n81074 = ~n48490 ;
  assign n48491 = n48148 & n81074 ;
  assign n48492 = n47927 | n48491 ;
  assign n48493 = n80978 & n48492 ;
  assign n48494 = n47799 & n80974 ;
  assign n48495 = n48237 & n48494 ;
  assign n48496 = n48493 | n48495 ;
  assign n48497 = n66043 & n48496 ;
  assign n81075 = ~n48495 ;
  assign n48631 = x75 & n81075 ;
  assign n81076 = ~n48493 ;
  assign n48632 = n81076 & n48631 ;
  assign n48633 = n48497 | n48632 ;
  assign n81077 = ~n48147 ;
  assign n48149 = n47921 & n81077 ;
  assign n48498 = n47816 | n47921 ;
  assign n81078 = ~n48498 ;
  assign n48499 = n47917 & n81078 ;
  assign n48500 = n48149 | n48499 ;
  assign n48501 = n80978 & n48500 ;
  assign n48502 = n47807 & n80974 ;
  assign n48503 = n48237 & n48502 ;
  assign n48504 = n48501 | n48503 ;
  assign n48505 = n65960 & n48504 ;
  assign n81079 = ~n47912 ;
  assign n47916 = n81079 & n47915 ;
  assign n48506 = n47824 | n47915 ;
  assign n81080 = ~n48506 ;
  assign n48507 = n48143 & n81080 ;
  assign n48508 = n47916 | n48507 ;
  assign n48509 = n80978 & n48508 ;
  assign n48510 = n47815 & n80974 ;
  assign n48511 = n48237 & n48510 ;
  assign n48512 = n48509 | n48511 ;
  assign n48513 = n65909 & n48512 ;
  assign n81081 = ~n48511 ;
  assign n48620 = x73 & n81081 ;
  assign n81082 = ~n48509 ;
  assign n48621 = n81082 & n48620 ;
  assign n48622 = n48513 | n48621 ;
  assign n81083 = ~n48142 ;
  assign n48144 = n47910 & n81083 ;
  assign n48514 = n47832 | n47910 ;
  assign n81084 = ~n48514 ;
  assign n48515 = n47906 & n81084 ;
  assign n48516 = n48144 | n48515 ;
  assign n48517 = n80978 & n48516 ;
  assign n48518 = n47823 & n80974 ;
  assign n48519 = n48237 & n48518 ;
  assign n48520 = n48517 | n48519 ;
  assign n48521 = n65877 & n48520 ;
  assign n81085 = ~n47901 ;
  assign n47905 = n81085 & n47904 ;
  assign n48522 = n47841 | n47904 ;
  assign n81086 = ~n48522 ;
  assign n48523 = n48139 & n81086 ;
  assign n48524 = n47905 | n48523 ;
  assign n48525 = n80978 & n48524 ;
  assign n48526 = n47831 & n80974 ;
  assign n48527 = n48237 & n48526 ;
  assign n48528 = n48525 | n48527 ;
  assign n48529 = n65820 & n48528 ;
  assign n81087 = ~n48527 ;
  assign n48609 = x71 & n81087 ;
  assign n81088 = ~n48525 ;
  assign n48610 = n81088 & n48609 ;
  assign n48611 = n48529 | n48610 ;
  assign n81089 = ~n48137 ;
  assign n48138 = n47899 & n81089 ;
  assign n48530 = n47850 | n47899 ;
  assign n81090 = ~n48530 ;
  assign n48531 = n47895 & n81090 ;
  assign n48532 = n48138 | n48531 ;
  assign n48533 = n80978 & n48532 ;
  assign n48534 = n47840 & n80974 ;
  assign n48535 = n48237 & n48534 ;
  assign n48536 = n48533 | n48535 ;
  assign n48537 = n65791 & n48536 ;
  assign n81091 = ~n47891 ;
  assign n48135 = n81091 & n47894 ;
  assign n48538 = n47889 | n48131 ;
  assign n48539 = n47858 | n47894 ;
  assign n81092 = ~n48539 ;
  assign n48540 = n48538 & n81092 ;
  assign n48541 = n48135 | n48540 ;
  assign n48542 = n80978 & n48541 ;
  assign n48543 = n47849 & n80974 ;
  assign n48544 = n48237 & n48543 ;
  assign n48545 = n48542 | n48544 ;
  assign n48546 = n65772 & n48545 ;
  assign n81093 = ~n48544 ;
  assign n48599 = x69 & n81093 ;
  assign n81094 = ~n48542 ;
  assign n48600 = n81094 & n48599 ;
  assign n48601 = n48546 | n48600 ;
  assign n81095 = ~n48131 ;
  assign n48133 = n47889 & n81095 ;
  assign n48547 = n47864 | n47889 ;
  assign n81096 = ~n48547 ;
  assign n48548 = n48130 & n81096 ;
  assign n48549 = n48133 | n48548 ;
  assign n48550 = n80978 & n48549 ;
  assign n48551 = n47857 & n80974 ;
  assign n48552 = n48237 & n48551 ;
  assign n48553 = n48550 | n48552 ;
  assign n48554 = n65746 & n48553 ;
  assign n81097 = ~n47882 ;
  assign n48129 = n81097 & n48128 ;
  assign n48555 = n47880 | n48128 ;
  assign n81098 = ~n48555 ;
  assign n48556 = n47881 & n81098 ;
  assign n48557 = n48129 | n48556 ;
  assign n48558 = n80978 & n48557 ;
  assign n48559 = n47863 & n80974 ;
  assign n48560 = n48237 & n48559 ;
  assign n48561 = n48558 | n48560 ;
  assign n48562 = n65721 & n48561 ;
  assign n81099 = ~n48560 ;
  assign n48589 = x67 & n81099 ;
  assign n81100 = ~n48558 ;
  assign n48590 = n81100 & n48589 ;
  assign n48591 = n48562 | n48590 ;
  assign n48563 = n15623 & n47878 ;
  assign n48564 = n80976 & n48563 ;
  assign n81101 = ~n48564 ;
  assign n48565 = n47881 & n81101 ;
  assign n48566 = n80978 & n48565 ;
  assign n48567 = n47875 & n80974 ;
  assign n48568 = n48237 & n48567 ;
  assign n48569 = n48566 | n48568 ;
  assign n48570 = n65686 & n48569 ;
  assign n48123 = n15623 & n80978 ;
  assign n48571 = n80974 & n48237 ;
  assign n81102 = ~n48571 ;
  assign n48572 = x64 & n81102 ;
  assign n81103 = ~n48572 ;
  assign n48573 = x20 & n81103 ;
  assign n48574 = n48123 | n48573 ;
  assign n48575 = x65 & n48574 ;
  assign n48122 = x64 & n80978 ;
  assign n81104 = ~n48122 ;
  assign n48576 = x20 & n81104 ;
  assign n48577 = n15623 & n81102 ;
  assign n48578 = x65 | n48577 ;
  assign n48579 = n48576 | n48578 ;
  assign n81105 = ~n48575 ;
  assign n48580 = n81105 & n48579 ;
  assign n48581 = n16327 | n48580 ;
  assign n48582 = n48123 | n48576 ;
  assign n48583 = n65670 & n48582 ;
  assign n81106 = ~n48583 ;
  assign n48584 = n48581 & n81106 ;
  assign n81107 = ~n48568 ;
  assign n48585 = x66 & n81107 ;
  assign n81108 = ~n48566 ;
  assign n48586 = n81108 & n48585 ;
  assign n48587 = n48570 | n48586 ;
  assign n48588 = n48584 | n48587 ;
  assign n81109 = ~n48570 ;
  assign n48592 = n81109 & n48588 ;
  assign n48593 = n48591 | n48592 ;
  assign n81110 = ~n48562 ;
  assign n48594 = n81110 & n48593 ;
  assign n81111 = ~n48552 ;
  assign n48595 = x68 & n81111 ;
  assign n81112 = ~n48550 ;
  assign n48596 = n81112 & n48595 ;
  assign n48597 = n48554 | n48596 ;
  assign n48598 = n48594 | n48597 ;
  assign n81113 = ~n48554 ;
  assign n48602 = n81113 & n48598 ;
  assign n48603 = n48601 | n48602 ;
  assign n81114 = ~n48546 ;
  assign n48604 = n81114 & n48603 ;
  assign n81115 = ~n48535 ;
  assign n48605 = x70 & n81115 ;
  assign n81116 = ~n48533 ;
  assign n48606 = n81116 & n48605 ;
  assign n48607 = n48537 | n48606 ;
  assign n48608 = n48604 | n48607 ;
  assign n81117 = ~n48537 ;
  assign n48613 = n81117 & n48608 ;
  assign n48614 = n48611 | n48613 ;
  assign n81118 = ~n48529 ;
  assign n48615 = n81118 & n48614 ;
  assign n81119 = ~n48519 ;
  assign n48616 = x72 & n81119 ;
  assign n81120 = ~n48517 ;
  assign n48617 = n81120 & n48616 ;
  assign n48618 = n48521 | n48617 ;
  assign n48619 = n48615 | n48618 ;
  assign n81121 = ~n48521 ;
  assign n48624 = n81121 & n48619 ;
  assign n48625 = n48622 | n48624 ;
  assign n81122 = ~n48513 ;
  assign n48626 = n81122 & n48625 ;
  assign n81123 = ~n48503 ;
  assign n48627 = x74 & n81123 ;
  assign n81124 = ~n48501 ;
  assign n48628 = n81124 & n48627 ;
  assign n48629 = n48505 | n48628 ;
  assign n48630 = n48626 | n48629 ;
  assign n81125 = ~n48505 ;
  assign n48634 = n81125 & n48630 ;
  assign n48635 = n48633 | n48634 ;
  assign n81126 = ~n48497 ;
  assign n48636 = n81126 & n48635 ;
  assign n81127 = ~n48487 ;
  assign n48637 = x76 & n81127 ;
  assign n81128 = ~n48485 ;
  assign n48638 = n81128 & n48637 ;
  assign n48639 = n48489 | n48638 ;
  assign n48640 = n48636 | n48639 ;
  assign n81129 = ~n48489 ;
  assign n48645 = n81129 & n48640 ;
  assign n48646 = n48643 | n48645 ;
  assign n81130 = ~n48481 ;
  assign n48647 = n81130 & n48646 ;
  assign n81131 = ~n48471 ;
  assign n48648 = x78 & n81131 ;
  assign n81132 = ~n48469 ;
  assign n48649 = n81132 & n48648 ;
  assign n48650 = n48473 | n48649 ;
  assign n48651 = n48647 | n48650 ;
  assign n81133 = ~n48473 ;
  assign n48655 = n81133 & n48651 ;
  assign n48656 = n48654 | n48655 ;
  assign n81134 = ~n48465 ;
  assign n48657 = n81134 & n48656 ;
  assign n81135 = ~n48455 ;
  assign n48658 = x80 & n81135 ;
  assign n81136 = ~n48453 ;
  assign n48659 = n81136 & n48658 ;
  assign n48660 = n48457 | n48659 ;
  assign n48661 = n48657 | n48660 ;
  assign n81137 = ~n48457 ;
  assign n48665 = n81137 & n48661 ;
  assign n48666 = n48664 | n48665 ;
  assign n81138 = ~n48449 ;
  assign n48667 = n81138 & n48666 ;
  assign n81139 = ~n48439 ;
  assign n48668 = x82 & n81139 ;
  assign n81140 = ~n48437 ;
  assign n48669 = n81140 & n48668 ;
  assign n48670 = n48441 | n48669 ;
  assign n48671 = n48667 | n48670 ;
  assign n81141 = ~n48441 ;
  assign n48675 = n81141 & n48671 ;
  assign n48676 = n48674 | n48675 ;
  assign n81142 = ~n48433 ;
  assign n48677 = n81142 & n48676 ;
  assign n81143 = ~n48423 ;
  assign n48678 = x84 & n81143 ;
  assign n81144 = ~n48421 ;
  assign n48679 = n81144 & n48678 ;
  assign n48680 = n48425 | n48679 ;
  assign n48681 = n48677 | n48680 ;
  assign n81145 = ~n48425 ;
  assign n48685 = n81145 & n48681 ;
  assign n48686 = n48684 | n48685 ;
  assign n81146 = ~n48417 ;
  assign n48687 = n81146 & n48686 ;
  assign n81147 = ~n48407 ;
  assign n48688 = x86 & n81147 ;
  assign n81148 = ~n48405 ;
  assign n48689 = n81148 & n48688 ;
  assign n48690 = n48409 | n48689 ;
  assign n48691 = n48687 | n48690 ;
  assign n81149 = ~n48409 ;
  assign n48695 = n81149 & n48691 ;
  assign n48696 = n48694 | n48695 ;
  assign n81150 = ~n48401 ;
  assign n48697 = n81150 & n48696 ;
  assign n81151 = ~n48391 ;
  assign n48698 = x88 & n81151 ;
  assign n81152 = ~n48389 ;
  assign n48699 = n81152 & n48698 ;
  assign n48700 = n48393 | n48699 ;
  assign n48701 = n48697 | n48700 ;
  assign n81153 = ~n48393 ;
  assign n48705 = n81153 & n48701 ;
  assign n48706 = n48704 | n48705 ;
  assign n81154 = ~n48385 ;
  assign n48707 = n81154 & n48706 ;
  assign n81155 = ~n48375 ;
  assign n48708 = x90 & n81155 ;
  assign n81156 = ~n48373 ;
  assign n48709 = n81156 & n48708 ;
  assign n48710 = n48377 | n48709 ;
  assign n48711 = n48707 | n48710 ;
  assign n81157 = ~n48377 ;
  assign n48715 = n81157 & n48711 ;
  assign n48716 = n48714 | n48715 ;
  assign n81158 = ~n48369 ;
  assign n48717 = n81158 & n48716 ;
  assign n81159 = ~n48359 ;
  assign n48718 = x92 & n81159 ;
  assign n81160 = ~n48357 ;
  assign n48719 = n81160 & n48718 ;
  assign n48720 = n48361 | n48719 ;
  assign n48721 = n48717 | n48720 ;
  assign n81161 = ~n48361 ;
  assign n48725 = n81161 & n48721 ;
  assign n48726 = n48724 | n48725 ;
  assign n81162 = ~n48353 ;
  assign n48727 = n81162 & n48726 ;
  assign n81163 = ~n48343 ;
  assign n48728 = x94 & n81163 ;
  assign n81164 = ~n48341 ;
  assign n48729 = n81164 & n48728 ;
  assign n48730 = n48345 | n48729 ;
  assign n48732 = n48727 | n48730 ;
  assign n81165 = ~n48345 ;
  assign n48736 = n81165 & n48732 ;
  assign n48737 = n48735 | n48736 ;
  assign n81166 = ~n48337 ;
  assign n48738 = n81166 & n48737 ;
  assign n81167 = ~n48327 ;
  assign n48739 = x96 & n81167 ;
  assign n81168 = ~n48325 ;
  assign n48740 = n81168 & n48739 ;
  assign n48741 = n48329 | n48740 ;
  assign n48742 = n48738 | n48741 ;
  assign n81169 = ~n48329 ;
  assign n48746 = n81169 & n48742 ;
  assign n48747 = n48745 | n48746 ;
  assign n81170 = ~n48321 ;
  assign n48748 = n81170 & n48747 ;
  assign n81171 = ~n48311 ;
  assign n48749 = x98 & n81171 ;
  assign n81172 = ~n48309 ;
  assign n48750 = n81172 & n48749 ;
  assign n48751 = n48313 | n48750 ;
  assign n48752 = n48748 | n48751 ;
  assign n81173 = ~n48313 ;
  assign n48756 = n81173 & n48752 ;
  assign n48757 = n48755 | n48756 ;
  assign n81174 = ~n48305 ;
  assign n48758 = n81174 & n48757 ;
  assign n81175 = ~n48295 ;
  assign n48759 = x100 & n81175 ;
  assign n81176 = ~n48293 ;
  assign n48760 = n81176 & n48759 ;
  assign n48761 = n48297 | n48760 ;
  assign n48762 = n48758 | n48761 ;
  assign n81177 = ~n48297 ;
  assign n48766 = n81177 & n48762 ;
  assign n48767 = n48765 | n48766 ;
  assign n81178 = ~n48289 ;
  assign n48768 = n81178 & n48767 ;
  assign n81179 = ~n48279 ;
  assign n48769 = x102 & n81179 ;
  assign n81180 = ~n48277 ;
  assign n48770 = n81180 & n48769 ;
  assign n48771 = n48281 | n48770 ;
  assign n48772 = n48768 | n48771 ;
  assign n81181 = ~n48281 ;
  assign n48777 = n81181 & n48772 ;
  assign n48778 = n48775 | n48777 ;
  assign n81182 = ~n48273 ;
  assign n48779 = n81182 & n48778 ;
  assign n81183 = ~n48263 ;
  assign n48780 = x104 & n81183 ;
  assign n81184 = ~n48261 ;
  assign n48781 = n81184 & n48780 ;
  assign n48782 = n48265 | n48781 ;
  assign n48783 = n48779 | n48782 ;
  assign n81185 = ~n48265 ;
  assign n48787 = n81185 & n48783 ;
  assign n48788 = n48786 | n48787 ;
  assign n81186 = ~n48257 ;
  assign n48789 = n81186 & n48788 ;
  assign n81187 = ~n48247 ;
  assign n48790 = x106 & n81187 ;
  assign n81188 = ~n48245 ;
  assign n48791 = n81188 & n48790 ;
  assign n48792 = n48249 | n48791 ;
  assign n48793 = n48789 | n48792 ;
  assign n81189 = ~n48249 ;
  assign n48797 = n81189 & n48793 ;
  assign n48798 = n48796 | n48797 ;
  assign n81190 = ~n48241 ;
  assign n48799 = n81190 & n48798 ;
  assign n48800 = n47544 | n48116 ;
  assign n48801 = n48112 | n48800 ;
  assign n81191 = ~n48801 ;
  assign n48802 = n48104 & n81191 ;
  assign n48803 = n48112 | n48116 ;
  assign n81192 = ~n48236 ;
  assign n48804 = n81192 & n48803 ;
  assign n48805 = n48802 | n48804 ;
  assign n48806 = n80978 & n48805 ;
  assign n48807 = n15167 & n46878 ;
  assign n48808 = n48237 & n48807 ;
  assign n48809 = n48806 | n48808 ;
  assign n48810 = n70927 & n48809 ;
  assign n81193 = ~n48808 ;
  assign n48811 = x108 & n81193 ;
  assign n81194 = ~n48806 ;
  assign n48812 = n81194 & n48811 ;
  assign n48813 = n16574 | n48812 ;
  assign n48814 = n48810 | n48813 ;
  assign n48815 = n48799 | n48814 ;
  assign n48816 = n70711 & n48809 ;
  assign n81195 = ~n48816 ;
  assign n48817 = n48815 & n81195 ;
  assign n81196 = ~n48797 ;
  assign n48906 = n48796 & n81196 ;
  assign n48819 = x65 & n48582 ;
  assign n81197 = ~n48819 ;
  assign n48820 = n48579 & n81197 ;
  assign n48821 = n16327 | n48820 ;
  assign n48823 = n81106 & n48821 ;
  assign n48824 = n48587 | n48823 ;
  assign n48825 = n81109 & n48824 ;
  assign n48826 = n48591 | n48825 ;
  assign n48827 = n81110 & n48826 ;
  assign n48828 = n48597 | n48827 ;
  assign n48829 = n81113 & n48828 ;
  assign n48830 = n48601 | n48829 ;
  assign n48831 = n81114 & n48830 ;
  assign n48832 = n48607 | n48831 ;
  assign n48833 = n81117 & n48832 ;
  assign n48834 = n48611 | n48833 ;
  assign n48835 = n81118 & n48834 ;
  assign n48836 = n48618 | n48835 ;
  assign n48837 = n81121 & n48836 ;
  assign n48838 = n48622 | n48837 ;
  assign n48839 = n81122 & n48838 ;
  assign n48840 = n48629 | n48839 ;
  assign n48841 = n81125 & n48840 ;
  assign n48842 = n48633 | n48841 ;
  assign n48843 = n81126 & n48842 ;
  assign n48844 = n48639 | n48843 ;
  assign n48845 = n81129 & n48844 ;
  assign n48846 = n48643 | n48845 ;
  assign n48847 = n81130 & n48846 ;
  assign n48848 = n48650 | n48847 ;
  assign n48849 = n81133 & n48848 ;
  assign n48850 = n48654 | n48849 ;
  assign n48851 = n81134 & n48850 ;
  assign n48852 = n48660 | n48851 ;
  assign n48853 = n81137 & n48852 ;
  assign n48854 = n48664 | n48853 ;
  assign n48855 = n81138 & n48854 ;
  assign n48856 = n48670 | n48855 ;
  assign n48857 = n81141 & n48856 ;
  assign n48858 = n48674 | n48857 ;
  assign n48859 = n81142 & n48858 ;
  assign n48860 = n48680 | n48859 ;
  assign n48861 = n81145 & n48860 ;
  assign n48862 = n48684 | n48861 ;
  assign n48863 = n81146 & n48862 ;
  assign n48864 = n48690 | n48863 ;
  assign n48865 = n81149 & n48864 ;
  assign n48866 = n48694 | n48865 ;
  assign n48867 = n81150 & n48866 ;
  assign n48868 = n48700 | n48867 ;
  assign n48869 = n81153 & n48868 ;
  assign n48870 = n48704 | n48869 ;
  assign n48871 = n81154 & n48870 ;
  assign n48872 = n48710 | n48871 ;
  assign n48873 = n81157 & n48872 ;
  assign n48874 = n48714 | n48873 ;
  assign n48875 = n81158 & n48874 ;
  assign n48876 = n48720 | n48875 ;
  assign n48877 = n81161 & n48876 ;
  assign n48878 = n48724 | n48877 ;
  assign n48879 = n81162 & n48878 ;
  assign n48880 = n48730 | n48879 ;
  assign n48881 = n81165 & n48880 ;
  assign n48882 = n48735 | n48881 ;
  assign n48883 = n81166 & n48882 ;
  assign n48884 = n48741 | n48883 ;
  assign n48885 = n81169 & n48884 ;
  assign n48886 = n48745 | n48885 ;
  assign n48887 = n81170 & n48886 ;
  assign n48888 = n48751 | n48887 ;
  assign n48889 = n81173 & n48888 ;
  assign n48890 = n48755 | n48889 ;
  assign n48891 = n81174 & n48890 ;
  assign n48892 = n48761 | n48891 ;
  assign n48893 = n81177 & n48892 ;
  assign n48894 = n48765 | n48893 ;
  assign n48895 = n81178 & n48894 ;
  assign n48896 = n48771 | n48895 ;
  assign n48897 = n81181 & n48896 ;
  assign n48898 = n48775 | n48897 ;
  assign n48899 = n81182 & n48898 ;
  assign n48900 = n48782 | n48899 ;
  assign n48901 = n81185 & n48900 ;
  assign n48902 = n48786 | n48901 ;
  assign n48903 = n81186 & n48902 ;
  assign n48904 = n48792 | n48903 ;
  assign n48907 = n48249 | n48796 ;
  assign n81198 = ~n48907 ;
  assign n48908 = n48904 & n81198 ;
  assign n48909 = n48906 | n48908 ;
  assign n81199 = ~n48817 ;
  assign n48910 = n81199 & n48909 ;
  assign n48911 = n48240 & n81195 ;
  assign n48912 = n48815 & n48911 ;
  assign n48913 = n48910 | n48912 ;
  assign n48914 = n48241 | n48812 ;
  assign n48915 = n48810 | n48914 ;
  assign n81200 = ~n48915 ;
  assign n48916 = n48798 & n81200 ;
  assign n48905 = n81189 & n48904 ;
  assign n48917 = n48796 | n48905 ;
  assign n48918 = n81190 & n48917 ;
  assign n48919 = n48810 | n48812 ;
  assign n81201 = ~n48918 ;
  assign n48920 = n81201 & n48919 ;
  assign n48921 = n48916 | n48920 ;
  assign n48922 = n81199 & n48921 ;
  assign n48923 = n15856 & n48809 ;
  assign n48924 = n48815 & n48923 ;
  assign n48925 = n48922 | n48924 ;
  assign n48926 = n70935 & n48925 ;
  assign n48927 = n70927 & n48913 ;
  assign n81202 = ~n48903 ;
  assign n48928 = n48792 & n81202 ;
  assign n48929 = n48257 | n48792 ;
  assign n81203 = ~n48929 ;
  assign n48930 = n48788 & n81203 ;
  assign n48931 = n48928 | n48930 ;
  assign n48932 = n81199 & n48931 ;
  assign n48933 = n48248 & n81195 ;
  assign n48934 = n48815 & n48933 ;
  assign n48935 = n48932 | n48934 ;
  assign n48936 = n70609 & n48935 ;
  assign n81204 = ~n48787 ;
  assign n48937 = n48786 & n81204 ;
  assign n48938 = n48265 | n48786 ;
  assign n81205 = ~n48938 ;
  assign n48939 = n48900 & n81205 ;
  assign n48940 = n48937 | n48939 ;
  assign n48941 = n81199 & n48940 ;
  assign n48942 = n48256 & n81195 ;
  assign n48943 = n48815 & n48942 ;
  assign n48944 = n48941 | n48943 ;
  assign n48945 = n70276 & n48944 ;
  assign n81206 = ~n48899 ;
  assign n48946 = n48782 & n81206 ;
  assign n48947 = n48273 | n48782 ;
  assign n81207 = ~n48947 ;
  assign n48948 = n48778 & n81207 ;
  assign n48949 = n48946 | n48948 ;
  assign n48950 = n81199 & n48949 ;
  assign n48951 = n48264 & n81195 ;
  assign n48952 = n48815 & n48951 ;
  assign n48953 = n48950 | n48952 ;
  assign n48954 = n70176 & n48953 ;
  assign n81208 = ~n48777 ;
  assign n48955 = n48775 & n81208 ;
  assign n48776 = n48281 | n48775 ;
  assign n81209 = ~n48776 ;
  assign n48956 = n48772 & n81209 ;
  assign n48957 = n48955 | n48956 ;
  assign n48958 = n81199 & n48957 ;
  assign n48959 = n48272 & n81195 ;
  assign n48960 = n48815 & n48959 ;
  assign n48961 = n48958 | n48960 ;
  assign n48962 = n69857 & n48961 ;
  assign n81210 = ~n48895 ;
  assign n48963 = n48771 & n81210 ;
  assign n48964 = n48289 | n48771 ;
  assign n81211 = ~n48964 ;
  assign n48965 = n48767 & n81211 ;
  assign n48966 = n48963 | n48965 ;
  assign n48967 = n81199 & n48966 ;
  assign n48968 = n48280 & n81195 ;
  assign n48969 = n48815 & n48968 ;
  assign n48970 = n48967 | n48969 ;
  assign n48971 = n69656 & n48970 ;
  assign n81212 = ~n48766 ;
  assign n48972 = n48765 & n81212 ;
  assign n48973 = n48297 | n48765 ;
  assign n81213 = ~n48973 ;
  assign n48974 = n48892 & n81213 ;
  assign n48975 = n48972 | n48974 ;
  assign n48976 = n81199 & n48975 ;
  assign n48977 = n48288 & n81195 ;
  assign n48978 = n48815 & n48977 ;
  assign n48979 = n48976 | n48978 ;
  assign n48980 = n69528 & n48979 ;
  assign n81214 = ~n48891 ;
  assign n48981 = n48761 & n81214 ;
  assign n48982 = n48305 | n48761 ;
  assign n81215 = ~n48982 ;
  assign n48983 = n48757 & n81215 ;
  assign n48984 = n48981 | n48983 ;
  assign n48985 = n81199 & n48984 ;
  assign n48986 = n48296 & n81195 ;
  assign n48987 = n48815 & n48986 ;
  assign n48988 = n48985 | n48987 ;
  assign n48989 = n69261 & n48988 ;
  assign n81216 = ~n48756 ;
  assign n48990 = n48755 & n81216 ;
  assign n48991 = n48313 | n48755 ;
  assign n81217 = ~n48991 ;
  assign n48992 = n48888 & n81217 ;
  assign n48993 = n48990 | n48992 ;
  assign n48994 = n81199 & n48993 ;
  assign n48995 = n48304 & n81195 ;
  assign n48996 = n48815 & n48995 ;
  assign n48997 = n48994 | n48996 ;
  assign n48998 = n69075 & n48997 ;
  assign n81218 = ~n48887 ;
  assign n48999 = n48751 & n81218 ;
  assign n49000 = n48321 | n48751 ;
  assign n81219 = ~n49000 ;
  assign n49001 = n48747 & n81219 ;
  assign n49002 = n48999 | n49001 ;
  assign n49003 = n81199 & n49002 ;
  assign n49004 = n48312 & n81195 ;
  assign n49005 = n48815 & n49004 ;
  assign n49006 = n49003 | n49005 ;
  assign n49007 = n68993 & n49006 ;
  assign n81220 = ~n48746 ;
  assign n49008 = n48745 & n81220 ;
  assign n49009 = n48329 | n48745 ;
  assign n81221 = ~n49009 ;
  assign n49010 = n48884 & n81221 ;
  assign n49011 = n49008 | n49010 ;
  assign n49012 = n81199 & n49011 ;
  assign n49013 = n48320 & n81195 ;
  assign n49014 = n48815 & n49013 ;
  assign n49015 = n49012 | n49014 ;
  assign n49016 = n68716 & n49015 ;
  assign n81222 = ~n48883 ;
  assign n49017 = n48741 & n81222 ;
  assign n49018 = n48337 | n48741 ;
  assign n81223 = ~n49018 ;
  assign n49019 = n48737 & n81223 ;
  assign n49020 = n49017 | n49019 ;
  assign n49021 = n81199 & n49020 ;
  assign n49022 = n48328 & n81195 ;
  assign n49023 = n48815 & n49022 ;
  assign n49024 = n49021 | n49023 ;
  assign n49025 = n68545 & n49024 ;
  assign n81224 = ~n48736 ;
  assign n49026 = n48735 & n81224 ;
  assign n49027 = n48345 | n48735 ;
  assign n81225 = ~n49027 ;
  assign n49028 = n48880 & n81225 ;
  assign n49029 = n49026 | n49028 ;
  assign n49030 = n81199 & n49029 ;
  assign n49031 = n48336 & n81195 ;
  assign n49032 = n48815 & n49031 ;
  assign n49033 = n49030 | n49032 ;
  assign n49034 = n68438 & n49033 ;
  assign n81226 = ~n48879 ;
  assign n49035 = n48730 & n81226 ;
  assign n48731 = n48353 | n48730 ;
  assign n81227 = ~n48731 ;
  assign n49036 = n81227 & n48878 ;
  assign n49037 = n49035 | n49036 ;
  assign n49038 = n81199 & n49037 ;
  assign n49039 = n48344 & n81195 ;
  assign n49040 = n48815 & n49039 ;
  assign n49041 = n49038 | n49040 ;
  assign n49042 = n68214 & n49041 ;
  assign n81228 = ~n48725 ;
  assign n49043 = n48724 & n81228 ;
  assign n49044 = n48361 | n48724 ;
  assign n81229 = ~n49044 ;
  assign n49045 = n48876 & n81229 ;
  assign n49046 = n49043 | n49045 ;
  assign n49047 = n81199 & n49046 ;
  assign n49048 = n48352 & n81195 ;
  assign n49049 = n48815 & n49048 ;
  assign n49050 = n49047 | n49049 ;
  assign n49051 = n68058 & n49050 ;
  assign n81230 = ~n48875 ;
  assign n49052 = n48720 & n81230 ;
  assign n49053 = n48369 | n48720 ;
  assign n81231 = ~n49053 ;
  assign n49054 = n48716 & n81231 ;
  assign n49055 = n49052 | n49054 ;
  assign n49056 = n81199 & n49055 ;
  assign n49057 = n48360 & n81195 ;
  assign n49058 = n48815 & n49057 ;
  assign n49059 = n49056 | n49058 ;
  assign n49060 = n67986 & n49059 ;
  assign n81232 = ~n48715 ;
  assign n49061 = n48714 & n81232 ;
  assign n49062 = n48377 | n48714 ;
  assign n81233 = ~n49062 ;
  assign n49063 = n48872 & n81233 ;
  assign n49064 = n49061 | n49063 ;
  assign n49065 = n81199 & n49064 ;
  assign n49066 = n48368 & n81195 ;
  assign n49067 = n48815 & n49066 ;
  assign n49068 = n49065 | n49067 ;
  assign n49069 = n67763 & n49068 ;
  assign n81234 = ~n48871 ;
  assign n49070 = n48710 & n81234 ;
  assign n49071 = n48385 | n48710 ;
  assign n81235 = ~n49071 ;
  assign n49072 = n48706 & n81235 ;
  assign n49073 = n49070 | n49072 ;
  assign n49074 = n81199 & n49073 ;
  assign n49075 = n48376 & n81195 ;
  assign n49076 = n48815 & n49075 ;
  assign n49077 = n49074 | n49076 ;
  assign n49078 = n67622 & n49077 ;
  assign n81236 = ~n48705 ;
  assign n49079 = n48704 & n81236 ;
  assign n49080 = n48393 | n48704 ;
  assign n81237 = ~n49080 ;
  assign n49081 = n48868 & n81237 ;
  assign n49082 = n49079 | n49081 ;
  assign n49083 = n81199 & n49082 ;
  assign n49084 = n48384 & n81195 ;
  assign n49085 = n48815 & n49084 ;
  assign n49086 = n49083 | n49085 ;
  assign n49087 = n67531 & n49086 ;
  assign n81238 = ~n48867 ;
  assign n49088 = n48700 & n81238 ;
  assign n49089 = n48401 | n48700 ;
  assign n81239 = ~n49089 ;
  assign n49090 = n48696 & n81239 ;
  assign n49091 = n49088 | n49090 ;
  assign n49092 = n81199 & n49091 ;
  assign n49093 = n48392 & n81195 ;
  assign n49094 = n48815 & n49093 ;
  assign n49095 = n49092 | n49094 ;
  assign n49096 = n67348 & n49095 ;
  assign n81240 = ~n48695 ;
  assign n49097 = n48694 & n81240 ;
  assign n49098 = n48409 | n48694 ;
  assign n81241 = ~n49098 ;
  assign n49099 = n48864 & n81241 ;
  assign n49100 = n49097 | n49099 ;
  assign n49101 = n81199 & n49100 ;
  assign n49102 = n48400 & n81195 ;
  assign n49103 = n48815 & n49102 ;
  assign n49104 = n49101 | n49103 ;
  assign n49105 = n67222 & n49104 ;
  assign n81242 = ~n48863 ;
  assign n49106 = n48690 & n81242 ;
  assign n49107 = n48417 | n48690 ;
  assign n81243 = ~n49107 ;
  assign n49108 = n48686 & n81243 ;
  assign n49109 = n49106 | n49108 ;
  assign n49110 = n81199 & n49109 ;
  assign n49111 = n48408 & n81195 ;
  assign n49112 = n48815 & n49111 ;
  assign n49113 = n49110 | n49112 ;
  assign n49114 = n67164 & n49113 ;
  assign n81244 = ~n48685 ;
  assign n49115 = n48684 & n81244 ;
  assign n49116 = n48425 | n48684 ;
  assign n81245 = ~n49116 ;
  assign n49117 = n48860 & n81245 ;
  assign n49118 = n49115 | n49117 ;
  assign n49119 = n81199 & n49118 ;
  assign n49120 = n48416 & n81195 ;
  assign n49121 = n48815 & n49120 ;
  assign n49122 = n49119 | n49121 ;
  assign n49123 = n66979 & n49122 ;
  assign n81246 = ~n48859 ;
  assign n49124 = n48680 & n81246 ;
  assign n49125 = n48433 | n48680 ;
  assign n81247 = ~n49125 ;
  assign n49126 = n48676 & n81247 ;
  assign n49127 = n49124 | n49126 ;
  assign n49128 = n81199 & n49127 ;
  assign n49129 = n48424 & n81195 ;
  assign n49130 = n48815 & n49129 ;
  assign n49131 = n49128 | n49130 ;
  assign n49132 = n66868 & n49131 ;
  assign n81248 = ~n48675 ;
  assign n49133 = n48674 & n81248 ;
  assign n49134 = n48441 | n48674 ;
  assign n81249 = ~n49134 ;
  assign n49135 = n48856 & n81249 ;
  assign n49136 = n49133 | n49135 ;
  assign n49137 = n81199 & n49136 ;
  assign n49138 = n48432 & n81195 ;
  assign n49139 = n48815 & n49138 ;
  assign n49140 = n49137 | n49139 ;
  assign n49141 = n66797 & n49140 ;
  assign n81250 = ~n48855 ;
  assign n49142 = n48670 & n81250 ;
  assign n49143 = n48449 | n48670 ;
  assign n81251 = ~n49143 ;
  assign n49144 = n48666 & n81251 ;
  assign n49145 = n49142 | n49144 ;
  assign n49146 = n81199 & n49145 ;
  assign n49147 = n48440 & n81195 ;
  assign n49148 = n48815 & n49147 ;
  assign n49149 = n49146 | n49148 ;
  assign n49150 = n66654 & n49149 ;
  assign n81252 = ~n48665 ;
  assign n49151 = n48664 & n81252 ;
  assign n49152 = n48457 | n48664 ;
  assign n81253 = ~n49152 ;
  assign n49153 = n48852 & n81253 ;
  assign n49154 = n49151 | n49153 ;
  assign n49155 = n81199 & n49154 ;
  assign n49156 = n48448 & n81195 ;
  assign n49157 = n48815 & n49156 ;
  assign n49158 = n49155 | n49157 ;
  assign n49159 = n66560 & n49158 ;
  assign n81254 = ~n48851 ;
  assign n49160 = n48660 & n81254 ;
  assign n49161 = n48465 | n48660 ;
  assign n81255 = ~n49161 ;
  assign n49162 = n48656 & n81255 ;
  assign n49163 = n49160 | n49162 ;
  assign n49164 = n81199 & n49163 ;
  assign n49165 = n48456 & n81195 ;
  assign n49166 = n48815 & n49165 ;
  assign n49167 = n49164 | n49166 ;
  assign n49168 = n66505 & n49167 ;
  assign n81256 = ~n48655 ;
  assign n49169 = n48654 & n81256 ;
  assign n49170 = n48473 | n48654 ;
  assign n81257 = ~n49170 ;
  assign n49171 = n48848 & n81257 ;
  assign n49172 = n49169 | n49171 ;
  assign n49173 = n81199 & n49172 ;
  assign n49174 = n48464 & n81195 ;
  assign n49175 = n48815 & n49174 ;
  assign n49176 = n49173 | n49175 ;
  assign n49177 = n66379 & n49176 ;
  assign n81258 = ~n48847 ;
  assign n49178 = n48650 & n81258 ;
  assign n49179 = n48481 | n48650 ;
  assign n81259 = ~n49179 ;
  assign n49180 = n48646 & n81259 ;
  assign n49181 = n49178 | n49180 ;
  assign n49182 = n81199 & n49181 ;
  assign n49183 = n48472 & n81195 ;
  assign n49184 = n48815 & n49183 ;
  assign n49185 = n49182 | n49184 ;
  assign n49186 = n66299 & n49185 ;
  assign n81260 = ~n48645 ;
  assign n49187 = n48643 & n81260 ;
  assign n48644 = n48489 | n48643 ;
  assign n81261 = ~n48644 ;
  assign n49188 = n48640 & n81261 ;
  assign n49189 = n49187 | n49188 ;
  assign n49190 = n81199 & n49189 ;
  assign n49191 = n48480 & n81195 ;
  assign n49192 = n48815 & n49191 ;
  assign n49193 = n49190 | n49192 ;
  assign n49194 = n66244 & n49193 ;
  assign n81262 = ~n48843 ;
  assign n49195 = n48639 & n81262 ;
  assign n49196 = n48497 | n48639 ;
  assign n81263 = ~n49196 ;
  assign n49197 = n48635 & n81263 ;
  assign n49198 = n49195 | n49197 ;
  assign n49199 = n81199 & n49198 ;
  assign n49200 = n48488 & n81195 ;
  assign n49201 = n48815 & n49200 ;
  assign n49202 = n49199 | n49201 ;
  assign n49203 = n66145 & n49202 ;
  assign n81264 = ~n48634 ;
  assign n49204 = n48633 & n81264 ;
  assign n49205 = n48505 | n48633 ;
  assign n81265 = ~n49205 ;
  assign n49206 = n48840 & n81265 ;
  assign n49207 = n49204 | n49206 ;
  assign n49208 = n81199 & n49207 ;
  assign n49209 = n48496 & n81195 ;
  assign n49210 = n48815 & n49209 ;
  assign n49211 = n49208 | n49210 ;
  assign n49212 = n66081 & n49211 ;
  assign n81266 = ~n48839 ;
  assign n49213 = n48629 & n81266 ;
  assign n49214 = n48513 | n48629 ;
  assign n81267 = ~n49214 ;
  assign n49215 = n48625 & n81267 ;
  assign n49216 = n49213 | n49215 ;
  assign n49217 = n81199 & n49216 ;
  assign n49218 = n48504 & n81195 ;
  assign n49219 = n48815 & n49218 ;
  assign n49220 = n49217 | n49219 ;
  assign n49221 = n66043 & n49220 ;
  assign n81268 = ~n48624 ;
  assign n49222 = n48622 & n81268 ;
  assign n48623 = n48521 | n48622 ;
  assign n81269 = ~n48623 ;
  assign n49223 = n48619 & n81269 ;
  assign n49224 = n49222 | n49223 ;
  assign n49225 = n81199 & n49224 ;
  assign n49226 = n48512 & n81195 ;
  assign n49227 = n48815 & n49226 ;
  assign n49228 = n49225 | n49227 ;
  assign n49229 = n65960 & n49228 ;
  assign n81270 = ~n48835 ;
  assign n49230 = n48618 & n81270 ;
  assign n49231 = n48529 | n48618 ;
  assign n81271 = ~n49231 ;
  assign n49232 = n48614 & n81271 ;
  assign n49233 = n49230 | n49232 ;
  assign n49234 = n81199 & n49233 ;
  assign n49235 = n48520 & n81195 ;
  assign n49236 = n48815 & n49235 ;
  assign n49237 = n49234 | n49236 ;
  assign n49238 = n65909 & n49237 ;
  assign n81272 = ~n48613 ;
  assign n49239 = n48611 & n81272 ;
  assign n48612 = n48537 | n48611 ;
  assign n81273 = ~n48612 ;
  assign n49240 = n48608 & n81273 ;
  assign n49241 = n49239 | n49240 ;
  assign n49242 = n81199 & n49241 ;
  assign n49243 = n48528 & n81195 ;
  assign n49244 = n48815 & n49243 ;
  assign n49245 = n49242 | n49244 ;
  assign n49246 = n65877 & n49245 ;
  assign n81274 = ~n48831 ;
  assign n49247 = n48607 & n81274 ;
  assign n49248 = n48546 | n48607 ;
  assign n81275 = ~n49248 ;
  assign n49249 = n48603 & n81275 ;
  assign n49250 = n49247 | n49249 ;
  assign n49251 = n81199 & n49250 ;
  assign n49252 = n48536 & n81195 ;
  assign n49253 = n48815 & n49252 ;
  assign n49254 = n49251 | n49253 ;
  assign n49255 = n65820 & n49254 ;
  assign n81276 = ~n48602 ;
  assign n49256 = n48601 & n81276 ;
  assign n49257 = n48554 | n48601 ;
  assign n81277 = ~n49257 ;
  assign n49258 = n48828 & n81277 ;
  assign n49259 = n49256 | n49258 ;
  assign n49260 = n81199 & n49259 ;
  assign n49261 = n48545 & n81195 ;
  assign n49262 = n48815 & n49261 ;
  assign n49263 = n49260 | n49262 ;
  assign n49264 = n65791 & n49263 ;
  assign n81278 = ~n48827 ;
  assign n49265 = n48597 & n81278 ;
  assign n49266 = n48562 | n48597 ;
  assign n81279 = ~n49266 ;
  assign n49267 = n48593 & n81279 ;
  assign n49268 = n49265 | n49267 ;
  assign n49269 = n81199 & n49268 ;
  assign n49270 = n48553 & n81195 ;
  assign n49271 = n48815 & n49270 ;
  assign n49272 = n49269 | n49271 ;
  assign n49273 = n65772 & n49272 ;
  assign n81280 = ~n48592 ;
  assign n49274 = n48591 & n81280 ;
  assign n49275 = n48570 | n48591 ;
  assign n81281 = ~n49275 ;
  assign n49276 = n48824 & n81281 ;
  assign n49277 = n49274 | n49276 ;
  assign n49278 = n81199 & n49277 ;
  assign n49279 = n48561 & n81195 ;
  assign n49280 = n48815 & n49279 ;
  assign n49281 = n49278 | n49280 ;
  assign n49282 = n65746 & n49281 ;
  assign n81282 = ~n48823 ;
  assign n49283 = n48587 & n81282 ;
  assign n48822 = n48583 | n48587 ;
  assign n81283 = ~n48822 ;
  assign n49284 = n48821 & n81283 ;
  assign n49285 = n49283 | n49284 ;
  assign n49286 = n81199 & n49285 ;
  assign n49287 = n48569 & n81195 ;
  assign n49288 = n48815 & n49287 ;
  assign n49289 = n49286 | n49288 ;
  assign n49290 = n65721 & n49289 ;
  assign n49291 = n16327 & n48579 ;
  assign n49292 = n81197 & n49291 ;
  assign n81284 = ~n49292 ;
  assign n49293 = n48821 & n81284 ;
  assign n49294 = n81199 & n49293 ;
  assign n49295 = n48582 & n81195 ;
  assign n49296 = n48815 & n49295 ;
  assign n49297 = n49294 | n49296 ;
  assign n49298 = n65686 & n49297 ;
  assign n48818 = n16327 & n81199 ;
  assign n49303 = x64 & n81199 ;
  assign n81285 = ~n49303 ;
  assign n49304 = x19 & n81285 ;
  assign n49305 = n48818 | n49304 ;
  assign n49307 = x65 & n49305 ;
  assign n49299 = n48814 | n48918 ;
  assign n49300 = n81195 & n49299 ;
  assign n81286 = ~n49300 ;
  assign n49301 = x64 & n81286 ;
  assign n81287 = ~n49301 ;
  assign n49302 = x19 & n81287 ;
  assign n49306 = x65 | n48818 ;
  assign n49308 = n49302 | n49306 ;
  assign n81288 = ~n49307 ;
  assign n49309 = n81288 & n49308 ;
  assign n49310 = n17058 | n49309 ;
  assign n49311 = n65670 & n49305 ;
  assign n81289 = ~n49311 ;
  assign n49312 = n49310 & n81289 ;
  assign n81290 = ~n49296 ;
  assign n49313 = x66 & n81290 ;
  assign n81291 = ~n49294 ;
  assign n49314 = n81291 & n49313 ;
  assign n49315 = n49298 | n49314 ;
  assign n49316 = n49312 | n49315 ;
  assign n81292 = ~n49298 ;
  assign n49317 = n81292 & n49316 ;
  assign n81293 = ~n49288 ;
  assign n49318 = x67 & n81293 ;
  assign n81294 = ~n49286 ;
  assign n49319 = n81294 & n49318 ;
  assign n49320 = n49317 | n49319 ;
  assign n81295 = ~n49290 ;
  assign n49321 = n81295 & n49320 ;
  assign n81296 = ~n49280 ;
  assign n49322 = x68 & n81296 ;
  assign n81297 = ~n49278 ;
  assign n49323 = n81297 & n49322 ;
  assign n49324 = n49282 | n49323 ;
  assign n49325 = n49321 | n49324 ;
  assign n81298 = ~n49282 ;
  assign n49326 = n81298 & n49325 ;
  assign n81299 = ~n49271 ;
  assign n49327 = x69 & n81299 ;
  assign n81300 = ~n49269 ;
  assign n49328 = n81300 & n49327 ;
  assign n49329 = n49326 | n49328 ;
  assign n81301 = ~n49273 ;
  assign n49330 = n81301 & n49329 ;
  assign n81302 = ~n49262 ;
  assign n49331 = x70 & n81302 ;
  assign n81303 = ~n49260 ;
  assign n49332 = n81303 & n49331 ;
  assign n49333 = n49264 | n49332 ;
  assign n49334 = n49330 | n49333 ;
  assign n81304 = ~n49264 ;
  assign n49335 = n81304 & n49334 ;
  assign n81305 = ~n49253 ;
  assign n49336 = x71 & n81305 ;
  assign n81306 = ~n49251 ;
  assign n49337 = n81306 & n49336 ;
  assign n49338 = n49255 | n49337 ;
  assign n49340 = n49335 | n49338 ;
  assign n81307 = ~n49255 ;
  assign n49341 = n81307 & n49340 ;
  assign n81308 = ~n49244 ;
  assign n49342 = x72 & n81308 ;
  assign n81309 = ~n49242 ;
  assign n49343 = n81309 & n49342 ;
  assign n49344 = n49246 | n49343 ;
  assign n49345 = n49341 | n49344 ;
  assign n81310 = ~n49246 ;
  assign n49346 = n81310 & n49345 ;
  assign n81311 = ~n49236 ;
  assign n49347 = x73 & n81311 ;
  assign n81312 = ~n49234 ;
  assign n49348 = n81312 & n49347 ;
  assign n49349 = n49238 | n49348 ;
  assign n49351 = n49346 | n49349 ;
  assign n81313 = ~n49238 ;
  assign n49352 = n81313 & n49351 ;
  assign n81314 = ~n49227 ;
  assign n49353 = x74 & n81314 ;
  assign n81315 = ~n49225 ;
  assign n49354 = n81315 & n49353 ;
  assign n49355 = n49229 | n49354 ;
  assign n49356 = n49352 | n49355 ;
  assign n81316 = ~n49229 ;
  assign n49357 = n81316 & n49356 ;
  assign n81317 = ~n49219 ;
  assign n49358 = x75 & n81317 ;
  assign n81318 = ~n49217 ;
  assign n49359 = n81318 & n49358 ;
  assign n49360 = n49221 | n49359 ;
  assign n49362 = n49357 | n49360 ;
  assign n81319 = ~n49221 ;
  assign n49363 = n81319 & n49362 ;
  assign n81320 = ~n49210 ;
  assign n49364 = x76 & n81320 ;
  assign n81321 = ~n49208 ;
  assign n49365 = n81321 & n49364 ;
  assign n49366 = n49212 | n49365 ;
  assign n49367 = n49363 | n49366 ;
  assign n81322 = ~n49212 ;
  assign n49368 = n81322 & n49367 ;
  assign n81323 = ~n49201 ;
  assign n49369 = x77 & n81323 ;
  assign n81324 = ~n49199 ;
  assign n49370 = n81324 & n49369 ;
  assign n49371 = n49203 | n49370 ;
  assign n49373 = n49368 | n49371 ;
  assign n81325 = ~n49203 ;
  assign n49374 = n81325 & n49373 ;
  assign n81326 = ~n49192 ;
  assign n49375 = x78 & n81326 ;
  assign n81327 = ~n49190 ;
  assign n49376 = n81327 & n49375 ;
  assign n49377 = n49194 | n49376 ;
  assign n49378 = n49374 | n49377 ;
  assign n81328 = ~n49194 ;
  assign n49379 = n81328 & n49378 ;
  assign n81329 = ~n49184 ;
  assign n49380 = x79 & n81329 ;
  assign n81330 = ~n49182 ;
  assign n49381 = n81330 & n49380 ;
  assign n49382 = n49186 | n49381 ;
  assign n49384 = n49379 | n49382 ;
  assign n81331 = ~n49186 ;
  assign n49385 = n81331 & n49384 ;
  assign n81332 = ~n49175 ;
  assign n49386 = x80 & n81332 ;
  assign n81333 = ~n49173 ;
  assign n49387 = n81333 & n49386 ;
  assign n49388 = n49177 | n49387 ;
  assign n49389 = n49385 | n49388 ;
  assign n81334 = ~n49177 ;
  assign n49390 = n81334 & n49389 ;
  assign n81335 = ~n49166 ;
  assign n49391 = x81 & n81335 ;
  assign n81336 = ~n49164 ;
  assign n49392 = n81336 & n49391 ;
  assign n49393 = n49168 | n49392 ;
  assign n49395 = n49390 | n49393 ;
  assign n81337 = ~n49168 ;
  assign n49396 = n81337 & n49395 ;
  assign n81338 = ~n49157 ;
  assign n49397 = x82 & n81338 ;
  assign n81339 = ~n49155 ;
  assign n49398 = n81339 & n49397 ;
  assign n49399 = n49159 | n49398 ;
  assign n49400 = n49396 | n49399 ;
  assign n81340 = ~n49159 ;
  assign n49401 = n81340 & n49400 ;
  assign n81341 = ~n49148 ;
  assign n49402 = x83 & n81341 ;
  assign n81342 = ~n49146 ;
  assign n49403 = n81342 & n49402 ;
  assign n49404 = n49150 | n49403 ;
  assign n49406 = n49401 | n49404 ;
  assign n81343 = ~n49150 ;
  assign n49407 = n81343 & n49406 ;
  assign n81344 = ~n49139 ;
  assign n49408 = x84 & n81344 ;
  assign n81345 = ~n49137 ;
  assign n49409 = n81345 & n49408 ;
  assign n49410 = n49141 | n49409 ;
  assign n49411 = n49407 | n49410 ;
  assign n81346 = ~n49141 ;
  assign n49412 = n81346 & n49411 ;
  assign n81347 = ~n49130 ;
  assign n49413 = x85 & n81347 ;
  assign n81348 = ~n49128 ;
  assign n49414 = n81348 & n49413 ;
  assign n49415 = n49132 | n49414 ;
  assign n49417 = n49412 | n49415 ;
  assign n81349 = ~n49132 ;
  assign n49418 = n81349 & n49417 ;
  assign n81350 = ~n49121 ;
  assign n49419 = x86 & n81350 ;
  assign n81351 = ~n49119 ;
  assign n49420 = n81351 & n49419 ;
  assign n49421 = n49123 | n49420 ;
  assign n49422 = n49418 | n49421 ;
  assign n81352 = ~n49123 ;
  assign n49423 = n81352 & n49422 ;
  assign n81353 = ~n49112 ;
  assign n49424 = x87 & n81353 ;
  assign n81354 = ~n49110 ;
  assign n49425 = n81354 & n49424 ;
  assign n49426 = n49114 | n49425 ;
  assign n49428 = n49423 | n49426 ;
  assign n81355 = ~n49114 ;
  assign n49429 = n81355 & n49428 ;
  assign n81356 = ~n49103 ;
  assign n49430 = x88 & n81356 ;
  assign n81357 = ~n49101 ;
  assign n49431 = n81357 & n49430 ;
  assign n49432 = n49105 | n49431 ;
  assign n49433 = n49429 | n49432 ;
  assign n81358 = ~n49105 ;
  assign n49434 = n81358 & n49433 ;
  assign n81359 = ~n49094 ;
  assign n49435 = x89 & n81359 ;
  assign n81360 = ~n49092 ;
  assign n49436 = n81360 & n49435 ;
  assign n49437 = n49096 | n49436 ;
  assign n49439 = n49434 | n49437 ;
  assign n81361 = ~n49096 ;
  assign n49440 = n81361 & n49439 ;
  assign n81362 = ~n49085 ;
  assign n49441 = x90 & n81362 ;
  assign n81363 = ~n49083 ;
  assign n49442 = n81363 & n49441 ;
  assign n49443 = n49087 | n49442 ;
  assign n49444 = n49440 | n49443 ;
  assign n81364 = ~n49087 ;
  assign n49445 = n81364 & n49444 ;
  assign n81365 = ~n49076 ;
  assign n49446 = x91 & n81365 ;
  assign n81366 = ~n49074 ;
  assign n49447 = n81366 & n49446 ;
  assign n49448 = n49078 | n49447 ;
  assign n49450 = n49445 | n49448 ;
  assign n81367 = ~n49078 ;
  assign n49451 = n81367 & n49450 ;
  assign n81368 = ~n49067 ;
  assign n49452 = x92 & n81368 ;
  assign n81369 = ~n49065 ;
  assign n49453 = n81369 & n49452 ;
  assign n49454 = n49069 | n49453 ;
  assign n49455 = n49451 | n49454 ;
  assign n81370 = ~n49069 ;
  assign n49456 = n81370 & n49455 ;
  assign n81371 = ~n49058 ;
  assign n49457 = x93 & n81371 ;
  assign n81372 = ~n49056 ;
  assign n49458 = n81372 & n49457 ;
  assign n49459 = n49060 | n49458 ;
  assign n49461 = n49456 | n49459 ;
  assign n81373 = ~n49060 ;
  assign n49462 = n81373 & n49461 ;
  assign n81374 = ~n49049 ;
  assign n49463 = x94 & n81374 ;
  assign n81375 = ~n49047 ;
  assign n49464 = n81375 & n49463 ;
  assign n49465 = n49051 | n49464 ;
  assign n49466 = n49462 | n49465 ;
  assign n81376 = ~n49051 ;
  assign n49467 = n81376 & n49466 ;
  assign n81377 = ~n49040 ;
  assign n49468 = x95 & n81377 ;
  assign n81378 = ~n49038 ;
  assign n49469 = n81378 & n49468 ;
  assign n49470 = n49042 | n49469 ;
  assign n49472 = n49467 | n49470 ;
  assign n81379 = ~n49042 ;
  assign n49473 = n81379 & n49472 ;
  assign n81380 = ~n49032 ;
  assign n49474 = x96 & n81380 ;
  assign n81381 = ~n49030 ;
  assign n49475 = n81381 & n49474 ;
  assign n49476 = n49034 | n49475 ;
  assign n49477 = n49473 | n49476 ;
  assign n81382 = ~n49034 ;
  assign n49478 = n81382 & n49477 ;
  assign n81383 = ~n49023 ;
  assign n49479 = x97 & n81383 ;
  assign n81384 = ~n49021 ;
  assign n49480 = n81384 & n49479 ;
  assign n49481 = n49025 | n49480 ;
  assign n49483 = n49478 | n49481 ;
  assign n81385 = ~n49025 ;
  assign n49484 = n81385 & n49483 ;
  assign n81386 = ~n49014 ;
  assign n49485 = x98 & n81386 ;
  assign n81387 = ~n49012 ;
  assign n49486 = n81387 & n49485 ;
  assign n49487 = n49016 | n49486 ;
  assign n49488 = n49484 | n49487 ;
  assign n81388 = ~n49016 ;
  assign n49489 = n81388 & n49488 ;
  assign n81389 = ~n49005 ;
  assign n49490 = x99 & n81389 ;
  assign n81390 = ~n49003 ;
  assign n49491 = n81390 & n49490 ;
  assign n49492 = n49007 | n49491 ;
  assign n49494 = n49489 | n49492 ;
  assign n81391 = ~n49007 ;
  assign n49495 = n81391 & n49494 ;
  assign n81392 = ~n48996 ;
  assign n49496 = x100 & n81392 ;
  assign n81393 = ~n48994 ;
  assign n49497 = n81393 & n49496 ;
  assign n49498 = n48998 | n49497 ;
  assign n49499 = n49495 | n49498 ;
  assign n81394 = ~n48998 ;
  assign n49500 = n81394 & n49499 ;
  assign n81395 = ~n48987 ;
  assign n49501 = x101 & n81395 ;
  assign n81396 = ~n48985 ;
  assign n49502 = n81396 & n49501 ;
  assign n49503 = n48989 | n49502 ;
  assign n49505 = n49500 | n49503 ;
  assign n81397 = ~n48989 ;
  assign n49506 = n81397 & n49505 ;
  assign n81398 = ~n48978 ;
  assign n49507 = x102 & n81398 ;
  assign n81399 = ~n48976 ;
  assign n49508 = n81399 & n49507 ;
  assign n49509 = n48980 | n49508 ;
  assign n49510 = n49506 | n49509 ;
  assign n81400 = ~n48980 ;
  assign n49511 = n81400 & n49510 ;
  assign n81401 = ~n48969 ;
  assign n49512 = x103 & n81401 ;
  assign n81402 = ~n48967 ;
  assign n49513 = n81402 & n49512 ;
  assign n49514 = n48971 | n49513 ;
  assign n49516 = n49511 | n49514 ;
  assign n81403 = ~n48971 ;
  assign n49517 = n81403 & n49516 ;
  assign n81404 = ~n48960 ;
  assign n49518 = x104 & n81404 ;
  assign n81405 = ~n48958 ;
  assign n49519 = n81405 & n49518 ;
  assign n49520 = n48962 | n49519 ;
  assign n49521 = n49517 | n49520 ;
  assign n81406 = ~n48962 ;
  assign n49522 = n81406 & n49521 ;
  assign n81407 = ~n48952 ;
  assign n49523 = x105 & n81407 ;
  assign n81408 = ~n48950 ;
  assign n49524 = n81408 & n49523 ;
  assign n49525 = n48954 | n49524 ;
  assign n49527 = n49522 | n49525 ;
  assign n81409 = ~n48954 ;
  assign n49528 = n81409 & n49527 ;
  assign n81410 = ~n48943 ;
  assign n49529 = x106 & n81410 ;
  assign n81411 = ~n48941 ;
  assign n49530 = n81411 & n49529 ;
  assign n49531 = n48945 | n49530 ;
  assign n49532 = n49528 | n49531 ;
  assign n81412 = ~n48945 ;
  assign n49533 = n81412 & n49532 ;
  assign n81413 = ~n48934 ;
  assign n49534 = x107 & n81413 ;
  assign n81414 = ~n48932 ;
  assign n49535 = n81414 & n49534 ;
  assign n49536 = n48936 | n49535 ;
  assign n49538 = n49533 | n49536 ;
  assign n81415 = ~n48936 ;
  assign n49539 = n81415 & n49538 ;
  assign n81416 = ~n48912 ;
  assign n49540 = x108 & n81416 ;
  assign n81417 = ~n48910 ;
  assign n49541 = n81417 & n49540 ;
  assign n49542 = n48927 | n49541 ;
  assign n49543 = n49539 | n49542 ;
  assign n81418 = ~n48927 ;
  assign n49544 = n81418 & n49543 ;
  assign n81419 = ~n48924 ;
  assign n49545 = x109 & n81419 ;
  assign n81420 = ~n48922 ;
  assign n49546 = n81420 & n49545 ;
  assign n49547 = n48926 | n49546 ;
  assign n49549 = n49544 | n49547 ;
  assign n81421 = ~n48926 ;
  assign n49550 = n81421 & n49549 ;
  assign n49551 = n17324 | n49550 ;
  assign n49552 = n48913 & n49551 ;
  assign n49553 = n48818 | n49302 ;
  assign n49554 = x65 & n49553 ;
  assign n81422 = ~n49554 ;
  assign n49555 = n49308 & n81422 ;
  assign n49556 = n17058 | n49555 ;
  assign n49557 = n81289 & n49556 ;
  assign n49558 = n49315 | n49557 ;
  assign n49559 = n81292 & n49558 ;
  assign n49560 = n49290 | n49319 ;
  assign n49562 = n49559 | n49560 ;
  assign n49563 = n81295 & n49562 ;
  assign n49564 = n49323 | n49563 ;
  assign n49566 = n81298 & n49564 ;
  assign n49567 = n49273 | n49328 ;
  assign n49569 = n49566 | n49567 ;
  assign n49570 = n81301 & n49569 ;
  assign n49571 = n49332 | n49570 ;
  assign n49573 = n81304 & n49571 ;
  assign n49574 = n49338 | n49573 ;
  assign n49575 = n81307 & n49574 ;
  assign n49576 = n49344 | n49575 ;
  assign n49578 = n81310 & n49576 ;
  assign n49579 = n49349 | n49578 ;
  assign n49580 = n81313 & n49579 ;
  assign n49581 = n49355 | n49580 ;
  assign n49583 = n81316 & n49581 ;
  assign n49584 = n49360 | n49583 ;
  assign n49585 = n81319 & n49584 ;
  assign n49586 = n49366 | n49585 ;
  assign n49588 = n81322 & n49586 ;
  assign n49589 = n49371 | n49588 ;
  assign n49590 = n81325 & n49589 ;
  assign n49591 = n49377 | n49590 ;
  assign n49593 = n81328 & n49591 ;
  assign n49594 = n49382 | n49593 ;
  assign n49595 = n81331 & n49594 ;
  assign n49596 = n49388 | n49595 ;
  assign n49598 = n81334 & n49596 ;
  assign n49599 = n49393 | n49598 ;
  assign n49600 = n81337 & n49599 ;
  assign n49601 = n49399 | n49600 ;
  assign n49603 = n81340 & n49601 ;
  assign n49604 = n49404 | n49603 ;
  assign n49605 = n81343 & n49604 ;
  assign n49606 = n49410 | n49605 ;
  assign n49608 = n81346 & n49606 ;
  assign n49609 = n49415 | n49608 ;
  assign n49610 = n81349 & n49609 ;
  assign n49611 = n49421 | n49610 ;
  assign n49613 = n81352 & n49611 ;
  assign n49614 = n49426 | n49613 ;
  assign n49615 = n81355 & n49614 ;
  assign n49616 = n49432 | n49615 ;
  assign n49618 = n81358 & n49616 ;
  assign n49619 = n49437 | n49618 ;
  assign n49620 = n81361 & n49619 ;
  assign n49621 = n49443 | n49620 ;
  assign n49623 = n81364 & n49621 ;
  assign n49624 = n49448 | n49623 ;
  assign n49625 = n81367 & n49624 ;
  assign n49626 = n49454 | n49625 ;
  assign n49628 = n81370 & n49626 ;
  assign n49629 = n49459 | n49628 ;
  assign n49630 = n81373 & n49629 ;
  assign n49631 = n49465 | n49630 ;
  assign n49633 = n81376 & n49631 ;
  assign n49634 = n49470 | n49633 ;
  assign n49635 = n81379 & n49634 ;
  assign n49636 = n49476 | n49635 ;
  assign n49638 = n81382 & n49636 ;
  assign n49639 = n49481 | n49638 ;
  assign n49640 = n81385 & n49639 ;
  assign n49641 = n49487 | n49640 ;
  assign n49643 = n81388 & n49641 ;
  assign n49644 = n49492 | n49643 ;
  assign n49645 = n81391 & n49644 ;
  assign n49646 = n49498 | n49645 ;
  assign n49648 = n81394 & n49646 ;
  assign n49649 = n49503 | n49648 ;
  assign n49650 = n81397 & n49649 ;
  assign n49651 = n49509 | n49650 ;
  assign n49653 = n81400 & n49651 ;
  assign n49654 = n49514 | n49653 ;
  assign n49655 = n81403 & n49654 ;
  assign n49656 = n49520 | n49655 ;
  assign n49658 = n81406 & n49656 ;
  assign n49659 = n49525 | n49658 ;
  assign n49660 = n81409 & n49659 ;
  assign n49661 = n49531 | n49660 ;
  assign n49663 = n81412 & n49661 ;
  assign n49664 = n49536 | n49663 ;
  assign n49665 = n81415 & n49664 ;
  assign n81423 = ~n49665 ;
  assign n49666 = n49542 & n81423 ;
  assign n49668 = n48936 | n49542 ;
  assign n81424 = ~n49668 ;
  assign n49669 = n49538 & n81424 ;
  assign n49670 = n49666 | n49669 ;
  assign n49671 = n71164 & n49670 ;
  assign n81425 = ~n49550 ;
  assign n49672 = n81425 & n49671 ;
  assign n49673 = n49552 | n49672 ;
  assign n49674 = n70935 & n49673 ;
  assign n81426 = ~n49672 ;
  assign n50259 = x109 & n81426 ;
  assign n81427 = ~n49552 ;
  assign n50260 = n81427 & n50259 ;
  assign n50261 = n49674 | n50260 ;
  assign n49675 = n48935 & n49551 ;
  assign n81428 = ~n49533 ;
  assign n49537 = n81428 & n49536 ;
  assign n49676 = n48945 | n49536 ;
  assign n81429 = ~n49676 ;
  assign n49677 = n49661 & n81429 ;
  assign n49678 = n49537 | n49677 ;
  assign n49679 = n71164 & n49678 ;
  assign n49680 = n81425 & n49679 ;
  assign n49681 = n49675 | n49680 ;
  assign n49682 = n70927 & n49681 ;
  assign n49683 = n48944 & n49551 ;
  assign n81430 = ~n49660 ;
  assign n49662 = n49531 & n81430 ;
  assign n49684 = n48954 | n49531 ;
  assign n81431 = ~n49684 ;
  assign n49685 = n49527 & n81431 ;
  assign n49686 = n49662 | n49685 ;
  assign n49687 = n71164 & n49686 ;
  assign n49688 = n81425 & n49687 ;
  assign n49689 = n49683 | n49688 ;
  assign n49690 = n70609 & n49689 ;
  assign n81432 = ~n49688 ;
  assign n50249 = x107 & n81432 ;
  assign n81433 = ~n49683 ;
  assign n50250 = n81433 & n50249 ;
  assign n50251 = n49690 | n50250 ;
  assign n49691 = n48953 & n49551 ;
  assign n81434 = ~n49522 ;
  assign n49526 = n81434 & n49525 ;
  assign n49692 = n48962 | n49525 ;
  assign n81435 = ~n49692 ;
  assign n49693 = n49656 & n81435 ;
  assign n49694 = n49526 | n49693 ;
  assign n49695 = n71164 & n49694 ;
  assign n49696 = n81425 & n49695 ;
  assign n49697 = n49691 | n49696 ;
  assign n49698 = n70276 & n49697 ;
  assign n49699 = n48961 & n49551 ;
  assign n81436 = ~n49655 ;
  assign n49657 = n49520 & n81436 ;
  assign n49700 = n48971 | n49520 ;
  assign n81437 = ~n49700 ;
  assign n49701 = n49516 & n81437 ;
  assign n49702 = n49657 | n49701 ;
  assign n49703 = n71164 & n49702 ;
  assign n49704 = n81425 & n49703 ;
  assign n49705 = n49699 | n49704 ;
  assign n49706 = n70176 & n49705 ;
  assign n81438 = ~n49704 ;
  assign n50239 = x105 & n81438 ;
  assign n81439 = ~n49699 ;
  assign n50240 = n81439 & n50239 ;
  assign n50241 = n49706 | n50240 ;
  assign n49707 = n48970 & n49551 ;
  assign n81440 = ~n49511 ;
  assign n49515 = n81440 & n49514 ;
  assign n49708 = n48980 | n49514 ;
  assign n81441 = ~n49708 ;
  assign n49709 = n49651 & n81441 ;
  assign n49710 = n49515 | n49709 ;
  assign n49711 = n71164 & n49710 ;
  assign n49712 = n81425 & n49711 ;
  assign n49713 = n49707 | n49712 ;
  assign n49714 = n69857 & n49713 ;
  assign n49715 = n48979 & n49551 ;
  assign n81442 = ~n49650 ;
  assign n49652 = n49509 & n81442 ;
  assign n49716 = n48989 | n49509 ;
  assign n81443 = ~n49716 ;
  assign n49717 = n49505 & n81443 ;
  assign n49718 = n49652 | n49717 ;
  assign n49719 = n71164 & n49718 ;
  assign n49720 = n81425 & n49719 ;
  assign n49721 = n49715 | n49720 ;
  assign n49722 = n69656 & n49721 ;
  assign n81444 = ~n49720 ;
  assign n50229 = x103 & n81444 ;
  assign n81445 = ~n49715 ;
  assign n50230 = n81445 & n50229 ;
  assign n50231 = n49722 | n50230 ;
  assign n49723 = n48988 & n49551 ;
  assign n81446 = ~n49500 ;
  assign n49504 = n81446 & n49503 ;
  assign n49724 = n48998 | n49503 ;
  assign n81447 = ~n49724 ;
  assign n49725 = n49646 & n81447 ;
  assign n49726 = n49504 | n49725 ;
  assign n49727 = n71164 & n49726 ;
  assign n49728 = n81425 & n49727 ;
  assign n49729 = n49723 | n49728 ;
  assign n49730 = n69528 & n49729 ;
  assign n49731 = n48997 & n49551 ;
  assign n81448 = ~n49645 ;
  assign n49647 = n49498 & n81448 ;
  assign n49732 = n49007 | n49498 ;
  assign n81449 = ~n49732 ;
  assign n49733 = n49494 & n81449 ;
  assign n49734 = n49647 | n49733 ;
  assign n49735 = n71164 & n49734 ;
  assign n49736 = n81425 & n49735 ;
  assign n49737 = n49731 | n49736 ;
  assign n49738 = n69261 & n49737 ;
  assign n81450 = ~n49736 ;
  assign n50219 = x101 & n81450 ;
  assign n81451 = ~n49731 ;
  assign n50220 = n81451 & n50219 ;
  assign n50221 = n49738 | n50220 ;
  assign n49739 = n49006 & n49551 ;
  assign n81452 = ~n49489 ;
  assign n49493 = n81452 & n49492 ;
  assign n49740 = n49016 | n49492 ;
  assign n81453 = ~n49740 ;
  assign n49741 = n49641 & n81453 ;
  assign n49742 = n49493 | n49741 ;
  assign n49743 = n71164 & n49742 ;
  assign n49744 = n81425 & n49743 ;
  assign n49745 = n49739 | n49744 ;
  assign n49746 = n69075 & n49745 ;
  assign n49747 = n49015 & n49551 ;
  assign n81454 = ~n49640 ;
  assign n49642 = n49487 & n81454 ;
  assign n49748 = n49025 | n49487 ;
  assign n81455 = ~n49748 ;
  assign n49749 = n49483 & n81455 ;
  assign n49750 = n49642 | n49749 ;
  assign n49751 = n71164 & n49750 ;
  assign n49752 = n81425 & n49751 ;
  assign n49753 = n49747 | n49752 ;
  assign n49754 = n68993 & n49753 ;
  assign n81456 = ~n49752 ;
  assign n50208 = x99 & n81456 ;
  assign n81457 = ~n49747 ;
  assign n50209 = n81457 & n50208 ;
  assign n50210 = n49754 | n50209 ;
  assign n49755 = n49024 & n49551 ;
  assign n81458 = ~n49478 ;
  assign n49482 = n81458 & n49481 ;
  assign n49756 = n49034 | n49481 ;
  assign n81459 = ~n49756 ;
  assign n49757 = n49636 & n81459 ;
  assign n49758 = n49482 | n49757 ;
  assign n49759 = n71164 & n49758 ;
  assign n49760 = n81425 & n49759 ;
  assign n49761 = n49755 | n49760 ;
  assign n49762 = n68716 & n49761 ;
  assign n49763 = n49033 & n49551 ;
  assign n81460 = ~n49635 ;
  assign n49637 = n49476 & n81460 ;
  assign n49764 = n49042 | n49476 ;
  assign n81461 = ~n49764 ;
  assign n49765 = n49472 & n81461 ;
  assign n49766 = n49637 | n49765 ;
  assign n49767 = n71164 & n49766 ;
  assign n49768 = n81425 & n49767 ;
  assign n49769 = n49763 | n49768 ;
  assign n49770 = n68545 & n49769 ;
  assign n81462 = ~n49768 ;
  assign n50198 = x97 & n81462 ;
  assign n81463 = ~n49763 ;
  assign n50199 = n81463 & n50198 ;
  assign n50200 = n49770 | n50199 ;
  assign n49771 = n49041 & n49551 ;
  assign n81464 = ~n49467 ;
  assign n49471 = n81464 & n49470 ;
  assign n49772 = n49051 | n49470 ;
  assign n81465 = ~n49772 ;
  assign n49773 = n49631 & n81465 ;
  assign n49774 = n49471 | n49773 ;
  assign n49775 = n71164 & n49774 ;
  assign n49776 = n81425 & n49775 ;
  assign n49777 = n49771 | n49776 ;
  assign n49778 = n68438 & n49777 ;
  assign n49779 = n49050 & n49551 ;
  assign n81466 = ~n49630 ;
  assign n49632 = n49465 & n81466 ;
  assign n49780 = n49060 | n49465 ;
  assign n81467 = ~n49780 ;
  assign n49781 = n49461 & n81467 ;
  assign n49782 = n49632 | n49781 ;
  assign n49783 = n71164 & n49782 ;
  assign n49784 = n81425 & n49783 ;
  assign n49785 = n49779 | n49784 ;
  assign n49786 = n68214 & n49785 ;
  assign n81468 = ~n49784 ;
  assign n50188 = x95 & n81468 ;
  assign n81469 = ~n49779 ;
  assign n50189 = n81469 & n50188 ;
  assign n50190 = n49786 | n50189 ;
  assign n49787 = n49059 & n49551 ;
  assign n81470 = ~n49456 ;
  assign n49460 = n81470 & n49459 ;
  assign n49788 = n49069 | n49459 ;
  assign n81471 = ~n49788 ;
  assign n49789 = n49626 & n81471 ;
  assign n49790 = n49460 | n49789 ;
  assign n49791 = n71164 & n49790 ;
  assign n49792 = n81425 & n49791 ;
  assign n49793 = n49787 | n49792 ;
  assign n49794 = n68058 & n49793 ;
  assign n49795 = n49068 & n49551 ;
  assign n81472 = ~n49625 ;
  assign n49627 = n49454 & n81472 ;
  assign n49796 = n49078 | n49454 ;
  assign n81473 = ~n49796 ;
  assign n49797 = n49450 & n81473 ;
  assign n49798 = n49627 | n49797 ;
  assign n49799 = n71164 & n49798 ;
  assign n49800 = n81425 & n49799 ;
  assign n49801 = n49795 | n49800 ;
  assign n49802 = n67986 & n49801 ;
  assign n81474 = ~n49800 ;
  assign n50178 = x93 & n81474 ;
  assign n81475 = ~n49795 ;
  assign n50179 = n81475 & n50178 ;
  assign n50180 = n49802 | n50179 ;
  assign n49803 = n49077 & n49551 ;
  assign n81476 = ~n49445 ;
  assign n49449 = n81476 & n49448 ;
  assign n49804 = n49087 | n49448 ;
  assign n81477 = ~n49804 ;
  assign n49805 = n49621 & n81477 ;
  assign n49806 = n49449 | n49805 ;
  assign n49807 = n71164 & n49806 ;
  assign n49808 = n81425 & n49807 ;
  assign n49809 = n49803 | n49808 ;
  assign n49810 = n67763 & n49809 ;
  assign n49811 = n49086 & n49551 ;
  assign n81478 = ~n49620 ;
  assign n49622 = n49443 & n81478 ;
  assign n49812 = n49096 | n49443 ;
  assign n81479 = ~n49812 ;
  assign n49813 = n49439 & n81479 ;
  assign n49814 = n49622 | n49813 ;
  assign n49815 = n71164 & n49814 ;
  assign n49816 = n81425 & n49815 ;
  assign n49817 = n49811 | n49816 ;
  assign n49818 = n67622 & n49817 ;
  assign n81480 = ~n49816 ;
  assign n50167 = x91 & n81480 ;
  assign n81481 = ~n49811 ;
  assign n50168 = n81481 & n50167 ;
  assign n50169 = n49818 | n50168 ;
  assign n49819 = n49095 & n49551 ;
  assign n81482 = ~n49434 ;
  assign n49438 = n81482 & n49437 ;
  assign n49820 = n49105 | n49437 ;
  assign n81483 = ~n49820 ;
  assign n49821 = n49616 & n81483 ;
  assign n49822 = n49438 | n49821 ;
  assign n49823 = n71164 & n49822 ;
  assign n49824 = n81425 & n49823 ;
  assign n49825 = n49819 | n49824 ;
  assign n49826 = n67531 & n49825 ;
  assign n49827 = n49104 & n49551 ;
  assign n81484 = ~n49615 ;
  assign n49617 = n49432 & n81484 ;
  assign n49828 = n49114 | n49432 ;
  assign n81485 = ~n49828 ;
  assign n49829 = n49428 & n81485 ;
  assign n49830 = n49617 | n49829 ;
  assign n49831 = n71164 & n49830 ;
  assign n49832 = n81425 & n49831 ;
  assign n49833 = n49827 | n49832 ;
  assign n49834 = n67348 & n49833 ;
  assign n81486 = ~n49832 ;
  assign n50157 = x89 & n81486 ;
  assign n81487 = ~n49827 ;
  assign n50158 = n81487 & n50157 ;
  assign n50159 = n49834 | n50158 ;
  assign n49835 = n49113 & n49551 ;
  assign n81488 = ~n49423 ;
  assign n49427 = n81488 & n49426 ;
  assign n49836 = n49123 | n49426 ;
  assign n81489 = ~n49836 ;
  assign n49837 = n49611 & n81489 ;
  assign n49838 = n49427 | n49837 ;
  assign n49839 = n71164 & n49838 ;
  assign n49840 = n81425 & n49839 ;
  assign n49841 = n49835 | n49840 ;
  assign n49842 = n67222 & n49841 ;
  assign n49843 = n49122 & n49551 ;
  assign n81490 = ~n49610 ;
  assign n49612 = n49421 & n81490 ;
  assign n49844 = n49132 | n49421 ;
  assign n81491 = ~n49844 ;
  assign n49845 = n49417 & n81491 ;
  assign n49846 = n49612 | n49845 ;
  assign n49847 = n71164 & n49846 ;
  assign n49848 = n81425 & n49847 ;
  assign n49849 = n49843 | n49848 ;
  assign n49850 = n67164 & n49849 ;
  assign n81492 = ~n49848 ;
  assign n50146 = x87 & n81492 ;
  assign n81493 = ~n49843 ;
  assign n50147 = n81493 & n50146 ;
  assign n50148 = n49850 | n50147 ;
  assign n49851 = n49131 & n49551 ;
  assign n81494 = ~n49412 ;
  assign n49416 = n81494 & n49415 ;
  assign n49852 = n49141 | n49415 ;
  assign n81495 = ~n49852 ;
  assign n49853 = n49606 & n81495 ;
  assign n49854 = n49416 | n49853 ;
  assign n49855 = n71164 & n49854 ;
  assign n49856 = n81425 & n49855 ;
  assign n49857 = n49851 | n49856 ;
  assign n49858 = n66979 & n49857 ;
  assign n49859 = n49140 & n49551 ;
  assign n81496 = ~n49605 ;
  assign n49607 = n49410 & n81496 ;
  assign n49860 = n49150 | n49410 ;
  assign n81497 = ~n49860 ;
  assign n49861 = n49406 & n81497 ;
  assign n49862 = n49607 | n49861 ;
  assign n49863 = n71164 & n49862 ;
  assign n49864 = n81425 & n49863 ;
  assign n49865 = n49859 | n49864 ;
  assign n49866 = n66868 & n49865 ;
  assign n81498 = ~n49864 ;
  assign n50136 = x85 & n81498 ;
  assign n81499 = ~n49859 ;
  assign n50137 = n81499 & n50136 ;
  assign n50138 = n49866 | n50137 ;
  assign n49867 = n49149 & n49551 ;
  assign n81500 = ~n49401 ;
  assign n49405 = n81500 & n49404 ;
  assign n49868 = n49159 | n49404 ;
  assign n81501 = ~n49868 ;
  assign n49869 = n49601 & n81501 ;
  assign n49870 = n49405 | n49869 ;
  assign n49871 = n71164 & n49870 ;
  assign n49872 = n81425 & n49871 ;
  assign n49873 = n49867 | n49872 ;
  assign n49874 = n66797 & n49873 ;
  assign n49875 = n49158 & n49551 ;
  assign n81502 = ~n49600 ;
  assign n49602 = n49399 & n81502 ;
  assign n49876 = n49168 | n49399 ;
  assign n81503 = ~n49876 ;
  assign n49877 = n49395 & n81503 ;
  assign n49878 = n49602 | n49877 ;
  assign n49879 = n71164 & n49878 ;
  assign n49880 = n81425 & n49879 ;
  assign n49881 = n49875 | n49880 ;
  assign n49882 = n66654 & n49881 ;
  assign n81504 = ~n49880 ;
  assign n50126 = x83 & n81504 ;
  assign n81505 = ~n49875 ;
  assign n50127 = n81505 & n50126 ;
  assign n50128 = n49882 | n50127 ;
  assign n49883 = n49167 & n49551 ;
  assign n81506 = ~n49390 ;
  assign n49394 = n81506 & n49393 ;
  assign n49884 = n49177 | n49393 ;
  assign n81507 = ~n49884 ;
  assign n49885 = n49596 & n81507 ;
  assign n49886 = n49394 | n49885 ;
  assign n49887 = n71164 & n49886 ;
  assign n49888 = n81425 & n49887 ;
  assign n49889 = n49883 | n49888 ;
  assign n49890 = n66560 & n49889 ;
  assign n49891 = n49176 & n49551 ;
  assign n81508 = ~n49595 ;
  assign n49597 = n49388 & n81508 ;
  assign n49892 = n49186 | n49388 ;
  assign n81509 = ~n49892 ;
  assign n49893 = n49384 & n81509 ;
  assign n49894 = n49597 | n49893 ;
  assign n49895 = n71164 & n49894 ;
  assign n49896 = n81425 & n49895 ;
  assign n49897 = n49891 | n49896 ;
  assign n49898 = n66505 & n49897 ;
  assign n81510 = ~n49896 ;
  assign n50116 = x81 & n81510 ;
  assign n81511 = ~n49891 ;
  assign n50117 = n81511 & n50116 ;
  assign n50118 = n49898 | n50117 ;
  assign n49899 = n49185 & n49551 ;
  assign n81512 = ~n49379 ;
  assign n49383 = n81512 & n49382 ;
  assign n49900 = n49194 | n49382 ;
  assign n81513 = ~n49900 ;
  assign n49901 = n49591 & n81513 ;
  assign n49902 = n49383 | n49901 ;
  assign n49903 = n71164 & n49902 ;
  assign n49904 = n81425 & n49903 ;
  assign n49905 = n49899 | n49904 ;
  assign n49906 = n66379 & n49905 ;
  assign n49907 = n49193 & n49551 ;
  assign n81514 = ~n49590 ;
  assign n49592 = n49377 & n81514 ;
  assign n49908 = n49203 | n49377 ;
  assign n81515 = ~n49908 ;
  assign n49909 = n49373 & n81515 ;
  assign n49910 = n49592 | n49909 ;
  assign n49911 = n71164 & n49910 ;
  assign n49912 = n81425 & n49911 ;
  assign n49913 = n49907 | n49912 ;
  assign n49914 = n66299 & n49913 ;
  assign n81516 = ~n49912 ;
  assign n50106 = x79 & n81516 ;
  assign n81517 = ~n49907 ;
  assign n50107 = n81517 & n50106 ;
  assign n50108 = n49914 | n50107 ;
  assign n49915 = n49202 & n49551 ;
  assign n81518 = ~n49368 ;
  assign n49372 = n81518 & n49371 ;
  assign n49916 = n49212 | n49371 ;
  assign n81519 = ~n49916 ;
  assign n49917 = n49586 & n81519 ;
  assign n49918 = n49372 | n49917 ;
  assign n49919 = n71164 & n49918 ;
  assign n49920 = n81425 & n49919 ;
  assign n49921 = n49915 | n49920 ;
  assign n49922 = n66244 & n49921 ;
  assign n49923 = n49211 & n49551 ;
  assign n81520 = ~n49585 ;
  assign n49587 = n49366 & n81520 ;
  assign n49924 = n49221 | n49366 ;
  assign n81521 = ~n49924 ;
  assign n49925 = n49362 & n81521 ;
  assign n49926 = n49587 | n49925 ;
  assign n49927 = n71164 & n49926 ;
  assign n49928 = n81425 & n49927 ;
  assign n49929 = n49923 | n49928 ;
  assign n49930 = n66145 & n49929 ;
  assign n81522 = ~n49928 ;
  assign n50096 = x77 & n81522 ;
  assign n81523 = ~n49923 ;
  assign n50097 = n81523 & n50096 ;
  assign n50098 = n49930 | n50097 ;
  assign n49931 = n49220 & n49551 ;
  assign n81524 = ~n49357 ;
  assign n49361 = n81524 & n49360 ;
  assign n49932 = n49229 | n49360 ;
  assign n81525 = ~n49932 ;
  assign n49933 = n49581 & n81525 ;
  assign n49934 = n49361 | n49933 ;
  assign n49935 = n71164 & n49934 ;
  assign n49936 = n81425 & n49935 ;
  assign n49937 = n49931 | n49936 ;
  assign n49938 = n66081 & n49937 ;
  assign n49939 = n49228 & n49551 ;
  assign n81526 = ~n49580 ;
  assign n49582 = n49355 & n81526 ;
  assign n49940 = n49238 | n49355 ;
  assign n81527 = ~n49940 ;
  assign n49941 = n49351 & n81527 ;
  assign n49942 = n49582 | n49941 ;
  assign n49943 = n71164 & n49942 ;
  assign n49944 = n81425 & n49943 ;
  assign n49945 = n49939 | n49944 ;
  assign n49946 = n66043 & n49945 ;
  assign n81528 = ~n49944 ;
  assign n50086 = x75 & n81528 ;
  assign n81529 = ~n49939 ;
  assign n50087 = n81529 & n50086 ;
  assign n50088 = n49946 | n50087 ;
  assign n49947 = n49237 & n49551 ;
  assign n81530 = ~n49346 ;
  assign n49350 = n81530 & n49349 ;
  assign n49948 = n49246 | n49349 ;
  assign n81531 = ~n49948 ;
  assign n49949 = n49576 & n81531 ;
  assign n49950 = n49350 | n49949 ;
  assign n49951 = n71164 & n49950 ;
  assign n49952 = n81425 & n49951 ;
  assign n49953 = n49947 | n49952 ;
  assign n49954 = n65960 & n49953 ;
  assign n49955 = n49245 & n49551 ;
  assign n81532 = ~n49575 ;
  assign n49577 = n49344 & n81532 ;
  assign n49956 = n49255 | n49344 ;
  assign n81533 = ~n49956 ;
  assign n49957 = n49340 & n81533 ;
  assign n49958 = n49577 | n49957 ;
  assign n49959 = n71164 & n49958 ;
  assign n49960 = n81425 & n49959 ;
  assign n49961 = n49955 | n49960 ;
  assign n49962 = n65909 & n49961 ;
  assign n81534 = ~n49960 ;
  assign n50076 = x73 & n81534 ;
  assign n81535 = ~n49955 ;
  assign n50077 = n81535 & n50076 ;
  assign n50078 = n49962 | n50077 ;
  assign n49963 = n49254 & n49551 ;
  assign n81536 = ~n49335 ;
  assign n49339 = n81536 & n49338 ;
  assign n49964 = n49333 | n49570 ;
  assign n49965 = n49264 | n49338 ;
  assign n81537 = ~n49965 ;
  assign n49966 = n49964 & n81537 ;
  assign n49967 = n49339 | n49966 ;
  assign n49968 = n71164 & n49967 ;
  assign n49969 = n81425 & n49968 ;
  assign n49970 = n49963 | n49969 ;
  assign n49971 = n65877 & n49970 ;
  assign n49972 = n49263 & n49551 ;
  assign n81538 = ~n49570 ;
  assign n49572 = n49333 & n81538 ;
  assign n49973 = n49326 | n49567 ;
  assign n49974 = n49273 | n49333 ;
  assign n81539 = ~n49974 ;
  assign n49975 = n49973 & n81539 ;
  assign n49976 = n49572 | n49975 ;
  assign n49977 = n71164 & n49976 ;
  assign n49978 = n81425 & n49977 ;
  assign n49979 = n49972 | n49978 ;
  assign n49980 = n65820 & n49979 ;
  assign n81540 = ~n49978 ;
  assign n50065 = x71 & n81540 ;
  assign n81541 = ~n49972 ;
  assign n50066 = n81541 & n50065 ;
  assign n50067 = n49980 | n50066 ;
  assign n49981 = n49272 & n49551 ;
  assign n81542 = ~n49326 ;
  assign n49568 = n81542 & n49567 ;
  assign n49982 = n49324 | n49563 ;
  assign n49983 = n49282 | n49567 ;
  assign n81543 = ~n49983 ;
  assign n49984 = n49982 & n81543 ;
  assign n49985 = n49568 | n49984 ;
  assign n49986 = n71164 & n49985 ;
  assign n49987 = n81425 & n49986 ;
  assign n49988 = n49981 | n49987 ;
  assign n49989 = n65791 & n49988 ;
  assign n49990 = n49281 & n49551 ;
  assign n81544 = ~n49563 ;
  assign n49565 = n49324 & n81544 ;
  assign n49991 = n49317 | n49560 ;
  assign n49992 = n49290 | n49324 ;
  assign n81545 = ~n49992 ;
  assign n49993 = n49991 & n81545 ;
  assign n49994 = n49565 | n49993 ;
  assign n49995 = n71164 & n49994 ;
  assign n49996 = n81425 & n49995 ;
  assign n49997 = n49990 | n49996 ;
  assign n49998 = n65772 & n49997 ;
  assign n81546 = ~n49996 ;
  assign n50055 = x69 & n81546 ;
  assign n81547 = ~n49990 ;
  assign n50056 = n81547 & n50055 ;
  assign n50057 = n49998 | n50056 ;
  assign n49999 = n49289 & n49551 ;
  assign n81548 = ~n49317 ;
  assign n49561 = n81548 & n49560 ;
  assign n50000 = n49298 | n49560 ;
  assign n81549 = ~n50000 ;
  assign n50001 = n49316 & n81549 ;
  assign n50002 = n49561 | n50001 ;
  assign n50003 = n71164 & n50002 ;
  assign n50004 = n81425 & n50003 ;
  assign n50005 = n49999 | n50004 ;
  assign n50006 = n65746 & n50005 ;
  assign n50007 = n49297 & n49551 ;
  assign n50008 = n49311 | n49315 ;
  assign n81550 = ~n50008 ;
  assign n50009 = n49556 & n81550 ;
  assign n81551 = ~n49557 ;
  assign n50010 = n49315 & n81551 ;
  assign n50011 = n50009 | n50010 ;
  assign n50012 = n71164 & n50011 ;
  assign n50013 = n81425 & n50012 ;
  assign n50014 = n50007 | n50013 ;
  assign n50015 = n65721 & n50014 ;
  assign n81552 = ~n50013 ;
  assign n50045 = x67 & n81552 ;
  assign n81553 = ~n50007 ;
  assign n50046 = n81553 & n50045 ;
  assign n50047 = n50015 | n50046 ;
  assign n50016 = n49551 & n49553 ;
  assign n50017 = n17058 & n49308 ;
  assign n50018 = n81288 & n50017 ;
  assign n50019 = n17324 | n50018 ;
  assign n81554 = ~n50019 ;
  assign n50020 = n49556 & n81554 ;
  assign n50021 = n81425 & n50020 ;
  assign n50022 = n50016 | n50021 ;
  assign n50023 = n65686 & n50022 ;
  assign n50024 = n17774 & n81425 ;
  assign n81555 = ~n50024 ;
  assign n50025 = x18 & n81555 ;
  assign n50026 = n17785 & n81425 ;
  assign n50027 = n50025 | n50026 ;
  assign n50028 = x65 & n50027 ;
  assign n49667 = n49542 | n49665 ;
  assign n50029 = n81418 & n49667 ;
  assign n50030 = n49547 | n50029 ;
  assign n50031 = n81421 & n50030 ;
  assign n81556 = ~n50031 ;
  assign n50032 = n17774 & n81556 ;
  assign n81557 = ~n50032 ;
  assign n50033 = x18 & n81557 ;
  assign n50034 = x65 | n50026 ;
  assign n50035 = n50033 | n50034 ;
  assign n81558 = ~n50028 ;
  assign n50036 = n81558 & n50035 ;
  assign n50037 = n17792 | n50036 ;
  assign n50038 = n50026 | n50033 ;
  assign n50039 = n65670 & n50038 ;
  assign n81559 = ~n50039 ;
  assign n50040 = n50037 & n81559 ;
  assign n81560 = ~n50021 ;
  assign n50041 = x66 & n81560 ;
  assign n81561 = ~n50016 ;
  assign n50042 = n81561 & n50041 ;
  assign n50043 = n50023 | n50042 ;
  assign n50044 = n50040 | n50043 ;
  assign n81562 = ~n50023 ;
  assign n50048 = n81562 & n50044 ;
  assign n50049 = n50047 | n50048 ;
  assign n81563 = ~n50015 ;
  assign n50050 = n81563 & n50049 ;
  assign n81564 = ~n50004 ;
  assign n50051 = x68 & n81564 ;
  assign n81565 = ~n49999 ;
  assign n50052 = n81565 & n50051 ;
  assign n50053 = n50006 | n50052 ;
  assign n50054 = n50050 | n50053 ;
  assign n81566 = ~n50006 ;
  assign n50058 = n81566 & n50054 ;
  assign n50059 = n50057 | n50058 ;
  assign n81567 = ~n49998 ;
  assign n50060 = n81567 & n50059 ;
  assign n81568 = ~n49987 ;
  assign n50061 = x70 & n81568 ;
  assign n81569 = ~n49981 ;
  assign n50062 = n81569 & n50061 ;
  assign n50063 = n49989 | n50062 ;
  assign n50064 = n50060 | n50063 ;
  assign n81570 = ~n49989 ;
  assign n50069 = n81570 & n50064 ;
  assign n50070 = n50067 | n50069 ;
  assign n81571 = ~n49980 ;
  assign n50071 = n81571 & n50070 ;
  assign n81572 = ~n49969 ;
  assign n50072 = x72 & n81572 ;
  assign n81573 = ~n49963 ;
  assign n50073 = n81573 & n50072 ;
  assign n50074 = n49971 | n50073 ;
  assign n50075 = n50071 | n50074 ;
  assign n81574 = ~n49971 ;
  assign n50079 = n81574 & n50075 ;
  assign n50080 = n50078 | n50079 ;
  assign n81575 = ~n49962 ;
  assign n50081 = n81575 & n50080 ;
  assign n81576 = ~n49952 ;
  assign n50082 = x74 & n81576 ;
  assign n81577 = ~n49947 ;
  assign n50083 = n81577 & n50082 ;
  assign n50084 = n49954 | n50083 ;
  assign n50085 = n50081 | n50084 ;
  assign n81578 = ~n49954 ;
  assign n50089 = n81578 & n50085 ;
  assign n50090 = n50088 | n50089 ;
  assign n81579 = ~n49946 ;
  assign n50091 = n81579 & n50090 ;
  assign n81580 = ~n49936 ;
  assign n50092 = x76 & n81580 ;
  assign n81581 = ~n49931 ;
  assign n50093 = n81581 & n50092 ;
  assign n50094 = n49938 | n50093 ;
  assign n50095 = n50091 | n50094 ;
  assign n81582 = ~n49938 ;
  assign n50099 = n81582 & n50095 ;
  assign n50100 = n50098 | n50099 ;
  assign n81583 = ~n49930 ;
  assign n50101 = n81583 & n50100 ;
  assign n81584 = ~n49920 ;
  assign n50102 = x78 & n81584 ;
  assign n81585 = ~n49915 ;
  assign n50103 = n81585 & n50102 ;
  assign n50104 = n49922 | n50103 ;
  assign n50105 = n50101 | n50104 ;
  assign n81586 = ~n49922 ;
  assign n50109 = n81586 & n50105 ;
  assign n50110 = n50108 | n50109 ;
  assign n81587 = ~n49914 ;
  assign n50111 = n81587 & n50110 ;
  assign n81588 = ~n49904 ;
  assign n50112 = x80 & n81588 ;
  assign n81589 = ~n49899 ;
  assign n50113 = n81589 & n50112 ;
  assign n50114 = n49906 | n50113 ;
  assign n50115 = n50111 | n50114 ;
  assign n81590 = ~n49906 ;
  assign n50119 = n81590 & n50115 ;
  assign n50120 = n50118 | n50119 ;
  assign n81591 = ~n49898 ;
  assign n50121 = n81591 & n50120 ;
  assign n81592 = ~n49888 ;
  assign n50122 = x82 & n81592 ;
  assign n81593 = ~n49883 ;
  assign n50123 = n81593 & n50122 ;
  assign n50124 = n49890 | n50123 ;
  assign n50125 = n50121 | n50124 ;
  assign n81594 = ~n49890 ;
  assign n50129 = n81594 & n50125 ;
  assign n50130 = n50128 | n50129 ;
  assign n81595 = ~n49882 ;
  assign n50131 = n81595 & n50130 ;
  assign n81596 = ~n49872 ;
  assign n50132 = x84 & n81596 ;
  assign n81597 = ~n49867 ;
  assign n50133 = n81597 & n50132 ;
  assign n50134 = n49874 | n50133 ;
  assign n50135 = n50131 | n50134 ;
  assign n81598 = ~n49874 ;
  assign n50139 = n81598 & n50135 ;
  assign n50140 = n50138 | n50139 ;
  assign n81599 = ~n49866 ;
  assign n50141 = n81599 & n50140 ;
  assign n81600 = ~n49856 ;
  assign n50142 = x86 & n81600 ;
  assign n81601 = ~n49851 ;
  assign n50143 = n81601 & n50142 ;
  assign n50144 = n49858 | n50143 ;
  assign n50145 = n50141 | n50144 ;
  assign n81602 = ~n49858 ;
  assign n50150 = n81602 & n50145 ;
  assign n50151 = n50148 | n50150 ;
  assign n81603 = ~n49850 ;
  assign n50152 = n81603 & n50151 ;
  assign n81604 = ~n49840 ;
  assign n50153 = x88 & n81604 ;
  assign n81605 = ~n49835 ;
  assign n50154 = n81605 & n50153 ;
  assign n50155 = n49842 | n50154 ;
  assign n50156 = n50152 | n50155 ;
  assign n81606 = ~n49842 ;
  assign n50160 = n81606 & n50156 ;
  assign n50161 = n50159 | n50160 ;
  assign n81607 = ~n49834 ;
  assign n50162 = n81607 & n50161 ;
  assign n81608 = ~n49824 ;
  assign n50163 = x90 & n81608 ;
  assign n81609 = ~n49819 ;
  assign n50164 = n81609 & n50163 ;
  assign n50165 = n49826 | n50164 ;
  assign n50166 = n50162 | n50165 ;
  assign n81610 = ~n49826 ;
  assign n50171 = n81610 & n50166 ;
  assign n50172 = n50169 | n50171 ;
  assign n81611 = ~n49818 ;
  assign n50173 = n81611 & n50172 ;
  assign n81612 = ~n49808 ;
  assign n50174 = x92 & n81612 ;
  assign n81613 = ~n49803 ;
  assign n50175 = n81613 & n50174 ;
  assign n50176 = n49810 | n50175 ;
  assign n50177 = n50173 | n50176 ;
  assign n81614 = ~n49810 ;
  assign n50181 = n81614 & n50177 ;
  assign n50182 = n50180 | n50181 ;
  assign n81615 = ~n49802 ;
  assign n50183 = n81615 & n50182 ;
  assign n81616 = ~n49792 ;
  assign n50184 = x94 & n81616 ;
  assign n81617 = ~n49787 ;
  assign n50185 = n81617 & n50184 ;
  assign n50186 = n49794 | n50185 ;
  assign n50187 = n50183 | n50186 ;
  assign n81618 = ~n49794 ;
  assign n50191 = n81618 & n50187 ;
  assign n50192 = n50190 | n50191 ;
  assign n81619 = ~n49786 ;
  assign n50193 = n81619 & n50192 ;
  assign n81620 = ~n49776 ;
  assign n50194 = x96 & n81620 ;
  assign n81621 = ~n49771 ;
  assign n50195 = n81621 & n50194 ;
  assign n50196 = n49778 | n50195 ;
  assign n50197 = n50193 | n50196 ;
  assign n81622 = ~n49778 ;
  assign n50201 = n81622 & n50197 ;
  assign n50202 = n50200 | n50201 ;
  assign n81623 = ~n49770 ;
  assign n50203 = n81623 & n50202 ;
  assign n81624 = ~n49760 ;
  assign n50204 = x98 & n81624 ;
  assign n81625 = ~n49755 ;
  assign n50205 = n81625 & n50204 ;
  assign n50206 = n49762 | n50205 ;
  assign n50207 = n50203 | n50206 ;
  assign n81626 = ~n49762 ;
  assign n50212 = n81626 & n50207 ;
  assign n50213 = n50210 | n50212 ;
  assign n81627 = ~n49754 ;
  assign n50214 = n81627 & n50213 ;
  assign n81628 = ~n49744 ;
  assign n50215 = x100 & n81628 ;
  assign n81629 = ~n49739 ;
  assign n50216 = n81629 & n50215 ;
  assign n50217 = n49746 | n50216 ;
  assign n50218 = n50214 | n50217 ;
  assign n81630 = ~n49746 ;
  assign n50222 = n81630 & n50218 ;
  assign n50223 = n50221 | n50222 ;
  assign n81631 = ~n49738 ;
  assign n50224 = n81631 & n50223 ;
  assign n81632 = ~n49728 ;
  assign n50225 = x102 & n81632 ;
  assign n81633 = ~n49723 ;
  assign n50226 = n81633 & n50225 ;
  assign n50227 = n49730 | n50226 ;
  assign n50228 = n50224 | n50227 ;
  assign n81634 = ~n49730 ;
  assign n50232 = n81634 & n50228 ;
  assign n50233 = n50231 | n50232 ;
  assign n81635 = ~n49722 ;
  assign n50234 = n81635 & n50233 ;
  assign n81636 = ~n49712 ;
  assign n50235 = x104 & n81636 ;
  assign n81637 = ~n49707 ;
  assign n50236 = n81637 & n50235 ;
  assign n50237 = n49714 | n50236 ;
  assign n50238 = n50234 | n50237 ;
  assign n81638 = ~n49714 ;
  assign n50242 = n81638 & n50238 ;
  assign n50243 = n50241 | n50242 ;
  assign n81639 = ~n49706 ;
  assign n50244 = n81639 & n50243 ;
  assign n81640 = ~n49696 ;
  assign n50245 = x106 & n81640 ;
  assign n81641 = ~n49691 ;
  assign n50246 = n81641 & n50245 ;
  assign n50247 = n49698 | n50246 ;
  assign n50248 = n50244 | n50247 ;
  assign n81642 = ~n49698 ;
  assign n50252 = n81642 & n50248 ;
  assign n50253 = n50251 | n50252 ;
  assign n81643 = ~n49690 ;
  assign n50254 = n81643 & n50253 ;
  assign n81644 = ~n49680 ;
  assign n50255 = x108 & n81644 ;
  assign n81645 = ~n49675 ;
  assign n50256 = n81645 & n50255 ;
  assign n50257 = n49682 | n50256 ;
  assign n50258 = n50254 | n50257 ;
  assign n81646 = ~n49682 ;
  assign n50263 = n81646 & n50258 ;
  assign n50264 = n50261 | n50263 ;
  assign n81647 = ~n49674 ;
  assign n50265 = n81647 & n50264 ;
  assign n81648 = ~n49544 ;
  assign n49548 = n81648 & n49547 ;
  assign n50266 = n48927 | n49547 ;
  assign n81649 = ~n50266 ;
  assign n50267 = n49667 & n81649 ;
  assign n50268 = n49548 | n50267 ;
  assign n50269 = n49551 | n50268 ;
  assign n81650 = ~n48925 ;
  assign n50270 = n81650 & n49551 ;
  assign n81651 = ~n50270 ;
  assign n50271 = n50269 & n81651 ;
  assign n50272 = n71253 & n50271 ;
  assign n81652 = ~n49551 ;
  assign n50273 = n81652 & n50268 ;
  assign n50274 = n48925 & n49551 ;
  assign n81653 = ~n50274 ;
  assign n50275 = x110 & n81653 ;
  assign n81654 = ~n50273 ;
  assign n50276 = n81654 & n50275 ;
  assign n50277 = n18047 | n50276 ;
  assign n50278 = n50272 | n50277 ;
  assign n50279 = n50265 | n50278 ;
  assign n50280 = n71164 & n50271 ;
  assign n81655 = ~n50280 ;
  assign n50281 = n50279 & n81655 ;
  assign n51035 = n49674 | n50276 ;
  assign n51036 = n50272 | n51035 ;
  assign n81656 = ~n51036 ;
  assign n51037 = n50264 & n81656 ;
  assign n50291 = x65 & n50038 ;
  assign n81657 = ~n50291 ;
  assign n50292 = n50035 & n81657 ;
  assign n50293 = n17792 | n50292 ;
  assign n50294 = n81559 & n50293 ;
  assign n50295 = n50043 | n50294 ;
  assign n50296 = n81562 & n50295 ;
  assign n50297 = n50047 | n50296 ;
  assign n50298 = n81563 & n50297 ;
  assign n50299 = n50053 | n50298 ;
  assign n50300 = n81566 & n50299 ;
  assign n50301 = n50057 | n50300 ;
  assign n50302 = n81567 & n50301 ;
  assign n50303 = n50063 | n50302 ;
  assign n50304 = n81570 & n50303 ;
  assign n50305 = n50067 | n50304 ;
  assign n50306 = n81571 & n50305 ;
  assign n50307 = n50074 | n50306 ;
  assign n50308 = n81574 & n50307 ;
  assign n50309 = n50078 | n50308 ;
  assign n50310 = n81575 & n50309 ;
  assign n50311 = n50084 | n50310 ;
  assign n50312 = n81578 & n50311 ;
  assign n50313 = n50088 | n50312 ;
  assign n50314 = n81579 & n50313 ;
  assign n50315 = n50094 | n50314 ;
  assign n50316 = n81582 & n50315 ;
  assign n50317 = n50098 | n50316 ;
  assign n50318 = n81583 & n50317 ;
  assign n50319 = n50104 | n50318 ;
  assign n50320 = n81586 & n50319 ;
  assign n50321 = n50108 | n50320 ;
  assign n50322 = n81587 & n50321 ;
  assign n50323 = n50114 | n50322 ;
  assign n50324 = n81590 & n50323 ;
  assign n50325 = n50118 | n50324 ;
  assign n50326 = n81591 & n50325 ;
  assign n50327 = n50124 | n50326 ;
  assign n50328 = n81594 & n50327 ;
  assign n50329 = n50128 | n50328 ;
  assign n50330 = n81595 & n50329 ;
  assign n50331 = n50134 | n50330 ;
  assign n50332 = n81598 & n50331 ;
  assign n50333 = n50138 | n50332 ;
  assign n50334 = n81599 & n50333 ;
  assign n50335 = n50144 | n50334 ;
  assign n50336 = n81602 & n50335 ;
  assign n50337 = n50148 | n50336 ;
  assign n50338 = n81603 & n50337 ;
  assign n50339 = n50155 | n50338 ;
  assign n50340 = n81606 & n50339 ;
  assign n50341 = n50159 | n50340 ;
  assign n50342 = n81607 & n50341 ;
  assign n50343 = n50165 | n50342 ;
  assign n50344 = n81610 & n50343 ;
  assign n50345 = n50169 | n50344 ;
  assign n50346 = n81611 & n50345 ;
  assign n50347 = n50176 | n50346 ;
  assign n50348 = n81614 & n50347 ;
  assign n50349 = n50180 | n50348 ;
  assign n50350 = n81615 & n50349 ;
  assign n50351 = n50186 | n50350 ;
  assign n50352 = n81618 & n50351 ;
  assign n50353 = n50190 | n50352 ;
  assign n50354 = n81619 & n50353 ;
  assign n50355 = n50196 | n50354 ;
  assign n50356 = n81622 & n50355 ;
  assign n50357 = n50200 | n50356 ;
  assign n50358 = n81623 & n50357 ;
  assign n50359 = n50206 | n50358 ;
  assign n50360 = n81626 & n50359 ;
  assign n50361 = n50210 | n50360 ;
  assign n50362 = n81627 & n50361 ;
  assign n50363 = n50217 | n50362 ;
  assign n50364 = n81630 & n50363 ;
  assign n50365 = n50221 | n50364 ;
  assign n50366 = n81631 & n50365 ;
  assign n50367 = n50227 | n50366 ;
  assign n50368 = n81634 & n50367 ;
  assign n50369 = n50231 | n50368 ;
  assign n50370 = n81635 & n50369 ;
  assign n50371 = n50237 | n50370 ;
  assign n50372 = n81638 & n50371 ;
  assign n50373 = n50241 | n50372 ;
  assign n50374 = n81639 & n50373 ;
  assign n50375 = n50247 | n50374 ;
  assign n50376 = n81642 & n50375 ;
  assign n50377 = n50251 | n50376 ;
  assign n50378 = n81643 & n50377 ;
  assign n50773 = n50257 | n50378 ;
  assign n50774 = n81646 & n50773 ;
  assign n50775 = n50261 | n50774 ;
  assign n50776 = n81647 & n50775 ;
  assign n51038 = n50272 | n50276 ;
  assign n81658 = ~n50776 ;
  assign n51039 = n81658 & n51038 ;
  assign n51040 = n51037 | n51039 ;
  assign n81659 = ~n50281 ;
  assign n51041 = n81659 & n51040 ;
  assign n51042 = n17324 & n48925 ;
  assign n51043 = n50279 & n51042 ;
  assign n51044 = n51041 | n51043 ;
  assign n51050 = n71636 & n51044 ;
  assign n81660 = ~n50263 ;
  assign n50283 = n50261 & n81660 ;
  assign n50262 = n49682 | n50261 ;
  assign n81661 = ~n50262 ;
  assign n50284 = n50258 & n81661 ;
  assign n50285 = n50283 | n50284 ;
  assign n50286 = n81659 & n50285 ;
  assign n50287 = n49673 & n81655 ;
  assign n50288 = n50279 & n50287 ;
  assign n50289 = n50286 | n50288 ;
  assign n50290 = n71253 & n50289 ;
  assign n81662 = ~n50378 ;
  assign n50379 = n50257 & n81662 ;
  assign n50380 = n49690 | n50257 ;
  assign n81663 = ~n50380 ;
  assign n50381 = n50253 & n81663 ;
  assign n50382 = n50379 | n50381 ;
  assign n50383 = n81659 & n50382 ;
  assign n50384 = n49681 & n81655 ;
  assign n50385 = n50279 & n50384 ;
  assign n50386 = n50383 | n50385 ;
  assign n50387 = n70935 & n50386 ;
  assign n81664 = ~n50252 ;
  assign n50388 = n50251 & n81664 ;
  assign n50389 = n49698 | n50251 ;
  assign n81665 = ~n50389 ;
  assign n50390 = n50375 & n81665 ;
  assign n50391 = n50388 | n50390 ;
  assign n50392 = n81659 & n50391 ;
  assign n50393 = n49689 & n81655 ;
  assign n50394 = n50279 & n50393 ;
  assign n50395 = n50392 | n50394 ;
  assign n50396 = n70927 & n50395 ;
  assign n81666 = ~n50374 ;
  assign n50397 = n50247 & n81666 ;
  assign n50398 = n49706 | n50247 ;
  assign n81667 = ~n50398 ;
  assign n50399 = n50243 & n81667 ;
  assign n50400 = n50397 | n50399 ;
  assign n50401 = n81659 & n50400 ;
  assign n50402 = n49697 & n81655 ;
  assign n50403 = n50279 & n50402 ;
  assign n50404 = n50401 | n50403 ;
  assign n50405 = n70609 & n50404 ;
  assign n81668 = ~n50242 ;
  assign n50406 = n50241 & n81668 ;
  assign n50407 = n49714 | n50241 ;
  assign n81669 = ~n50407 ;
  assign n50408 = n50371 & n81669 ;
  assign n50409 = n50406 | n50408 ;
  assign n50410 = n81659 & n50409 ;
  assign n50411 = n49705 & n81655 ;
  assign n50412 = n50279 & n50411 ;
  assign n50413 = n50410 | n50412 ;
  assign n50414 = n70276 & n50413 ;
  assign n81670 = ~n50370 ;
  assign n50415 = n50237 & n81670 ;
  assign n50416 = n49722 | n50237 ;
  assign n81671 = ~n50416 ;
  assign n50417 = n50233 & n81671 ;
  assign n50418 = n50415 | n50417 ;
  assign n50419 = n81659 & n50418 ;
  assign n50420 = n49713 & n81655 ;
  assign n50421 = n50279 & n50420 ;
  assign n50422 = n50419 | n50421 ;
  assign n50423 = n70176 & n50422 ;
  assign n81672 = ~n50232 ;
  assign n50424 = n50231 & n81672 ;
  assign n50425 = n49730 | n50231 ;
  assign n81673 = ~n50425 ;
  assign n50426 = n50367 & n81673 ;
  assign n50427 = n50424 | n50426 ;
  assign n50428 = n81659 & n50427 ;
  assign n50429 = n49721 & n81655 ;
  assign n50430 = n50279 & n50429 ;
  assign n50431 = n50428 | n50430 ;
  assign n50432 = n69857 & n50431 ;
  assign n81674 = ~n50366 ;
  assign n50433 = n50227 & n81674 ;
  assign n50434 = n49738 | n50227 ;
  assign n81675 = ~n50434 ;
  assign n50435 = n50223 & n81675 ;
  assign n50436 = n50433 | n50435 ;
  assign n50437 = n81659 & n50436 ;
  assign n50438 = n49729 & n81655 ;
  assign n50439 = n50279 & n50438 ;
  assign n50440 = n50437 | n50439 ;
  assign n50441 = n69656 & n50440 ;
  assign n81676 = ~n50222 ;
  assign n50442 = n50221 & n81676 ;
  assign n50443 = n49746 | n50221 ;
  assign n81677 = ~n50443 ;
  assign n50444 = n50363 & n81677 ;
  assign n50445 = n50442 | n50444 ;
  assign n50446 = n81659 & n50445 ;
  assign n50447 = n49737 & n81655 ;
  assign n50448 = n50279 & n50447 ;
  assign n50449 = n50446 | n50448 ;
  assign n50450 = n69528 & n50449 ;
  assign n81678 = ~n50362 ;
  assign n50451 = n50217 & n81678 ;
  assign n50452 = n49754 | n50217 ;
  assign n81679 = ~n50452 ;
  assign n50453 = n50213 & n81679 ;
  assign n50454 = n50451 | n50453 ;
  assign n50455 = n81659 & n50454 ;
  assign n50456 = n49745 & n81655 ;
  assign n50457 = n50279 & n50456 ;
  assign n50458 = n50455 | n50457 ;
  assign n50459 = n69261 & n50458 ;
  assign n81680 = ~n50212 ;
  assign n50460 = n50210 & n81680 ;
  assign n50211 = n49762 | n50210 ;
  assign n81681 = ~n50211 ;
  assign n50461 = n50207 & n81681 ;
  assign n50462 = n50460 | n50461 ;
  assign n50463 = n81659 & n50462 ;
  assign n50464 = n49753 & n81655 ;
  assign n50465 = n50279 & n50464 ;
  assign n50466 = n50463 | n50465 ;
  assign n50467 = n69075 & n50466 ;
  assign n81682 = ~n50358 ;
  assign n50468 = n50206 & n81682 ;
  assign n50469 = n49770 | n50206 ;
  assign n81683 = ~n50469 ;
  assign n50470 = n50202 & n81683 ;
  assign n50471 = n50468 | n50470 ;
  assign n50472 = n81659 & n50471 ;
  assign n50473 = n49761 & n81655 ;
  assign n50474 = n50279 & n50473 ;
  assign n50475 = n50472 | n50474 ;
  assign n50476 = n68993 & n50475 ;
  assign n81684 = ~n50201 ;
  assign n50477 = n50200 & n81684 ;
  assign n50478 = n49778 | n50200 ;
  assign n81685 = ~n50478 ;
  assign n50479 = n50355 & n81685 ;
  assign n50480 = n50477 | n50479 ;
  assign n50481 = n81659 & n50480 ;
  assign n50482 = n49769 & n81655 ;
  assign n50483 = n50279 & n50482 ;
  assign n50484 = n50481 | n50483 ;
  assign n50485 = n68716 & n50484 ;
  assign n81686 = ~n50354 ;
  assign n50486 = n50196 & n81686 ;
  assign n50487 = n49786 | n50196 ;
  assign n81687 = ~n50487 ;
  assign n50488 = n50192 & n81687 ;
  assign n50489 = n50486 | n50488 ;
  assign n50490 = n81659 & n50489 ;
  assign n50491 = n49777 & n81655 ;
  assign n50492 = n50279 & n50491 ;
  assign n50493 = n50490 | n50492 ;
  assign n50494 = n68545 & n50493 ;
  assign n81688 = ~n50191 ;
  assign n50495 = n50190 & n81688 ;
  assign n50496 = n49794 | n50190 ;
  assign n81689 = ~n50496 ;
  assign n50497 = n50351 & n81689 ;
  assign n50498 = n50495 | n50497 ;
  assign n50499 = n81659 & n50498 ;
  assign n50500 = n49785 & n81655 ;
  assign n50501 = n50279 & n50500 ;
  assign n50502 = n50499 | n50501 ;
  assign n50503 = n68438 & n50502 ;
  assign n81690 = ~n50350 ;
  assign n50504 = n50186 & n81690 ;
  assign n50505 = n49802 | n50186 ;
  assign n81691 = ~n50505 ;
  assign n50506 = n50182 & n81691 ;
  assign n50507 = n50504 | n50506 ;
  assign n50508 = n81659 & n50507 ;
  assign n50509 = n49793 & n81655 ;
  assign n50510 = n50279 & n50509 ;
  assign n50511 = n50508 | n50510 ;
  assign n50512 = n68214 & n50511 ;
  assign n81692 = ~n50181 ;
  assign n50513 = n50180 & n81692 ;
  assign n50514 = n49810 | n50180 ;
  assign n81693 = ~n50514 ;
  assign n50515 = n50347 & n81693 ;
  assign n50516 = n50513 | n50515 ;
  assign n50517 = n81659 & n50516 ;
  assign n50518 = n49801 & n81655 ;
  assign n50519 = n50279 & n50518 ;
  assign n50520 = n50517 | n50519 ;
  assign n50521 = n68058 & n50520 ;
  assign n81694 = ~n50346 ;
  assign n50522 = n50176 & n81694 ;
  assign n50523 = n49818 | n50176 ;
  assign n81695 = ~n50523 ;
  assign n50524 = n50172 & n81695 ;
  assign n50525 = n50522 | n50524 ;
  assign n50526 = n81659 & n50525 ;
  assign n50527 = n49809 & n81655 ;
  assign n50528 = n50279 & n50527 ;
  assign n50529 = n50526 | n50528 ;
  assign n50530 = n67986 & n50529 ;
  assign n81696 = ~n50171 ;
  assign n50531 = n50169 & n81696 ;
  assign n50170 = n49826 | n50169 ;
  assign n81697 = ~n50170 ;
  assign n50532 = n50166 & n81697 ;
  assign n50533 = n50531 | n50532 ;
  assign n50534 = n81659 & n50533 ;
  assign n50535 = n49817 & n81655 ;
  assign n50536 = n50279 & n50535 ;
  assign n50537 = n50534 | n50536 ;
  assign n50538 = n67763 & n50537 ;
  assign n81698 = ~n50342 ;
  assign n50539 = n50165 & n81698 ;
  assign n50540 = n49834 | n50165 ;
  assign n81699 = ~n50540 ;
  assign n50541 = n50161 & n81699 ;
  assign n50542 = n50539 | n50541 ;
  assign n50543 = n81659 & n50542 ;
  assign n50544 = n49825 & n81655 ;
  assign n50545 = n50279 & n50544 ;
  assign n50546 = n50543 | n50545 ;
  assign n50547 = n67622 & n50546 ;
  assign n81700 = ~n50160 ;
  assign n50548 = n50159 & n81700 ;
  assign n50549 = n49842 | n50159 ;
  assign n81701 = ~n50549 ;
  assign n50550 = n50339 & n81701 ;
  assign n50551 = n50548 | n50550 ;
  assign n50552 = n81659 & n50551 ;
  assign n50553 = n49833 & n81655 ;
  assign n50554 = n50279 & n50553 ;
  assign n50555 = n50552 | n50554 ;
  assign n50556 = n67531 & n50555 ;
  assign n81702 = ~n50338 ;
  assign n50557 = n50155 & n81702 ;
  assign n50558 = n49850 | n50155 ;
  assign n81703 = ~n50558 ;
  assign n50559 = n50151 & n81703 ;
  assign n50560 = n50557 | n50559 ;
  assign n50561 = n81659 & n50560 ;
  assign n50562 = n49841 & n81655 ;
  assign n50563 = n50279 & n50562 ;
  assign n50564 = n50561 | n50563 ;
  assign n50565 = n67348 & n50564 ;
  assign n81704 = ~n50150 ;
  assign n50566 = n50148 & n81704 ;
  assign n50149 = n49858 | n50148 ;
  assign n81705 = ~n50149 ;
  assign n50567 = n50145 & n81705 ;
  assign n50568 = n50566 | n50567 ;
  assign n50569 = n81659 & n50568 ;
  assign n50570 = n49849 & n81655 ;
  assign n50571 = n50279 & n50570 ;
  assign n50572 = n50569 | n50571 ;
  assign n50573 = n67222 & n50572 ;
  assign n81706 = ~n50334 ;
  assign n50574 = n50144 & n81706 ;
  assign n50575 = n49866 | n50144 ;
  assign n81707 = ~n50575 ;
  assign n50576 = n50140 & n81707 ;
  assign n50577 = n50574 | n50576 ;
  assign n50578 = n81659 & n50577 ;
  assign n50579 = n49857 & n81655 ;
  assign n50580 = n50279 & n50579 ;
  assign n50581 = n50578 | n50580 ;
  assign n50582 = n67164 & n50581 ;
  assign n81708 = ~n50139 ;
  assign n50583 = n50138 & n81708 ;
  assign n50584 = n49874 | n50138 ;
  assign n81709 = ~n50584 ;
  assign n50585 = n50331 & n81709 ;
  assign n50586 = n50583 | n50585 ;
  assign n50587 = n81659 & n50586 ;
  assign n50588 = n49865 & n81655 ;
  assign n50589 = n50279 & n50588 ;
  assign n50590 = n50587 | n50589 ;
  assign n50591 = n66979 & n50590 ;
  assign n81710 = ~n50330 ;
  assign n50592 = n50134 & n81710 ;
  assign n50593 = n49882 | n50134 ;
  assign n81711 = ~n50593 ;
  assign n50594 = n50130 & n81711 ;
  assign n50595 = n50592 | n50594 ;
  assign n50596 = n81659 & n50595 ;
  assign n50597 = n49873 & n81655 ;
  assign n50598 = n50279 & n50597 ;
  assign n50599 = n50596 | n50598 ;
  assign n50600 = n66868 & n50599 ;
  assign n81712 = ~n50129 ;
  assign n50601 = n50128 & n81712 ;
  assign n50602 = n49890 | n50128 ;
  assign n81713 = ~n50602 ;
  assign n50603 = n50327 & n81713 ;
  assign n50604 = n50601 | n50603 ;
  assign n50605 = n81659 & n50604 ;
  assign n50606 = n49881 & n81655 ;
  assign n50607 = n50279 & n50606 ;
  assign n50608 = n50605 | n50607 ;
  assign n50609 = n66797 & n50608 ;
  assign n81714 = ~n50326 ;
  assign n50610 = n50124 & n81714 ;
  assign n50611 = n49898 | n50124 ;
  assign n81715 = ~n50611 ;
  assign n50612 = n50120 & n81715 ;
  assign n50613 = n50610 | n50612 ;
  assign n50614 = n81659 & n50613 ;
  assign n50615 = n49889 & n81655 ;
  assign n50616 = n50279 & n50615 ;
  assign n50617 = n50614 | n50616 ;
  assign n50618 = n66654 & n50617 ;
  assign n81716 = ~n50119 ;
  assign n50619 = n50118 & n81716 ;
  assign n50620 = n49906 | n50118 ;
  assign n81717 = ~n50620 ;
  assign n50621 = n50323 & n81717 ;
  assign n50622 = n50619 | n50621 ;
  assign n50623 = n81659 & n50622 ;
  assign n50624 = n49897 & n81655 ;
  assign n50625 = n50279 & n50624 ;
  assign n50626 = n50623 | n50625 ;
  assign n50627 = n66560 & n50626 ;
  assign n81718 = ~n50322 ;
  assign n50628 = n50114 & n81718 ;
  assign n50629 = n49914 | n50114 ;
  assign n81719 = ~n50629 ;
  assign n50630 = n50110 & n81719 ;
  assign n50631 = n50628 | n50630 ;
  assign n50632 = n81659 & n50631 ;
  assign n50633 = n49905 & n81655 ;
  assign n50634 = n50279 & n50633 ;
  assign n50635 = n50632 | n50634 ;
  assign n50636 = n66505 & n50635 ;
  assign n81720 = ~n50109 ;
  assign n50637 = n50108 & n81720 ;
  assign n50638 = n49922 | n50108 ;
  assign n81721 = ~n50638 ;
  assign n50639 = n50319 & n81721 ;
  assign n50640 = n50637 | n50639 ;
  assign n50641 = n81659 & n50640 ;
  assign n50642 = n49913 & n81655 ;
  assign n50643 = n50279 & n50642 ;
  assign n50644 = n50641 | n50643 ;
  assign n50645 = n66379 & n50644 ;
  assign n81722 = ~n50318 ;
  assign n50646 = n50104 & n81722 ;
  assign n50647 = n49930 | n50104 ;
  assign n81723 = ~n50647 ;
  assign n50648 = n50100 & n81723 ;
  assign n50649 = n50646 | n50648 ;
  assign n50650 = n81659 & n50649 ;
  assign n50651 = n49921 & n81655 ;
  assign n50652 = n50279 & n50651 ;
  assign n50653 = n50650 | n50652 ;
  assign n50654 = n66299 & n50653 ;
  assign n81724 = ~n50099 ;
  assign n50655 = n50098 & n81724 ;
  assign n50656 = n49938 | n50098 ;
  assign n81725 = ~n50656 ;
  assign n50657 = n50315 & n81725 ;
  assign n50658 = n50655 | n50657 ;
  assign n50659 = n81659 & n50658 ;
  assign n50660 = n49929 & n81655 ;
  assign n50661 = n50279 & n50660 ;
  assign n50662 = n50659 | n50661 ;
  assign n50663 = n66244 & n50662 ;
  assign n81726 = ~n50314 ;
  assign n50664 = n50094 & n81726 ;
  assign n50665 = n49946 | n50094 ;
  assign n81727 = ~n50665 ;
  assign n50666 = n50090 & n81727 ;
  assign n50667 = n50664 | n50666 ;
  assign n50668 = n81659 & n50667 ;
  assign n50669 = n49937 & n81655 ;
  assign n50670 = n50279 & n50669 ;
  assign n50671 = n50668 | n50670 ;
  assign n50672 = n66145 & n50671 ;
  assign n81728 = ~n50089 ;
  assign n50673 = n50088 & n81728 ;
  assign n50674 = n49954 | n50088 ;
  assign n81729 = ~n50674 ;
  assign n50675 = n50311 & n81729 ;
  assign n50676 = n50673 | n50675 ;
  assign n50677 = n81659 & n50676 ;
  assign n50678 = n49945 & n81655 ;
  assign n50679 = n50279 & n50678 ;
  assign n50680 = n50677 | n50679 ;
  assign n50681 = n66081 & n50680 ;
  assign n81730 = ~n50310 ;
  assign n50682 = n50084 & n81730 ;
  assign n50683 = n49962 | n50084 ;
  assign n81731 = ~n50683 ;
  assign n50684 = n50080 & n81731 ;
  assign n50685 = n50682 | n50684 ;
  assign n50686 = n81659 & n50685 ;
  assign n50687 = n49953 & n81655 ;
  assign n50688 = n50279 & n50687 ;
  assign n50689 = n50686 | n50688 ;
  assign n50690 = n66043 & n50689 ;
  assign n81732 = ~n50079 ;
  assign n50691 = n50078 & n81732 ;
  assign n50692 = n49971 | n50078 ;
  assign n81733 = ~n50692 ;
  assign n50693 = n50307 & n81733 ;
  assign n50694 = n50691 | n50693 ;
  assign n50695 = n81659 & n50694 ;
  assign n50696 = n49961 & n81655 ;
  assign n50697 = n50279 & n50696 ;
  assign n50698 = n50695 | n50697 ;
  assign n50699 = n65960 & n50698 ;
  assign n81734 = ~n50306 ;
  assign n50700 = n50074 & n81734 ;
  assign n50701 = n49980 | n50074 ;
  assign n81735 = ~n50701 ;
  assign n50702 = n50070 & n81735 ;
  assign n50703 = n50700 | n50702 ;
  assign n50704 = n81659 & n50703 ;
  assign n50705 = n49970 & n81655 ;
  assign n50706 = n50279 & n50705 ;
  assign n50707 = n50704 | n50706 ;
  assign n50708 = n65909 & n50707 ;
  assign n81736 = ~n50069 ;
  assign n50709 = n50067 & n81736 ;
  assign n50068 = n49989 | n50067 ;
  assign n81737 = ~n50068 ;
  assign n50710 = n50064 & n81737 ;
  assign n50711 = n50709 | n50710 ;
  assign n50712 = n81659 & n50711 ;
  assign n50713 = n49979 & n81655 ;
  assign n50714 = n50279 & n50713 ;
  assign n50715 = n50712 | n50714 ;
  assign n50716 = n65877 & n50715 ;
  assign n81738 = ~n50302 ;
  assign n50717 = n50063 & n81738 ;
  assign n50718 = n49998 | n50063 ;
  assign n81739 = ~n50718 ;
  assign n50719 = n50059 & n81739 ;
  assign n50720 = n50717 | n50719 ;
  assign n50721 = n81659 & n50720 ;
  assign n50722 = n49988 & n81655 ;
  assign n50723 = n50279 & n50722 ;
  assign n50724 = n50721 | n50723 ;
  assign n50725 = n65820 & n50724 ;
  assign n81740 = ~n50058 ;
  assign n50727 = n50057 & n81740 ;
  assign n50726 = n50006 | n50057 ;
  assign n81741 = ~n50726 ;
  assign n50728 = n50054 & n81741 ;
  assign n50729 = n50727 | n50728 ;
  assign n50730 = n81659 & n50729 ;
  assign n50731 = n49997 & n81655 ;
  assign n50732 = n50279 & n50731 ;
  assign n50733 = n50730 | n50732 ;
  assign n50734 = n65791 & n50733 ;
  assign n81742 = ~n50298 ;
  assign n50736 = n50053 & n81742 ;
  assign n50735 = n50015 | n50053 ;
  assign n81743 = ~n50735 ;
  assign n50737 = n50297 & n81743 ;
  assign n50738 = n50736 | n50737 ;
  assign n50739 = n81659 & n50738 ;
  assign n50740 = n50005 & n81655 ;
  assign n50741 = n50279 & n50740 ;
  assign n50742 = n50739 | n50741 ;
  assign n50743 = n65772 & n50742 ;
  assign n81744 = ~n50048 ;
  assign n50745 = n50047 & n81744 ;
  assign n50744 = n50023 | n50047 ;
  assign n81745 = ~n50744 ;
  assign n50746 = n50044 & n81745 ;
  assign n50747 = n50745 | n50746 ;
  assign n50748 = n81659 & n50747 ;
  assign n50749 = n50014 & n81655 ;
  assign n50750 = n50279 & n50749 ;
  assign n50751 = n50748 | n50750 ;
  assign n50752 = n65746 & n50751 ;
  assign n81746 = ~n50294 ;
  assign n50754 = n50043 & n81746 ;
  assign n50753 = n50039 | n50043 ;
  assign n81747 = ~n50753 ;
  assign n50755 = n50293 & n81747 ;
  assign n50756 = n50754 | n50755 ;
  assign n50757 = n81659 & n50756 ;
  assign n50758 = n50022 & n81655 ;
  assign n50759 = n50279 & n50758 ;
  assign n50760 = n50757 | n50759 ;
  assign n50761 = n65721 & n50760 ;
  assign n50762 = n17792 & n50035 ;
  assign n50763 = n81657 & n50762 ;
  assign n81748 = ~n50763 ;
  assign n50764 = n50293 & n81748 ;
  assign n50765 = n81659 & n50764 ;
  assign n50766 = n50038 & n81655 ;
  assign n50767 = n50279 & n50766 ;
  assign n50768 = n50765 | n50767 ;
  assign n50769 = n65686 & n50768 ;
  assign n50282 = n17792 & n81659 ;
  assign n50770 = x64 & n81659 ;
  assign n81749 = ~n50770 ;
  assign n50771 = x17 & n81749 ;
  assign n50772 = n50282 | n50771 ;
  assign n50786 = n65670 & n50772 ;
  assign n50777 = n50278 | n50776 ;
  assign n50778 = n81655 & n50777 ;
  assign n81750 = ~n50778 ;
  assign n50779 = x64 & n81750 ;
  assign n81751 = ~n50779 ;
  assign n50780 = x17 & n81751 ;
  assign n50781 = n50282 | n50780 ;
  assign n50782 = x65 & n50781 ;
  assign n50783 = x65 | n50282 ;
  assign n50784 = n50780 | n50783 ;
  assign n81752 = ~n50782 ;
  assign n50785 = n81752 & n50784 ;
  assign n50787 = n18543 | n50785 ;
  assign n81753 = ~n50786 ;
  assign n50788 = n81753 & n50787 ;
  assign n81754 = ~n50767 ;
  assign n50789 = x66 & n81754 ;
  assign n81755 = ~n50765 ;
  assign n50790 = n81755 & n50789 ;
  assign n50791 = n50769 | n50790 ;
  assign n50792 = n50788 | n50791 ;
  assign n81756 = ~n50769 ;
  assign n50793 = n81756 & n50792 ;
  assign n81757 = ~n50759 ;
  assign n50794 = x67 & n81757 ;
  assign n81758 = ~n50757 ;
  assign n50795 = n81758 & n50794 ;
  assign n50796 = n50761 | n50795 ;
  assign n50797 = n50793 | n50796 ;
  assign n81759 = ~n50761 ;
  assign n50798 = n81759 & n50797 ;
  assign n81760 = ~n50750 ;
  assign n50799 = x68 & n81760 ;
  assign n81761 = ~n50748 ;
  assign n50800 = n81761 & n50799 ;
  assign n50801 = n50752 | n50800 ;
  assign n50802 = n50798 | n50801 ;
  assign n81762 = ~n50752 ;
  assign n50803 = n81762 & n50802 ;
  assign n81763 = ~n50741 ;
  assign n50804 = x69 & n81763 ;
  assign n81764 = ~n50739 ;
  assign n50805 = n81764 & n50804 ;
  assign n50806 = n50743 | n50805 ;
  assign n50807 = n50803 | n50806 ;
  assign n81765 = ~n50743 ;
  assign n50808 = n81765 & n50807 ;
  assign n81766 = ~n50732 ;
  assign n50809 = x70 & n81766 ;
  assign n81767 = ~n50730 ;
  assign n50810 = n81767 & n50809 ;
  assign n50811 = n50734 | n50810 ;
  assign n50813 = n50808 | n50811 ;
  assign n81768 = ~n50734 ;
  assign n50814 = n81768 & n50813 ;
  assign n81769 = ~n50723 ;
  assign n50815 = x71 & n81769 ;
  assign n81770 = ~n50721 ;
  assign n50816 = n81770 & n50815 ;
  assign n50817 = n50725 | n50816 ;
  assign n50818 = n50814 | n50817 ;
  assign n81771 = ~n50725 ;
  assign n50819 = n81771 & n50818 ;
  assign n81772 = ~n50714 ;
  assign n50820 = x72 & n81772 ;
  assign n81773 = ~n50712 ;
  assign n50821 = n81773 & n50820 ;
  assign n50822 = n50716 | n50821 ;
  assign n50824 = n50819 | n50822 ;
  assign n81774 = ~n50716 ;
  assign n50825 = n81774 & n50824 ;
  assign n81775 = ~n50706 ;
  assign n50826 = x73 & n81775 ;
  assign n81776 = ~n50704 ;
  assign n50827 = n81776 & n50826 ;
  assign n50828 = n50708 | n50827 ;
  assign n50829 = n50825 | n50828 ;
  assign n81777 = ~n50708 ;
  assign n50830 = n81777 & n50829 ;
  assign n81778 = ~n50697 ;
  assign n50831 = x74 & n81778 ;
  assign n81779 = ~n50695 ;
  assign n50832 = n81779 & n50831 ;
  assign n50833 = n50699 | n50832 ;
  assign n50835 = n50830 | n50833 ;
  assign n81780 = ~n50699 ;
  assign n50836 = n81780 & n50835 ;
  assign n81781 = ~n50688 ;
  assign n50837 = x75 & n81781 ;
  assign n81782 = ~n50686 ;
  assign n50838 = n81782 & n50837 ;
  assign n50839 = n50690 | n50838 ;
  assign n50840 = n50836 | n50839 ;
  assign n81783 = ~n50690 ;
  assign n50841 = n81783 & n50840 ;
  assign n81784 = ~n50679 ;
  assign n50842 = x76 & n81784 ;
  assign n81785 = ~n50677 ;
  assign n50843 = n81785 & n50842 ;
  assign n50844 = n50681 | n50843 ;
  assign n50846 = n50841 | n50844 ;
  assign n81786 = ~n50681 ;
  assign n50847 = n81786 & n50846 ;
  assign n81787 = ~n50670 ;
  assign n50848 = x77 & n81787 ;
  assign n81788 = ~n50668 ;
  assign n50849 = n81788 & n50848 ;
  assign n50850 = n50672 | n50849 ;
  assign n50851 = n50847 | n50850 ;
  assign n81789 = ~n50672 ;
  assign n50852 = n81789 & n50851 ;
  assign n81790 = ~n50661 ;
  assign n50853 = x78 & n81790 ;
  assign n81791 = ~n50659 ;
  assign n50854 = n81791 & n50853 ;
  assign n50855 = n50663 | n50854 ;
  assign n50857 = n50852 | n50855 ;
  assign n81792 = ~n50663 ;
  assign n50858 = n81792 & n50857 ;
  assign n81793 = ~n50652 ;
  assign n50859 = x79 & n81793 ;
  assign n81794 = ~n50650 ;
  assign n50860 = n81794 & n50859 ;
  assign n50861 = n50654 | n50860 ;
  assign n50862 = n50858 | n50861 ;
  assign n81795 = ~n50654 ;
  assign n50863 = n81795 & n50862 ;
  assign n81796 = ~n50643 ;
  assign n50864 = x80 & n81796 ;
  assign n81797 = ~n50641 ;
  assign n50865 = n81797 & n50864 ;
  assign n50866 = n50645 | n50865 ;
  assign n50868 = n50863 | n50866 ;
  assign n81798 = ~n50645 ;
  assign n50869 = n81798 & n50868 ;
  assign n81799 = ~n50634 ;
  assign n50870 = x81 & n81799 ;
  assign n81800 = ~n50632 ;
  assign n50871 = n81800 & n50870 ;
  assign n50872 = n50636 | n50871 ;
  assign n50873 = n50869 | n50872 ;
  assign n81801 = ~n50636 ;
  assign n50874 = n81801 & n50873 ;
  assign n81802 = ~n50625 ;
  assign n50875 = x82 & n81802 ;
  assign n81803 = ~n50623 ;
  assign n50876 = n81803 & n50875 ;
  assign n50877 = n50627 | n50876 ;
  assign n50879 = n50874 | n50877 ;
  assign n81804 = ~n50627 ;
  assign n50880 = n81804 & n50879 ;
  assign n81805 = ~n50616 ;
  assign n50881 = x83 & n81805 ;
  assign n81806 = ~n50614 ;
  assign n50882 = n81806 & n50881 ;
  assign n50883 = n50618 | n50882 ;
  assign n50884 = n50880 | n50883 ;
  assign n81807 = ~n50618 ;
  assign n50885 = n81807 & n50884 ;
  assign n81808 = ~n50607 ;
  assign n50886 = x84 & n81808 ;
  assign n81809 = ~n50605 ;
  assign n50887 = n81809 & n50886 ;
  assign n50888 = n50609 | n50887 ;
  assign n50890 = n50885 | n50888 ;
  assign n81810 = ~n50609 ;
  assign n50891 = n81810 & n50890 ;
  assign n81811 = ~n50598 ;
  assign n50892 = x85 & n81811 ;
  assign n81812 = ~n50596 ;
  assign n50893 = n81812 & n50892 ;
  assign n50894 = n50600 | n50893 ;
  assign n50895 = n50891 | n50894 ;
  assign n81813 = ~n50600 ;
  assign n50896 = n81813 & n50895 ;
  assign n81814 = ~n50589 ;
  assign n50897 = x86 & n81814 ;
  assign n81815 = ~n50587 ;
  assign n50898 = n81815 & n50897 ;
  assign n50899 = n50591 | n50898 ;
  assign n50901 = n50896 | n50899 ;
  assign n81816 = ~n50591 ;
  assign n50902 = n81816 & n50901 ;
  assign n81817 = ~n50580 ;
  assign n50903 = x87 & n81817 ;
  assign n81818 = ~n50578 ;
  assign n50904 = n81818 & n50903 ;
  assign n50905 = n50582 | n50904 ;
  assign n50906 = n50902 | n50905 ;
  assign n81819 = ~n50582 ;
  assign n50907 = n81819 & n50906 ;
  assign n81820 = ~n50571 ;
  assign n50908 = x88 & n81820 ;
  assign n81821 = ~n50569 ;
  assign n50909 = n81821 & n50908 ;
  assign n50910 = n50573 | n50909 ;
  assign n50912 = n50907 | n50910 ;
  assign n81822 = ~n50573 ;
  assign n50913 = n81822 & n50912 ;
  assign n81823 = ~n50563 ;
  assign n50914 = x89 & n81823 ;
  assign n81824 = ~n50561 ;
  assign n50915 = n81824 & n50914 ;
  assign n50916 = n50565 | n50915 ;
  assign n50917 = n50913 | n50916 ;
  assign n81825 = ~n50565 ;
  assign n50918 = n81825 & n50917 ;
  assign n81826 = ~n50554 ;
  assign n50919 = x90 & n81826 ;
  assign n81827 = ~n50552 ;
  assign n50920 = n81827 & n50919 ;
  assign n50921 = n50556 | n50920 ;
  assign n50923 = n50918 | n50921 ;
  assign n81828 = ~n50556 ;
  assign n50924 = n81828 & n50923 ;
  assign n81829 = ~n50545 ;
  assign n50925 = x91 & n81829 ;
  assign n81830 = ~n50543 ;
  assign n50926 = n81830 & n50925 ;
  assign n50927 = n50547 | n50926 ;
  assign n50928 = n50924 | n50927 ;
  assign n81831 = ~n50547 ;
  assign n50929 = n81831 & n50928 ;
  assign n81832 = ~n50536 ;
  assign n50930 = x92 & n81832 ;
  assign n81833 = ~n50534 ;
  assign n50931 = n81833 & n50930 ;
  assign n50932 = n50538 | n50931 ;
  assign n50934 = n50929 | n50932 ;
  assign n81834 = ~n50538 ;
  assign n50935 = n81834 & n50934 ;
  assign n81835 = ~n50528 ;
  assign n50936 = x93 & n81835 ;
  assign n81836 = ~n50526 ;
  assign n50937 = n81836 & n50936 ;
  assign n50938 = n50530 | n50937 ;
  assign n50939 = n50935 | n50938 ;
  assign n81837 = ~n50530 ;
  assign n50940 = n81837 & n50939 ;
  assign n81838 = ~n50519 ;
  assign n50941 = x94 & n81838 ;
  assign n81839 = ~n50517 ;
  assign n50942 = n81839 & n50941 ;
  assign n50943 = n50521 | n50942 ;
  assign n50945 = n50940 | n50943 ;
  assign n81840 = ~n50521 ;
  assign n50946 = n81840 & n50945 ;
  assign n81841 = ~n50510 ;
  assign n50947 = x95 & n81841 ;
  assign n81842 = ~n50508 ;
  assign n50948 = n81842 & n50947 ;
  assign n50949 = n50512 | n50948 ;
  assign n50950 = n50946 | n50949 ;
  assign n81843 = ~n50512 ;
  assign n50951 = n81843 & n50950 ;
  assign n81844 = ~n50501 ;
  assign n50952 = x96 & n81844 ;
  assign n81845 = ~n50499 ;
  assign n50953 = n81845 & n50952 ;
  assign n50954 = n50503 | n50953 ;
  assign n50956 = n50951 | n50954 ;
  assign n81846 = ~n50503 ;
  assign n50957 = n81846 & n50956 ;
  assign n81847 = ~n50492 ;
  assign n50958 = x97 & n81847 ;
  assign n81848 = ~n50490 ;
  assign n50959 = n81848 & n50958 ;
  assign n50960 = n50494 | n50959 ;
  assign n50961 = n50957 | n50960 ;
  assign n81849 = ~n50494 ;
  assign n50962 = n81849 & n50961 ;
  assign n81850 = ~n50483 ;
  assign n50963 = x98 & n81850 ;
  assign n81851 = ~n50481 ;
  assign n50964 = n81851 & n50963 ;
  assign n50965 = n50485 | n50964 ;
  assign n50967 = n50962 | n50965 ;
  assign n81852 = ~n50485 ;
  assign n50968 = n81852 & n50967 ;
  assign n81853 = ~n50474 ;
  assign n50969 = x99 & n81853 ;
  assign n81854 = ~n50472 ;
  assign n50970 = n81854 & n50969 ;
  assign n50971 = n50476 | n50970 ;
  assign n50972 = n50968 | n50971 ;
  assign n81855 = ~n50476 ;
  assign n50973 = n81855 & n50972 ;
  assign n81856 = ~n50465 ;
  assign n50974 = x100 & n81856 ;
  assign n81857 = ~n50463 ;
  assign n50975 = n81857 & n50974 ;
  assign n50976 = n50467 | n50975 ;
  assign n50978 = n50973 | n50976 ;
  assign n81858 = ~n50467 ;
  assign n50979 = n81858 & n50978 ;
  assign n81859 = ~n50457 ;
  assign n50980 = x101 & n81859 ;
  assign n81860 = ~n50455 ;
  assign n50981 = n81860 & n50980 ;
  assign n50982 = n50459 | n50981 ;
  assign n50983 = n50979 | n50982 ;
  assign n81861 = ~n50459 ;
  assign n50984 = n81861 & n50983 ;
  assign n81862 = ~n50448 ;
  assign n50985 = x102 & n81862 ;
  assign n81863 = ~n50446 ;
  assign n50986 = n81863 & n50985 ;
  assign n50987 = n50450 | n50986 ;
  assign n50989 = n50984 | n50987 ;
  assign n81864 = ~n50450 ;
  assign n50990 = n81864 & n50989 ;
  assign n81865 = ~n50439 ;
  assign n50991 = x103 & n81865 ;
  assign n81866 = ~n50437 ;
  assign n50992 = n81866 & n50991 ;
  assign n50993 = n50441 | n50992 ;
  assign n50994 = n50990 | n50993 ;
  assign n81867 = ~n50441 ;
  assign n50995 = n81867 & n50994 ;
  assign n81868 = ~n50430 ;
  assign n50996 = x104 & n81868 ;
  assign n81869 = ~n50428 ;
  assign n50997 = n81869 & n50996 ;
  assign n50998 = n50432 | n50997 ;
  assign n51000 = n50995 | n50998 ;
  assign n81870 = ~n50432 ;
  assign n51001 = n81870 & n51000 ;
  assign n81871 = ~n50421 ;
  assign n51002 = x105 & n81871 ;
  assign n81872 = ~n50419 ;
  assign n51003 = n81872 & n51002 ;
  assign n51004 = n50423 | n51003 ;
  assign n51005 = n51001 | n51004 ;
  assign n81873 = ~n50423 ;
  assign n51006 = n81873 & n51005 ;
  assign n81874 = ~n50412 ;
  assign n51007 = x106 & n81874 ;
  assign n81875 = ~n50410 ;
  assign n51008 = n81875 & n51007 ;
  assign n51009 = n50414 | n51008 ;
  assign n51011 = n51006 | n51009 ;
  assign n81876 = ~n50414 ;
  assign n51012 = n81876 & n51011 ;
  assign n81877 = ~n50403 ;
  assign n51013 = x107 & n81877 ;
  assign n81878 = ~n50401 ;
  assign n51014 = n81878 & n51013 ;
  assign n51015 = n50405 | n51014 ;
  assign n51016 = n51012 | n51015 ;
  assign n81879 = ~n50405 ;
  assign n51017 = n81879 & n51016 ;
  assign n81880 = ~n50394 ;
  assign n51018 = x108 & n81880 ;
  assign n81881 = ~n50392 ;
  assign n51019 = n81881 & n51018 ;
  assign n51020 = n50396 | n51019 ;
  assign n51022 = n51017 | n51020 ;
  assign n81882 = ~n50396 ;
  assign n51023 = n81882 & n51022 ;
  assign n81883 = ~n50385 ;
  assign n51024 = x109 & n81883 ;
  assign n81884 = ~n50383 ;
  assign n51025 = n81884 & n51024 ;
  assign n51026 = n50387 | n51025 ;
  assign n51027 = n51023 | n51026 ;
  assign n81885 = ~n50387 ;
  assign n51028 = n81885 & n51027 ;
  assign n81886 = ~n50288 ;
  assign n51029 = x110 & n81886 ;
  assign n81887 = ~n50286 ;
  assign n51030 = n81887 & n51029 ;
  assign n51031 = n50290 | n51030 ;
  assign n51033 = n51028 | n51031 ;
  assign n81888 = ~n50290 ;
  assign n51034 = n81888 & n51033 ;
  assign n51045 = n71633 & n51044 ;
  assign n81889 = ~n51043 ;
  assign n51046 = x111 & n81889 ;
  assign n81890 = ~n51041 ;
  assign n51047 = n81890 & n51046 ;
  assign n51048 = n66858 | n51047 ;
  assign n51049 = n51045 | n51048 ;
  assign n51051 = n51034 | n51049 ;
  assign n81891 = ~n51050 ;
  assign n51052 = n81891 & n51051 ;
  assign n51180 = n50290 | n51047 ;
  assign n51181 = n51045 | n51180 ;
  assign n81892 = ~n51181 ;
  assign n51182 = n51033 & n81892 ;
  assign n51055 = x65 & n50772 ;
  assign n81893 = ~n51055 ;
  assign n51056 = n50784 & n81893 ;
  assign n51057 = n18543 | n51056 ;
  assign n51058 = n81753 & n51057 ;
  assign n51059 = n50791 | n51058 ;
  assign n51060 = n81756 & n51059 ;
  assign n51062 = n50796 | n51060 ;
  assign n51063 = n81759 & n51062 ;
  assign n51065 = n50801 | n51063 ;
  assign n51066 = n81762 & n51065 ;
  assign n51067 = n50806 | n51066 ;
  assign n51069 = n81765 & n51067 ;
  assign n51070 = n50811 | n51069 ;
  assign n51071 = n81768 & n51070 ;
  assign n51072 = n50817 | n51071 ;
  assign n51074 = n81771 & n51072 ;
  assign n51075 = n50822 | n51074 ;
  assign n51076 = n81774 & n51075 ;
  assign n51077 = n50828 | n51076 ;
  assign n51079 = n81777 & n51077 ;
  assign n51080 = n50833 | n51079 ;
  assign n51081 = n81780 & n51080 ;
  assign n51082 = n50839 | n51081 ;
  assign n51084 = n81783 & n51082 ;
  assign n51085 = n50844 | n51084 ;
  assign n51086 = n81786 & n51085 ;
  assign n51087 = n50850 | n51086 ;
  assign n51089 = n81789 & n51087 ;
  assign n51090 = n50855 | n51089 ;
  assign n51091 = n81792 & n51090 ;
  assign n51092 = n50861 | n51091 ;
  assign n51094 = n81795 & n51092 ;
  assign n51095 = n50866 | n51094 ;
  assign n51096 = n81798 & n51095 ;
  assign n51097 = n50872 | n51096 ;
  assign n51099 = n81801 & n51097 ;
  assign n51100 = n50877 | n51099 ;
  assign n51101 = n81804 & n51100 ;
  assign n51102 = n50883 | n51101 ;
  assign n51104 = n81807 & n51102 ;
  assign n51105 = n50888 | n51104 ;
  assign n51106 = n81810 & n51105 ;
  assign n51107 = n50894 | n51106 ;
  assign n51109 = n81813 & n51107 ;
  assign n51110 = n50899 | n51109 ;
  assign n51111 = n81816 & n51110 ;
  assign n51112 = n50905 | n51111 ;
  assign n51114 = n81819 & n51112 ;
  assign n51115 = n50910 | n51114 ;
  assign n51116 = n81822 & n51115 ;
  assign n51117 = n50916 | n51116 ;
  assign n51119 = n81825 & n51117 ;
  assign n51120 = n50921 | n51119 ;
  assign n51121 = n81828 & n51120 ;
  assign n51122 = n50927 | n51121 ;
  assign n51124 = n81831 & n51122 ;
  assign n51125 = n50932 | n51124 ;
  assign n51126 = n81834 & n51125 ;
  assign n51127 = n50938 | n51126 ;
  assign n51129 = n81837 & n51127 ;
  assign n51130 = n50943 | n51129 ;
  assign n51131 = n81840 & n51130 ;
  assign n51132 = n50949 | n51131 ;
  assign n51134 = n81843 & n51132 ;
  assign n51135 = n50954 | n51134 ;
  assign n51136 = n81846 & n51135 ;
  assign n51137 = n50960 | n51136 ;
  assign n51139 = n81849 & n51137 ;
  assign n51140 = n50965 | n51139 ;
  assign n51141 = n81852 & n51140 ;
  assign n51142 = n50971 | n51141 ;
  assign n51144 = n81855 & n51142 ;
  assign n51145 = n50976 | n51144 ;
  assign n51146 = n81858 & n51145 ;
  assign n51147 = n50982 | n51146 ;
  assign n51149 = n81861 & n51147 ;
  assign n51150 = n50987 | n51149 ;
  assign n51151 = n81864 & n51150 ;
  assign n51152 = n50993 | n51151 ;
  assign n51154 = n81867 & n51152 ;
  assign n51155 = n50998 | n51154 ;
  assign n51156 = n81870 & n51155 ;
  assign n51157 = n51004 | n51156 ;
  assign n51159 = n81873 & n51157 ;
  assign n51160 = n51009 | n51159 ;
  assign n51161 = n81876 & n51160 ;
  assign n51162 = n51015 | n51161 ;
  assign n51164 = n81879 & n51162 ;
  assign n51165 = n51020 | n51164 ;
  assign n51166 = n81882 & n51165 ;
  assign n51167 = n51026 | n51166 ;
  assign n51173 = n81885 & n51167 ;
  assign n51174 = n51031 | n51173 ;
  assign n51175 = n81888 & n51174 ;
  assign n51183 = n51045 | n51047 ;
  assign n81894 = ~n51175 ;
  assign n51184 = n81894 & n51183 ;
  assign n51185 = n51182 | n51184 ;
  assign n81895 = ~n51052 ;
  assign n51186 = n81895 & n51185 ;
  assign n51176 = n51049 | n51175 ;
  assign n51187 = n18047 & n51044 ;
  assign n51188 = n51176 & n51187 ;
  assign n51189 = n51186 | n51188 ;
  assign n51190 = n71645 & n51189 ;
  assign n81896 = ~n51188 ;
  assign n51837 = x112 & n81896 ;
  assign n81897 = ~n51186 ;
  assign n51838 = n81897 & n51837 ;
  assign n51839 = n51190 | n51838 ;
  assign n81898 = ~n51028 ;
  assign n51032 = n81898 & n51031 ;
  assign n51169 = n50387 | n51031 ;
  assign n81899 = ~n51169 ;
  assign n51170 = n51167 & n81899 ;
  assign n51171 = n51032 | n51170 ;
  assign n51172 = n81895 & n51171 ;
  assign n51177 = n50289 & n81891 ;
  assign n51178 = n51176 & n51177 ;
  assign n51179 = n51172 | n51178 ;
  assign n51191 = n71633 & n51179 ;
  assign n81900 = ~n51166 ;
  assign n51168 = n51026 & n81900 ;
  assign n51192 = n50396 | n51026 ;
  assign n81901 = ~n51192 ;
  assign n51193 = n51022 & n81901 ;
  assign n51194 = n51168 | n51193 ;
  assign n51195 = n81895 & n51194 ;
  assign n51196 = n50386 & n81891 ;
  assign n51197 = n51176 & n51196 ;
  assign n51198 = n51195 | n51197 ;
  assign n51199 = n71253 & n51198 ;
  assign n81902 = ~n51197 ;
  assign n51825 = x110 & n81902 ;
  assign n81903 = ~n51195 ;
  assign n51826 = n81903 & n51825 ;
  assign n51827 = n51199 | n51826 ;
  assign n81904 = ~n51017 ;
  assign n51021 = n81904 & n51020 ;
  assign n51200 = n50405 | n51020 ;
  assign n81905 = ~n51200 ;
  assign n51201 = n51162 & n81905 ;
  assign n51202 = n51021 | n51201 ;
  assign n51203 = n81895 & n51202 ;
  assign n51204 = n50395 & n81891 ;
  assign n51205 = n51176 & n51204 ;
  assign n51206 = n51203 | n51205 ;
  assign n51207 = n70935 & n51206 ;
  assign n81906 = ~n51161 ;
  assign n51163 = n51015 & n81906 ;
  assign n51208 = n50414 | n51015 ;
  assign n81907 = ~n51208 ;
  assign n51209 = n51011 & n81907 ;
  assign n51210 = n51163 | n51209 ;
  assign n51211 = n81895 & n51210 ;
  assign n51212 = n50404 & n81891 ;
  assign n51213 = n51176 & n51212 ;
  assign n51214 = n51211 | n51213 ;
  assign n51215 = n70927 & n51214 ;
  assign n81908 = ~n51213 ;
  assign n51813 = x108 & n81908 ;
  assign n81909 = ~n51211 ;
  assign n51814 = n81909 & n51813 ;
  assign n51815 = n51215 | n51814 ;
  assign n81910 = ~n51006 ;
  assign n51010 = n81910 & n51009 ;
  assign n51216 = n50423 | n51009 ;
  assign n81911 = ~n51216 ;
  assign n51217 = n51157 & n81911 ;
  assign n51218 = n51010 | n51217 ;
  assign n51219 = n81895 & n51218 ;
  assign n51220 = n50413 & n81891 ;
  assign n51221 = n51176 & n51220 ;
  assign n51222 = n51219 | n51221 ;
  assign n51223 = n70609 & n51222 ;
  assign n81912 = ~n51156 ;
  assign n51158 = n51004 & n81912 ;
  assign n51224 = n50432 | n51004 ;
  assign n81913 = ~n51224 ;
  assign n51225 = n51000 & n81913 ;
  assign n51226 = n51158 | n51225 ;
  assign n51227 = n81895 & n51226 ;
  assign n51228 = n50422 & n81891 ;
  assign n51229 = n51176 & n51228 ;
  assign n51230 = n51227 | n51229 ;
  assign n51231 = n70276 & n51230 ;
  assign n81914 = ~n51229 ;
  assign n51801 = x106 & n81914 ;
  assign n81915 = ~n51227 ;
  assign n51802 = n81915 & n51801 ;
  assign n51803 = n51231 | n51802 ;
  assign n81916 = ~n50995 ;
  assign n50999 = n81916 & n50998 ;
  assign n51232 = n50441 | n50998 ;
  assign n81917 = ~n51232 ;
  assign n51233 = n51152 & n81917 ;
  assign n51234 = n50999 | n51233 ;
  assign n51235 = n81895 & n51234 ;
  assign n51236 = n50431 & n81891 ;
  assign n51237 = n51176 & n51236 ;
  assign n51238 = n51235 | n51237 ;
  assign n51239 = n70176 & n51238 ;
  assign n81918 = ~n51151 ;
  assign n51153 = n50993 & n81918 ;
  assign n51240 = n50450 | n50993 ;
  assign n81919 = ~n51240 ;
  assign n51241 = n50989 & n81919 ;
  assign n51242 = n51153 | n51241 ;
  assign n51243 = n81895 & n51242 ;
  assign n51244 = n50440 & n81891 ;
  assign n51245 = n51176 & n51244 ;
  assign n51246 = n51243 | n51245 ;
  assign n51247 = n69857 & n51246 ;
  assign n81920 = ~n51245 ;
  assign n51789 = x104 & n81920 ;
  assign n81921 = ~n51243 ;
  assign n51790 = n81921 & n51789 ;
  assign n51791 = n51247 | n51790 ;
  assign n81922 = ~n50984 ;
  assign n50988 = n81922 & n50987 ;
  assign n51248 = n50459 | n50987 ;
  assign n81923 = ~n51248 ;
  assign n51249 = n51147 & n81923 ;
  assign n51250 = n50988 | n51249 ;
  assign n51251 = n81895 & n51250 ;
  assign n51252 = n50449 & n81891 ;
  assign n51253 = n51176 & n51252 ;
  assign n51254 = n51251 | n51253 ;
  assign n51255 = n69656 & n51254 ;
  assign n81924 = ~n51146 ;
  assign n51148 = n50982 & n81924 ;
  assign n51256 = n50467 | n50982 ;
  assign n81925 = ~n51256 ;
  assign n51257 = n50978 & n81925 ;
  assign n51258 = n51148 | n51257 ;
  assign n51259 = n81895 & n51258 ;
  assign n51260 = n50458 & n81891 ;
  assign n51261 = n51176 & n51260 ;
  assign n51262 = n51259 | n51261 ;
  assign n51263 = n69528 & n51262 ;
  assign n81926 = ~n51261 ;
  assign n51777 = x102 & n81926 ;
  assign n81927 = ~n51259 ;
  assign n51778 = n81927 & n51777 ;
  assign n51779 = n51263 | n51778 ;
  assign n81928 = ~n50973 ;
  assign n50977 = n81928 & n50976 ;
  assign n51264 = n50476 | n50976 ;
  assign n81929 = ~n51264 ;
  assign n51265 = n51142 & n81929 ;
  assign n51266 = n50977 | n51265 ;
  assign n51267 = n81895 & n51266 ;
  assign n51268 = n50466 & n81891 ;
  assign n51269 = n51176 & n51268 ;
  assign n51270 = n51267 | n51269 ;
  assign n51271 = n69261 & n51270 ;
  assign n81930 = ~n51141 ;
  assign n51143 = n50971 & n81930 ;
  assign n51272 = n50485 | n50971 ;
  assign n81931 = ~n51272 ;
  assign n51273 = n50967 & n81931 ;
  assign n51274 = n51143 | n51273 ;
  assign n51275 = n81895 & n51274 ;
  assign n51276 = n50475 & n81891 ;
  assign n51277 = n51176 & n51276 ;
  assign n51278 = n51275 | n51277 ;
  assign n51279 = n69075 & n51278 ;
  assign n81932 = ~n51277 ;
  assign n51765 = x100 & n81932 ;
  assign n81933 = ~n51275 ;
  assign n51766 = n81933 & n51765 ;
  assign n51767 = n51279 | n51766 ;
  assign n81934 = ~n50962 ;
  assign n50966 = n81934 & n50965 ;
  assign n51280 = n50494 | n50965 ;
  assign n81935 = ~n51280 ;
  assign n51281 = n51137 & n81935 ;
  assign n51282 = n50966 | n51281 ;
  assign n51283 = n81895 & n51282 ;
  assign n51284 = n50484 & n81891 ;
  assign n51285 = n51176 & n51284 ;
  assign n51286 = n51283 | n51285 ;
  assign n51287 = n68993 & n51286 ;
  assign n81936 = ~n51136 ;
  assign n51138 = n50960 & n81936 ;
  assign n51288 = n50503 | n50960 ;
  assign n81937 = ~n51288 ;
  assign n51289 = n50956 & n81937 ;
  assign n51290 = n51138 | n51289 ;
  assign n51291 = n81895 & n51290 ;
  assign n51292 = n50493 & n81891 ;
  assign n51293 = n51176 & n51292 ;
  assign n51294 = n51291 | n51293 ;
  assign n51295 = n68716 & n51294 ;
  assign n81938 = ~n51293 ;
  assign n51753 = x98 & n81938 ;
  assign n81939 = ~n51291 ;
  assign n51754 = n81939 & n51753 ;
  assign n51755 = n51295 | n51754 ;
  assign n81940 = ~n50951 ;
  assign n50955 = n81940 & n50954 ;
  assign n51296 = n50512 | n50954 ;
  assign n81941 = ~n51296 ;
  assign n51297 = n51132 & n81941 ;
  assign n51298 = n50955 | n51297 ;
  assign n51299 = n81895 & n51298 ;
  assign n51300 = n50502 & n81891 ;
  assign n51301 = n51176 & n51300 ;
  assign n51302 = n51299 | n51301 ;
  assign n51303 = n68545 & n51302 ;
  assign n81942 = ~n51131 ;
  assign n51133 = n50949 & n81942 ;
  assign n51304 = n50521 | n50949 ;
  assign n81943 = ~n51304 ;
  assign n51305 = n50945 & n81943 ;
  assign n51306 = n51133 | n51305 ;
  assign n51307 = n81895 & n51306 ;
  assign n51308 = n50511 & n81891 ;
  assign n51309 = n51176 & n51308 ;
  assign n51310 = n51307 | n51309 ;
  assign n51311 = n68438 & n51310 ;
  assign n81944 = ~n51309 ;
  assign n51741 = x96 & n81944 ;
  assign n81945 = ~n51307 ;
  assign n51742 = n81945 & n51741 ;
  assign n51743 = n51311 | n51742 ;
  assign n81946 = ~n50940 ;
  assign n50944 = n81946 & n50943 ;
  assign n51312 = n50530 | n50943 ;
  assign n81947 = ~n51312 ;
  assign n51313 = n51127 & n81947 ;
  assign n51314 = n50944 | n51313 ;
  assign n51315 = n81895 & n51314 ;
  assign n51316 = n50520 & n81891 ;
  assign n51317 = n51176 & n51316 ;
  assign n51318 = n51315 | n51317 ;
  assign n51319 = n68214 & n51318 ;
  assign n81948 = ~n51126 ;
  assign n51128 = n50938 & n81948 ;
  assign n51320 = n50538 | n50938 ;
  assign n81949 = ~n51320 ;
  assign n51321 = n50934 & n81949 ;
  assign n51322 = n51128 | n51321 ;
  assign n51323 = n81895 & n51322 ;
  assign n51324 = n50529 & n81891 ;
  assign n51325 = n51176 & n51324 ;
  assign n51326 = n51323 | n51325 ;
  assign n51327 = n68058 & n51326 ;
  assign n81950 = ~n51325 ;
  assign n51729 = x94 & n81950 ;
  assign n81951 = ~n51323 ;
  assign n51730 = n81951 & n51729 ;
  assign n51731 = n51327 | n51730 ;
  assign n81952 = ~n50929 ;
  assign n50933 = n81952 & n50932 ;
  assign n51328 = n50547 | n50932 ;
  assign n81953 = ~n51328 ;
  assign n51329 = n51122 & n81953 ;
  assign n51330 = n50933 | n51329 ;
  assign n51331 = n81895 & n51330 ;
  assign n51332 = n50537 & n81891 ;
  assign n51333 = n51176 & n51332 ;
  assign n51334 = n51331 | n51333 ;
  assign n51335 = n67986 & n51334 ;
  assign n81954 = ~n51121 ;
  assign n51123 = n50927 & n81954 ;
  assign n51336 = n50556 | n50927 ;
  assign n81955 = ~n51336 ;
  assign n51337 = n50923 & n81955 ;
  assign n51338 = n51123 | n51337 ;
  assign n51339 = n81895 & n51338 ;
  assign n51340 = n50546 & n81891 ;
  assign n51341 = n51176 & n51340 ;
  assign n51342 = n51339 | n51341 ;
  assign n51343 = n67763 & n51342 ;
  assign n81956 = ~n51341 ;
  assign n51717 = x92 & n81956 ;
  assign n81957 = ~n51339 ;
  assign n51718 = n81957 & n51717 ;
  assign n51719 = n51343 | n51718 ;
  assign n81958 = ~n50918 ;
  assign n50922 = n81958 & n50921 ;
  assign n51344 = n50565 | n50921 ;
  assign n81959 = ~n51344 ;
  assign n51345 = n51117 & n81959 ;
  assign n51346 = n50922 | n51345 ;
  assign n51347 = n81895 & n51346 ;
  assign n51348 = n50555 & n81891 ;
  assign n51349 = n51176 & n51348 ;
  assign n51350 = n51347 | n51349 ;
  assign n51351 = n67622 & n51350 ;
  assign n81960 = ~n51116 ;
  assign n51118 = n50916 & n81960 ;
  assign n51352 = n50573 | n50916 ;
  assign n81961 = ~n51352 ;
  assign n51353 = n50912 & n81961 ;
  assign n51354 = n51118 | n51353 ;
  assign n51355 = n81895 & n51354 ;
  assign n51356 = n50564 & n81891 ;
  assign n51357 = n51176 & n51356 ;
  assign n51358 = n51355 | n51357 ;
  assign n51359 = n67531 & n51358 ;
  assign n81962 = ~n51357 ;
  assign n51705 = x90 & n81962 ;
  assign n81963 = ~n51355 ;
  assign n51706 = n81963 & n51705 ;
  assign n51707 = n51359 | n51706 ;
  assign n81964 = ~n50907 ;
  assign n50911 = n81964 & n50910 ;
  assign n51360 = n50582 | n50910 ;
  assign n81965 = ~n51360 ;
  assign n51361 = n51112 & n81965 ;
  assign n51362 = n50911 | n51361 ;
  assign n51363 = n81895 & n51362 ;
  assign n51364 = n50572 & n81891 ;
  assign n51365 = n51176 & n51364 ;
  assign n51366 = n51363 | n51365 ;
  assign n51367 = n67348 & n51366 ;
  assign n81966 = ~n51111 ;
  assign n51113 = n50905 & n81966 ;
  assign n51368 = n50591 | n50905 ;
  assign n81967 = ~n51368 ;
  assign n51369 = n50901 & n81967 ;
  assign n51370 = n51113 | n51369 ;
  assign n51371 = n81895 & n51370 ;
  assign n51372 = n50581 & n81891 ;
  assign n51373 = n51176 & n51372 ;
  assign n51374 = n51371 | n51373 ;
  assign n51375 = n67222 & n51374 ;
  assign n81968 = ~n51373 ;
  assign n51693 = x88 & n81968 ;
  assign n81969 = ~n51371 ;
  assign n51694 = n81969 & n51693 ;
  assign n51695 = n51375 | n51694 ;
  assign n81970 = ~n50896 ;
  assign n50900 = n81970 & n50899 ;
  assign n51376 = n50600 | n50899 ;
  assign n81971 = ~n51376 ;
  assign n51377 = n51107 & n81971 ;
  assign n51378 = n50900 | n51377 ;
  assign n51379 = n81895 & n51378 ;
  assign n51380 = n50590 & n81891 ;
  assign n51381 = n51176 & n51380 ;
  assign n51382 = n51379 | n51381 ;
  assign n51383 = n67164 & n51382 ;
  assign n81972 = ~n51106 ;
  assign n51108 = n50894 & n81972 ;
  assign n51384 = n50609 | n50894 ;
  assign n81973 = ~n51384 ;
  assign n51385 = n50890 & n81973 ;
  assign n51386 = n51108 | n51385 ;
  assign n51387 = n81895 & n51386 ;
  assign n51388 = n50599 & n81891 ;
  assign n51389 = n51176 & n51388 ;
  assign n51390 = n51387 | n51389 ;
  assign n51391 = n66979 & n51390 ;
  assign n81974 = ~n51389 ;
  assign n51681 = x86 & n81974 ;
  assign n81975 = ~n51387 ;
  assign n51682 = n81975 & n51681 ;
  assign n51683 = n51391 | n51682 ;
  assign n81976 = ~n50885 ;
  assign n50889 = n81976 & n50888 ;
  assign n51392 = n50618 | n50888 ;
  assign n81977 = ~n51392 ;
  assign n51393 = n51102 & n81977 ;
  assign n51394 = n50889 | n51393 ;
  assign n51395 = n81895 & n51394 ;
  assign n51396 = n50608 & n81891 ;
  assign n51397 = n51176 & n51396 ;
  assign n51398 = n51395 | n51397 ;
  assign n51399 = n66868 & n51398 ;
  assign n81978 = ~n51101 ;
  assign n51103 = n50883 & n81978 ;
  assign n51400 = n50627 | n50883 ;
  assign n81979 = ~n51400 ;
  assign n51401 = n50879 & n81979 ;
  assign n51402 = n51103 | n51401 ;
  assign n51403 = n81895 & n51402 ;
  assign n51404 = n50617 & n81891 ;
  assign n51405 = n51176 & n51404 ;
  assign n51406 = n51403 | n51405 ;
  assign n51407 = n66797 & n51406 ;
  assign n81980 = ~n51405 ;
  assign n51669 = x84 & n81980 ;
  assign n81981 = ~n51403 ;
  assign n51670 = n81981 & n51669 ;
  assign n51671 = n51407 | n51670 ;
  assign n81982 = ~n50874 ;
  assign n50878 = n81982 & n50877 ;
  assign n51408 = n50636 | n50877 ;
  assign n81983 = ~n51408 ;
  assign n51409 = n51097 & n81983 ;
  assign n51410 = n50878 | n51409 ;
  assign n51411 = n81895 & n51410 ;
  assign n51412 = n50626 & n81891 ;
  assign n51413 = n51176 & n51412 ;
  assign n51414 = n51411 | n51413 ;
  assign n51415 = n66654 & n51414 ;
  assign n81984 = ~n51096 ;
  assign n51098 = n50872 & n81984 ;
  assign n51416 = n50645 | n50872 ;
  assign n81985 = ~n51416 ;
  assign n51417 = n50868 & n81985 ;
  assign n51418 = n51098 | n51417 ;
  assign n51419 = n81895 & n51418 ;
  assign n51420 = n50635 & n81891 ;
  assign n51421 = n51176 & n51420 ;
  assign n51422 = n51419 | n51421 ;
  assign n51423 = n66560 & n51422 ;
  assign n81986 = ~n51421 ;
  assign n51657 = x82 & n81986 ;
  assign n81987 = ~n51419 ;
  assign n51658 = n81987 & n51657 ;
  assign n51659 = n51423 | n51658 ;
  assign n81988 = ~n50863 ;
  assign n50867 = n81988 & n50866 ;
  assign n51424 = n50654 | n50866 ;
  assign n81989 = ~n51424 ;
  assign n51425 = n51092 & n81989 ;
  assign n51426 = n50867 | n51425 ;
  assign n51427 = n81895 & n51426 ;
  assign n51428 = n50644 & n81891 ;
  assign n51429 = n51176 & n51428 ;
  assign n51430 = n51427 | n51429 ;
  assign n51431 = n66505 & n51430 ;
  assign n81990 = ~n51091 ;
  assign n51093 = n50861 & n81990 ;
  assign n51432 = n50663 | n50861 ;
  assign n81991 = ~n51432 ;
  assign n51433 = n50857 & n81991 ;
  assign n51434 = n51093 | n51433 ;
  assign n51435 = n81895 & n51434 ;
  assign n51436 = n50653 & n81891 ;
  assign n51437 = n51176 & n51436 ;
  assign n51438 = n51435 | n51437 ;
  assign n51439 = n66379 & n51438 ;
  assign n81992 = ~n51437 ;
  assign n51645 = x80 & n81992 ;
  assign n81993 = ~n51435 ;
  assign n51646 = n81993 & n51645 ;
  assign n51647 = n51439 | n51646 ;
  assign n81994 = ~n50852 ;
  assign n50856 = n81994 & n50855 ;
  assign n51440 = n50672 | n50855 ;
  assign n81995 = ~n51440 ;
  assign n51441 = n51087 & n81995 ;
  assign n51442 = n50856 | n51441 ;
  assign n51443 = n81895 & n51442 ;
  assign n51444 = n50662 & n81891 ;
  assign n51445 = n51176 & n51444 ;
  assign n51446 = n51443 | n51445 ;
  assign n51447 = n66299 & n51446 ;
  assign n81996 = ~n51086 ;
  assign n51088 = n50850 & n81996 ;
  assign n51448 = n50681 | n50850 ;
  assign n81997 = ~n51448 ;
  assign n51449 = n50846 & n81997 ;
  assign n51450 = n51088 | n51449 ;
  assign n51451 = n81895 & n51450 ;
  assign n51452 = n50671 & n81891 ;
  assign n51453 = n51176 & n51452 ;
  assign n51454 = n51451 | n51453 ;
  assign n51455 = n66244 & n51454 ;
  assign n81998 = ~n51453 ;
  assign n51633 = x78 & n81998 ;
  assign n81999 = ~n51451 ;
  assign n51634 = n81999 & n51633 ;
  assign n51635 = n51455 | n51634 ;
  assign n82000 = ~n50841 ;
  assign n50845 = n82000 & n50844 ;
  assign n51456 = n50690 | n50844 ;
  assign n82001 = ~n51456 ;
  assign n51457 = n51082 & n82001 ;
  assign n51458 = n50845 | n51457 ;
  assign n51459 = n81895 & n51458 ;
  assign n51460 = n50680 & n81891 ;
  assign n51461 = n51176 & n51460 ;
  assign n51462 = n51459 | n51461 ;
  assign n51463 = n66145 & n51462 ;
  assign n82002 = ~n51081 ;
  assign n51083 = n50839 & n82002 ;
  assign n51464 = n50699 | n50839 ;
  assign n82003 = ~n51464 ;
  assign n51465 = n50835 & n82003 ;
  assign n51466 = n51083 | n51465 ;
  assign n51467 = n81895 & n51466 ;
  assign n51468 = n50689 & n81891 ;
  assign n51469 = n51176 & n51468 ;
  assign n51470 = n51467 | n51469 ;
  assign n51471 = n66081 & n51470 ;
  assign n82004 = ~n51469 ;
  assign n51621 = x76 & n82004 ;
  assign n82005 = ~n51467 ;
  assign n51622 = n82005 & n51621 ;
  assign n51623 = n51471 | n51622 ;
  assign n82006 = ~n50830 ;
  assign n50834 = n82006 & n50833 ;
  assign n51472 = n50708 | n50833 ;
  assign n82007 = ~n51472 ;
  assign n51473 = n51077 & n82007 ;
  assign n51474 = n50834 | n51473 ;
  assign n51475 = n81895 & n51474 ;
  assign n51476 = n50698 & n81891 ;
  assign n51477 = n51176 & n51476 ;
  assign n51478 = n51475 | n51477 ;
  assign n51479 = n66043 & n51478 ;
  assign n82008 = ~n51076 ;
  assign n51078 = n50828 & n82008 ;
  assign n51480 = n50716 | n50828 ;
  assign n82009 = ~n51480 ;
  assign n51481 = n50824 & n82009 ;
  assign n51482 = n51078 | n51481 ;
  assign n51483 = n81895 & n51482 ;
  assign n51484 = n50707 & n81891 ;
  assign n51485 = n51176 & n51484 ;
  assign n51486 = n51483 | n51485 ;
  assign n51487 = n65960 & n51486 ;
  assign n82010 = ~n51485 ;
  assign n51609 = x74 & n82010 ;
  assign n82011 = ~n51483 ;
  assign n51610 = n82011 & n51609 ;
  assign n51611 = n51487 | n51610 ;
  assign n82012 = ~n50819 ;
  assign n50823 = n82012 & n50822 ;
  assign n51488 = n50725 | n50822 ;
  assign n82013 = ~n51488 ;
  assign n51489 = n51072 & n82013 ;
  assign n51490 = n50823 | n51489 ;
  assign n51491 = n81895 & n51490 ;
  assign n51492 = n50715 & n81891 ;
  assign n51493 = n51176 & n51492 ;
  assign n51494 = n51491 | n51493 ;
  assign n51495 = n65909 & n51494 ;
  assign n82014 = ~n51071 ;
  assign n51073 = n50817 & n82014 ;
  assign n51496 = n50734 | n50817 ;
  assign n82015 = ~n51496 ;
  assign n51497 = n50813 & n82015 ;
  assign n51498 = n51073 | n51497 ;
  assign n51499 = n81895 & n51498 ;
  assign n51500 = n50724 & n81891 ;
  assign n51501 = n51176 & n51500 ;
  assign n51502 = n51499 | n51501 ;
  assign n51503 = n65877 & n51502 ;
  assign n82016 = ~n51501 ;
  assign n51597 = x72 & n82016 ;
  assign n82017 = ~n51499 ;
  assign n51598 = n82017 & n51597 ;
  assign n51599 = n51503 | n51598 ;
  assign n82018 = ~n50808 ;
  assign n50812 = n82018 & n50811 ;
  assign n51504 = n50743 | n50811 ;
  assign n82019 = ~n51504 ;
  assign n51505 = n51067 & n82019 ;
  assign n51506 = n50812 | n51505 ;
  assign n51507 = n81895 & n51506 ;
  assign n51508 = n50733 & n81891 ;
  assign n51509 = n51176 & n51508 ;
  assign n51510 = n51507 | n51509 ;
  assign n51511 = n65820 & n51510 ;
  assign n82020 = ~n51066 ;
  assign n51068 = n50806 & n82020 ;
  assign n51512 = n50752 | n50806 ;
  assign n82021 = ~n51512 ;
  assign n51513 = n50802 & n82021 ;
  assign n51514 = n51068 | n51513 ;
  assign n51515 = n81895 & n51514 ;
  assign n51516 = n50742 & n81891 ;
  assign n51517 = n51176 & n51516 ;
  assign n51518 = n51515 | n51517 ;
  assign n51519 = n65791 & n51518 ;
  assign n82022 = ~n51517 ;
  assign n51585 = x70 & n82022 ;
  assign n82023 = ~n51515 ;
  assign n51586 = n82023 & n51585 ;
  assign n51587 = n51519 | n51586 ;
  assign n82024 = ~n50798 ;
  assign n51064 = n82024 & n50801 ;
  assign n51520 = n50761 | n50801 ;
  assign n82025 = ~n51520 ;
  assign n51521 = n51062 & n82025 ;
  assign n51522 = n51064 | n51521 ;
  assign n51523 = n81895 & n51522 ;
  assign n51524 = n50751 & n81891 ;
  assign n51525 = n51176 & n51524 ;
  assign n51526 = n51523 | n51525 ;
  assign n51527 = n65772 & n51526 ;
  assign n82026 = ~n51060 ;
  assign n51061 = n50796 & n82026 ;
  assign n51528 = n50769 | n50796 ;
  assign n82027 = ~n51528 ;
  assign n51529 = n51059 & n82027 ;
  assign n51530 = n51061 | n51529 ;
  assign n51531 = n81895 & n51530 ;
  assign n51532 = n50760 & n81891 ;
  assign n51533 = n51176 & n51532 ;
  assign n51534 = n51531 | n51533 ;
  assign n51535 = n65746 & n51534 ;
  assign n82028 = ~n51533 ;
  assign n51574 = x68 & n82028 ;
  assign n82029 = ~n51531 ;
  assign n51575 = n82029 & n51574 ;
  assign n51576 = n51535 | n51575 ;
  assign n82030 = ~n51058 ;
  assign n51537 = n50791 & n82030 ;
  assign n51536 = n50786 | n50791 ;
  assign n82031 = ~n51536 ;
  assign n51538 = n50787 & n82031 ;
  assign n51539 = n51537 | n51538 ;
  assign n51540 = n81895 & n51539 ;
  assign n51541 = n50768 & n81891 ;
  assign n51542 = n51176 & n51541 ;
  assign n51543 = n51540 | n51542 ;
  assign n51544 = n65721 & n51543 ;
  assign n51545 = n18543 & n50784 ;
  assign n51546 = n81893 & n51545 ;
  assign n82032 = ~n51546 ;
  assign n51547 = n50787 & n82032 ;
  assign n51548 = n81895 & n51547 ;
  assign n51549 = n50772 & n81891 ;
  assign n51550 = n51176 & n51549 ;
  assign n51551 = n51548 | n51550 ;
  assign n51552 = n65686 & n51551 ;
  assign n82033 = ~n51550 ;
  assign n51564 = x66 & n82033 ;
  assign n82034 = ~n51548 ;
  assign n51565 = n82034 & n51564 ;
  assign n51566 = n51552 | n51565 ;
  assign n51054 = n18543 & n81895 ;
  assign n51053 = x64 & n81895 ;
  assign n82035 = ~n51053 ;
  assign n51553 = x16 & n82035 ;
  assign n51554 = n51054 | n51553 ;
  assign n51555 = x65 & n51554 ;
  assign n51556 = n81891 & n51176 ;
  assign n82036 = ~n51556 ;
  assign n51557 = n18543 & n82036 ;
  assign n51558 = x65 | n51557 ;
  assign n51559 = n51553 | n51558 ;
  assign n82037 = ~n51555 ;
  assign n51560 = n82037 & n51559 ;
  assign n51562 = n19324 | n51560 ;
  assign n51563 = n65670 & n51554 ;
  assign n82038 = ~n51563 ;
  assign n51567 = n51562 & n82038 ;
  assign n51568 = n51566 | n51567 ;
  assign n82039 = ~n51552 ;
  assign n51569 = n82039 & n51568 ;
  assign n82040 = ~n51542 ;
  assign n51570 = x67 & n82040 ;
  assign n82041 = ~n51540 ;
  assign n51571 = n82041 & n51570 ;
  assign n51572 = n51544 | n51571 ;
  assign n51573 = n51569 | n51572 ;
  assign n82042 = ~n51544 ;
  assign n51577 = n82042 & n51573 ;
  assign n51578 = n51576 | n51577 ;
  assign n82043 = ~n51535 ;
  assign n51579 = n82043 & n51578 ;
  assign n82044 = ~n51525 ;
  assign n51580 = x69 & n82044 ;
  assign n82045 = ~n51523 ;
  assign n51581 = n82045 & n51580 ;
  assign n51582 = n51527 | n51581 ;
  assign n51584 = n51579 | n51582 ;
  assign n82046 = ~n51527 ;
  assign n51589 = n82046 & n51584 ;
  assign n51590 = n51587 | n51589 ;
  assign n82047 = ~n51519 ;
  assign n51591 = n82047 & n51590 ;
  assign n82048 = ~n51509 ;
  assign n51592 = x71 & n82048 ;
  assign n82049 = ~n51507 ;
  assign n51593 = n82049 & n51592 ;
  assign n51594 = n51511 | n51593 ;
  assign n51596 = n51591 | n51594 ;
  assign n82050 = ~n51511 ;
  assign n51601 = n82050 & n51596 ;
  assign n51602 = n51599 | n51601 ;
  assign n82051 = ~n51503 ;
  assign n51603 = n82051 & n51602 ;
  assign n82052 = ~n51493 ;
  assign n51604 = x73 & n82052 ;
  assign n82053 = ~n51491 ;
  assign n51605 = n82053 & n51604 ;
  assign n51606 = n51495 | n51605 ;
  assign n51608 = n51603 | n51606 ;
  assign n82054 = ~n51495 ;
  assign n51613 = n82054 & n51608 ;
  assign n51614 = n51611 | n51613 ;
  assign n82055 = ~n51487 ;
  assign n51615 = n82055 & n51614 ;
  assign n82056 = ~n51477 ;
  assign n51616 = x75 & n82056 ;
  assign n82057 = ~n51475 ;
  assign n51617 = n82057 & n51616 ;
  assign n51618 = n51479 | n51617 ;
  assign n51620 = n51615 | n51618 ;
  assign n82058 = ~n51479 ;
  assign n51625 = n82058 & n51620 ;
  assign n51626 = n51623 | n51625 ;
  assign n82059 = ~n51471 ;
  assign n51627 = n82059 & n51626 ;
  assign n82060 = ~n51461 ;
  assign n51628 = x77 & n82060 ;
  assign n82061 = ~n51459 ;
  assign n51629 = n82061 & n51628 ;
  assign n51630 = n51463 | n51629 ;
  assign n51632 = n51627 | n51630 ;
  assign n82062 = ~n51463 ;
  assign n51637 = n82062 & n51632 ;
  assign n51638 = n51635 | n51637 ;
  assign n82063 = ~n51455 ;
  assign n51639 = n82063 & n51638 ;
  assign n82064 = ~n51445 ;
  assign n51640 = x79 & n82064 ;
  assign n82065 = ~n51443 ;
  assign n51641 = n82065 & n51640 ;
  assign n51642 = n51447 | n51641 ;
  assign n51644 = n51639 | n51642 ;
  assign n82066 = ~n51447 ;
  assign n51649 = n82066 & n51644 ;
  assign n51650 = n51647 | n51649 ;
  assign n82067 = ~n51439 ;
  assign n51651 = n82067 & n51650 ;
  assign n82068 = ~n51429 ;
  assign n51652 = x81 & n82068 ;
  assign n82069 = ~n51427 ;
  assign n51653 = n82069 & n51652 ;
  assign n51654 = n51431 | n51653 ;
  assign n51656 = n51651 | n51654 ;
  assign n82070 = ~n51431 ;
  assign n51661 = n82070 & n51656 ;
  assign n51662 = n51659 | n51661 ;
  assign n82071 = ~n51423 ;
  assign n51663 = n82071 & n51662 ;
  assign n82072 = ~n51413 ;
  assign n51664 = x83 & n82072 ;
  assign n82073 = ~n51411 ;
  assign n51665 = n82073 & n51664 ;
  assign n51666 = n51415 | n51665 ;
  assign n51668 = n51663 | n51666 ;
  assign n82074 = ~n51415 ;
  assign n51673 = n82074 & n51668 ;
  assign n51674 = n51671 | n51673 ;
  assign n82075 = ~n51407 ;
  assign n51675 = n82075 & n51674 ;
  assign n82076 = ~n51397 ;
  assign n51676 = x85 & n82076 ;
  assign n82077 = ~n51395 ;
  assign n51677 = n82077 & n51676 ;
  assign n51678 = n51399 | n51677 ;
  assign n51680 = n51675 | n51678 ;
  assign n82078 = ~n51399 ;
  assign n51685 = n82078 & n51680 ;
  assign n51686 = n51683 | n51685 ;
  assign n82079 = ~n51391 ;
  assign n51687 = n82079 & n51686 ;
  assign n82080 = ~n51381 ;
  assign n51688 = x87 & n82080 ;
  assign n82081 = ~n51379 ;
  assign n51689 = n82081 & n51688 ;
  assign n51690 = n51383 | n51689 ;
  assign n51692 = n51687 | n51690 ;
  assign n82082 = ~n51383 ;
  assign n51697 = n82082 & n51692 ;
  assign n51698 = n51695 | n51697 ;
  assign n82083 = ~n51375 ;
  assign n51699 = n82083 & n51698 ;
  assign n82084 = ~n51365 ;
  assign n51700 = x89 & n82084 ;
  assign n82085 = ~n51363 ;
  assign n51701 = n82085 & n51700 ;
  assign n51702 = n51367 | n51701 ;
  assign n51704 = n51699 | n51702 ;
  assign n82086 = ~n51367 ;
  assign n51709 = n82086 & n51704 ;
  assign n51710 = n51707 | n51709 ;
  assign n82087 = ~n51359 ;
  assign n51711 = n82087 & n51710 ;
  assign n82088 = ~n51349 ;
  assign n51712 = x91 & n82088 ;
  assign n82089 = ~n51347 ;
  assign n51713 = n82089 & n51712 ;
  assign n51714 = n51351 | n51713 ;
  assign n51716 = n51711 | n51714 ;
  assign n82090 = ~n51351 ;
  assign n51721 = n82090 & n51716 ;
  assign n51722 = n51719 | n51721 ;
  assign n82091 = ~n51343 ;
  assign n51723 = n82091 & n51722 ;
  assign n82092 = ~n51333 ;
  assign n51724 = x93 & n82092 ;
  assign n82093 = ~n51331 ;
  assign n51725 = n82093 & n51724 ;
  assign n51726 = n51335 | n51725 ;
  assign n51728 = n51723 | n51726 ;
  assign n82094 = ~n51335 ;
  assign n51733 = n82094 & n51728 ;
  assign n51734 = n51731 | n51733 ;
  assign n82095 = ~n51327 ;
  assign n51735 = n82095 & n51734 ;
  assign n82096 = ~n51317 ;
  assign n51736 = x95 & n82096 ;
  assign n82097 = ~n51315 ;
  assign n51737 = n82097 & n51736 ;
  assign n51738 = n51319 | n51737 ;
  assign n51740 = n51735 | n51738 ;
  assign n82098 = ~n51319 ;
  assign n51745 = n82098 & n51740 ;
  assign n51746 = n51743 | n51745 ;
  assign n82099 = ~n51311 ;
  assign n51747 = n82099 & n51746 ;
  assign n82100 = ~n51301 ;
  assign n51748 = x97 & n82100 ;
  assign n82101 = ~n51299 ;
  assign n51749 = n82101 & n51748 ;
  assign n51750 = n51303 | n51749 ;
  assign n51752 = n51747 | n51750 ;
  assign n82102 = ~n51303 ;
  assign n51757 = n82102 & n51752 ;
  assign n51758 = n51755 | n51757 ;
  assign n82103 = ~n51295 ;
  assign n51759 = n82103 & n51758 ;
  assign n82104 = ~n51285 ;
  assign n51760 = x99 & n82104 ;
  assign n82105 = ~n51283 ;
  assign n51761 = n82105 & n51760 ;
  assign n51762 = n51287 | n51761 ;
  assign n51764 = n51759 | n51762 ;
  assign n82106 = ~n51287 ;
  assign n51769 = n82106 & n51764 ;
  assign n51770 = n51767 | n51769 ;
  assign n82107 = ~n51279 ;
  assign n51771 = n82107 & n51770 ;
  assign n82108 = ~n51269 ;
  assign n51772 = x101 & n82108 ;
  assign n82109 = ~n51267 ;
  assign n51773 = n82109 & n51772 ;
  assign n51774 = n51271 | n51773 ;
  assign n51776 = n51771 | n51774 ;
  assign n82110 = ~n51271 ;
  assign n51781 = n82110 & n51776 ;
  assign n51782 = n51779 | n51781 ;
  assign n82111 = ~n51263 ;
  assign n51783 = n82111 & n51782 ;
  assign n82112 = ~n51253 ;
  assign n51784 = x103 & n82112 ;
  assign n82113 = ~n51251 ;
  assign n51785 = n82113 & n51784 ;
  assign n51786 = n51255 | n51785 ;
  assign n51788 = n51783 | n51786 ;
  assign n82114 = ~n51255 ;
  assign n51793 = n82114 & n51788 ;
  assign n51794 = n51791 | n51793 ;
  assign n82115 = ~n51247 ;
  assign n51795 = n82115 & n51794 ;
  assign n82116 = ~n51237 ;
  assign n51796 = x105 & n82116 ;
  assign n82117 = ~n51235 ;
  assign n51797 = n82117 & n51796 ;
  assign n51798 = n51239 | n51797 ;
  assign n51800 = n51795 | n51798 ;
  assign n82118 = ~n51239 ;
  assign n51805 = n82118 & n51800 ;
  assign n51806 = n51803 | n51805 ;
  assign n82119 = ~n51231 ;
  assign n51807 = n82119 & n51806 ;
  assign n82120 = ~n51221 ;
  assign n51808 = x107 & n82120 ;
  assign n82121 = ~n51219 ;
  assign n51809 = n82121 & n51808 ;
  assign n51810 = n51223 | n51809 ;
  assign n51812 = n51807 | n51810 ;
  assign n82122 = ~n51223 ;
  assign n51817 = n82122 & n51812 ;
  assign n51818 = n51815 | n51817 ;
  assign n82123 = ~n51215 ;
  assign n51819 = n82123 & n51818 ;
  assign n82124 = ~n51205 ;
  assign n51820 = x109 & n82124 ;
  assign n82125 = ~n51203 ;
  assign n51821 = n82125 & n51820 ;
  assign n51822 = n51207 | n51821 ;
  assign n51824 = n51819 | n51822 ;
  assign n82126 = ~n51207 ;
  assign n51829 = n82126 & n51824 ;
  assign n51830 = n51827 | n51829 ;
  assign n82127 = ~n51199 ;
  assign n51831 = n82127 & n51830 ;
  assign n82128 = ~n51178 ;
  assign n51832 = x111 & n82128 ;
  assign n82129 = ~n51172 ;
  assign n51833 = n82129 & n51832 ;
  assign n51834 = n51191 | n51833 ;
  assign n51836 = n51831 | n51834 ;
  assign n82130 = ~n51191 ;
  assign n51840 = n82130 & n51836 ;
  assign n51841 = n51839 | n51840 ;
  assign n82131 = ~n51190 ;
  assign n51842 = n82131 & n51841 ;
  assign n51843 = n279 | n51842 ;
  assign n82132 = ~n51189 ;
  assign n51845 = n82132 & n51843 ;
  assign n82133 = ~n51840 ;
  assign n52594 = n51839 & n82133 ;
  assign n51847 = x64 & n82036 ;
  assign n82134 = ~n51847 ;
  assign n51848 = x16 & n82134 ;
  assign n51849 = n51054 | n51848 ;
  assign n51850 = x65 & n51849 ;
  assign n82135 = ~n51850 ;
  assign n51851 = n51559 & n82135 ;
  assign n51852 = n19324 | n51851 ;
  assign n51853 = n82038 & n51852 ;
  assign n51855 = n51566 | n51853 ;
  assign n51856 = n82039 & n51855 ;
  assign n51857 = n51572 | n51856 ;
  assign n51858 = n82042 & n51857 ;
  assign n51859 = n51576 | n51858 ;
  assign n51860 = n82043 & n51859 ;
  assign n51861 = n51582 | n51860 ;
  assign n51862 = n82046 & n51861 ;
  assign n51863 = n51587 | n51862 ;
  assign n51864 = n82047 & n51863 ;
  assign n51865 = n51594 | n51864 ;
  assign n51866 = n82050 & n51865 ;
  assign n51867 = n51599 | n51866 ;
  assign n51868 = n82051 & n51867 ;
  assign n51869 = n51606 | n51868 ;
  assign n51870 = n82054 & n51869 ;
  assign n51871 = n51611 | n51870 ;
  assign n51872 = n82055 & n51871 ;
  assign n51873 = n51618 | n51872 ;
  assign n51874 = n82058 & n51873 ;
  assign n51875 = n51623 | n51874 ;
  assign n51876 = n82059 & n51875 ;
  assign n51877 = n51630 | n51876 ;
  assign n51878 = n82062 & n51877 ;
  assign n51879 = n51635 | n51878 ;
  assign n51880 = n82063 & n51879 ;
  assign n51881 = n51642 | n51880 ;
  assign n51882 = n82066 & n51881 ;
  assign n51883 = n51647 | n51882 ;
  assign n51884 = n82067 & n51883 ;
  assign n51885 = n51654 | n51884 ;
  assign n51886 = n82070 & n51885 ;
  assign n51887 = n51659 | n51886 ;
  assign n51888 = n82071 & n51887 ;
  assign n51889 = n51666 | n51888 ;
  assign n51890 = n82074 & n51889 ;
  assign n51891 = n51671 | n51890 ;
  assign n51892 = n82075 & n51891 ;
  assign n51893 = n51678 | n51892 ;
  assign n51894 = n82078 & n51893 ;
  assign n51895 = n51683 | n51894 ;
  assign n51896 = n82079 & n51895 ;
  assign n51897 = n51690 | n51896 ;
  assign n51898 = n82082 & n51897 ;
  assign n51899 = n51695 | n51898 ;
  assign n51900 = n82083 & n51899 ;
  assign n51901 = n51702 | n51900 ;
  assign n51902 = n82086 & n51901 ;
  assign n51903 = n51707 | n51902 ;
  assign n51904 = n82087 & n51903 ;
  assign n51905 = n51714 | n51904 ;
  assign n51906 = n82090 & n51905 ;
  assign n51907 = n51719 | n51906 ;
  assign n51908 = n82091 & n51907 ;
  assign n51909 = n51726 | n51908 ;
  assign n51910 = n82094 & n51909 ;
  assign n51911 = n51731 | n51910 ;
  assign n51912 = n82095 & n51911 ;
  assign n51913 = n51738 | n51912 ;
  assign n51914 = n82098 & n51913 ;
  assign n51915 = n51743 | n51914 ;
  assign n51916 = n82099 & n51915 ;
  assign n51917 = n51750 | n51916 ;
  assign n51918 = n82102 & n51917 ;
  assign n51919 = n51755 | n51918 ;
  assign n51920 = n82103 & n51919 ;
  assign n51921 = n51762 | n51920 ;
  assign n51922 = n82106 & n51921 ;
  assign n51923 = n51767 | n51922 ;
  assign n51924 = n82107 & n51923 ;
  assign n51925 = n51774 | n51924 ;
  assign n51926 = n82110 & n51925 ;
  assign n51927 = n51779 | n51926 ;
  assign n51928 = n82111 & n51927 ;
  assign n51929 = n51786 | n51928 ;
  assign n51930 = n82114 & n51929 ;
  assign n51931 = n51791 | n51930 ;
  assign n51932 = n82115 & n51931 ;
  assign n51933 = n51798 | n51932 ;
  assign n51934 = n82118 & n51933 ;
  assign n51935 = n51803 | n51934 ;
  assign n51936 = n82119 & n51935 ;
  assign n51937 = n51810 | n51936 ;
  assign n51938 = n82122 & n51937 ;
  assign n51939 = n51815 | n51938 ;
  assign n51940 = n82123 & n51939 ;
  assign n51941 = n51822 | n51940 ;
  assign n51942 = n82126 & n51941 ;
  assign n51943 = n51827 | n51942 ;
  assign n51945 = n82127 & n51943 ;
  assign n52321 = n51834 | n51945 ;
  assign n52595 = n51191 | n51839 ;
  assign n82136 = ~n52595 ;
  assign n52596 = n52321 & n82136 ;
  assign n52597 = n52594 | n52596 ;
  assign n52598 = n51843 | n52597 ;
  assign n82137 = ~n51845 ;
  assign n52599 = n82137 & n52598 ;
  assign n52607 = n66715 & n52599 ;
  assign n51846 = n51179 & n51843 ;
  assign n51835 = n51199 | n51834 ;
  assign n82138 = ~n51835 ;
  assign n51944 = n82138 & n51943 ;
  assign n82139 = ~n51945 ;
  assign n51946 = n51834 & n82139 ;
  assign n51947 = n51944 | n51946 ;
  assign n51948 = n66715 & n51947 ;
  assign n82140 = ~n51842 ;
  assign n51949 = n82140 & n51948 ;
  assign n51950 = n51846 | n51949 ;
  assign n51951 = n71645 & n51950 ;
  assign n51952 = n51198 & n51843 ;
  assign n51828 = n51207 | n51827 ;
  assign n82141 = ~n51828 ;
  assign n51953 = n51824 & n82141 ;
  assign n82142 = ~n51829 ;
  assign n51954 = n51827 & n82142 ;
  assign n51955 = n51953 | n51954 ;
  assign n51956 = n66715 & n51955 ;
  assign n51957 = n82140 & n51956 ;
  assign n51958 = n51952 | n51957 ;
  assign n51959 = n71633 & n51958 ;
  assign n51960 = n51206 & n51843 ;
  assign n51823 = n51215 | n51822 ;
  assign n82143 = ~n51823 ;
  assign n51961 = n82143 & n51939 ;
  assign n82144 = ~n51940 ;
  assign n51962 = n51822 & n82144 ;
  assign n51963 = n51961 | n51962 ;
  assign n51964 = n66715 & n51963 ;
  assign n51965 = n82140 & n51964 ;
  assign n51966 = n51960 | n51965 ;
  assign n51967 = n71253 & n51966 ;
  assign n51968 = n51214 & n51843 ;
  assign n51816 = n51223 | n51815 ;
  assign n82145 = ~n51816 ;
  assign n51969 = n51812 & n82145 ;
  assign n82146 = ~n51817 ;
  assign n51970 = n51815 & n82146 ;
  assign n51971 = n51969 | n51970 ;
  assign n51972 = n66715 & n51971 ;
  assign n51973 = n82140 & n51972 ;
  assign n51974 = n51968 | n51973 ;
  assign n51975 = n70935 & n51974 ;
  assign n51976 = n51222 & n51843 ;
  assign n51811 = n51231 | n51810 ;
  assign n82147 = ~n51811 ;
  assign n51977 = n82147 & n51935 ;
  assign n82148 = ~n51936 ;
  assign n51978 = n51810 & n82148 ;
  assign n51979 = n51977 | n51978 ;
  assign n51980 = n66715 & n51979 ;
  assign n51981 = n82140 & n51980 ;
  assign n51982 = n51976 | n51981 ;
  assign n51983 = n70927 & n51982 ;
  assign n51984 = n51230 & n51843 ;
  assign n51804 = n51239 | n51803 ;
  assign n82149 = ~n51804 ;
  assign n51985 = n51800 & n82149 ;
  assign n82150 = ~n51805 ;
  assign n51986 = n51803 & n82150 ;
  assign n51987 = n51985 | n51986 ;
  assign n51988 = n66715 & n51987 ;
  assign n51989 = n82140 & n51988 ;
  assign n51990 = n51984 | n51989 ;
  assign n51991 = n70609 & n51990 ;
  assign n51992 = n51238 & n51843 ;
  assign n51799 = n51247 | n51798 ;
  assign n82151 = ~n51799 ;
  assign n51993 = n82151 & n51931 ;
  assign n82152 = ~n51932 ;
  assign n51994 = n51798 & n82152 ;
  assign n51995 = n51993 | n51994 ;
  assign n51996 = n66715 & n51995 ;
  assign n51997 = n82140 & n51996 ;
  assign n51998 = n51992 | n51997 ;
  assign n51999 = n70276 & n51998 ;
  assign n52000 = n51246 & n51843 ;
  assign n51792 = n51255 | n51791 ;
  assign n82153 = ~n51792 ;
  assign n52001 = n51788 & n82153 ;
  assign n82154 = ~n51793 ;
  assign n52002 = n51791 & n82154 ;
  assign n52003 = n52001 | n52002 ;
  assign n52004 = n66715 & n52003 ;
  assign n52005 = n82140 & n52004 ;
  assign n52006 = n52000 | n52005 ;
  assign n52007 = n70176 & n52006 ;
  assign n52008 = n51254 & n51843 ;
  assign n51787 = n51263 | n51786 ;
  assign n82155 = ~n51787 ;
  assign n52009 = n82155 & n51927 ;
  assign n82156 = ~n51928 ;
  assign n52010 = n51786 & n82156 ;
  assign n52011 = n52009 | n52010 ;
  assign n52012 = n66715 & n52011 ;
  assign n52013 = n82140 & n52012 ;
  assign n52014 = n52008 | n52013 ;
  assign n52015 = n69857 & n52014 ;
  assign n52016 = n51262 & n51843 ;
  assign n51780 = n51271 | n51779 ;
  assign n82157 = ~n51780 ;
  assign n52017 = n51776 & n82157 ;
  assign n82158 = ~n51781 ;
  assign n52018 = n51779 & n82158 ;
  assign n52019 = n52017 | n52018 ;
  assign n52020 = n66715 & n52019 ;
  assign n52021 = n82140 & n52020 ;
  assign n52022 = n52016 | n52021 ;
  assign n52023 = n69656 & n52022 ;
  assign n52024 = n51270 & n51843 ;
  assign n51775 = n51279 | n51774 ;
  assign n82159 = ~n51775 ;
  assign n52025 = n82159 & n51923 ;
  assign n82160 = ~n51924 ;
  assign n52026 = n51774 & n82160 ;
  assign n52027 = n52025 | n52026 ;
  assign n52028 = n66715 & n52027 ;
  assign n52029 = n82140 & n52028 ;
  assign n52030 = n52024 | n52029 ;
  assign n52031 = n69528 & n52030 ;
  assign n52032 = n51278 & n51843 ;
  assign n51768 = n51287 | n51767 ;
  assign n82161 = ~n51768 ;
  assign n52033 = n51764 & n82161 ;
  assign n82162 = ~n51769 ;
  assign n52034 = n51767 & n82162 ;
  assign n52035 = n52033 | n52034 ;
  assign n52036 = n66715 & n52035 ;
  assign n52037 = n82140 & n52036 ;
  assign n52038 = n52032 | n52037 ;
  assign n52039 = n69261 & n52038 ;
  assign n52040 = n51286 & n51843 ;
  assign n51763 = n51295 | n51762 ;
  assign n82163 = ~n51763 ;
  assign n52041 = n82163 & n51919 ;
  assign n82164 = ~n51920 ;
  assign n52042 = n51762 & n82164 ;
  assign n52043 = n52041 | n52042 ;
  assign n52044 = n66715 & n52043 ;
  assign n52045 = n82140 & n52044 ;
  assign n52046 = n52040 | n52045 ;
  assign n52047 = n69075 & n52046 ;
  assign n52048 = n51294 & n51843 ;
  assign n51756 = n51303 | n51755 ;
  assign n82165 = ~n51756 ;
  assign n52049 = n51752 & n82165 ;
  assign n82166 = ~n51757 ;
  assign n52050 = n51755 & n82166 ;
  assign n52051 = n52049 | n52050 ;
  assign n52052 = n66715 & n52051 ;
  assign n52053 = n82140 & n52052 ;
  assign n52054 = n52048 | n52053 ;
  assign n52055 = n68993 & n52054 ;
  assign n52056 = n51302 & n51843 ;
  assign n51751 = n51311 | n51750 ;
  assign n82167 = ~n51751 ;
  assign n52057 = n82167 & n51915 ;
  assign n82168 = ~n51916 ;
  assign n52058 = n51750 & n82168 ;
  assign n52059 = n52057 | n52058 ;
  assign n52060 = n66715 & n52059 ;
  assign n52061 = n82140 & n52060 ;
  assign n52062 = n52056 | n52061 ;
  assign n52063 = n68716 & n52062 ;
  assign n52064 = n51310 & n51843 ;
  assign n51744 = n51319 | n51743 ;
  assign n82169 = ~n51744 ;
  assign n52065 = n51740 & n82169 ;
  assign n82170 = ~n51745 ;
  assign n52066 = n51743 & n82170 ;
  assign n52067 = n52065 | n52066 ;
  assign n52068 = n66715 & n52067 ;
  assign n52069 = n82140 & n52068 ;
  assign n52070 = n52064 | n52069 ;
  assign n52071 = n68545 & n52070 ;
  assign n52072 = n51318 & n51843 ;
  assign n51739 = n51327 | n51738 ;
  assign n82171 = ~n51739 ;
  assign n52073 = n82171 & n51911 ;
  assign n82172 = ~n51912 ;
  assign n52074 = n51738 & n82172 ;
  assign n52075 = n52073 | n52074 ;
  assign n52076 = n66715 & n52075 ;
  assign n52077 = n82140 & n52076 ;
  assign n52078 = n52072 | n52077 ;
  assign n52079 = n68438 & n52078 ;
  assign n52080 = n51326 & n51843 ;
  assign n51732 = n51335 | n51731 ;
  assign n82173 = ~n51732 ;
  assign n52081 = n51728 & n82173 ;
  assign n82174 = ~n51733 ;
  assign n52082 = n51731 & n82174 ;
  assign n52083 = n52081 | n52082 ;
  assign n52084 = n66715 & n52083 ;
  assign n52085 = n82140 & n52084 ;
  assign n52086 = n52080 | n52085 ;
  assign n52087 = n68214 & n52086 ;
  assign n52088 = n51334 & n51843 ;
  assign n51727 = n51343 | n51726 ;
  assign n82175 = ~n51727 ;
  assign n52089 = n82175 & n51907 ;
  assign n82176 = ~n51908 ;
  assign n52090 = n51726 & n82176 ;
  assign n52091 = n52089 | n52090 ;
  assign n52092 = n66715 & n52091 ;
  assign n52093 = n82140 & n52092 ;
  assign n52094 = n52088 | n52093 ;
  assign n52095 = n68058 & n52094 ;
  assign n52096 = n51342 & n51843 ;
  assign n51720 = n51351 | n51719 ;
  assign n82177 = ~n51720 ;
  assign n52097 = n51716 & n82177 ;
  assign n82178 = ~n51721 ;
  assign n52098 = n51719 & n82178 ;
  assign n52099 = n52097 | n52098 ;
  assign n52100 = n66715 & n52099 ;
  assign n52101 = n82140 & n52100 ;
  assign n52102 = n52096 | n52101 ;
  assign n52103 = n67986 & n52102 ;
  assign n52104 = n51350 & n51843 ;
  assign n51715 = n51359 | n51714 ;
  assign n82179 = ~n51715 ;
  assign n52105 = n82179 & n51903 ;
  assign n82180 = ~n51904 ;
  assign n52106 = n51714 & n82180 ;
  assign n52107 = n52105 | n52106 ;
  assign n52108 = n66715 & n52107 ;
  assign n52109 = n82140 & n52108 ;
  assign n52110 = n52104 | n52109 ;
  assign n52111 = n67763 & n52110 ;
  assign n52112 = n51358 & n51843 ;
  assign n51708 = n51367 | n51707 ;
  assign n82181 = ~n51708 ;
  assign n52113 = n51704 & n82181 ;
  assign n82182 = ~n51709 ;
  assign n52114 = n51707 & n82182 ;
  assign n52115 = n52113 | n52114 ;
  assign n52116 = n66715 & n52115 ;
  assign n52117 = n82140 & n52116 ;
  assign n52118 = n52112 | n52117 ;
  assign n52119 = n67622 & n52118 ;
  assign n52120 = n51366 & n51843 ;
  assign n51703 = n51375 | n51702 ;
  assign n82183 = ~n51703 ;
  assign n52121 = n82183 & n51899 ;
  assign n82184 = ~n51900 ;
  assign n52122 = n51702 & n82184 ;
  assign n52123 = n52121 | n52122 ;
  assign n52124 = n66715 & n52123 ;
  assign n52125 = n82140 & n52124 ;
  assign n52126 = n52120 | n52125 ;
  assign n52127 = n67531 & n52126 ;
  assign n52128 = n51374 & n51843 ;
  assign n51696 = n51383 | n51695 ;
  assign n82185 = ~n51696 ;
  assign n52129 = n51692 & n82185 ;
  assign n82186 = ~n51697 ;
  assign n52130 = n51695 & n82186 ;
  assign n52131 = n52129 | n52130 ;
  assign n52132 = n66715 & n52131 ;
  assign n52133 = n82140 & n52132 ;
  assign n52134 = n52128 | n52133 ;
  assign n52135 = n67348 & n52134 ;
  assign n52136 = n51382 & n51843 ;
  assign n51691 = n51391 | n51690 ;
  assign n82187 = ~n51691 ;
  assign n52137 = n82187 & n51895 ;
  assign n82188 = ~n51896 ;
  assign n52138 = n51690 & n82188 ;
  assign n52139 = n52137 | n52138 ;
  assign n52140 = n66715 & n52139 ;
  assign n52141 = n82140 & n52140 ;
  assign n52142 = n52136 | n52141 ;
  assign n52143 = n67222 & n52142 ;
  assign n52144 = n51390 & n51843 ;
  assign n51684 = n51399 | n51683 ;
  assign n82189 = ~n51684 ;
  assign n52145 = n51680 & n82189 ;
  assign n82190 = ~n51685 ;
  assign n52146 = n51683 & n82190 ;
  assign n52147 = n52145 | n52146 ;
  assign n52148 = n66715 & n52147 ;
  assign n52149 = n82140 & n52148 ;
  assign n52150 = n52144 | n52149 ;
  assign n52151 = n67164 & n52150 ;
  assign n52152 = n51398 & n51843 ;
  assign n51679 = n51407 | n51678 ;
  assign n82191 = ~n51679 ;
  assign n52153 = n82191 & n51891 ;
  assign n82192 = ~n51892 ;
  assign n52154 = n51678 & n82192 ;
  assign n52155 = n52153 | n52154 ;
  assign n52156 = n66715 & n52155 ;
  assign n52157 = n82140 & n52156 ;
  assign n52158 = n52152 | n52157 ;
  assign n52159 = n66979 & n52158 ;
  assign n52160 = n51406 & n51843 ;
  assign n51672 = n51415 | n51671 ;
  assign n82193 = ~n51672 ;
  assign n52161 = n51668 & n82193 ;
  assign n82194 = ~n51673 ;
  assign n52162 = n51671 & n82194 ;
  assign n52163 = n52161 | n52162 ;
  assign n52164 = n66715 & n52163 ;
  assign n52165 = n82140 & n52164 ;
  assign n52166 = n52160 | n52165 ;
  assign n52167 = n66868 & n52166 ;
  assign n52168 = n51414 & n51843 ;
  assign n51667 = n51423 | n51666 ;
  assign n82195 = ~n51667 ;
  assign n52169 = n82195 & n51887 ;
  assign n82196 = ~n51888 ;
  assign n52170 = n51666 & n82196 ;
  assign n52171 = n52169 | n52170 ;
  assign n52172 = n66715 & n52171 ;
  assign n52173 = n82140 & n52172 ;
  assign n52174 = n52168 | n52173 ;
  assign n52175 = n66797 & n52174 ;
  assign n52176 = n51422 & n51843 ;
  assign n51660 = n51431 | n51659 ;
  assign n82197 = ~n51660 ;
  assign n52177 = n51656 & n82197 ;
  assign n82198 = ~n51661 ;
  assign n52178 = n51659 & n82198 ;
  assign n52179 = n52177 | n52178 ;
  assign n52180 = n66715 & n52179 ;
  assign n52181 = n82140 & n52180 ;
  assign n52182 = n52176 | n52181 ;
  assign n52183 = n66654 & n52182 ;
  assign n52184 = n51430 & n51843 ;
  assign n51655 = n51439 | n51654 ;
  assign n82199 = ~n51655 ;
  assign n52185 = n82199 & n51883 ;
  assign n82200 = ~n51884 ;
  assign n52186 = n51654 & n82200 ;
  assign n52187 = n52185 | n52186 ;
  assign n52188 = n66715 & n52187 ;
  assign n52189 = n82140 & n52188 ;
  assign n52190 = n52184 | n52189 ;
  assign n52191 = n66560 & n52190 ;
  assign n52192 = n51438 & n51843 ;
  assign n51648 = n51447 | n51647 ;
  assign n82201 = ~n51648 ;
  assign n52193 = n51644 & n82201 ;
  assign n82202 = ~n51649 ;
  assign n52194 = n51647 & n82202 ;
  assign n52195 = n52193 | n52194 ;
  assign n52196 = n66715 & n52195 ;
  assign n52197 = n82140 & n52196 ;
  assign n52198 = n52192 | n52197 ;
  assign n52199 = n66505 & n52198 ;
  assign n52200 = n51446 & n51843 ;
  assign n51643 = n51455 | n51642 ;
  assign n82203 = ~n51643 ;
  assign n52201 = n82203 & n51879 ;
  assign n82204 = ~n51880 ;
  assign n52202 = n51642 & n82204 ;
  assign n52203 = n52201 | n52202 ;
  assign n52204 = n66715 & n52203 ;
  assign n52205 = n82140 & n52204 ;
  assign n52206 = n52200 | n52205 ;
  assign n52207 = n66379 & n52206 ;
  assign n52208 = n51454 & n51843 ;
  assign n51636 = n51463 | n51635 ;
  assign n82205 = ~n51636 ;
  assign n52209 = n51632 & n82205 ;
  assign n82206 = ~n51637 ;
  assign n52210 = n51635 & n82206 ;
  assign n52211 = n52209 | n52210 ;
  assign n52212 = n66715 & n52211 ;
  assign n52213 = n82140 & n52212 ;
  assign n52214 = n52208 | n52213 ;
  assign n52215 = n66299 & n52214 ;
  assign n52216 = n51462 & n51843 ;
  assign n51631 = n51471 | n51630 ;
  assign n82207 = ~n51631 ;
  assign n52217 = n82207 & n51875 ;
  assign n82208 = ~n51876 ;
  assign n52218 = n51630 & n82208 ;
  assign n52219 = n52217 | n52218 ;
  assign n52220 = n66715 & n52219 ;
  assign n52221 = n82140 & n52220 ;
  assign n52222 = n52216 | n52221 ;
  assign n52223 = n66244 & n52222 ;
  assign n52224 = n51470 & n51843 ;
  assign n51624 = n51479 | n51623 ;
  assign n82209 = ~n51624 ;
  assign n52225 = n51620 & n82209 ;
  assign n82210 = ~n51625 ;
  assign n52226 = n51623 & n82210 ;
  assign n52227 = n52225 | n52226 ;
  assign n52228 = n66715 & n52227 ;
  assign n52229 = n82140 & n52228 ;
  assign n52230 = n52224 | n52229 ;
  assign n52231 = n66145 & n52230 ;
  assign n52232 = n51478 & n51843 ;
  assign n51619 = n51487 | n51618 ;
  assign n82211 = ~n51619 ;
  assign n52233 = n82211 & n51871 ;
  assign n82212 = ~n51872 ;
  assign n52234 = n51618 & n82212 ;
  assign n52235 = n52233 | n52234 ;
  assign n52236 = n66715 & n52235 ;
  assign n52237 = n82140 & n52236 ;
  assign n52238 = n52232 | n52237 ;
  assign n52239 = n66081 & n52238 ;
  assign n52240 = n51486 & n51843 ;
  assign n51612 = n51495 | n51611 ;
  assign n82213 = ~n51612 ;
  assign n52241 = n51608 & n82213 ;
  assign n82214 = ~n51613 ;
  assign n52242 = n51611 & n82214 ;
  assign n52243 = n52241 | n52242 ;
  assign n52244 = n66715 & n52243 ;
  assign n52245 = n82140 & n52244 ;
  assign n52246 = n52240 | n52245 ;
  assign n52247 = n66043 & n52246 ;
  assign n52248 = n51494 & n51843 ;
  assign n51607 = n51503 | n51606 ;
  assign n82215 = ~n51607 ;
  assign n52249 = n82215 & n51867 ;
  assign n82216 = ~n51868 ;
  assign n52250 = n51606 & n82216 ;
  assign n52251 = n52249 | n52250 ;
  assign n52252 = n66715 & n52251 ;
  assign n52253 = n82140 & n52252 ;
  assign n52254 = n52248 | n52253 ;
  assign n52255 = n65960 & n52254 ;
  assign n52256 = n51502 & n51843 ;
  assign n51600 = n51511 | n51599 ;
  assign n82217 = ~n51600 ;
  assign n52257 = n51596 & n82217 ;
  assign n82218 = ~n51601 ;
  assign n52258 = n51599 & n82218 ;
  assign n52259 = n52257 | n52258 ;
  assign n52260 = n66715 & n52259 ;
  assign n52261 = n82140 & n52260 ;
  assign n52262 = n52256 | n52261 ;
  assign n52263 = n65909 & n52262 ;
  assign n52264 = n51510 & n51843 ;
  assign n51595 = n51519 | n51594 ;
  assign n82219 = ~n51595 ;
  assign n52265 = n82219 & n51863 ;
  assign n82220 = ~n51864 ;
  assign n52266 = n51594 & n82220 ;
  assign n52267 = n52265 | n52266 ;
  assign n52268 = n66715 & n52267 ;
  assign n52269 = n82140 & n52268 ;
  assign n52270 = n52264 | n52269 ;
  assign n52271 = n65877 & n52270 ;
  assign n52272 = n51518 & n51843 ;
  assign n51588 = n51527 | n51587 ;
  assign n82221 = ~n51588 ;
  assign n52273 = n51584 & n82221 ;
  assign n82222 = ~n51589 ;
  assign n52274 = n51587 & n82222 ;
  assign n52275 = n52273 | n52274 ;
  assign n52276 = n66715 & n52275 ;
  assign n52277 = n82140 & n52276 ;
  assign n52278 = n52272 | n52277 ;
  assign n52279 = n65820 & n52278 ;
  assign n52280 = n51526 & n51843 ;
  assign n51583 = n51535 | n51582 ;
  assign n82223 = ~n51583 ;
  assign n52281 = n82223 & n51859 ;
  assign n82224 = ~n51860 ;
  assign n52282 = n51582 & n82224 ;
  assign n52283 = n52281 | n52282 ;
  assign n52284 = n66715 & n52283 ;
  assign n52285 = n82140 & n52284 ;
  assign n52286 = n52280 | n52285 ;
  assign n52287 = n65791 & n52286 ;
  assign n52288 = n51534 & n51843 ;
  assign n52289 = n51544 | n51576 ;
  assign n82225 = ~n52289 ;
  assign n52290 = n51573 & n82225 ;
  assign n82226 = ~n51577 ;
  assign n52291 = n51576 & n82226 ;
  assign n52292 = n52290 | n52291 ;
  assign n52293 = n66715 & n52292 ;
  assign n52294 = n82140 & n52293 ;
  assign n52295 = n52288 | n52294 ;
  assign n52296 = n65772 & n52295 ;
  assign n52297 = n51543 & n51843 ;
  assign n52298 = n51552 | n51572 ;
  assign n82227 = ~n52298 ;
  assign n52299 = n51568 & n82227 ;
  assign n82228 = ~n51856 ;
  assign n52300 = n51572 & n82228 ;
  assign n52301 = n52299 | n52300 ;
  assign n52302 = n66715 & n52301 ;
  assign n52303 = n82140 & n52302 ;
  assign n52304 = n52297 | n52303 ;
  assign n52305 = n65746 & n52304 ;
  assign n52306 = n51551 & n51843 ;
  assign n51854 = n51563 | n51566 ;
  assign n82229 = ~n51854 ;
  assign n52307 = n51852 & n82229 ;
  assign n82230 = ~n51567 ;
  assign n52308 = n51566 & n82230 ;
  assign n52309 = n52307 | n52308 ;
  assign n52310 = n66715 & n52309 ;
  assign n52311 = n82140 & n52310 ;
  assign n52312 = n52306 | n52311 ;
  assign n52313 = n65721 & n52312 ;
  assign n51844 = n51554 & n51843 ;
  assign n51561 = n19324 & n51559 ;
  assign n52314 = n51561 & n82135 ;
  assign n52315 = n279 | n52314 ;
  assign n82231 = ~n52315 ;
  assign n52316 = n51852 & n82231 ;
  assign n52317 = n82140 & n52316 ;
  assign n52318 = n51844 | n52317 ;
  assign n52319 = n65686 & n52318 ;
  assign n52320 = n20095 & n82140 ;
  assign n52322 = n82130 & n52321 ;
  assign n52323 = n51839 | n52322 ;
  assign n52324 = n82131 & n52323 ;
  assign n82232 = ~n52324 ;
  assign n52325 = n20091 & n82232 ;
  assign n82233 = ~n52325 ;
  assign n52326 = x15 & n82233 ;
  assign n52327 = n52320 | n52326 ;
  assign n52335 = n65670 & n52327 ;
  assign n52328 = n20091 & n82140 ;
  assign n82234 = ~n52328 ;
  assign n52329 = x15 & n82234 ;
  assign n52330 = n52320 | n52329 ;
  assign n52331 = x65 & n52330 ;
  assign n52332 = x65 | n52320 ;
  assign n52333 = n52329 | n52332 ;
  assign n82235 = ~n52331 ;
  assign n52334 = n82235 & n52333 ;
  assign n52336 = n20102 | n52334 ;
  assign n82236 = ~n52335 ;
  assign n52337 = n82236 & n52336 ;
  assign n82237 = ~n52317 ;
  assign n52338 = x66 & n82237 ;
  assign n82238 = ~n51844 ;
  assign n52339 = n82238 & n52338 ;
  assign n52340 = n52337 | n52339 ;
  assign n82239 = ~n52319 ;
  assign n52341 = n82239 & n52340 ;
  assign n82240 = ~n52311 ;
  assign n52342 = x67 & n82240 ;
  assign n82241 = ~n52306 ;
  assign n52343 = n82241 & n52342 ;
  assign n52344 = n52313 | n52343 ;
  assign n52345 = n52341 | n52344 ;
  assign n82242 = ~n52313 ;
  assign n52346 = n82242 & n52345 ;
  assign n82243 = ~n52303 ;
  assign n52347 = x68 & n82243 ;
  assign n82244 = ~n52297 ;
  assign n52348 = n82244 & n52347 ;
  assign n52349 = n52305 | n52348 ;
  assign n52350 = n52346 | n52349 ;
  assign n82245 = ~n52305 ;
  assign n52351 = n82245 & n52350 ;
  assign n82246 = ~n52294 ;
  assign n52352 = x69 & n82246 ;
  assign n82247 = ~n52288 ;
  assign n52353 = n82247 & n52352 ;
  assign n52354 = n52296 | n52353 ;
  assign n52355 = n52351 | n52354 ;
  assign n82248 = ~n52296 ;
  assign n52356 = n82248 & n52355 ;
  assign n82249 = ~n52285 ;
  assign n52357 = x70 & n82249 ;
  assign n82250 = ~n52280 ;
  assign n52358 = n82250 & n52357 ;
  assign n52359 = n52287 | n52358 ;
  assign n52361 = n52356 | n52359 ;
  assign n82251 = ~n52287 ;
  assign n52362 = n82251 & n52361 ;
  assign n82252 = ~n52277 ;
  assign n52363 = x71 & n82252 ;
  assign n82253 = ~n52272 ;
  assign n52364 = n82253 & n52363 ;
  assign n52365 = n52279 | n52364 ;
  assign n52366 = n52362 | n52365 ;
  assign n82254 = ~n52279 ;
  assign n52367 = n82254 & n52366 ;
  assign n82255 = ~n52269 ;
  assign n52368 = x72 & n82255 ;
  assign n82256 = ~n52264 ;
  assign n52369 = n82256 & n52368 ;
  assign n52370 = n52271 | n52369 ;
  assign n52372 = n52367 | n52370 ;
  assign n82257 = ~n52271 ;
  assign n52373 = n82257 & n52372 ;
  assign n82258 = ~n52261 ;
  assign n52374 = x73 & n82258 ;
  assign n82259 = ~n52256 ;
  assign n52375 = n82259 & n52374 ;
  assign n52376 = n52263 | n52375 ;
  assign n52377 = n52373 | n52376 ;
  assign n82260 = ~n52263 ;
  assign n52378 = n82260 & n52377 ;
  assign n82261 = ~n52253 ;
  assign n52379 = x74 & n82261 ;
  assign n82262 = ~n52248 ;
  assign n52380 = n82262 & n52379 ;
  assign n52381 = n52255 | n52380 ;
  assign n52383 = n52378 | n52381 ;
  assign n82263 = ~n52255 ;
  assign n52384 = n82263 & n52383 ;
  assign n82264 = ~n52245 ;
  assign n52385 = x75 & n82264 ;
  assign n82265 = ~n52240 ;
  assign n52386 = n82265 & n52385 ;
  assign n52387 = n52247 | n52386 ;
  assign n52388 = n52384 | n52387 ;
  assign n82266 = ~n52247 ;
  assign n52389 = n82266 & n52388 ;
  assign n82267 = ~n52237 ;
  assign n52390 = x76 & n82267 ;
  assign n82268 = ~n52232 ;
  assign n52391 = n82268 & n52390 ;
  assign n52392 = n52239 | n52391 ;
  assign n52394 = n52389 | n52392 ;
  assign n82269 = ~n52239 ;
  assign n52395 = n82269 & n52394 ;
  assign n82270 = ~n52229 ;
  assign n52396 = x77 & n82270 ;
  assign n82271 = ~n52224 ;
  assign n52397 = n82271 & n52396 ;
  assign n52398 = n52231 | n52397 ;
  assign n52399 = n52395 | n52398 ;
  assign n82272 = ~n52231 ;
  assign n52400 = n82272 & n52399 ;
  assign n82273 = ~n52221 ;
  assign n52401 = x78 & n82273 ;
  assign n82274 = ~n52216 ;
  assign n52402 = n82274 & n52401 ;
  assign n52403 = n52223 | n52402 ;
  assign n52405 = n52400 | n52403 ;
  assign n82275 = ~n52223 ;
  assign n52406 = n82275 & n52405 ;
  assign n82276 = ~n52213 ;
  assign n52407 = x79 & n82276 ;
  assign n82277 = ~n52208 ;
  assign n52408 = n82277 & n52407 ;
  assign n52409 = n52215 | n52408 ;
  assign n52410 = n52406 | n52409 ;
  assign n82278 = ~n52215 ;
  assign n52411 = n82278 & n52410 ;
  assign n82279 = ~n52205 ;
  assign n52412 = x80 & n82279 ;
  assign n82280 = ~n52200 ;
  assign n52413 = n82280 & n52412 ;
  assign n52414 = n52207 | n52413 ;
  assign n52416 = n52411 | n52414 ;
  assign n82281 = ~n52207 ;
  assign n52417 = n82281 & n52416 ;
  assign n82282 = ~n52197 ;
  assign n52418 = x81 & n82282 ;
  assign n82283 = ~n52192 ;
  assign n52419 = n82283 & n52418 ;
  assign n52420 = n52199 | n52419 ;
  assign n52421 = n52417 | n52420 ;
  assign n82284 = ~n52199 ;
  assign n52422 = n82284 & n52421 ;
  assign n82285 = ~n52189 ;
  assign n52423 = x82 & n82285 ;
  assign n82286 = ~n52184 ;
  assign n52424 = n82286 & n52423 ;
  assign n52425 = n52191 | n52424 ;
  assign n52427 = n52422 | n52425 ;
  assign n82287 = ~n52191 ;
  assign n52428 = n82287 & n52427 ;
  assign n82288 = ~n52181 ;
  assign n52429 = x83 & n82288 ;
  assign n82289 = ~n52176 ;
  assign n52430 = n82289 & n52429 ;
  assign n52431 = n52183 | n52430 ;
  assign n52432 = n52428 | n52431 ;
  assign n82290 = ~n52183 ;
  assign n52433 = n82290 & n52432 ;
  assign n82291 = ~n52173 ;
  assign n52434 = x84 & n82291 ;
  assign n82292 = ~n52168 ;
  assign n52435 = n82292 & n52434 ;
  assign n52436 = n52175 | n52435 ;
  assign n52438 = n52433 | n52436 ;
  assign n82293 = ~n52175 ;
  assign n52439 = n82293 & n52438 ;
  assign n82294 = ~n52165 ;
  assign n52440 = x85 & n82294 ;
  assign n82295 = ~n52160 ;
  assign n52441 = n82295 & n52440 ;
  assign n52442 = n52167 | n52441 ;
  assign n52443 = n52439 | n52442 ;
  assign n82296 = ~n52167 ;
  assign n52444 = n82296 & n52443 ;
  assign n82297 = ~n52157 ;
  assign n52445 = x86 & n82297 ;
  assign n82298 = ~n52152 ;
  assign n52446 = n82298 & n52445 ;
  assign n52447 = n52159 | n52446 ;
  assign n52449 = n52444 | n52447 ;
  assign n82299 = ~n52159 ;
  assign n52450 = n82299 & n52449 ;
  assign n82300 = ~n52149 ;
  assign n52451 = x87 & n82300 ;
  assign n82301 = ~n52144 ;
  assign n52452 = n82301 & n52451 ;
  assign n52453 = n52151 | n52452 ;
  assign n52454 = n52450 | n52453 ;
  assign n82302 = ~n52151 ;
  assign n52455 = n82302 & n52454 ;
  assign n82303 = ~n52141 ;
  assign n52456 = x88 & n82303 ;
  assign n82304 = ~n52136 ;
  assign n52457 = n82304 & n52456 ;
  assign n52458 = n52143 | n52457 ;
  assign n52460 = n52455 | n52458 ;
  assign n82305 = ~n52143 ;
  assign n52461 = n82305 & n52460 ;
  assign n82306 = ~n52133 ;
  assign n52462 = x89 & n82306 ;
  assign n82307 = ~n52128 ;
  assign n52463 = n82307 & n52462 ;
  assign n52464 = n52135 | n52463 ;
  assign n52465 = n52461 | n52464 ;
  assign n82308 = ~n52135 ;
  assign n52466 = n82308 & n52465 ;
  assign n82309 = ~n52125 ;
  assign n52467 = x90 & n82309 ;
  assign n82310 = ~n52120 ;
  assign n52468 = n82310 & n52467 ;
  assign n52469 = n52127 | n52468 ;
  assign n52471 = n52466 | n52469 ;
  assign n82311 = ~n52127 ;
  assign n52472 = n82311 & n52471 ;
  assign n82312 = ~n52117 ;
  assign n52473 = x91 & n82312 ;
  assign n82313 = ~n52112 ;
  assign n52474 = n82313 & n52473 ;
  assign n52475 = n52119 | n52474 ;
  assign n52476 = n52472 | n52475 ;
  assign n82314 = ~n52119 ;
  assign n52477 = n82314 & n52476 ;
  assign n82315 = ~n52109 ;
  assign n52478 = x92 & n82315 ;
  assign n82316 = ~n52104 ;
  assign n52479 = n82316 & n52478 ;
  assign n52480 = n52111 | n52479 ;
  assign n52482 = n52477 | n52480 ;
  assign n82317 = ~n52111 ;
  assign n52483 = n82317 & n52482 ;
  assign n82318 = ~n52101 ;
  assign n52484 = x93 & n82318 ;
  assign n82319 = ~n52096 ;
  assign n52485 = n82319 & n52484 ;
  assign n52486 = n52103 | n52485 ;
  assign n52487 = n52483 | n52486 ;
  assign n82320 = ~n52103 ;
  assign n52488 = n82320 & n52487 ;
  assign n82321 = ~n52093 ;
  assign n52489 = x94 & n82321 ;
  assign n82322 = ~n52088 ;
  assign n52490 = n82322 & n52489 ;
  assign n52491 = n52095 | n52490 ;
  assign n52493 = n52488 | n52491 ;
  assign n82323 = ~n52095 ;
  assign n52494 = n82323 & n52493 ;
  assign n82324 = ~n52085 ;
  assign n52495 = x95 & n82324 ;
  assign n82325 = ~n52080 ;
  assign n52496 = n82325 & n52495 ;
  assign n52497 = n52087 | n52496 ;
  assign n52498 = n52494 | n52497 ;
  assign n82326 = ~n52087 ;
  assign n52499 = n82326 & n52498 ;
  assign n82327 = ~n52077 ;
  assign n52500 = x96 & n82327 ;
  assign n82328 = ~n52072 ;
  assign n52501 = n82328 & n52500 ;
  assign n52502 = n52079 | n52501 ;
  assign n52504 = n52499 | n52502 ;
  assign n82329 = ~n52079 ;
  assign n52505 = n82329 & n52504 ;
  assign n82330 = ~n52069 ;
  assign n52506 = x97 & n82330 ;
  assign n82331 = ~n52064 ;
  assign n52507 = n82331 & n52506 ;
  assign n52508 = n52071 | n52507 ;
  assign n52509 = n52505 | n52508 ;
  assign n82332 = ~n52071 ;
  assign n52510 = n82332 & n52509 ;
  assign n82333 = ~n52061 ;
  assign n52511 = x98 & n82333 ;
  assign n82334 = ~n52056 ;
  assign n52512 = n82334 & n52511 ;
  assign n52513 = n52063 | n52512 ;
  assign n52515 = n52510 | n52513 ;
  assign n82335 = ~n52063 ;
  assign n52516 = n82335 & n52515 ;
  assign n82336 = ~n52053 ;
  assign n52517 = x99 & n82336 ;
  assign n82337 = ~n52048 ;
  assign n52518 = n82337 & n52517 ;
  assign n52519 = n52055 | n52518 ;
  assign n52520 = n52516 | n52519 ;
  assign n82338 = ~n52055 ;
  assign n52521 = n82338 & n52520 ;
  assign n82339 = ~n52045 ;
  assign n52522 = x100 & n82339 ;
  assign n82340 = ~n52040 ;
  assign n52523 = n82340 & n52522 ;
  assign n52524 = n52047 | n52523 ;
  assign n52526 = n52521 | n52524 ;
  assign n82341 = ~n52047 ;
  assign n52527 = n82341 & n52526 ;
  assign n82342 = ~n52037 ;
  assign n52528 = x101 & n82342 ;
  assign n82343 = ~n52032 ;
  assign n52529 = n82343 & n52528 ;
  assign n52530 = n52039 | n52529 ;
  assign n52531 = n52527 | n52530 ;
  assign n82344 = ~n52039 ;
  assign n52532 = n82344 & n52531 ;
  assign n82345 = ~n52029 ;
  assign n52533 = x102 & n82345 ;
  assign n82346 = ~n52024 ;
  assign n52534 = n82346 & n52533 ;
  assign n52535 = n52031 | n52534 ;
  assign n52537 = n52532 | n52535 ;
  assign n82347 = ~n52031 ;
  assign n52538 = n82347 & n52537 ;
  assign n82348 = ~n52021 ;
  assign n52539 = x103 & n82348 ;
  assign n82349 = ~n52016 ;
  assign n52540 = n82349 & n52539 ;
  assign n52541 = n52023 | n52540 ;
  assign n52542 = n52538 | n52541 ;
  assign n82350 = ~n52023 ;
  assign n52543 = n82350 & n52542 ;
  assign n82351 = ~n52013 ;
  assign n52544 = x104 & n82351 ;
  assign n82352 = ~n52008 ;
  assign n52545 = n82352 & n52544 ;
  assign n52546 = n52015 | n52545 ;
  assign n52548 = n52543 | n52546 ;
  assign n82353 = ~n52015 ;
  assign n52549 = n82353 & n52548 ;
  assign n82354 = ~n52005 ;
  assign n52550 = x105 & n82354 ;
  assign n82355 = ~n52000 ;
  assign n52551 = n82355 & n52550 ;
  assign n52552 = n52007 | n52551 ;
  assign n52553 = n52549 | n52552 ;
  assign n82356 = ~n52007 ;
  assign n52554 = n82356 & n52553 ;
  assign n82357 = ~n51997 ;
  assign n52555 = x106 & n82357 ;
  assign n82358 = ~n51992 ;
  assign n52556 = n82358 & n52555 ;
  assign n52557 = n51999 | n52556 ;
  assign n52559 = n52554 | n52557 ;
  assign n82359 = ~n51999 ;
  assign n52560 = n82359 & n52559 ;
  assign n82360 = ~n51989 ;
  assign n52561 = x107 & n82360 ;
  assign n82361 = ~n51984 ;
  assign n52562 = n82361 & n52561 ;
  assign n52563 = n51991 | n52562 ;
  assign n52564 = n52560 | n52563 ;
  assign n82362 = ~n51991 ;
  assign n52565 = n82362 & n52564 ;
  assign n82363 = ~n51981 ;
  assign n52566 = x108 & n82363 ;
  assign n82364 = ~n51976 ;
  assign n52567 = n82364 & n52566 ;
  assign n52568 = n51983 | n52567 ;
  assign n52570 = n52565 | n52568 ;
  assign n82365 = ~n51983 ;
  assign n52571 = n82365 & n52570 ;
  assign n82366 = ~n51973 ;
  assign n52572 = x109 & n82366 ;
  assign n82367 = ~n51968 ;
  assign n52573 = n82367 & n52572 ;
  assign n52574 = n51975 | n52573 ;
  assign n52575 = n52571 | n52574 ;
  assign n82368 = ~n51975 ;
  assign n52576 = n82368 & n52575 ;
  assign n82369 = ~n51965 ;
  assign n52577 = x110 & n82369 ;
  assign n82370 = ~n51960 ;
  assign n52578 = n82370 & n52577 ;
  assign n52579 = n51967 | n52578 ;
  assign n52581 = n52576 | n52579 ;
  assign n82371 = ~n51967 ;
  assign n52582 = n82371 & n52581 ;
  assign n82372 = ~n51957 ;
  assign n52583 = x111 & n82372 ;
  assign n82373 = ~n51952 ;
  assign n52584 = n82373 & n52583 ;
  assign n52585 = n51959 | n52584 ;
  assign n52586 = n52582 | n52585 ;
  assign n82374 = ~n51959 ;
  assign n52587 = n82374 & n52586 ;
  assign n82375 = ~n51949 ;
  assign n52588 = x112 & n82375 ;
  assign n82376 = ~n51846 ;
  assign n52589 = n82376 & n52588 ;
  assign n52590 = n51951 | n52589 ;
  assign n52592 = n52587 | n52590 ;
  assign n82377 = ~n51951 ;
  assign n52593 = n82377 & n52592 ;
  assign n52600 = n72025 & n52599 ;
  assign n82378 = ~n51843 ;
  assign n52601 = n82378 & n52597 ;
  assign n52602 = n51189 & n51843 ;
  assign n82379 = ~n52602 ;
  assign n52603 = x113 & n82379 ;
  assign n82380 = ~n52601 ;
  assign n52604 = n82380 & n52603 ;
  assign n52605 = n20358 | n52604 ;
  assign n52606 = n52600 | n52605 ;
  assign n52608 = n52593 | n52606 ;
  assign n82381 = ~n52607 ;
  assign n52609 = n82381 & n52608 ;
  assign n82382 = ~n52587 ;
  assign n52591 = n82382 & n52590 ;
  assign n52612 = x65 & n52327 ;
  assign n82383 = ~n52612 ;
  assign n52613 = n52333 & n82383 ;
  assign n52614 = n20102 | n52613 ;
  assign n52615 = n82236 & n52614 ;
  assign n52616 = n52319 | n52339 ;
  assign n52618 = n52615 | n52616 ;
  assign n52619 = n82239 & n52618 ;
  assign n52620 = n52343 | n52619 ;
  assign n52622 = n82242 & n52620 ;
  assign n52624 = n52349 | n52622 ;
  assign n52625 = n82245 & n52624 ;
  assign n52627 = n52354 | n52625 ;
  assign n52628 = n82248 & n52627 ;
  assign n52629 = n52359 | n52628 ;
  assign n52630 = n82251 & n52629 ;
  assign n52631 = n52365 | n52630 ;
  assign n52633 = n82254 & n52631 ;
  assign n52634 = n52370 | n52633 ;
  assign n52635 = n82257 & n52634 ;
  assign n52636 = n52376 | n52635 ;
  assign n52638 = n82260 & n52636 ;
  assign n52639 = n52381 | n52638 ;
  assign n52640 = n82263 & n52639 ;
  assign n52641 = n52387 | n52640 ;
  assign n52643 = n82266 & n52641 ;
  assign n52644 = n52392 | n52643 ;
  assign n52645 = n82269 & n52644 ;
  assign n52646 = n52398 | n52645 ;
  assign n52648 = n82272 & n52646 ;
  assign n52649 = n52403 | n52648 ;
  assign n52650 = n82275 & n52649 ;
  assign n52651 = n52409 | n52650 ;
  assign n52653 = n82278 & n52651 ;
  assign n52654 = n52414 | n52653 ;
  assign n52655 = n82281 & n52654 ;
  assign n52656 = n52420 | n52655 ;
  assign n52658 = n82284 & n52656 ;
  assign n52659 = n52425 | n52658 ;
  assign n52660 = n82287 & n52659 ;
  assign n52661 = n52431 | n52660 ;
  assign n52663 = n82290 & n52661 ;
  assign n52664 = n52436 | n52663 ;
  assign n52665 = n82293 & n52664 ;
  assign n52666 = n52442 | n52665 ;
  assign n52668 = n82296 & n52666 ;
  assign n52669 = n52447 | n52668 ;
  assign n52670 = n82299 & n52669 ;
  assign n52671 = n52453 | n52670 ;
  assign n52673 = n82302 & n52671 ;
  assign n52674 = n52458 | n52673 ;
  assign n52675 = n82305 & n52674 ;
  assign n52676 = n52464 | n52675 ;
  assign n52678 = n82308 & n52676 ;
  assign n52679 = n52469 | n52678 ;
  assign n52680 = n82311 & n52679 ;
  assign n52681 = n52475 | n52680 ;
  assign n52683 = n82314 & n52681 ;
  assign n52684 = n52480 | n52683 ;
  assign n52685 = n82317 & n52684 ;
  assign n52686 = n52486 | n52685 ;
  assign n52688 = n82320 & n52686 ;
  assign n52689 = n52491 | n52688 ;
  assign n52690 = n82323 & n52689 ;
  assign n52691 = n52497 | n52690 ;
  assign n52693 = n82326 & n52691 ;
  assign n52694 = n52502 | n52693 ;
  assign n52695 = n82329 & n52694 ;
  assign n52696 = n52508 | n52695 ;
  assign n52698 = n82332 & n52696 ;
  assign n52699 = n52513 | n52698 ;
  assign n52700 = n82335 & n52699 ;
  assign n52701 = n52519 | n52700 ;
  assign n52703 = n82338 & n52701 ;
  assign n52704 = n52524 | n52703 ;
  assign n52705 = n82341 & n52704 ;
  assign n52706 = n52530 | n52705 ;
  assign n52708 = n82344 & n52706 ;
  assign n52709 = n52535 | n52708 ;
  assign n52710 = n82347 & n52709 ;
  assign n52711 = n52541 | n52710 ;
  assign n52713 = n82350 & n52711 ;
  assign n52714 = n52546 | n52713 ;
  assign n52715 = n82353 & n52714 ;
  assign n52716 = n52552 | n52715 ;
  assign n52718 = n82356 & n52716 ;
  assign n52719 = n52557 | n52718 ;
  assign n52720 = n82359 & n52719 ;
  assign n52721 = n52563 | n52720 ;
  assign n52723 = n82362 & n52721 ;
  assign n52724 = n52568 | n52723 ;
  assign n52725 = n82365 & n52724 ;
  assign n52726 = n52574 | n52725 ;
  assign n52728 = n82368 & n52726 ;
  assign n52729 = n52579 | n52728 ;
  assign n52730 = n82371 & n52729 ;
  assign n52731 = n52585 | n52730 ;
  assign n52733 = n51959 | n52590 ;
  assign n82384 = ~n52733 ;
  assign n52734 = n52731 & n82384 ;
  assign n52735 = n52591 | n52734 ;
  assign n82385 = ~n52609 ;
  assign n52736 = n82385 & n52735 ;
  assign n52737 = n82374 & n52731 ;
  assign n52738 = n52590 | n52737 ;
  assign n52739 = n82377 & n52738 ;
  assign n52740 = n52606 | n52739 ;
  assign n52741 = n51950 & n82381 ;
  assign n52742 = n52740 & n52741 ;
  assign n52743 = n52736 | n52742 ;
  assign n52744 = n72025 & n52743 ;
  assign n82386 = ~n52742 ;
  assign n53374 = x113 & n82386 ;
  assign n82387 = ~n52736 ;
  assign n53375 = n82387 & n53374 ;
  assign n53376 = n52744 | n53375 ;
  assign n82388 = ~n52730 ;
  assign n52732 = n52585 & n82388 ;
  assign n52745 = n51967 | n52585 ;
  assign n82389 = ~n52745 ;
  assign n52746 = n52581 & n82389 ;
  assign n52747 = n52732 | n52746 ;
  assign n52748 = n82385 & n52747 ;
  assign n52749 = n51958 & n82381 ;
  assign n52750 = n52740 & n52749 ;
  assign n52751 = n52748 | n52750 ;
  assign n52752 = n71645 & n52751 ;
  assign n82390 = ~n52576 ;
  assign n52580 = n82390 & n52579 ;
  assign n52753 = n51975 | n52579 ;
  assign n82391 = ~n52753 ;
  assign n52754 = n52726 & n82391 ;
  assign n52755 = n52580 | n52754 ;
  assign n52756 = n82385 & n52755 ;
  assign n52757 = n51966 & n82381 ;
  assign n52758 = n52740 & n52757 ;
  assign n52759 = n52756 | n52758 ;
  assign n52760 = n71633 & n52759 ;
  assign n82392 = ~n52758 ;
  assign n53364 = x111 & n82392 ;
  assign n82393 = ~n52756 ;
  assign n53365 = n82393 & n53364 ;
  assign n53366 = n52760 | n53365 ;
  assign n82394 = ~n52725 ;
  assign n52727 = n52574 & n82394 ;
  assign n52761 = n51983 | n52574 ;
  assign n82395 = ~n52761 ;
  assign n52762 = n52570 & n82395 ;
  assign n52763 = n52727 | n52762 ;
  assign n52764 = n82385 & n52763 ;
  assign n52765 = n51974 & n82381 ;
  assign n52766 = n52740 & n52765 ;
  assign n52767 = n52764 | n52766 ;
  assign n52768 = n71253 & n52767 ;
  assign n82396 = ~n52565 ;
  assign n52569 = n82396 & n52568 ;
  assign n52769 = n51991 | n52568 ;
  assign n82397 = ~n52769 ;
  assign n52770 = n52721 & n82397 ;
  assign n52771 = n52569 | n52770 ;
  assign n52772 = n82385 & n52771 ;
  assign n52773 = n51982 & n82381 ;
  assign n52774 = n52740 & n52773 ;
  assign n52775 = n52772 | n52774 ;
  assign n52776 = n70935 & n52775 ;
  assign n82398 = ~n52774 ;
  assign n53354 = x109 & n82398 ;
  assign n82399 = ~n52772 ;
  assign n53355 = n82399 & n53354 ;
  assign n53356 = n52776 | n53355 ;
  assign n82400 = ~n52720 ;
  assign n52722 = n52563 & n82400 ;
  assign n52777 = n51999 | n52563 ;
  assign n82401 = ~n52777 ;
  assign n52778 = n52559 & n82401 ;
  assign n52779 = n52722 | n52778 ;
  assign n52780 = n82385 & n52779 ;
  assign n52781 = n51990 & n82381 ;
  assign n52782 = n52740 & n52781 ;
  assign n52783 = n52780 | n52782 ;
  assign n52784 = n70927 & n52783 ;
  assign n82402 = ~n52554 ;
  assign n52558 = n82402 & n52557 ;
  assign n52785 = n52007 | n52557 ;
  assign n82403 = ~n52785 ;
  assign n52786 = n52716 & n82403 ;
  assign n52787 = n52558 | n52786 ;
  assign n52788 = n82385 & n52787 ;
  assign n52789 = n51998 & n82381 ;
  assign n52790 = n52740 & n52789 ;
  assign n52791 = n52788 | n52790 ;
  assign n52792 = n70609 & n52791 ;
  assign n82404 = ~n52790 ;
  assign n53344 = x107 & n82404 ;
  assign n82405 = ~n52788 ;
  assign n53345 = n82405 & n53344 ;
  assign n53346 = n52792 | n53345 ;
  assign n82406 = ~n52715 ;
  assign n52717 = n52552 & n82406 ;
  assign n52793 = n52015 | n52552 ;
  assign n82407 = ~n52793 ;
  assign n52794 = n52548 & n82407 ;
  assign n52795 = n52717 | n52794 ;
  assign n52796 = n82385 & n52795 ;
  assign n52797 = n52006 & n82381 ;
  assign n52798 = n52740 & n52797 ;
  assign n52799 = n52796 | n52798 ;
  assign n52800 = n70276 & n52799 ;
  assign n82408 = ~n52543 ;
  assign n52547 = n82408 & n52546 ;
  assign n52801 = n52023 | n52546 ;
  assign n82409 = ~n52801 ;
  assign n52802 = n52711 & n82409 ;
  assign n52803 = n52547 | n52802 ;
  assign n52804 = n82385 & n52803 ;
  assign n52805 = n52014 & n82381 ;
  assign n52806 = n52740 & n52805 ;
  assign n52807 = n52804 | n52806 ;
  assign n52808 = n70176 & n52807 ;
  assign n82410 = ~n52806 ;
  assign n53334 = x105 & n82410 ;
  assign n82411 = ~n52804 ;
  assign n53335 = n82411 & n53334 ;
  assign n53336 = n52808 | n53335 ;
  assign n82412 = ~n52710 ;
  assign n52712 = n52541 & n82412 ;
  assign n52809 = n52031 | n52541 ;
  assign n82413 = ~n52809 ;
  assign n52810 = n52537 & n82413 ;
  assign n52811 = n52712 | n52810 ;
  assign n52812 = n82385 & n52811 ;
  assign n52813 = n52022 & n82381 ;
  assign n52814 = n52740 & n52813 ;
  assign n52815 = n52812 | n52814 ;
  assign n52816 = n69857 & n52815 ;
  assign n82414 = ~n52532 ;
  assign n52536 = n82414 & n52535 ;
  assign n52817 = n52039 | n52535 ;
  assign n82415 = ~n52817 ;
  assign n52818 = n52706 & n82415 ;
  assign n52819 = n52536 | n52818 ;
  assign n52820 = n82385 & n52819 ;
  assign n52821 = n52030 & n82381 ;
  assign n52822 = n52740 & n52821 ;
  assign n52823 = n52820 | n52822 ;
  assign n52824 = n69656 & n52823 ;
  assign n82416 = ~n52822 ;
  assign n53324 = x103 & n82416 ;
  assign n82417 = ~n52820 ;
  assign n53325 = n82417 & n53324 ;
  assign n53326 = n52824 | n53325 ;
  assign n82418 = ~n52705 ;
  assign n52707 = n52530 & n82418 ;
  assign n52825 = n52047 | n52530 ;
  assign n82419 = ~n52825 ;
  assign n52826 = n52526 & n82419 ;
  assign n52827 = n52707 | n52826 ;
  assign n52828 = n82385 & n52827 ;
  assign n52829 = n52038 & n82381 ;
  assign n52830 = n52740 & n52829 ;
  assign n52831 = n52828 | n52830 ;
  assign n52832 = n69528 & n52831 ;
  assign n82420 = ~n52521 ;
  assign n52525 = n82420 & n52524 ;
  assign n52833 = n52055 | n52524 ;
  assign n82421 = ~n52833 ;
  assign n52834 = n52701 & n82421 ;
  assign n52835 = n52525 | n52834 ;
  assign n52836 = n82385 & n52835 ;
  assign n52837 = n52046 & n82381 ;
  assign n52838 = n52740 & n52837 ;
  assign n52839 = n52836 | n52838 ;
  assign n52840 = n69261 & n52839 ;
  assign n82422 = ~n52838 ;
  assign n53314 = x101 & n82422 ;
  assign n82423 = ~n52836 ;
  assign n53315 = n82423 & n53314 ;
  assign n53316 = n52840 | n53315 ;
  assign n82424 = ~n52700 ;
  assign n52702 = n52519 & n82424 ;
  assign n52841 = n52063 | n52519 ;
  assign n82425 = ~n52841 ;
  assign n52842 = n52515 & n82425 ;
  assign n52843 = n52702 | n52842 ;
  assign n52844 = n82385 & n52843 ;
  assign n52845 = n52054 & n82381 ;
  assign n52846 = n52740 & n52845 ;
  assign n52847 = n52844 | n52846 ;
  assign n52848 = n69075 & n52847 ;
  assign n82426 = ~n52510 ;
  assign n52514 = n82426 & n52513 ;
  assign n52849 = n52071 | n52513 ;
  assign n82427 = ~n52849 ;
  assign n52850 = n52696 & n82427 ;
  assign n52851 = n52514 | n52850 ;
  assign n52852 = n82385 & n52851 ;
  assign n52853 = n52062 & n82381 ;
  assign n52854 = n52740 & n52853 ;
  assign n52855 = n52852 | n52854 ;
  assign n52856 = n68993 & n52855 ;
  assign n82428 = ~n52854 ;
  assign n53304 = x99 & n82428 ;
  assign n82429 = ~n52852 ;
  assign n53305 = n82429 & n53304 ;
  assign n53306 = n52856 | n53305 ;
  assign n82430 = ~n52695 ;
  assign n52697 = n52508 & n82430 ;
  assign n52857 = n52079 | n52508 ;
  assign n82431 = ~n52857 ;
  assign n52858 = n52504 & n82431 ;
  assign n52859 = n52697 | n52858 ;
  assign n52860 = n82385 & n52859 ;
  assign n52861 = n52070 & n82381 ;
  assign n52862 = n52740 & n52861 ;
  assign n52863 = n52860 | n52862 ;
  assign n52864 = n68716 & n52863 ;
  assign n82432 = ~n52499 ;
  assign n52503 = n82432 & n52502 ;
  assign n52865 = n52087 | n52502 ;
  assign n82433 = ~n52865 ;
  assign n52866 = n52691 & n82433 ;
  assign n52867 = n52503 | n52866 ;
  assign n52868 = n82385 & n52867 ;
  assign n52869 = n52078 & n82381 ;
  assign n52870 = n52740 & n52869 ;
  assign n52871 = n52868 | n52870 ;
  assign n52872 = n68545 & n52871 ;
  assign n82434 = ~n52870 ;
  assign n53294 = x97 & n82434 ;
  assign n82435 = ~n52868 ;
  assign n53295 = n82435 & n53294 ;
  assign n53296 = n52872 | n53295 ;
  assign n82436 = ~n52690 ;
  assign n52692 = n52497 & n82436 ;
  assign n52873 = n52095 | n52497 ;
  assign n82437 = ~n52873 ;
  assign n52874 = n52493 & n82437 ;
  assign n52875 = n52692 | n52874 ;
  assign n52876 = n82385 & n52875 ;
  assign n52877 = n52086 & n82381 ;
  assign n52878 = n52740 & n52877 ;
  assign n52879 = n52876 | n52878 ;
  assign n52880 = n68438 & n52879 ;
  assign n82438 = ~n52488 ;
  assign n52492 = n82438 & n52491 ;
  assign n52881 = n52103 | n52491 ;
  assign n82439 = ~n52881 ;
  assign n52882 = n52686 & n82439 ;
  assign n52883 = n52492 | n52882 ;
  assign n52884 = n82385 & n52883 ;
  assign n52885 = n52094 & n82381 ;
  assign n52886 = n52740 & n52885 ;
  assign n52887 = n52884 | n52886 ;
  assign n52888 = n68214 & n52887 ;
  assign n82440 = ~n52886 ;
  assign n53284 = x95 & n82440 ;
  assign n82441 = ~n52884 ;
  assign n53285 = n82441 & n53284 ;
  assign n53286 = n52888 | n53285 ;
  assign n82442 = ~n52685 ;
  assign n52687 = n52486 & n82442 ;
  assign n52889 = n52111 | n52486 ;
  assign n82443 = ~n52889 ;
  assign n52890 = n52482 & n82443 ;
  assign n52891 = n52687 | n52890 ;
  assign n52892 = n82385 & n52891 ;
  assign n52893 = n52102 & n82381 ;
  assign n52894 = n52740 & n52893 ;
  assign n52895 = n52892 | n52894 ;
  assign n52896 = n68058 & n52895 ;
  assign n82444 = ~n52477 ;
  assign n52481 = n82444 & n52480 ;
  assign n52897 = n52119 | n52480 ;
  assign n82445 = ~n52897 ;
  assign n52898 = n52681 & n82445 ;
  assign n52899 = n52481 | n52898 ;
  assign n52900 = n82385 & n52899 ;
  assign n52901 = n52110 & n82381 ;
  assign n52902 = n52740 & n52901 ;
  assign n52903 = n52900 | n52902 ;
  assign n52904 = n67986 & n52903 ;
  assign n82446 = ~n52902 ;
  assign n53274 = x93 & n82446 ;
  assign n82447 = ~n52900 ;
  assign n53275 = n82447 & n53274 ;
  assign n53276 = n52904 | n53275 ;
  assign n82448 = ~n52680 ;
  assign n52682 = n52475 & n82448 ;
  assign n52905 = n52127 | n52475 ;
  assign n82449 = ~n52905 ;
  assign n52906 = n52471 & n82449 ;
  assign n52907 = n52682 | n52906 ;
  assign n52908 = n82385 & n52907 ;
  assign n52909 = n52118 & n82381 ;
  assign n52910 = n52740 & n52909 ;
  assign n52911 = n52908 | n52910 ;
  assign n52912 = n67763 & n52911 ;
  assign n82450 = ~n52466 ;
  assign n52470 = n82450 & n52469 ;
  assign n52913 = n52135 | n52469 ;
  assign n82451 = ~n52913 ;
  assign n52914 = n52676 & n82451 ;
  assign n52915 = n52470 | n52914 ;
  assign n52916 = n82385 & n52915 ;
  assign n52917 = n52126 & n82381 ;
  assign n52918 = n52740 & n52917 ;
  assign n52919 = n52916 | n52918 ;
  assign n52920 = n67622 & n52919 ;
  assign n82452 = ~n52918 ;
  assign n53264 = x91 & n82452 ;
  assign n82453 = ~n52916 ;
  assign n53265 = n82453 & n53264 ;
  assign n53266 = n52920 | n53265 ;
  assign n82454 = ~n52675 ;
  assign n52677 = n52464 & n82454 ;
  assign n52921 = n52143 | n52464 ;
  assign n82455 = ~n52921 ;
  assign n52922 = n52460 & n82455 ;
  assign n52923 = n52677 | n52922 ;
  assign n52924 = n82385 & n52923 ;
  assign n52925 = n52134 & n82381 ;
  assign n52926 = n52740 & n52925 ;
  assign n52927 = n52924 | n52926 ;
  assign n52928 = n67531 & n52927 ;
  assign n82456 = ~n52455 ;
  assign n52459 = n82456 & n52458 ;
  assign n52929 = n52151 | n52458 ;
  assign n82457 = ~n52929 ;
  assign n52930 = n52671 & n82457 ;
  assign n52931 = n52459 | n52930 ;
  assign n52932 = n82385 & n52931 ;
  assign n52933 = n52142 & n82381 ;
  assign n52934 = n52740 & n52933 ;
  assign n52935 = n52932 | n52934 ;
  assign n52936 = n67348 & n52935 ;
  assign n82458 = ~n52934 ;
  assign n53254 = x89 & n82458 ;
  assign n82459 = ~n52932 ;
  assign n53255 = n82459 & n53254 ;
  assign n53256 = n52936 | n53255 ;
  assign n82460 = ~n52670 ;
  assign n52672 = n52453 & n82460 ;
  assign n52937 = n52159 | n52453 ;
  assign n82461 = ~n52937 ;
  assign n52938 = n52449 & n82461 ;
  assign n52939 = n52672 | n52938 ;
  assign n52940 = n82385 & n52939 ;
  assign n52941 = n52150 & n82381 ;
  assign n52942 = n52740 & n52941 ;
  assign n52943 = n52940 | n52942 ;
  assign n52944 = n67222 & n52943 ;
  assign n82462 = ~n52444 ;
  assign n52448 = n82462 & n52447 ;
  assign n52945 = n52167 | n52447 ;
  assign n82463 = ~n52945 ;
  assign n52946 = n52666 & n82463 ;
  assign n52947 = n52448 | n52946 ;
  assign n52948 = n82385 & n52947 ;
  assign n52949 = n52158 & n82381 ;
  assign n52950 = n52740 & n52949 ;
  assign n52951 = n52948 | n52950 ;
  assign n52952 = n67164 & n52951 ;
  assign n82464 = ~n52950 ;
  assign n53243 = x87 & n82464 ;
  assign n82465 = ~n52948 ;
  assign n53244 = n82465 & n53243 ;
  assign n53245 = n52952 | n53244 ;
  assign n82466 = ~n52665 ;
  assign n52667 = n52442 & n82466 ;
  assign n52953 = n52175 | n52442 ;
  assign n82467 = ~n52953 ;
  assign n52954 = n52438 & n82467 ;
  assign n52955 = n52667 | n52954 ;
  assign n52956 = n82385 & n52955 ;
  assign n52957 = n52166 & n82381 ;
  assign n52958 = n52740 & n52957 ;
  assign n52959 = n52956 | n52958 ;
  assign n52960 = n66979 & n52959 ;
  assign n82468 = ~n52433 ;
  assign n52437 = n82468 & n52436 ;
  assign n52961 = n52183 | n52436 ;
  assign n82469 = ~n52961 ;
  assign n52962 = n52661 & n82469 ;
  assign n52963 = n52437 | n52962 ;
  assign n52964 = n82385 & n52963 ;
  assign n52965 = n52174 & n82381 ;
  assign n52966 = n52740 & n52965 ;
  assign n52967 = n52964 | n52966 ;
  assign n52968 = n66868 & n52967 ;
  assign n82470 = ~n52966 ;
  assign n53233 = x85 & n82470 ;
  assign n82471 = ~n52964 ;
  assign n53234 = n82471 & n53233 ;
  assign n53235 = n52968 | n53234 ;
  assign n82472 = ~n52660 ;
  assign n52662 = n52431 & n82472 ;
  assign n52969 = n52191 | n52431 ;
  assign n82473 = ~n52969 ;
  assign n52970 = n52427 & n82473 ;
  assign n52971 = n52662 | n52970 ;
  assign n52972 = n82385 & n52971 ;
  assign n52973 = n52182 & n82381 ;
  assign n52974 = n52740 & n52973 ;
  assign n52975 = n52972 | n52974 ;
  assign n52976 = n66797 & n52975 ;
  assign n82474 = ~n52422 ;
  assign n52426 = n82474 & n52425 ;
  assign n52977 = n52199 | n52425 ;
  assign n82475 = ~n52977 ;
  assign n52978 = n52656 & n82475 ;
  assign n52979 = n52426 | n52978 ;
  assign n52980 = n82385 & n52979 ;
  assign n52981 = n52190 & n82381 ;
  assign n52982 = n52740 & n52981 ;
  assign n52983 = n52980 | n52982 ;
  assign n52984 = n66654 & n52983 ;
  assign n82476 = ~n52982 ;
  assign n53222 = x83 & n82476 ;
  assign n82477 = ~n52980 ;
  assign n53223 = n82477 & n53222 ;
  assign n53224 = n52984 | n53223 ;
  assign n82478 = ~n52655 ;
  assign n52657 = n52420 & n82478 ;
  assign n52985 = n52207 | n52420 ;
  assign n82479 = ~n52985 ;
  assign n52986 = n52416 & n82479 ;
  assign n52987 = n52657 | n52986 ;
  assign n52988 = n82385 & n52987 ;
  assign n52989 = n52198 & n82381 ;
  assign n52990 = n52740 & n52989 ;
  assign n52991 = n52988 | n52990 ;
  assign n52992 = n66560 & n52991 ;
  assign n82480 = ~n52411 ;
  assign n52415 = n82480 & n52414 ;
  assign n52993 = n52215 | n52414 ;
  assign n82481 = ~n52993 ;
  assign n52994 = n52651 & n82481 ;
  assign n52995 = n52415 | n52994 ;
  assign n52996 = n82385 & n52995 ;
  assign n52997 = n52206 & n82381 ;
  assign n52998 = n52740 & n52997 ;
  assign n52999 = n52996 | n52998 ;
  assign n53000 = n66505 & n52999 ;
  assign n82482 = ~n52998 ;
  assign n53212 = x81 & n82482 ;
  assign n82483 = ~n52996 ;
  assign n53213 = n82483 & n53212 ;
  assign n53214 = n53000 | n53213 ;
  assign n82484 = ~n52650 ;
  assign n52652 = n52409 & n82484 ;
  assign n53001 = n52223 | n52409 ;
  assign n82485 = ~n53001 ;
  assign n53002 = n52405 & n82485 ;
  assign n53003 = n52652 | n53002 ;
  assign n53004 = n82385 & n53003 ;
  assign n53005 = n52214 & n82381 ;
  assign n53006 = n52740 & n53005 ;
  assign n53007 = n53004 | n53006 ;
  assign n53008 = n66379 & n53007 ;
  assign n82486 = ~n52400 ;
  assign n52404 = n82486 & n52403 ;
  assign n53009 = n52231 | n52403 ;
  assign n82487 = ~n53009 ;
  assign n53010 = n52646 & n82487 ;
  assign n53011 = n52404 | n53010 ;
  assign n53012 = n82385 & n53011 ;
  assign n53013 = n52222 & n82381 ;
  assign n53014 = n52740 & n53013 ;
  assign n53015 = n53012 | n53014 ;
  assign n53016 = n66299 & n53015 ;
  assign n82488 = ~n53014 ;
  assign n53202 = x79 & n82488 ;
  assign n82489 = ~n53012 ;
  assign n53203 = n82489 & n53202 ;
  assign n53204 = n53016 | n53203 ;
  assign n82490 = ~n52645 ;
  assign n52647 = n52398 & n82490 ;
  assign n53017 = n52239 | n52398 ;
  assign n82491 = ~n53017 ;
  assign n53018 = n52394 & n82491 ;
  assign n53019 = n52647 | n53018 ;
  assign n53020 = n82385 & n53019 ;
  assign n53021 = n52230 & n82381 ;
  assign n53022 = n52740 & n53021 ;
  assign n53023 = n53020 | n53022 ;
  assign n53024 = n66244 & n53023 ;
  assign n82492 = ~n52389 ;
  assign n52393 = n82492 & n52392 ;
  assign n53025 = n52247 | n52392 ;
  assign n82493 = ~n53025 ;
  assign n53026 = n52641 & n82493 ;
  assign n53027 = n52393 | n53026 ;
  assign n53028 = n82385 & n53027 ;
  assign n53029 = n52238 & n82381 ;
  assign n53030 = n52740 & n53029 ;
  assign n53031 = n53028 | n53030 ;
  assign n53032 = n66145 & n53031 ;
  assign n82494 = ~n53030 ;
  assign n53191 = x77 & n82494 ;
  assign n82495 = ~n53028 ;
  assign n53192 = n82495 & n53191 ;
  assign n53193 = n53032 | n53192 ;
  assign n82496 = ~n52640 ;
  assign n52642 = n52387 & n82496 ;
  assign n53033 = n52255 | n52387 ;
  assign n82497 = ~n53033 ;
  assign n53034 = n52383 & n82497 ;
  assign n53035 = n52642 | n53034 ;
  assign n53036 = n82385 & n53035 ;
  assign n53037 = n52246 & n82381 ;
  assign n53038 = n52740 & n53037 ;
  assign n53039 = n53036 | n53038 ;
  assign n53040 = n66081 & n53039 ;
  assign n82498 = ~n52378 ;
  assign n52382 = n82498 & n52381 ;
  assign n53041 = n52263 | n52381 ;
  assign n82499 = ~n53041 ;
  assign n53042 = n52636 & n82499 ;
  assign n53043 = n52382 | n53042 ;
  assign n53044 = n82385 & n53043 ;
  assign n53045 = n52254 & n82381 ;
  assign n53046 = n52740 & n53045 ;
  assign n53047 = n53044 | n53046 ;
  assign n53048 = n66043 & n53047 ;
  assign n82500 = ~n53046 ;
  assign n53181 = x75 & n82500 ;
  assign n82501 = ~n53044 ;
  assign n53182 = n82501 & n53181 ;
  assign n53183 = n53048 | n53182 ;
  assign n82502 = ~n52635 ;
  assign n52637 = n52376 & n82502 ;
  assign n53049 = n52271 | n52376 ;
  assign n82503 = ~n53049 ;
  assign n53050 = n52372 & n82503 ;
  assign n53051 = n52637 | n53050 ;
  assign n53052 = n82385 & n53051 ;
  assign n53053 = n52262 & n82381 ;
  assign n53054 = n52740 & n53053 ;
  assign n53055 = n53052 | n53054 ;
  assign n53056 = n65960 & n53055 ;
  assign n82504 = ~n52367 ;
  assign n52371 = n82504 & n52370 ;
  assign n53057 = n52279 | n52370 ;
  assign n82505 = ~n53057 ;
  assign n53058 = n52631 & n82505 ;
  assign n53059 = n52371 | n53058 ;
  assign n53060 = n82385 & n53059 ;
  assign n53061 = n52270 & n82381 ;
  assign n53062 = n52740 & n53061 ;
  assign n53063 = n53060 | n53062 ;
  assign n53064 = n65909 & n53063 ;
  assign n82506 = ~n53062 ;
  assign n53170 = x73 & n82506 ;
  assign n82507 = ~n53060 ;
  assign n53171 = n82507 & n53170 ;
  assign n53172 = n53064 | n53171 ;
  assign n82508 = ~n52630 ;
  assign n52632 = n52365 & n82508 ;
  assign n53065 = n52287 | n52365 ;
  assign n82509 = ~n53065 ;
  assign n53066 = n52361 & n82509 ;
  assign n53067 = n52632 | n53066 ;
  assign n53068 = n82385 & n53067 ;
  assign n53069 = n52278 & n82381 ;
  assign n53070 = n52740 & n53069 ;
  assign n53071 = n53068 | n53070 ;
  assign n53072 = n65877 & n53071 ;
  assign n82510 = ~n52356 ;
  assign n52360 = n82510 & n52359 ;
  assign n53073 = n52296 | n52359 ;
  assign n82511 = ~n53073 ;
  assign n53074 = n52627 & n82511 ;
  assign n53075 = n52360 | n53074 ;
  assign n53076 = n82385 & n53075 ;
  assign n53077 = n52286 & n82381 ;
  assign n53078 = n52740 & n53077 ;
  assign n53079 = n53076 | n53078 ;
  assign n53080 = n65820 & n53079 ;
  assign n82512 = ~n53078 ;
  assign n53160 = x71 & n82512 ;
  assign n82513 = ~n53076 ;
  assign n53161 = n82513 & n53160 ;
  assign n53162 = n53080 | n53161 ;
  assign n82514 = ~n52625 ;
  assign n52626 = n52354 & n82514 ;
  assign n53081 = n52305 | n52354 ;
  assign n82515 = ~n53081 ;
  assign n53082 = n52350 & n82515 ;
  assign n53083 = n52626 | n53082 ;
  assign n53084 = n82385 & n53083 ;
  assign n53085 = n52295 & n82381 ;
  assign n53086 = n52740 & n53085 ;
  assign n53087 = n53084 | n53086 ;
  assign n53088 = n65791 & n53087 ;
  assign n82516 = ~n52346 ;
  assign n52623 = n82516 & n52349 ;
  assign n53089 = n52344 | n52619 ;
  assign n53090 = n52313 | n52349 ;
  assign n82517 = ~n53090 ;
  assign n53091 = n53089 & n82517 ;
  assign n53092 = n52623 | n53091 ;
  assign n53093 = n82385 & n53092 ;
  assign n53094 = n52304 & n82381 ;
  assign n53095 = n52740 & n53094 ;
  assign n53096 = n53093 | n53095 ;
  assign n53097 = n65772 & n53096 ;
  assign n82518 = ~n53095 ;
  assign n53150 = x69 & n82518 ;
  assign n82519 = ~n53093 ;
  assign n53151 = n82519 & n53150 ;
  assign n53152 = n53097 | n53151 ;
  assign n82520 = ~n52619 ;
  assign n52621 = n52344 & n82520 ;
  assign n53098 = n52319 | n52344 ;
  assign n82521 = ~n53098 ;
  assign n53099 = n52618 & n82521 ;
  assign n53100 = n52621 | n53099 ;
  assign n53101 = n82385 & n53100 ;
  assign n53102 = n52312 & n82381 ;
  assign n53103 = n52740 & n53102 ;
  assign n53104 = n53101 | n53103 ;
  assign n53105 = n65746 & n53104 ;
  assign n82522 = ~n52337 ;
  assign n52617 = n82522 & n52616 ;
  assign n53106 = n52335 | n52616 ;
  assign n82523 = ~n53106 ;
  assign n53107 = n52336 & n82523 ;
  assign n53108 = n52617 | n53107 ;
  assign n53109 = n82385 & n53108 ;
  assign n53110 = n52318 & n82381 ;
  assign n53111 = n52740 & n53110 ;
  assign n53112 = n53109 | n53111 ;
  assign n53113 = n65721 & n53112 ;
  assign n82524 = ~n53111 ;
  assign n53140 = x67 & n82524 ;
  assign n82525 = ~n53109 ;
  assign n53141 = n82525 & n53140 ;
  assign n53142 = n53113 | n53141 ;
  assign n53114 = n20102 & n52333 ;
  assign n53115 = n82383 & n53114 ;
  assign n82526 = ~n53115 ;
  assign n53116 = n52336 & n82526 ;
  assign n53117 = n82385 & n53116 ;
  assign n53118 = n52330 & n82381 ;
  assign n53119 = n52740 & n53118 ;
  assign n53120 = n53117 | n53119 ;
  assign n53121 = n65686 & n53120 ;
  assign n52611 = n20102 & n82385 ;
  assign n53122 = n82381 & n52740 ;
  assign n82527 = ~n53122 ;
  assign n53123 = x64 & n82527 ;
  assign n82528 = ~n53123 ;
  assign n53124 = x14 & n82528 ;
  assign n53125 = n52611 | n53124 ;
  assign n53126 = x65 & n53125 ;
  assign n52610 = x64 & n82385 ;
  assign n82529 = ~n52610 ;
  assign n53127 = x14 & n82529 ;
  assign n53128 = n20102 & n82527 ;
  assign n53129 = x65 | n53128 ;
  assign n53130 = n53127 | n53129 ;
  assign n82530 = ~n53126 ;
  assign n53131 = n82530 & n53130 ;
  assign n53132 = n20903 | n53131 ;
  assign n53133 = n52611 | n53127 ;
  assign n53134 = n65670 & n53133 ;
  assign n82531 = ~n53134 ;
  assign n53135 = n53132 & n82531 ;
  assign n82532 = ~n53119 ;
  assign n53136 = x66 & n82532 ;
  assign n82533 = ~n53117 ;
  assign n53137 = n82533 & n53136 ;
  assign n53138 = n53121 | n53137 ;
  assign n53139 = n53135 | n53138 ;
  assign n82534 = ~n53121 ;
  assign n53143 = n82534 & n53139 ;
  assign n53144 = n53142 | n53143 ;
  assign n82535 = ~n53113 ;
  assign n53145 = n82535 & n53144 ;
  assign n82536 = ~n53103 ;
  assign n53146 = x68 & n82536 ;
  assign n82537 = ~n53101 ;
  assign n53147 = n82537 & n53146 ;
  assign n53148 = n53105 | n53147 ;
  assign n53149 = n53145 | n53148 ;
  assign n82538 = ~n53105 ;
  assign n53153 = n82538 & n53149 ;
  assign n53154 = n53152 | n53153 ;
  assign n82539 = ~n53097 ;
  assign n53155 = n82539 & n53154 ;
  assign n82540 = ~n53086 ;
  assign n53156 = x70 & n82540 ;
  assign n82541 = ~n53084 ;
  assign n53157 = n82541 & n53156 ;
  assign n53158 = n53088 | n53157 ;
  assign n53159 = n53155 | n53158 ;
  assign n82542 = ~n53088 ;
  assign n53163 = n82542 & n53159 ;
  assign n53164 = n53162 | n53163 ;
  assign n82543 = ~n53080 ;
  assign n53165 = n82543 & n53164 ;
  assign n82544 = ~n53070 ;
  assign n53166 = x72 & n82544 ;
  assign n82545 = ~n53068 ;
  assign n53167 = n82545 & n53166 ;
  assign n53168 = n53072 | n53167 ;
  assign n53169 = n53165 | n53168 ;
  assign n82546 = ~n53072 ;
  assign n53173 = n82546 & n53169 ;
  assign n53174 = n53172 | n53173 ;
  assign n82547 = ~n53064 ;
  assign n53175 = n82547 & n53174 ;
  assign n82548 = ~n53054 ;
  assign n53176 = x74 & n82548 ;
  assign n82549 = ~n53052 ;
  assign n53177 = n82549 & n53176 ;
  assign n53178 = n53056 | n53177 ;
  assign n53180 = n53175 | n53178 ;
  assign n82550 = ~n53056 ;
  assign n53184 = n82550 & n53180 ;
  assign n53185 = n53183 | n53184 ;
  assign n82551 = ~n53048 ;
  assign n53186 = n82551 & n53185 ;
  assign n82552 = ~n53038 ;
  assign n53187 = x76 & n82552 ;
  assign n82553 = ~n53036 ;
  assign n53188 = n82553 & n53187 ;
  assign n53189 = n53040 | n53188 ;
  assign n53190 = n53186 | n53189 ;
  assign n82554 = ~n53040 ;
  assign n53195 = n82554 & n53190 ;
  assign n53196 = n53193 | n53195 ;
  assign n82555 = ~n53032 ;
  assign n53197 = n82555 & n53196 ;
  assign n82556 = ~n53022 ;
  assign n53198 = x78 & n82556 ;
  assign n82557 = ~n53020 ;
  assign n53199 = n82557 & n53198 ;
  assign n53200 = n53024 | n53199 ;
  assign n53201 = n53197 | n53200 ;
  assign n82558 = ~n53024 ;
  assign n53205 = n82558 & n53201 ;
  assign n53206 = n53204 | n53205 ;
  assign n82559 = ~n53016 ;
  assign n53207 = n82559 & n53206 ;
  assign n82560 = ~n53006 ;
  assign n53208 = x80 & n82560 ;
  assign n82561 = ~n53004 ;
  assign n53209 = n82561 & n53208 ;
  assign n53210 = n53008 | n53209 ;
  assign n53211 = n53207 | n53210 ;
  assign n82562 = ~n53008 ;
  assign n53215 = n82562 & n53211 ;
  assign n53216 = n53214 | n53215 ;
  assign n82563 = ~n53000 ;
  assign n53217 = n82563 & n53216 ;
  assign n82564 = ~n52990 ;
  assign n53218 = x82 & n82564 ;
  assign n82565 = ~n52988 ;
  assign n53219 = n82565 & n53218 ;
  assign n53220 = n52992 | n53219 ;
  assign n53221 = n53217 | n53220 ;
  assign n82566 = ~n52992 ;
  assign n53226 = n82566 & n53221 ;
  assign n53227 = n53224 | n53226 ;
  assign n82567 = ~n52984 ;
  assign n53228 = n82567 & n53227 ;
  assign n82568 = ~n52974 ;
  assign n53229 = x84 & n82568 ;
  assign n82569 = ~n52972 ;
  assign n53230 = n82569 & n53229 ;
  assign n53231 = n52976 | n53230 ;
  assign n53232 = n53228 | n53231 ;
  assign n82570 = ~n52976 ;
  assign n53236 = n82570 & n53232 ;
  assign n53237 = n53235 | n53236 ;
  assign n82571 = ~n52968 ;
  assign n53238 = n82571 & n53237 ;
  assign n82572 = ~n52958 ;
  assign n53239 = x86 & n82572 ;
  assign n82573 = ~n52956 ;
  assign n53240 = n82573 & n53239 ;
  assign n53241 = n52960 | n53240 ;
  assign n53242 = n53238 | n53241 ;
  assign n82574 = ~n52960 ;
  assign n53246 = n82574 & n53242 ;
  assign n53247 = n53245 | n53246 ;
  assign n82575 = ~n52952 ;
  assign n53248 = n82575 & n53247 ;
  assign n82576 = ~n52942 ;
  assign n53249 = x88 & n82576 ;
  assign n82577 = ~n52940 ;
  assign n53250 = n82577 & n53249 ;
  assign n53251 = n52944 | n53250 ;
  assign n53253 = n53248 | n53251 ;
  assign n82578 = ~n52944 ;
  assign n53257 = n82578 & n53253 ;
  assign n53258 = n53256 | n53257 ;
  assign n82579 = ~n52936 ;
  assign n53259 = n82579 & n53258 ;
  assign n82580 = ~n52926 ;
  assign n53260 = x90 & n82580 ;
  assign n82581 = ~n52924 ;
  assign n53261 = n82581 & n53260 ;
  assign n53262 = n52928 | n53261 ;
  assign n53263 = n53259 | n53262 ;
  assign n82582 = ~n52928 ;
  assign n53267 = n82582 & n53263 ;
  assign n53268 = n53266 | n53267 ;
  assign n82583 = ~n52920 ;
  assign n53269 = n82583 & n53268 ;
  assign n82584 = ~n52910 ;
  assign n53270 = x92 & n82584 ;
  assign n82585 = ~n52908 ;
  assign n53271 = n82585 & n53270 ;
  assign n53272 = n52912 | n53271 ;
  assign n53273 = n53269 | n53272 ;
  assign n82586 = ~n52912 ;
  assign n53277 = n82586 & n53273 ;
  assign n53278 = n53276 | n53277 ;
  assign n82587 = ~n52904 ;
  assign n53279 = n82587 & n53278 ;
  assign n82588 = ~n52894 ;
  assign n53280 = x94 & n82588 ;
  assign n82589 = ~n52892 ;
  assign n53281 = n82589 & n53280 ;
  assign n53282 = n52896 | n53281 ;
  assign n53283 = n53279 | n53282 ;
  assign n82590 = ~n52896 ;
  assign n53287 = n82590 & n53283 ;
  assign n53288 = n53286 | n53287 ;
  assign n82591 = ~n52888 ;
  assign n53289 = n82591 & n53288 ;
  assign n82592 = ~n52878 ;
  assign n53290 = x96 & n82592 ;
  assign n82593 = ~n52876 ;
  assign n53291 = n82593 & n53290 ;
  assign n53292 = n52880 | n53291 ;
  assign n53293 = n53289 | n53292 ;
  assign n82594 = ~n52880 ;
  assign n53297 = n82594 & n53293 ;
  assign n53298 = n53296 | n53297 ;
  assign n82595 = ~n52872 ;
  assign n53299 = n82595 & n53298 ;
  assign n82596 = ~n52862 ;
  assign n53300 = x98 & n82596 ;
  assign n82597 = ~n52860 ;
  assign n53301 = n82597 & n53300 ;
  assign n53302 = n52864 | n53301 ;
  assign n53303 = n53299 | n53302 ;
  assign n82598 = ~n52864 ;
  assign n53307 = n82598 & n53303 ;
  assign n53308 = n53306 | n53307 ;
  assign n82599 = ~n52856 ;
  assign n53309 = n82599 & n53308 ;
  assign n82600 = ~n52846 ;
  assign n53310 = x100 & n82600 ;
  assign n82601 = ~n52844 ;
  assign n53311 = n82601 & n53310 ;
  assign n53312 = n52848 | n53311 ;
  assign n53313 = n53309 | n53312 ;
  assign n82602 = ~n52848 ;
  assign n53317 = n82602 & n53313 ;
  assign n53318 = n53316 | n53317 ;
  assign n82603 = ~n52840 ;
  assign n53319 = n82603 & n53318 ;
  assign n82604 = ~n52830 ;
  assign n53320 = x102 & n82604 ;
  assign n82605 = ~n52828 ;
  assign n53321 = n82605 & n53320 ;
  assign n53322 = n52832 | n53321 ;
  assign n53323 = n53319 | n53322 ;
  assign n82606 = ~n52832 ;
  assign n53327 = n82606 & n53323 ;
  assign n53328 = n53326 | n53327 ;
  assign n82607 = ~n52824 ;
  assign n53329 = n82607 & n53328 ;
  assign n82608 = ~n52814 ;
  assign n53330 = x104 & n82608 ;
  assign n82609 = ~n52812 ;
  assign n53331 = n82609 & n53330 ;
  assign n53332 = n52816 | n53331 ;
  assign n53333 = n53329 | n53332 ;
  assign n82610 = ~n52816 ;
  assign n53337 = n82610 & n53333 ;
  assign n53338 = n53336 | n53337 ;
  assign n82611 = ~n52808 ;
  assign n53339 = n82611 & n53338 ;
  assign n82612 = ~n52798 ;
  assign n53340 = x106 & n82612 ;
  assign n82613 = ~n52796 ;
  assign n53341 = n82613 & n53340 ;
  assign n53342 = n52800 | n53341 ;
  assign n53343 = n53339 | n53342 ;
  assign n82614 = ~n52800 ;
  assign n53347 = n82614 & n53343 ;
  assign n53348 = n53346 | n53347 ;
  assign n82615 = ~n52792 ;
  assign n53349 = n82615 & n53348 ;
  assign n82616 = ~n52782 ;
  assign n53350 = x108 & n82616 ;
  assign n82617 = ~n52780 ;
  assign n53351 = n82617 & n53350 ;
  assign n53352 = n52784 | n53351 ;
  assign n53353 = n53349 | n53352 ;
  assign n82618 = ~n52784 ;
  assign n53357 = n82618 & n53353 ;
  assign n53358 = n53356 | n53357 ;
  assign n82619 = ~n52776 ;
  assign n53359 = n82619 & n53358 ;
  assign n82620 = ~n52766 ;
  assign n53360 = x110 & n82620 ;
  assign n82621 = ~n52764 ;
  assign n53361 = n82621 & n53360 ;
  assign n53362 = n52768 | n53361 ;
  assign n53363 = n53359 | n53362 ;
  assign n82622 = ~n52768 ;
  assign n53367 = n82622 & n53363 ;
  assign n53368 = n53366 | n53367 ;
  assign n82623 = ~n52760 ;
  assign n53369 = n82623 & n53368 ;
  assign n82624 = ~n52750 ;
  assign n53370 = x112 & n82624 ;
  assign n82625 = ~n52748 ;
  assign n53371 = n82625 & n53370 ;
  assign n53372 = n52752 | n53371 ;
  assign n53373 = n53369 | n53372 ;
  assign n82626 = ~n52752 ;
  assign n53377 = n82626 & n53373 ;
  assign n53378 = n53376 | n53377 ;
  assign n82627 = ~n52744 ;
  assign n53379 = n82627 & n53378 ;
  assign n53380 = n51951 | n52604 ;
  assign n53381 = n52600 | n53380 ;
  assign n82628 = ~n53381 ;
  assign n53382 = n52592 & n82628 ;
  assign n53383 = n52600 | n52604 ;
  assign n82629 = ~n52739 ;
  assign n53384 = n82629 & n53383 ;
  assign n53385 = n53382 | n53384 ;
  assign n53386 = n82385 & n53385 ;
  assign n53387 = n279 & n51189 ;
  assign n53388 = n52740 & n53387 ;
  assign n53389 = n53386 | n53388 ;
  assign n53390 = n72385 & n53389 ;
  assign n82630 = ~n53388 ;
  assign n53391 = x114 & n82630 ;
  assign n82631 = ~n53386 ;
  assign n53392 = n82631 & n53391 ;
  assign n53393 = n21184 | n53392 ;
  assign n53394 = n53390 | n53393 ;
  assign n53395 = n53379 | n53394 ;
  assign n53396 = n72139 & n53389 ;
  assign n82632 = ~n53396 ;
  assign n53397 = n53395 & n82632 ;
  assign n82633 = ~n53377 ;
  assign n53497 = n53376 & n82633 ;
  assign n53398 = x65 & n53133 ;
  assign n82634 = ~n53398 ;
  assign n53399 = n53130 & n82634 ;
  assign n53400 = n20903 | n53399 ;
  assign n53402 = n82531 & n53400 ;
  assign n53403 = n53138 | n53402 ;
  assign n53404 = n82534 & n53403 ;
  assign n53405 = n53142 | n53404 ;
  assign n53406 = n82535 & n53405 ;
  assign n53407 = n53148 | n53406 ;
  assign n53408 = n82538 & n53407 ;
  assign n53409 = n53152 | n53408 ;
  assign n53410 = n82539 & n53409 ;
  assign n53411 = n53158 | n53410 ;
  assign n53412 = n82542 & n53411 ;
  assign n53413 = n53162 | n53412 ;
  assign n53414 = n82543 & n53413 ;
  assign n53415 = n53168 | n53414 ;
  assign n53416 = n82546 & n53415 ;
  assign n53417 = n53172 | n53416 ;
  assign n53418 = n82547 & n53417 ;
  assign n53419 = n53178 | n53418 ;
  assign n53420 = n82550 & n53419 ;
  assign n53421 = n53183 | n53420 ;
  assign n53422 = n82551 & n53421 ;
  assign n53423 = n53189 | n53422 ;
  assign n53424 = n82554 & n53423 ;
  assign n53425 = n53193 | n53424 ;
  assign n53426 = n82555 & n53425 ;
  assign n53427 = n53200 | n53426 ;
  assign n53428 = n82558 & n53427 ;
  assign n53429 = n53204 | n53428 ;
  assign n53430 = n82559 & n53429 ;
  assign n53431 = n53210 | n53430 ;
  assign n53432 = n82562 & n53431 ;
  assign n53433 = n53214 | n53432 ;
  assign n53434 = n82563 & n53433 ;
  assign n53435 = n53220 | n53434 ;
  assign n53436 = n82566 & n53435 ;
  assign n53437 = n53224 | n53436 ;
  assign n53438 = n82567 & n53437 ;
  assign n53439 = n53231 | n53438 ;
  assign n53440 = n82570 & n53439 ;
  assign n53441 = n53235 | n53440 ;
  assign n53442 = n82571 & n53441 ;
  assign n53443 = n53241 | n53442 ;
  assign n53444 = n82574 & n53443 ;
  assign n53445 = n53245 | n53444 ;
  assign n53446 = n82575 & n53445 ;
  assign n53447 = n53251 | n53446 ;
  assign n53448 = n82578 & n53447 ;
  assign n53449 = n53256 | n53448 ;
  assign n53450 = n82579 & n53449 ;
  assign n53451 = n53262 | n53450 ;
  assign n53452 = n82582 & n53451 ;
  assign n53453 = n53266 | n53452 ;
  assign n53454 = n82583 & n53453 ;
  assign n53455 = n53272 | n53454 ;
  assign n53456 = n82586 & n53455 ;
  assign n53457 = n53276 | n53456 ;
  assign n53458 = n82587 & n53457 ;
  assign n53459 = n53282 | n53458 ;
  assign n53460 = n82590 & n53459 ;
  assign n53461 = n53286 | n53460 ;
  assign n53462 = n82591 & n53461 ;
  assign n53463 = n53292 | n53462 ;
  assign n53464 = n82594 & n53463 ;
  assign n53465 = n53296 | n53464 ;
  assign n53466 = n82595 & n53465 ;
  assign n53467 = n53302 | n53466 ;
  assign n53468 = n82598 & n53467 ;
  assign n53469 = n53306 | n53468 ;
  assign n53470 = n82599 & n53469 ;
  assign n53471 = n53312 | n53470 ;
  assign n53472 = n82602 & n53471 ;
  assign n53473 = n53316 | n53472 ;
  assign n53474 = n82603 & n53473 ;
  assign n53475 = n53322 | n53474 ;
  assign n53476 = n82606 & n53475 ;
  assign n53477 = n53326 | n53476 ;
  assign n53478 = n82607 & n53477 ;
  assign n53479 = n53332 | n53478 ;
  assign n53480 = n82610 & n53479 ;
  assign n53481 = n53336 | n53480 ;
  assign n53482 = n82611 & n53481 ;
  assign n53483 = n53342 | n53482 ;
  assign n53484 = n82614 & n53483 ;
  assign n53485 = n53346 | n53484 ;
  assign n53486 = n82615 & n53485 ;
  assign n53487 = n53352 | n53486 ;
  assign n53488 = n82618 & n53487 ;
  assign n53489 = n53356 | n53488 ;
  assign n53490 = n82619 & n53489 ;
  assign n53491 = n53362 | n53490 ;
  assign n53492 = n82622 & n53491 ;
  assign n53493 = n53366 | n53492 ;
  assign n53494 = n82623 & n53493 ;
  assign n53495 = n53372 | n53494 ;
  assign n53498 = n52752 | n53376 ;
  assign n82635 = ~n53498 ;
  assign n53499 = n53495 & n82635 ;
  assign n53500 = n53497 | n53499 ;
  assign n82636 = ~n53397 ;
  assign n53501 = n82636 & n53500 ;
  assign n53502 = n52743 & n82632 ;
  assign n53503 = n53395 & n53502 ;
  assign n53504 = n53501 | n53503 ;
  assign n53505 = n52744 | n53392 ;
  assign n53506 = n53390 | n53505 ;
  assign n82637 = ~n53506 ;
  assign n53507 = n53378 & n82637 ;
  assign n53496 = n82626 & n53495 ;
  assign n53508 = n53376 | n53496 ;
  assign n53509 = n82627 & n53508 ;
  assign n53510 = n53390 | n53392 ;
  assign n82638 = ~n53509 ;
  assign n53511 = n82638 & n53510 ;
  assign n53512 = n53507 | n53511 ;
  assign n53513 = n82636 & n53512 ;
  assign n53514 = n20358 & n53389 ;
  assign n53515 = n53395 & n53514 ;
  assign n53516 = n53513 | n53515 ;
  assign n53517 = n72393 & n53516 ;
  assign n53518 = n72385 & n53504 ;
  assign n82639 = ~n53494 ;
  assign n53519 = n53372 & n82639 ;
  assign n53520 = n52760 | n53372 ;
  assign n82640 = ~n53520 ;
  assign n53521 = n53368 & n82640 ;
  assign n53522 = n53519 | n53521 ;
  assign n53523 = n82636 & n53522 ;
  assign n53524 = n52751 & n82632 ;
  assign n53525 = n53395 & n53524 ;
  assign n53526 = n53523 | n53525 ;
  assign n53527 = n72025 & n53526 ;
  assign n82641 = ~n53367 ;
  assign n53528 = n53366 & n82641 ;
  assign n53529 = n52768 | n53366 ;
  assign n82642 = ~n53529 ;
  assign n53530 = n53491 & n82642 ;
  assign n53531 = n53528 | n53530 ;
  assign n53532 = n82636 & n53531 ;
  assign n53533 = n52759 & n82632 ;
  assign n53534 = n53395 & n53533 ;
  assign n53535 = n53532 | n53534 ;
  assign n53536 = n71645 & n53535 ;
  assign n82643 = ~n53490 ;
  assign n53537 = n53362 & n82643 ;
  assign n53538 = n52776 | n53362 ;
  assign n82644 = ~n53538 ;
  assign n53539 = n53358 & n82644 ;
  assign n53540 = n53537 | n53539 ;
  assign n53541 = n82636 & n53540 ;
  assign n53542 = n52767 & n82632 ;
  assign n53543 = n53395 & n53542 ;
  assign n53544 = n53541 | n53543 ;
  assign n53545 = n71633 & n53544 ;
  assign n82645 = ~n53357 ;
  assign n53546 = n53356 & n82645 ;
  assign n53547 = n52784 | n53356 ;
  assign n82646 = ~n53547 ;
  assign n53548 = n53487 & n82646 ;
  assign n53549 = n53546 | n53548 ;
  assign n53550 = n82636 & n53549 ;
  assign n53551 = n52775 & n82632 ;
  assign n53552 = n53395 & n53551 ;
  assign n53553 = n53550 | n53552 ;
  assign n53554 = n71253 & n53553 ;
  assign n82647 = ~n53486 ;
  assign n53555 = n53352 & n82647 ;
  assign n53556 = n52792 | n53352 ;
  assign n82648 = ~n53556 ;
  assign n53557 = n53348 & n82648 ;
  assign n53558 = n53555 | n53557 ;
  assign n53559 = n82636 & n53558 ;
  assign n53560 = n52783 & n82632 ;
  assign n53561 = n53395 & n53560 ;
  assign n53562 = n53559 | n53561 ;
  assign n53563 = n70935 & n53562 ;
  assign n82649 = ~n53347 ;
  assign n53564 = n53346 & n82649 ;
  assign n53565 = n52800 | n53346 ;
  assign n82650 = ~n53565 ;
  assign n53566 = n53483 & n82650 ;
  assign n53567 = n53564 | n53566 ;
  assign n53568 = n82636 & n53567 ;
  assign n53569 = n52791 & n82632 ;
  assign n53570 = n53395 & n53569 ;
  assign n53571 = n53568 | n53570 ;
  assign n53572 = n70927 & n53571 ;
  assign n82651 = ~n53482 ;
  assign n53573 = n53342 & n82651 ;
  assign n53574 = n52808 | n53342 ;
  assign n82652 = ~n53574 ;
  assign n53575 = n53338 & n82652 ;
  assign n53576 = n53573 | n53575 ;
  assign n53577 = n82636 & n53576 ;
  assign n53578 = n52799 & n82632 ;
  assign n53579 = n53395 & n53578 ;
  assign n53580 = n53577 | n53579 ;
  assign n53581 = n70609 & n53580 ;
  assign n82653 = ~n53337 ;
  assign n53582 = n53336 & n82653 ;
  assign n53583 = n52816 | n53336 ;
  assign n82654 = ~n53583 ;
  assign n53584 = n53479 & n82654 ;
  assign n53585 = n53582 | n53584 ;
  assign n53586 = n82636 & n53585 ;
  assign n53587 = n52807 & n82632 ;
  assign n53588 = n53395 & n53587 ;
  assign n53589 = n53586 | n53588 ;
  assign n53590 = n70276 & n53589 ;
  assign n82655 = ~n53478 ;
  assign n53591 = n53332 & n82655 ;
  assign n53592 = n52824 | n53332 ;
  assign n82656 = ~n53592 ;
  assign n53593 = n53328 & n82656 ;
  assign n53594 = n53591 | n53593 ;
  assign n53595 = n82636 & n53594 ;
  assign n53596 = n52815 & n82632 ;
  assign n53597 = n53395 & n53596 ;
  assign n53598 = n53595 | n53597 ;
  assign n53599 = n70176 & n53598 ;
  assign n82657 = ~n53327 ;
  assign n53600 = n53326 & n82657 ;
  assign n53601 = n52832 | n53326 ;
  assign n82658 = ~n53601 ;
  assign n53602 = n53475 & n82658 ;
  assign n53603 = n53600 | n53602 ;
  assign n53604 = n82636 & n53603 ;
  assign n53605 = n52823 & n82632 ;
  assign n53606 = n53395 & n53605 ;
  assign n53607 = n53604 | n53606 ;
  assign n53608 = n69857 & n53607 ;
  assign n82659 = ~n53474 ;
  assign n53609 = n53322 & n82659 ;
  assign n53610 = n52840 | n53322 ;
  assign n82660 = ~n53610 ;
  assign n53611 = n53318 & n82660 ;
  assign n53612 = n53609 | n53611 ;
  assign n53613 = n82636 & n53612 ;
  assign n53614 = n52831 & n82632 ;
  assign n53615 = n53395 & n53614 ;
  assign n53616 = n53613 | n53615 ;
  assign n53617 = n69656 & n53616 ;
  assign n82661 = ~n53317 ;
  assign n53618 = n53316 & n82661 ;
  assign n53619 = n52848 | n53316 ;
  assign n82662 = ~n53619 ;
  assign n53620 = n53471 & n82662 ;
  assign n53621 = n53618 | n53620 ;
  assign n53622 = n82636 & n53621 ;
  assign n53623 = n52839 & n82632 ;
  assign n53624 = n53395 & n53623 ;
  assign n53625 = n53622 | n53624 ;
  assign n53626 = n69528 & n53625 ;
  assign n82663 = ~n53470 ;
  assign n53627 = n53312 & n82663 ;
  assign n53628 = n52856 | n53312 ;
  assign n82664 = ~n53628 ;
  assign n53629 = n53308 & n82664 ;
  assign n53630 = n53627 | n53629 ;
  assign n53631 = n82636 & n53630 ;
  assign n53632 = n52847 & n82632 ;
  assign n53633 = n53395 & n53632 ;
  assign n53634 = n53631 | n53633 ;
  assign n53635 = n69261 & n53634 ;
  assign n82665 = ~n53307 ;
  assign n53636 = n53306 & n82665 ;
  assign n53637 = n52864 | n53306 ;
  assign n82666 = ~n53637 ;
  assign n53638 = n53467 & n82666 ;
  assign n53639 = n53636 | n53638 ;
  assign n53640 = n82636 & n53639 ;
  assign n53641 = n52855 & n82632 ;
  assign n53642 = n53395 & n53641 ;
  assign n53643 = n53640 | n53642 ;
  assign n53644 = n69075 & n53643 ;
  assign n82667 = ~n53466 ;
  assign n53645 = n53302 & n82667 ;
  assign n53646 = n52872 | n53302 ;
  assign n82668 = ~n53646 ;
  assign n53647 = n53298 & n82668 ;
  assign n53648 = n53645 | n53647 ;
  assign n53649 = n82636 & n53648 ;
  assign n53650 = n52863 & n82632 ;
  assign n53651 = n53395 & n53650 ;
  assign n53652 = n53649 | n53651 ;
  assign n53653 = n68993 & n53652 ;
  assign n82669 = ~n53297 ;
  assign n53654 = n53296 & n82669 ;
  assign n53655 = n52880 | n53296 ;
  assign n82670 = ~n53655 ;
  assign n53656 = n53463 & n82670 ;
  assign n53657 = n53654 | n53656 ;
  assign n53658 = n82636 & n53657 ;
  assign n53659 = n52871 & n82632 ;
  assign n53660 = n53395 & n53659 ;
  assign n53661 = n53658 | n53660 ;
  assign n53662 = n68716 & n53661 ;
  assign n82671 = ~n53462 ;
  assign n53663 = n53292 & n82671 ;
  assign n53664 = n52888 | n53292 ;
  assign n82672 = ~n53664 ;
  assign n53665 = n53288 & n82672 ;
  assign n53666 = n53663 | n53665 ;
  assign n53667 = n82636 & n53666 ;
  assign n53668 = n52879 & n82632 ;
  assign n53669 = n53395 & n53668 ;
  assign n53670 = n53667 | n53669 ;
  assign n53671 = n68545 & n53670 ;
  assign n82673 = ~n53287 ;
  assign n53672 = n53286 & n82673 ;
  assign n53673 = n52896 | n53286 ;
  assign n82674 = ~n53673 ;
  assign n53674 = n53459 & n82674 ;
  assign n53675 = n53672 | n53674 ;
  assign n53676 = n82636 & n53675 ;
  assign n53677 = n52887 & n82632 ;
  assign n53678 = n53395 & n53677 ;
  assign n53679 = n53676 | n53678 ;
  assign n53680 = n68438 & n53679 ;
  assign n82675 = ~n53458 ;
  assign n53681 = n53282 & n82675 ;
  assign n53682 = n52904 | n53282 ;
  assign n82676 = ~n53682 ;
  assign n53683 = n53278 & n82676 ;
  assign n53684 = n53681 | n53683 ;
  assign n53685 = n82636 & n53684 ;
  assign n53686 = n52895 & n82632 ;
  assign n53687 = n53395 & n53686 ;
  assign n53688 = n53685 | n53687 ;
  assign n53689 = n68214 & n53688 ;
  assign n82677 = ~n53277 ;
  assign n53690 = n53276 & n82677 ;
  assign n53691 = n52912 | n53276 ;
  assign n82678 = ~n53691 ;
  assign n53692 = n53455 & n82678 ;
  assign n53693 = n53690 | n53692 ;
  assign n53694 = n82636 & n53693 ;
  assign n53695 = n52903 & n82632 ;
  assign n53696 = n53395 & n53695 ;
  assign n53697 = n53694 | n53696 ;
  assign n53698 = n68058 & n53697 ;
  assign n82679 = ~n53454 ;
  assign n53699 = n53272 & n82679 ;
  assign n53700 = n52920 | n53272 ;
  assign n82680 = ~n53700 ;
  assign n53701 = n53268 & n82680 ;
  assign n53702 = n53699 | n53701 ;
  assign n53703 = n82636 & n53702 ;
  assign n53704 = n52911 & n82632 ;
  assign n53705 = n53395 & n53704 ;
  assign n53706 = n53703 | n53705 ;
  assign n53707 = n67986 & n53706 ;
  assign n82681 = ~n53267 ;
  assign n53708 = n53266 & n82681 ;
  assign n53709 = n52928 | n53266 ;
  assign n82682 = ~n53709 ;
  assign n53710 = n53451 & n82682 ;
  assign n53711 = n53708 | n53710 ;
  assign n53712 = n82636 & n53711 ;
  assign n53713 = n52919 & n82632 ;
  assign n53714 = n53395 & n53713 ;
  assign n53715 = n53712 | n53714 ;
  assign n53716 = n67763 & n53715 ;
  assign n82683 = ~n53450 ;
  assign n53717 = n53262 & n82683 ;
  assign n53718 = n52936 | n53262 ;
  assign n82684 = ~n53718 ;
  assign n53719 = n53258 & n82684 ;
  assign n53720 = n53717 | n53719 ;
  assign n53721 = n82636 & n53720 ;
  assign n53722 = n52927 & n82632 ;
  assign n53723 = n53395 & n53722 ;
  assign n53724 = n53721 | n53723 ;
  assign n53725 = n67622 & n53724 ;
  assign n82685 = ~n53257 ;
  assign n53726 = n53256 & n82685 ;
  assign n53727 = n52944 | n53256 ;
  assign n82686 = ~n53727 ;
  assign n53728 = n53447 & n82686 ;
  assign n53729 = n53726 | n53728 ;
  assign n53730 = n82636 & n53729 ;
  assign n53731 = n52935 & n82632 ;
  assign n53732 = n53395 & n53731 ;
  assign n53733 = n53730 | n53732 ;
  assign n53734 = n67531 & n53733 ;
  assign n82687 = ~n53446 ;
  assign n53736 = n53251 & n82687 ;
  assign n53252 = n52952 | n53251 ;
  assign n82688 = ~n53252 ;
  assign n53737 = n82688 & n53445 ;
  assign n53738 = n53736 | n53737 ;
  assign n53739 = n82636 & n53738 ;
  assign n53740 = n52943 & n82632 ;
  assign n53741 = n53395 & n53740 ;
  assign n53742 = n53739 | n53741 ;
  assign n53743 = n67348 & n53742 ;
  assign n82689 = ~n53246 ;
  assign n53744 = n53245 & n82689 ;
  assign n53745 = n52960 | n53245 ;
  assign n82690 = ~n53745 ;
  assign n53746 = n53443 & n82690 ;
  assign n53747 = n53744 | n53746 ;
  assign n53748 = n82636 & n53747 ;
  assign n53749 = n52951 & n82632 ;
  assign n53750 = n53395 & n53749 ;
  assign n53751 = n53748 | n53750 ;
  assign n53752 = n67222 & n53751 ;
  assign n82691 = ~n53442 ;
  assign n53753 = n53241 & n82691 ;
  assign n53754 = n52968 | n53241 ;
  assign n82692 = ~n53754 ;
  assign n53755 = n53237 & n82692 ;
  assign n53756 = n53753 | n53755 ;
  assign n53757 = n82636 & n53756 ;
  assign n53758 = n52959 & n82632 ;
  assign n53759 = n53395 & n53758 ;
  assign n53760 = n53757 | n53759 ;
  assign n53761 = n67164 & n53760 ;
  assign n82693 = ~n53236 ;
  assign n53762 = n53235 & n82693 ;
  assign n53763 = n52976 | n53235 ;
  assign n82694 = ~n53763 ;
  assign n53764 = n53439 & n82694 ;
  assign n53765 = n53762 | n53764 ;
  assign n53766 = n82636 & n53765 ;
  assign n53767 = n52967 & n82632 ;
  assign n53768 = n53395 & n53767 ;
  assign n53769 = n53766 | n53768 ;
  assign n53770 = n66979 & n53769 ;
  assign n82695 = ~n53438 ;
  assign n53771 = n53231 & n82695 ;
  assign n53772 = n52984 | n53231 ;
  assign n82696 = ~n53772 ;
  assign n53773 = n53227 & n82696 ;
  assign n53774 = n53771 | n53773 ;
  assign n53775 = n82636 & n53774 ;
  assign n53776 = n52975 & n82632 ;
  assign n53777 = n53395 & n53776 ;
  assign n53778 = n53775 | n53777 ;
  assign n53779 = n66868 & n53778 ;
  assign n82697 = ~n53226 ;
  assign n53780 = n53224 & n82697 ;
  assign n53225 = n52992 | n53224 ;
  assign n82698 = ~n53225 ;
  assign n53781 = n53221 & n82698 ;
  assign n53782 = n53780 | n53781 ;
  assign n53783 = n82636 & n53782 ;
  assign n53784 = n52983 & n82632 ;
  assign n53785 = n53395 & n53784 ;
  assign n53786 = n53783 | n53785 ;
  assign n53787 = n66797 & n53786 ;
  assign n82699 = ~n53434 ;
  assign n53788 = n53220 & n82699 ;
  assign n53789 = n53000 | n53220 ;
  assign n82700 = ~n53789 ;
  assign n53790 = n53216 & n82700 ;
  assign n53791 = n53788 | n53790 ;
  assign n53792 = n82636 & n53791 ;
  assign n53793 = n52991 & n82632 ;
  assign n53794 = n53395 & n53793 ;
  assign n53795 = n53792 | n53794 ;
  assign n53796 = n66654 & n53795 ;
  assign n82701 = ~n53215 ;
  assign n53797 = n53214 & n82701 ;
  assign n53798 = n53008 | n53214 ;
  assign n82702 = ~n53798 ;
  assign n53799 = n53431 & n82702 ;
  assign n53800 = n53797 | n53799 ;
  assign n53801 = n82636 & n53800 ;
  assign n53802 = n52999 & n82632 ;
  assign n53803 = n53395 & n53802 ;
  assign n53804 = n53801 | n53803 ;
  assign n53805 = n66560 & n53804 ;
  assign n82703 = ~n53430 ;
  assign n53806 = n53210 & n82703 ;
  assign n53807 = n53016 | n53210 ;
  assign n82704 = ~n53807 ;
  assign n53808 = n53206 & n82704 ;
  assign n53809 = n53806 | n53808 ;
  assign n53810 = n82636 & n53809 ;
  assign n53811 = n53007 & n82632 ;
  assign n53812 = n53395 & n53811 ;
  assign n53813 = n53810 | n53812 ;
  assign n53814 = n66505 & n53813 ;
  assign n82705 = ~n53205 ;
  assign n53815 = n53204 & n82705 ;
  assign n53816 = n53024 | n53204 ;
  assign n82706 = ~n53816 ;
  assign n53817 = n53427 & n82706 ;
  assign n53818 = n53815 | n53817 ;
  assign n53819 = n82636 & n53818 ;
  assign n53820 = n53015 & n82632 ;
  assign n53821 = n53395 & n53820 ;
  assign n53822 = n53819 | n53821 ;
  assign n53823 = n66379 & n53822 ;
  assign n82707 = ~n53426 ;
  assign n53824 = n53200 & n82707 ;
  assign n53825 = n53032 | n53200 ;
  assign n82708 = ~n53825 ;
  assign n53826 = n53196 & n82708 ;
  assign n53827 = n53824 | n53826 ;
  assign n53828 = n82636 & n53827 ;
  assign n53829 = n53023 & n82632 ;
  assign n53830 = n53395 & n53829 ;
  assign n53831 = n53828 | n53830 ;
  assign n53832 = n66299 & n53831 ;
  assign n82709 = ~n53195 ;
  assign n53833 = n53193 & n82709 ;
  assign n53194 = n53040 | n53193 ;
  assign n82710 = ~n53194 ;
  assign n53834 = n53190 & n82710 ;
  assign n53835 = n53833 | n53834 ;
  assign n53836 = n82636 & n53835 ;
  assign n53837 = n53031 & n82632 ;
  assign n53838 = n53395 & n53837 ;
  assign n53839 = n53836 | n53838 ;
  assign n53840 = n66244 & n53839 ;
  assign n82711 = ~n53422 ;
  assign n53841 = n53189 & n82711 ;
  assign n53842 = n53048 | n53189 ;
  assign n82712 = ~n53842 ;
  assign n53843 = n53185 & n82712 ;
  assign n53844 = n53841 | n53843 ;
  assign n53845 = n82636 & n53844 ;
  assign n53846 = n53039 & n82632 ;
  assign n53847 = n53395 & n53846 ;
  assign n53848 = n53845 | n53847 ;
  assign n53849 = n66145 & n53848 ;
  assign n82713 = ~n53184 ;
  assign n53850 = n53183 & n82713 ;
  assign n53851 = n53056 | n53183 ;
  assign n82714 = ~n53851 ;
  assign n53852 = n53419 & n82714 ;
  assign n53853 = n53850 | n53852 ;
  assign n53854 = n82636 & n53853 ;
  assign n53855 = n53047 & n82632 ;
  assign n53856 = n53395 & n53855 ;
  assign n53857 = n53854 | n53856 ;
  assign n53858 = n66081 & n53857 ;
  assign n82715 = ~n53418 ;
  assign n53859 = n53178 & n82715 ;
  assign n53179 = n53064 | n53178 ;
  assign n82716 = ~n53179 ;
  assign n53860 = n82716 & n53417 ;
  assign n53861 = n53859 | n53860 ;
  assign n53862 = n82636 & n53861 ;
  assign n53863 = n53055 & n82632 ;
  assign n53864 = n53395 & n53863 ;
  assign n53865 = n53862 | n53864 ;
  assign n53866 = n66043 & n53865 ;
  assign n82717 = ~n53173 ;
  assign n53867 = n53172 & n82717 ;
  assign n53868 = n53072 | n53172 ;
  assign n82718 = ~n53868 ;
  assign n53869 = n53415 & n82718 ;
  assign n53870 = n53867 | n53869 ;
  assign n53871 = n82636 & n53870 ;
  assign n53872 = n53063 & n82632 ;
  assign n53873 = n53395 & n53872 ;
  assign n53874 = n53871 | n53873 ;
  assign n53875 = n65960 & n53874 ;
  assign n82719 = ~n53414 ;
  assign n53876 = n53168 & n82719 ;
  assign n53877 = n53080 | n53168 ;
  assign n82720 = ~n53877 ;
  assign n53878 = n53164 & n82720 ;
  assign n53879 = n53876 | n53878 ;
  assign n53880 = n82636 & n53879 ;
  assign n53881 = n53071 & n82632 ;
  assign n53882 = n53395 & n53881 ;
  assign n53883 = n53880 | n53882 ;
  assign n53884 = n65909 & n53883 ;
  assign n82721 = ~n53163 ;
  assign n53885 = n53162 & n82721 ;
  assign n53886 = n53088 | n53162 ;
  assign n82722 = ~n53886 ;
  assign n53887 = n53411 & n82722 ;
  assign n53888 = n53885 | n53887 ;
  assign n53889 = n82636 & n53888 ;
  assign n53890 = n53079 & n82632 ;
  assign n53891 = n53395 & n53890 ;
  assign n53892 = n53889 | n53891 ;
  assign n53893 = n65877 & n53892 ;
  assign n82723 = ~n53410 ;
  assign n53894 = n53158 & n82723 ;
  assign n53895 = n53097 | n53158 ;
  assign n82724 = ~n53895 ;
  assign n53896 = n53154 & n82724 ;
  assign n53897 = n53894 | n53896 ;
  assign n53898 = n82636 & n53897 ;
  assign n53899 = n53087 & n82632 ;
  assign n53900 = n53395 & n53899 ;
  assign n53901 = n53898 | n53900 ;
  assign n53902 = n65820 & n53901 ;
  assign n82725 = ~n53153 ;
  assign n53903 = n53152 & n82725 ;
  assign n53904 = n53105 | n53152 ;
  assign n82726 = ~n53904 ;
  assign n53905 = n53407 & n82726 ;
  assign n53906 = n53903 | n53905 ;
  assign n53907 = n82636 & n53906 ;
  assign n53908 = n53096 & n82632 ;
  assign n53909 = n53395 & n53908 ;
  assign n53910 = n53907 | n53909 ;
  assign n53911 = n65791 & n53910 ;
  assign n82727 = ~n53406 ;
  assign n53912 = n53148 & n82727 ;
  assign n53913 = n53113 | n53148 ;
  assign n82728 = ~n53913 ;
  assign n53914 = n53144 & n82728 ;
  assign n53915 = n53912 | n53914 ;
  assign n53916 = n82636 & n53915 ;
  assign n53917 = n53104 & n82632 ;
  assign n53918 = n53395 & n53917 ;
  assign n53919 = n53916 | n53918 ;
  assign n53920 = n65772 & n53919 ;
  assign n82729 = ~n53143 ;
  assign n53922 = n53142 & n82729 ;
  assign n53921 = n53121 | n53142 ;
  assign n82730 = ~n53921 ;
  assign n53923 = n53139 & n82730 ;
  assign n53924 = n53922 | n53923 ;
  assign n53925 = n82636 & n53924 ;
  assign n53926 = n53112 & n82632 ;
  assign n53927 = n53395 & n53926 ;
  assign n53928 = n53925 | n53927 ;
  assign n53929 = n65746 & n53928 ;
  assign n82731 = ~n53402 ;
  assign n53930 = n53138 & n82731 ;
  assign n53401 = n53134 | n53138 ;
  assign n82732 = ~n53401 ;
  assign n53931 = n53400 & n82732 ;
  assign n53932 = n53930 | n53931 ;
  assign n53933 = n82636 & n53932 ;
  assign n53934 = n53120 & n82632 ;
  assign n53935 = n53395 & n53934 ;
  assign n53936 = n53933 | n53935 ;
  assign n53937 = n65721 & n53936 ;
  assign n53938 = n20903 & n53130 ;
  assign n53939 = n82634 & n53938 ;
  assign n82733 = ~n53939 ;
  assign n53940 = n53400 & n82733 ;
  assign n53941 = n82636 & n53940 ;
  assign n53942 = n53133 & n82632 ;
  assign n53943 = n53395 & n53942 ;
  assign n53944 = n53941 | n53943 ;
  assign n53945 = n65686 & n53944 ;
  assign n53735 = n20903 & n82636 ;
  assign n53950 = x64 & n82636 ;
  assign n82734 = ~n53950 ;
  assign n53951 = x13 & n82734 ;
  assign n53952 = n53735 | n53951 ;
  assign n53954 = x65 & n53952 ;
  assign n53946 = n53394 | n53509 ;
  assign n53947 = n82632 & n53946 ;
  assign n82735 = ~n53947 ;
  assign n53948 = x64 & n82735 ;
  assign n82736 = ~n53948 ;
  assign n53949 = x13 & n82736 ;
  assign n53953 = x65 | n53735 ;
  assign n53955 = n53949 | n53953 ;
  assign n82737 = ~n53954 ;
  assign n53956 = n82737 & n53955 ;
  assign n53957 = n21731 | n53956 ;
  assign n53958 = n65670 & n53952 ;
  assign n82738 = ~n53958 ;
  assign n53959 = n53957 & n82738 ;
  assign n82739 = ~n53943 ;
  assign n53960 = x66 & n82739 ;
  assign n82740 = ~n53941 ;
  assign n53961 = n82740 & n53960 ;
  assign n53962 = n53945 | n53961 ;
  assign n53963 = n53959 | n53962 ;
  assign n82741 = ~n53945 ;
  assign n53964 = n82741 & n53963 ;
  assign n82742 = ~n53935 ;
  assign n53965 = x67 & n82742 ;
  assign n82743 = ~n53933 ;
  assign n53966 = n82743 & n53965 ;
  assign n53967 = n53964 | n53966 ;
  assign n82744 = ~n53937 ;
  assign n53968 = n82744 & n53967 ;
  assign n82745 = ~n53927 ;
  assign n53969 = x68 & n82745 ;
  assign n82746 = ~n53925 ;
  assign n53970 = n82746 & n53969 ;
  assign n53971 = n53929 | n53970 ;
  assign n53972 = n53968 | n53971 ;
  assign n82747 = ~n53929 ;
  assign n53973 = n82747 & n53972 ;
  assign n82748 = ~n53918 ;
  assign n53974 = x69 & n82748 ;
  assign n82749 = ~n53916 ;
  assign n53975 = n82749 & n53974 ;
  assign n53976 = n53973 | n53975 ;
  assign n82750 = ~n53920 ;
  assign n53977 = n82750 & n53976 ;
  assign n82751 = ~n53909 ;
  assign n53978 = x70 & n82751 ;
  assign n82752 = ~n53907 ;
  assign n53979 = n82752 & n53978 ;
  assign n53980 = n53911 | n53979 ;
  assign n53981 = n53977 | n53980 ;
  assign n82753 = ~n53911 ;
  assign n53982 = n82753 & n53981 ;
  assign n82754 = ~n53900 ;
  assign n53983 = x71 & n82754 ;
  assign n82755 = ~n53898 ;
  assign n53984 = n82755 & n53983 ;
  assign n53985 = n53902 | n53984 ;
  assign n53987 = n53982 | n53985 ;
  assign n82756 = ~n53902 ;
  assign n53988 = n82756 & n53987 ;
  assign n82757 = ~n53891 ;
  assign n53989 = x72 & n82757 ;
  assign n82758 = ~n53889 ;
  assign n53990 = n82758 & n53989 ;
  assign n53991 = n53893 | n53990 ;
  assign n53992 = n53988 | n53991 ;
  assign n82759 = ~n53893 ;
  assign n53993 = n82759 & n53992 ;
  assign n82760 = ~n53882 ;
  assign n53994 = x73 & n82760 ;
  assign n82761 = ~n53880 ;
  assign n53995 = n82761 & n53994 ;
  assign n53996 = n53884 | n53995 ;
  assign n53998 = n53993 | n53996 ;
  assign n82762 = ~n53884 ;
  assign n53999 = n82762 & n53998 ;
  assign n82763 = ~n53873 ;
  assign n54000 = x74 & n82763 ;
  assign n82764 = ~n53871 ;
  assign n54001 = n82764 & n54000 ;
  assign n54002 = n53875 | n54001 ;
  assign n54003 = n53999 | n54002 ;
  assign n82765 = ~n53875 ;
  assign n54004 = n82765 & n54003 ;
  assign n82766 = ~n53864 ;
  assign n54005 = x75 & n82766 ;
  assign n82767 = ~n53862 ;
  assign n54006 = n82767 & n54005 ;
  assign n54007 = n53866 | n54006 ;
  assign n54009 = n54004 | n54007 ;
  assign n82768 = ~n53866 ;
  assign n54010 = n82768 & n54009 ;
  assign n82769 = ~n53856 ;
  assign n54011 = x76 & n82769 ;
  assign n82770 = ~n53854 ;
  assign n54012 = n82770 & n54011 ;
  assign n54013 = n53858 | n54012 ;
  assign n54014 = n54010 | n54013 ;
  assign n82771 = ~n53858 ;
  assign n54015 = n82771 & n54014 ;
  assign n82772 = ~n53847 ;
  assign n54016 = x77 & n82772 ;
  assign n82773 = ~n53845 ;
  assign n54017 = n82773 & n54016 ;
  assign n54018 = n53849 | n54017 ;
  assign n54020 = n54015 | n54018 ;
  assign n82774 = ~n53849 ;
  assign n54021 = n82774 & n54020 ;
  assign n82775 = ~n53838 ;
  assign n54022 = x78 & n82775 ;
  assign n82776 = ~n53836 ;
  assign n54023 = n82776 & n54022 ;
  assign n54024 = n53840 | n54023 ;
  assign n54025 = n54021 | n54024 ;
  assign n82777 = ~n53840 ;
  assign n54026 = n82777 & n54025 ;
  assign n82778 = ~n53830 ;
  assign n54027 = x79 & n82778 ;
  assign n82779 = ~n53828 ;
  assign n54028 = n82779 & n54027 ;
  assign n54029 = n53832 | n54028 ;
  assign n54031 = n54026 | n54029 ;
  assign n82780 = ~n53832 ;
  assign n54032 = n82780 & n54031 ;
  assign n82781 = ~n53821 ;
  assign n54033 = x80 & n82781 ;
  assign n82782 = ~n53819 ;
  assign n54034 = n82782 & n54033 ;
  assign n54035 = n53823 | n54034 ;
  assign n54036 = n54032 | n54035 ;
  assign n82783 = ~n53823 ;
  assign n54037 = n82783 & n54036 ;
  assign n82784 = ~n53812 ;
  assign n54038 = x81 & n82784 ;
  assign n82785 = ~n53810 ;
  assign n54039 = n82785 & n54038 ;
  assign n54040 = n53814 | n54039 ;
  assign n54042 = n54037 | n54040 ;
  assign n82786 = ~n53814 ;
  assign n54043 = n82786 & n54042 ;
  assign n82787 = ~n53803 ;
  assign n54044 = x82 & n82787 ;
  assign n82788 = ~n53801 ;
  assign n54045 = n82788 & n54044 ;
  assign n54046 = n53805 | n54045 ;
  assign n54047 = n54043 | n54046 ;
  assign n82789 = ~n53805 ;
  assign n54048 = n82789 & n54047 ;
  assign n82790 = ~n53794 ;
  assign n54049 = x83 & n82790 ;
  assign n82791 = ~n53792 ;
  assign n54050 = n82791 & n54049 ;
  assign n54051 = n53796 | n54050 ;
  assign n54053 = n54048 | n54051 ;
  assign n82792 = ~n53796 ;
  assign n54054 = n82792 & n54053 ;
  assign n82793 = ~n53785 ;
  assign n54055 = x84 & n82793 ;
  assign n82794 = ~n53783 ;
  assign n54056 = n82794 & n54055 ;
  assign n54057 = n53787 | n54056 ;
  assign n54058 = n54054 | n54057 ;
  assign n82795 = ~n53787 ;
  assign n54059 = n82795 & n54058 ;
  assign n82796 = ~n53777 ;
  assign n54060 = x85 & n82796 ;
  assign n82797 = ~n53775 ;
  assign n54061 = n82797 & n54060 ;
  assign n54062 = n53779 | n54061 ;
  assign n54064 = n54059 | n54062 ;
  assign n82798 = ~n53779 ;
  assign n54065 = n82798 & n54064 ;
  assign n82799 = ~n53768 ;
  assign n54066 = x86 & n82799 ;
  assign n82800 = ~n53766 ;
  assign n54067 = n82800 & n54066 ;
  assign n54068 = n53770 | n54067 ;
  assign n54069 = n54065 | n54068 ;
  assign n82801 = ~n53770 ;
  assign n54070 = n82801 & n54069 ;
  assign n82802 = ~n53759 ;
  assign n54071 = x87 & n82802 ;
  assign n82803 = ~n53757 ;
  assign n54072 = n82803 & n54071 ;
  assign n54073 = n53761 | n54072 ;
  assign n54075 = n54070 | n54073 ;
  assign n82804 = ~n53761 ;
  assign n54076 = n82804 & n54075 ;
  assign n82805 = ~n53750 ;
  assign n54077 = x88 & n82805 ;
  assign n82806 = ~n53748 ;
  assign n54078 = n82806 & n54077 ;
  assign n54079 = n53752 | n54078 ;
  assign n54080 = n54076 | n54079 ;
  assign n82807 = ~n53752 ;
  assign n54081 = n82807 & n54080 ;
  assign n82808 = ~n53741 ;
  assign n54082 = x89 & n82808 ;
  assign n82809 = ~n53739 ;
  assign n54083 = n82809 & n54082 ;
  assign n54084 = n53743 | n54083 ;
  assign n54086 = n54081 | n54084 ;
  assign n82810 = ~n53743 ;
  assign n54087 = n82810 & n54086 ;
  assign n82811 = ~n53732 ;
  assign n54088 = x90 & n82811 ;
  assign n82812 = ~n53730 ;
  assign n54089 = n82812 & n54088 ;
  assign n54090 = n53734 | n54089 ;
  assign n54091 = n54087 | n54090 ;
  assign n82813 = ~n53734 ;
  assign n54092 = n82813 & n54091 ;
  assign n82814 = ~n53723 ;
  assign n54093 = x91 & n82814 ;
  assign n82815 = ~n53721 ;
  assign n54094 = n82815 & n54093 ;
  assign n54095 = n53725 | n54094 ;
  assign n54097 = n54092 | n54095 ;
  assign n82816 = ~n53725 ;
  assign n54098 = n82816 & n54097 ;
  assign n82817 = ~n53714 ;
  assign n54099 = x92 & n82817 ;
  assign n82818 = ~n53712 ;
  assign n54100 = n82818 & n54099 ;
  assign n54101 = n53716 | n54100 ;
  assign n54102 = n54098 | n54101 ;
  assign n82819 = ~n53716 ;
  assign n54103 = n82819 & n54102 ;
  assign n82820 = ~n53705 ;
  assign n54104 = x93 & n82820 ;
  assign n82821 = ~n53703 ;
  assign n54105 = n82821 & n54104 ;
  assign n54106 = n53707 | n54105 ;
  assign n54108 = n54103 | n54106 ;
  assign n82822 = ~n53707 ;
  assign n54109 = n82822 & n54108 ;
  assign n82823 = ~n53696 ;
  assign n54110 = x94 & n82823 ;
  assign n82824 = ~n53694 ;
  assign n54111 = n82824 & n54110 ;
  assign n54112 = n53698 | n54111 ;
  assign n54113 = n54109 | n54112 ;
  assign n82825 = ~n53698 ;
  assign n54114 = n82825 & n54113 ;
  assign n82826 = ~n53687 ;
  assign n54115 = x95 & n82826 ;
  assign n82827 = ~n53685 ;
  assign n54116 = n82827 & n54115 ;
  assign n54117 = n53689 | n54116 ;
  assign n54119 = n54114 | n54117 ;
  assign n82828 = ~n53689 ;
  assign n54120 = n82828 & n54119 ;
  assign n82829 = ~n53678 ;
  assign n54121 = x96 & n82829 ;
  assign n82830 = ~n53676 ;
  assign n54122 = n82830 & n54121 ;
  assign n54123 = n53680 | n54122 ;
  assign n54124 = n54120 | n54123 ;
  assign n82831 = ~n53680 ;
  assign n54125 = n82831 & n54124 ;
  assign n82832 = ~n53669 ;
  assign n54126 = x97 & n82832 ;
  assign n82833 = ~n53667 ;
  assign n54127 = n82833 & n54126 ;
  assign n54128 = n53671 | n54127 ;
  assign n54130 = n54125 | n54128 ;
  assign n82834 = ~n53671 ;
  assign n54131 = n82834 & n54130 ;
  assign n82835 = ~n53660 ;
  assign n54132 = x98 & n82835 ;
  assign n82836 = ~n53658 ;
  assign n54133 = n82836 & n54132 ;
  assign n54134 = n53662 | n54133 ;
  assign n54135 = n54131 | n54134 ;
  assign n82837 = ~n53662 ;
  assign n54136 = n82837 & n54135 ;
  assign n82838 = ~n53651 ;
  assign n54137 = x99 & n82838 ;
  assign n82839 = ~n53649 ;
  assign n54138 = n82839 & n54137 ;
  assign n54139 = n53653 | n54138 ;
  assign n54141 = n54136 | n54139 ;
  assign n82840 = ~n53653 ;
  assign n54142 = n82840 & n54141 ;
  assign n82841 = ~n53642 ;
  assign n54143 = x100 & n82841 ;
  assign n82842 = ~n53640 ;
  assign n54144 = n82842 & n54143 ;
  assign n54145 = n53644 | n54144 ;
  assign n54146 = n54142 | n54145 ;
  assign n82843 = ~n53644 ;
  assign n54147 = n82843 & n54146 ;
  assign n82844 = ~n53633 ;
  assign n54148 = x101 & n82844 ;
  assign n82845 = ~n53631 ;
  assign n54149 = n82845 & n54148 ;
  assign n54150 = n53635 | n54149 ;
  assign n54152 = n54147 | n54150 ;
  assign n82846 = ~n53635 ;
  assign n54153 = n82846 & n54152 ;
  assign n82847 = ~n53624 ;
  assign n54154 = x102 & n82847 ;
  assign n82848 = ~n53622 ;
  assign n54155 = n82848 & n54154 ;
  assign n54156 = n53626 | n54155 ;
  assign n54157 = n54153 | n54156 ;
  assign n82849 = ~n53626 ;
  assign n54158 = n82849 & n54157 ;
  assign n82850 = ~n53615 ;
  assign n54159 = x103 & n82850 ;
  assign n82851 = ~n53613 ;
  assign n54160 = n82851 & n54159 ;
  assign n54161 = n53617 | n54160 ;
  assign n54163 = n54158 | n54161 ;
  assign n82852 = ~n53617 ;
  assign n54164 = n82852 & n54163 ;
  assign n82853 = ~n53606 ;
  assign n54165 = x104 & n82853 ;
  assign n82854 = ~n53604 ;
  assign n54166 = n82854 & n54165 ;
  assign n54167 = n53608 | n54166 ;
  assign n54168 = n54164 | n54167 ;
  assign n82855 = ~n53608 ;
  assign n54169 = n82855 & n54168 ;
  assign n82856 = ~n53597 ;
  assign n54170 = x105 & n82856 ;
  assign n82857 = ~n53595 ;
  assign n54171 = n82857 & n54170 ;
  assign n54172 = n53599 | n54171 ;
  assign n54174 = n54169 | n54172 ;
  assign n82858 = ~n53599 ;
  assign n54175 = n82858 & n54174 ;
  assign n82859 = ~n53588 ;
  assign n54176 = x106 & n82859 ;
  assign n82860 = ~n53586 ;
  assign n54177 = n82860 & n54176 ;
  assign n54178 = n53590 | n54177 ;
  assign n54179 = n54175 | n54178 ;
  assign n82861 = ~n53590 ;
  assign n54180 = n82861 & n54179 ;
  assign n82862 = ~n53579 ;
  assign n54181 = x107 & n82862 ;
  assign n82863 = ~n53577 ;
  assign n54182 = n82863 & n54181 ;
  assign n54183 = n53581 | n54182 ;
  assign n54185 = n54180 | n54183 ;
  assign n82864 = ~n53581 ;
  assign n54186 = n82864 & n54185 ;
  assign n82865 = ~n53570 ;
  assign n54187 = x108 & n82865 ;
  assign n82866 = ~n53568 ;
  assign n54188 = n82866 & n54187 ;
  assign n54189 = n53572 | n54188 ;
  assign n54190 = n54186 | n54189 ;
  assign n82867 = ~n53572 ;
  assign n54191 = n82867 & n54190 ;
  assign n82868 = ~n53561 ;
  assign n54192 = x109 & n82868 ;
  assign n82869 = ~n53559 ;
  assign n54193 = n82869 & n54192 ;
  assign n54194 = n53563 | n54193 ;
  assign n54196 = n54191 | n54194 ;
  assign n82870 = ~n53563 ;
  assign n54197 = n82870 & n54196 ;
  assign n82871 = ~n53552 ;
  assign n54198 = x110 & n82871 ;
  assign n82872 = ~n53550 ;
  assign n54199 = n82872 & n54198 ;
  assign n54200 = n53554 | n54199 ;
  assign n54201 = n54197 | n54200 ;
  assign n82873 = ~n53554 ;
  assign n54202 = n82873 & n54201 ;
  assign n82874 = ~n53543 ;
  assign n54203 = x111 & n82874 ;
  assign n82875 = ~n53541 ;
  assign n54204 = n82875 & n54203 ;
  assign n54205 = n53545 | n54204 ;
  assign n54207 = n54202 | n54205 ;
  assign n82876 = ~n53545 ;
  assign n54208 = n82876 & n54207 ;
  assign n82877 = ~n53534 ;
  assign n54209 = x112 & n82877 ;
  assign n82878 = ~n53532 ;
  assign n54210 = n82878 & n54209 ;
  assign n54211 = n53536 | n54210 ;
  assign n54212 = n54208 | n54211 ;
  assign n82879 = ~n53536 ;
  assign n54213 = n82879 & n54212 ;
  assign n82880 = ~n53525 ;
  assign n54214 = x113 & n82880 ;
  assign n82881 = ~n53523 ;
  assign n54215 = n82881 & n54214 ;
  assign n54216 = n53527 | n54215 ;
  assign n54218 = n54213 | n54216 ;
  assign n82882 = ~n53527 ;
  assign n54219 = n82882 & n54218 ;
  assign n82883 = ~n53503 ;
  assign n54220 = x114 & n82883 ;
  assign n82884 = ~n53501 ;
  assign n54221 = n82884 & n54220 ;
  assign n54222 = n53518 | n54221 ;
  assign n54223 = n54219 | n54222 ;
  assign n82885 = ~n53518 ;
  assign n54224 = n82885 & n54223 ;
  assign n82886 = ~n53515 ;
  assign n54225 = x115 & n82886 ;
  assign n82887 = ~n53513 ;
  assign n54226 = n82887 & n54225 ;
  assign n54227 = n53517 | n54226 ;
  assign n54229 = n54224 | n54227 ;
  assign n82888 = ~n53517 ;
  assign n54230 = n82888 & n54229 ;
  assign n54231 = n65429 | n54230 ;
  assign n54232 = n53504 & n54231 ;
  assign n54233 = n53735 | n53949 ;
  assign n54234 = x65 & n54233 ;
  assign n82889 = ~n54234 ;
  assign n54235 = n53955 & n82889 ;
  assign n54236 = n21731 | n54235 ;
  assign n54237 = n82738 & n54236 ;
  assign n54238 = n53962 | n54237 ;
  assign n54239 = n82741 & n54238 ;
  assign n54240 = n53937 | n53966 ;
  assign n54242 = n54239 | n54240 ;
  assign n54243 = n82744 & n54242 ;
  assign n54245 = n53971 | n54243 ;
  assign n54246 = n82747 & n54245 ;
  assign n54247 = n53920 | n53975 ;
  assign n54249 = n54246 | n54247 ;
  assign n54250 = n82750 & n54249 ;
  assign n54251 = n53979 | n54250 ;
  assign n54253 = n82753 & n54251 ;
  assign n54254 = n53985 | n54253 ;
  assign n54255 = n82756 & n54254 ;
  assign n54256 = n53991 | n54255 ;
  assign n54258 = n82759 & n54256 ;
  assign n54259 = n53996 | n54258 ;
  assign n54260 = n82762 & n54259 ;
  assign n54261 = n54002 | n54260 ;
  assign n54263 = n82765 & n54261 ;
  assign n54264 = n54007 | n54263 ;
  assign n54265 = n82768 & n54264 ;
  assign n54266 = n54013 | n54265 ;
  assign n54268 = n82771 & n54266 ;
  assign n54269 = n54018 | n54268 ;
  assign n54270 = n82774 & n54269 ;
  assign n54271 = n54024 | n54270 ;
  assign n54273 = n82777 & n54271 ;
  assign n54274 = n54029 | n54273 ;
  assign n54275 = n82780 & n54274 ;
  assign n54276 = n54035 | n54275 ;
  assign n54278 = n82783 & n54276 ;
  assign n54279 = n54040 | n54278 ;
  assign n54280 = n82786 & n54279 ;
  assign n54281 = n54046 | n54280 ;
  assign n54283 = n82789 & n54281 ;
  assign n54284 = n54051 | n54283 ;
  assign n54285 = n82792 & n54284 ;
  assign n54286 = n54057 | n54285 ;
  assign n54288 = n82795 & n54286 ;
  assign n54289 = n54062 | n54288 ;
  assign n54290 = n82798 & n54289 ;
  assign n54291 = n54068 | n54290 ;
  assign n54293 = n82801 & n54291 ;
  assign n54294 = n54073 | n54293 ;
  assign n54295 = n82804 & n54294 ;
  assign n54296 = n54079 | n54295 ;
  assign n54298 = n82807 & n54296 ;
  assign n54299 = n54084 | n54298 ;
  assign n54300 = n82810 & n54299 ;
  assign n54301 = n54090 | n54300 ;
  assign n54303 = n82813 & n54301 ;
  assign n54304 = n54095 | n54303 ;
  assign n54305 = n82816 & n54304 ;
  assign n54306 = n54101 | n54305 ;
  assign n54308 = n82819 & n54306 ;
  assign n54309 = n54106 | n54308 ;
  assign n54310 = n82822 & n54309 ;
  assign n54311 = n54112 | n54310 ;
  assign n54313 = n82825 & n54311 ;
  assign n54314 = n54117 | n54313 ;
  assign n54315 = n82828 & n54314 ;
  assign n54316 = n54123 | n54315 ;
  assign n54318 = n82831 & n54316 ;
  assign n54319 = n54128 | n54318 ;
  assign n54320 = n82834 & n54319 ;
  assign n54321 = n54134 | n54320 ;
  assign n54323 = n82837 & n54321 ;
  assign n54324 = n54139 | n54323 ;
  assign n54325 = n82840 & n54324 ;
  assign n54326 = n54145 | n54325 ;
  assign n54328 = n82843 & n54326 ;
  assign n54329 = n54150 | n54328 ;
  assign n54330 = n82846 & n54329 ;
  assign n54331 = n54156 | n54330 ;
  assign n54333 = n82849 & n54331 ;
  assign n54334 = n54161 | n54333 ;
  assign n54335 = n82852 & n54334 ;
  assign n54336 = n54167 | n54335 ;
  assign n54338 = n82855 & n54336 ;
  assign n54339 = n54172 | n54338 ;
  assign n54340 = n82858 & n54339 ;
  assign n54341 = n54178 | n54340 ;
  assign n54343 = n82861 & n54341 ;
  assign n54344 = n54183 | n54343 ;
  assign n54345 = n82864 & n54344 ;
  assign n54346 = n54189 | n54345 ;
  assign n54348 = n82867 & n54346 ;
  assign n54349 = n54194 | n54348 ;
  assign n54350 = n82870 & n54349 ;
  assign n54351 = n54200 | n54350 ;
  assign n54353 = n82873 & n54351 ;
  assign n54354 = n54205 | n54353 ;
  assign n54355 = n82876 & n54354 ;
  assign n54356 = n54211 | n54355 ;
  assign n54358 = n82879 & n54356 ;
  assign n54359 = n54216 | n54358 ;
  assign n54360 = n82882 & n54359 ;
  assign n82890 = ~n54360 ;
  assign n54361 = n54222 & n82890 ;
  assign n54363 = n53527 | n54222 ;
  assign n82891 = ~n54363 ;
  assign n54364 = n54218 & n82891 ;
  assign n54365 = n54361 | n54364 ;
  assign n54366 = n67021 & n54365 ;
  assign n82892 = ~n54230 ;
  assign n54367 = n82892 & n54366 ;
  assign n54368 = n54232 | n54367 ;
  assign n54369 = n72393 & n54368 ;
  assign n82893 = ~n54367 ;
  assign n55039 = x115 & n82893 ;
  assign n82894 = ~n54232 ;
  assign n55040 = n82894 & n55039 ;
  assign n55041 = n54369 | n55040 ;
  assign n54370 = n53526 & n54231 ;
  assign n82895 = ~n54213 ;
  assign n54217 = n82895 & n54216 ;
  assign n54371 = n53536 | n54216 ;
  assign n82896 = ~n54371 ;
  assign n54372 = n54356 & n82896 ;
  assign n54373 = n54217 | n54372 ;
  assign n54374 = n67021 & n54373 ;
  assign n54375 = n82892 & n54374 ;
  assign n54376 = n54370 | n54375 ;
  assign n54377 = n72385 & n54376 ;
  assign n54378 = n53535 & n54231 ;
  assign n82897 = ~n54355 ;
  assign n54357 = n54211 & n82897 ;
  assign n54379 = n53545 | n54211 ;
  assign n82898 = ~n54379 ;
  assign n54380 = n54207 & n82898 ;
  assign n54381 = n54357 | n54380 ;
  assign n54382 = n67021 & n54381 ;
  assign n54383 = n82892 & n54382 ;
  assign n54384 = n54378 | n54383 ;
  assign n54385 = n72025 & n54384 ;
  assign n82899 = ~n54383 ;
  assign n55029 = x113 & n82899 ;
  assign n82900 = ~n54378 ;
  assign n55030 = n82900 & n55029 ;
  assign n55031 = n54385 | n55030 ;
  assign n54386 = n53544 & n54231 ;
  assign n82901 = ~n54202 ;
  assign n54206 = n82901 & n54205 ;
  assign n54387 = n53554 | n54205 ;
  assign n82902 = ~n54387 ;
  assign n54388 = n54351 & n82902 ;
  assign n54389 = n54206 | n54388 ;
  assign n54390 = n67021 & n54389 ;
  assign n54391 = n82892 & n54390 ;
  assign n54392 = n54386 | n54391 ;
  assign n54393 = n71645 & n54392 ;
  assign n54394 = n53553 & n54231 ;
  assign n82903 = ~n54350 ;
  assign n54352 = n54200 & n82903 ;
  assign n54395 = n53563 | n54200 ;
  assign n82904 = ~n54395 ;
  assign n54396 = n54196 & n82904 ;
  assign n54397 = n54352 | n54396 ;
  assign n54398 = n67021 & n54397 ;
  assign n54399 = n82892 & n54398 ;
  assign n54400 = n54394 | n54399 ;
  assign n54401 = n71633 & n54400 ;
  assign n82905 = ~n54399 ;
  assign n55019 = x111 & n82905 ;
  assign n82906 = ~n54394 ;
  assign n55020 = n82906 & n55019 ;
  assign n55021 = n54401 | n55020 ;
  assign n54402 = n53562 & n54231 ;
  assign n82907 = ~n54191 ;
  assign n54195 = n82907 & n54194 ;
  assign n54403 = n53572 | n54194 ;
  assign n82908 = ~n54403 ;
  assign n54404 = n54346 & n82908 ;
  assign n54405 = n54195 | n54404 ;
  assign n54406 = n67021 & n54405 ;
  assign n54407 = n82892 & n54406 ;
  assign n54408 = n54402 | n54407 ;
  assign n54409 = n71253 & n54408 ;
  assign n54410 = n53571 & n54231 ;
  assign n82909 = ~n54345 ;
  assign n54347 = n54189 & n82909 ;
  assign n54411 = n53581 | n54189 ;
  assign n82910 = ~n54411 ;
  assign n54412 = n54185 & n82910 ;
  assign n54413 = n54347 | n54412 ;
  assign n54414 = n67021 & n54413 ;
  assign n54415 = n82892 & n54414 ;
  assign n54416 = n54410 | n54415 ;
  assign n54417 = n70935 & n54416 ;
  assign n82911 = ~n54415 ;
  assign n55009 = x109 & n82911 ;
  assign n82912 = ~n54410 ;
  assign n55010 = n82912 & n55009 ;
  assign n55011 = n54417 | n55010 ;
  assign n54418 = n53580 & n54231 ;
  assign n82913 = ~n54180 ;
  assign n54184 = n82913 & n54183 ;
  assign n54419 = n53590 | n54183 ;
  assign n82914 = ~n54419 ;
  assign n54420 = n54341 & n82914 ;
  assign n54421 = n54184 | n54420 ;
  assign n54422 = n67021 & n54421 ;
  assign n54423 = n82892 & n54422 ;
  assign n54424 = n54418 | n54423 ;
  assign n54425 = n70927 & n54424 ;
  assign n54426 = n53589 & n54231 ;
  assign n82915 = ~n54340 ;
  assign n54342 = n54178 & n82915 ;
  assign n54427 = n53599 | n54178 ;
  assign n82916 = ~n54427 ;
  assign n54428 = n54174 & n82916 ;
  assign n54429 = n54342 | n54428 ;
  assign n54430 = n67021 & n54429 ;
  assign n54431 = n82892 & n54430 ;
  assign n54432 = n54426 | n54431 ;
  assign n54433 = n70609 & n54432 ;
  assign n82917 = ~n54431 ;
  assign n54998 = x107 & n82917 ;
  assign n82918 = ~n54426 ;
  assign n54999 = n82918 & n54998 ;
  assign n55000 = n54433 | n54999 ;
  assign n54434 = n53598 & n54231 ;
  assign n82919 = ~n54169 ;
  assign n54173 = n82919 & n54172 ;
  assign n54435 = n53608 | n54172 ;
  assign n82920 = ~n54435 ;
  assign n54436 = n54336 & n82920 ;
  assign n54437 = n54173 | n54436 ;
  assign n54438 = n67021 & n54437 ;
  assign n54439 = n82892 & n54438 ;
  assign n54440 = n54434 | n54439 ;
  assign n54441 = n70276 & n54440 ;
  assign n54442 = n53607 & n54231 ;
  assign n82921 = ~n54335 ;
  assign n54337 = n54167 & n82921 ;
  assign n54443 = n53617 | n54167 ;
  assign n82922 = ~n54443 ;
  assign n54444 = n54163 & n82922 ;
  assign n54445 = n54337 | n54444 ;
  assign n54446 = n67021 & n54445 ;
  assign n54447 = n82892 & n54446 ;
  assign n54448 = n54442 | n54447 ;
  assign n54449 = n70176 & n54448 ;
  assign n82923 = ~n54447 ;
  assign n54988 = x105 & n82923 ;
  assign n82924 = ~n54442 ;
  assign n54989 = n82924 & n54988 ;
  assign n54990 = n54449 | n54989 ;
  assign n54450 = n53616 & n54231 ;
  assign n82925 = ~n54158 ;
  assign n54162 = n82925 & n54161 ;
  assign n54451 = n53626 | n54161 ;
  assign n82926 = ~n54451 ;
  assign n54452 = n54331 & n82926 ;
  assign n54453 = n54162 | n54452 ;
  assign n54454 = n67021 & n54453 ;
  assign n54455 = n82892 & n54454 ;
  assign n54456 = n54450 | n54455 ;
  assign n54457 = n69857 & n54456 ;
  assign n54458 = n53625 & n54231 ;
  assign n82927 = ~n54330 ;
  assign n54332 = n54156 & n82927 ;
  assign n54459 = n53635 | n54156 ;
  assign n82928 = ~n54459 ;
  assign n54460 = n54152 & n82928 ;
  assign n54461 = n54332 | n54460 ;
  assign n54462 = n67021 & n54461 ;
  assign n54463 = n82892 & n54462 ;
  assign n54464 = n54458 | n54463 ;
  assign n54465 = n69656 & n54464 ;
  assign n82929 = ~n54463 ;
  assign n54977 = x103 & n82929 ;
  assign n82930 = ~n54458 ;
  assign n54978 = n82930 & n54977 ;
  assign n54979 = n54465 | n54978 ;
  assign n54466 = n53634 & n54231 ;
  assign n82931 = ~n54147 ;
  assign n54151 = n82931 & n54150 ;
  assign n54467 = n53644 | n54150 ;
  assign n82932 = ~n54467 ;
  assign n54468 = n54326 & n82932 ;
  assign n54469 = n54151 | n54468 ;
  assign n54470 = n67021 & n54469 ;
  assign n54471 = n82892 & n54470 ;
  assign n54472 = n54466 | n54471 ;
  assign n54473 = n69528 & n54472 ;
  assign n54474 = n53643 & n54231 ;
  assign n82933 = ~n54325 ;
  assign n54327 = n54145 & n82933 ;
  assign n54475 = n53653 | n54145 ;
  assign n82934 = ~n54475 ;
  assign n54476 = n54141 & n82934 ;
  assign n54477 = n54327 | n54476 ;
  assign n54478 = n67021 & n54477 ;
  assign n54479 = n82892 & n54478 ;
  assign n54480 = n54474 | n54479 ;
  assign n54481 = n69261 & n54480 ;
  assign n82935 = ~n54479 ;
  assign n54966 = x101 & n82935 ;
  assign n82936 = ~n54474 ;
  assign n54967 = n82936 & n54966 ;
  assign n54968 = n54481 | n54967 ;
  assign n54482 = n53652 & n54231 ;
  assign n82937 = ~n54136 ;
  assign n54140 = n82937 & n54139 ;
  assign n54483 = n53662 | n54139 ;
  assign n82938 = ~n54483 ;
  assign n54484 = n54321 & n82938 ;
  assign n54485 = n54140 | n54484 ;
  assign n54486 = n67021 & n54485 ;
  assign n54487 = n82892 & n54486 ;
  assign n54488 = n54482 | n54487 ;
  assign n54489 = n69075 & n54488 ;
  assign n54490 = n53661 & n54231 ;
  assign n82939 = ~n54320 ;
  assign n54322 = n54134 & n82939 ;
  assign n54491 = n53671 | n54134 ;
  assign n82940 = ~n54491 ;
  assign n54492 = n54130 & n82940 ;
  assign n54493 = n54322 | n54492 ;
  assign n54494 = n67021 & n54493 ;
  assign n54495 = n82892 & n54494 ;
  assign n54496 = n54490 | n54495 ;
  assign n54497 = n68993 & n54496 ;
  assign n82941 = ~n54495 ;
  assign n54956 = x99 & n82941 ;
  assign n82942 = ~n54490 ;
  assign n54957 = n82942 & n54956 ;
  assign n54958 = n54497 | n54957 ;
  assign n54498 = n53670 & n54231 ;
  assign n82943 = ~n54125 ;
  assign n54129 = n82943 & n54128 ;
  assign n54499 = n53680 | n54128 ;
  assign n82944 = ~n54499 ;
  assign n54500 = n54316 & n82944 ;
  assign n54501 = n54129 | n54500 ;
  assign n54502 = n67021 & n54501 ;
  assign n54503 = n82892 & n54502 ;
  assign n54504 = n54498 | n54503 ;
  assign n54505 = n68716 & n54504 ;
  assign n54506 = n53679 & n54231 ;
  assign n82945 = ~n54315 ;
  assign n54317 = n54123 & n82945 ;
  assign n54507 = n53689 | n54123 ;
  assign n82946 = ~n54507 ;
  assign n54508 = n54119 & n82946 ;
  assign n54509 = n54317 | n54508 ;
  assign n54510 = n67021 & n54509 ;
  assign n54511 = n82892 & n54510 ;
  assign n54512 = n54506 | n54511 ;
  assign n54513 = n68545 & n54512 ;
  assign n82947 = ~n54511 ;
  assign n54946 = x97 & n82947 ;
  assign n82948 = ~n54506 ;
  assign n54947 = n82948 & n54946 ;
  assign n54948 = n54513 | n54947 ;
  assign n54514 = n53688 & n54231 ;
  assign n82949 = ~n54114 ;
  assign n54118 = n82949 & n54117 ;
  assign n54515 = n53698 | n54117 ;
  assign n82950 = ~n54515 ;
  assign n54516 = n54311 & n82950 ;
  assign n54517 = n54118 | n54516 ;
  assign n54518 = n67021 & n54517 ;
  assign n54519 = n82892 & n54518 ;
  assign n54520 = n54514 | n54519 ;
  assign n54521 = n68438 & n54520 ;
  assign n54522 = n53697 & n54231 ;
  assign n82951 = ~n54310 ;
  assign n54312 = n54112 & n82951 ;
  assign n54523 = n53707 | n54112 ;
  assign n82952 = ~n54523 ;
  assign n54524 = n54108 & n82952 ;
  assign n54525 = n54312 | n54524 ;
  assign n54526 = n67021 & n54525 ;
  assign n54527 = n82892 & n54526 ;
  assign n54528 = n54522 | n54527 ;
  assign n54529 = n68214 & n54528 ;
  assign n82953 = ~n54527 ;
  assign n54936 = x95 & n82953 ;
  assign n82954 = ~n54522 ;
  assign n54937 = n82954 & n54936 ;
  assign n54938 = n54529 | n54937 ;
  assign n54530 = n53706 & n54231 ;
  assign n82955 = ~n54103 ;
  assign n54107 = n82955 & n54106 ;
  assign n54531 = n53716 | n54106 ;
  assign n82956 = ~n54531 ;
  assign n54532 = n54306 & n82956 ;
  assign n54533 = n54107 | n54532 ;
  assign n54534 = n67021 & n54533 ;
  assign n54535 = n82892 & n54534 ;
  assign n54536 = n54530 | n54535 ;
  assign n54537 = n68058 & n54536 ;
  assign n54538 = n53715 & n54231 ;
  assign n82957 = ~n54305 ;
  assign n54307 = n54101 & n82957 ;
  assign n54539 = n53725 | n54101 ;
  assign n82958 = ~n54539 ;
  assign n54540 = n54097 & n82958 ;
  assign n54541 = n54307 | n54540 ;
  assign n54542 = n67021 & n54541 ;
  assign n54543 = n82892 & n54542 ;
  assign n54544 = n54538 | n54543 ;
  assign n54545 = n67986 & n54544 ;
  assign n82959 = ~n54543 ;
  assign n54925 = x93 & n82959 ;
  assign n82960 = ~n54538 ;
  assign n54926 = n82960 & n54925 ;
  assign n54927 = n54545 | n54926 ;
  assign n54546 = n53724 & n54231 ;
  assign n82961 = ~n54092 ;
  assign n54096 = n82961 & n54095 ;
  assign n54547 = n53734 | n54095 ;
  assign n82962 = ~n54547 ;
  assign n54548 = n54301 & n82962 ;
  assign n54549 = n54096 | n54548 ;
  assign n54550 = n67021 & n54549 ;
  assign n54551 = n82892 & n54550 ;
  assign n54552 = n54546 | n54551 ;
  assign n54553 = n67763 & n54552 ;
  assign n54554 = n53733 & n54231 ;
  assign n82963 = ~n54300 ;
  assign n54302 = n54090 & n82963 ;
  assign n54555 = n53743 | n54090 ;
  assign n82964 = ~n54555 ;
  assign n54556 = n54086 & n82964 ;
  assign n54557 = n54302 | n54556 ;
  assign n54558 = n67021 & n54557 ;
  assign n54559 = n82892 & n54558 ;
  assign n54560 = n54554 | n54559 ;
  assign n54561 = n67622 & n54560 ;
  assign n82965 = ~n54559 ;
  assign n54915 = x91 & n82965 ;
  assign n82966 = ~n54554 ;
  assign n54916 = n82966 & n54915 ;
  assign n54917 = n54561 | n54916 ;
  assign n54562 = n53742 & n54231 ;
  assign n82967 = ~n54081 ;
  assign n54085 = n82967 & n54084 ;
  assign n54563 = n53752 | n54084 ;
  assign n82968 = ~n54563 ;
  assign n54564 = n54296 & n82968 ;
  assign n54565 = n54085 | n54564 ;
  assign n54566 = n67021 & n54565 ;
  assign n54567 = n82892 & n54566 ;
  assign n54568 = n54562 | n54567 ;
  assign n54569 = n67531 & n54568 ;
  assign n54570 = n53751 & n54231 ;
  assign n82969 = ~n54295 ;
  assign n54297 = n54079 & n82969 ;
  assign n54571 = n53761 | n54079 ;
  assign n82970 = ~n54571 ;
  assign n54572 = n54075 & n82970 ;
  assign n54573 = n54297 | n54572 ;
  assign n54574 = n67021 & n54573 ;
  assign n54575 = n82892 & n54574 ;
  assign n54576 = n54570 | n54575 ;
  assign n54577 = n67348 & n54576 ;
  assign n82971 = ~n54575 ;
  assign n54905 = x89 & n82971 ;
  assign n82972 = ~n54570 ;
  assign n54906 = n82972 & n54905 ;
  assign n54907 = n54577 | n54906 ;
  assign n54578 = n53760 & n54231 ;
  assign n82973 = ~n54070 ;
  assign n54074 = n82973 & n54073 ;
  assign n54579 = n53770 | n54073 ;
  assign n82974 = ~n54579 ;
  assign n54580 = n54291 & n82974 ;
  assign n54581 = n54074 | n54580 ;
  assign n54582 = n67021 & n54581 ;
  assign n54583 = n82892 & n54582 ;
  assign n54584 = n54578 | n54583 ;
  assign n54585 = n67222 & n54584 ;
  assign n54586 = n53769 & n54231 ;
  assign n82975 = ~n54290 ;
  assign n54292 = n54068 & n82975 ;
  assign n54587 = n53779 | n54068 ;
  assign n82976 = ~n54587 ;
  assign n54588 = n54064 & n82976 ;
  assign n54589 = n54292 | n54588 ;
  assign n54590 = n67021 & n54589 ;
  assign n54591 = n82892 & n54590 ;
  assign n54592 = n54586 | n54591 ;
  assign n54593 = n67164 & n54592 ;
  assign n82977 = ~n54591 ;
  assign n54895 = x87 & n82977 ;
  assign n82978 = ~n54586 ;
  assign n54896 = n82978 & n54895 ;
  assign n54897 = n54593 | n54896 ;
  assign n54594 = n53778 & n54231 ;
  assign n82979 = ~n54059 ;
  assign n54063 = n82979 & n54062 ;
  assign n54595 = n53787 | n54062 ;
  assign n82980 = ~n54595 ;
  assign n54596 = n54286 & n82980 ;
  assign n54597 = n54063 | n54596 ;
  assign n54598 = n67021 & n54597 ;
  assign n54599 = n82892 & n54598 ;
  assign n54600 = n54594 | n54599 ;
  assign n54601 = n66979 & n54600 ;
  assign n54602 = n53786 & n54231 ;
  assign n82981 = ~n54285 ;
  assign n54287 = n54057 & n82981 ;
  assign n54603 = n53796 | n54057 ;
  assign n82982 = ~n54603 ;
  assign n54604 = n54053 & n82982 ;
  assign n54605 = n54287 | n54604 ;
  assign n54606 = n67021 & n54605 ;
  assign n54607 = n82892 & n54606 ;
  assign n54608 = n54602 | n54607 ;
  assign n54609 = n66868 & n54608 ;
  assign n82983 = ~n54607 ;
  assign n54885 = x85 & n82983 ;
  assign n82984 = ~n54602 ;
  assign n54886 = n82984 & n54885 ;
  assign n54887 = n54609 | n54886 ;
  assign n54610 = n53795 & n54231 ;
  assign n82985 = ~n54048 ;
  assign n54052 = n82985 & n54051 ;
  assign n54611 = n53805 | n54051 ;
  assign n82986 = ~n54611 ;
  assign n54612 = n54281 & n82986 ;
  assign n54613 = n54052 | n54612 ;
  assign n54614 = n67021 & n54613 ;
  assign n54615 = n82892 & n54614 ;
  assign n54616 = n54610 | n54615 ;
  assign n54617 = n66797 & n54616 ;
  assign n54618 = n53804 & n54231 ;
  assign n82987 = ~n54280 ;
  assign n54282 = n54046 & n82987 ;
  assign n54619 = n53814 | n54046 ;
  assign n82988 = ~n54619 ;
  assign n54620 = n54042 & n82988 ;
  assign n54621 = n54282 | n54620 ;
  assign n54622 = n67021 & n54621 ;
  assign n54623 = n82892 & n54622 ;
  assign n54624 = n54618 | n54623 ;
  assign n54625 = n66654 & n54624 ;
  assign n82989 = ~n54623 ;
  assign n54874 = x83 & n82989 ;
  assign n82990 = ~n54618 ;
  assign n54875 = n82990 & n54874 ;
  assign n54876 = n54625 | n54875 ;
  assign n54626 = n53813 & n54231 ;
  assign n82991 = ~n54037 ;
  assign n54041 = n82991 & n54040 ;
  assign n54627 = n53823 | n54040 ;
  assign n82992 = ~n54627 ;
  assign n54628 = n54276 & n82992 ;
  assign n54629 = n54041 | n54628 ;
  assign n54630 = n67021 & n54629 ;
  assign n54631 = n82892 & n54630 ;
  assign n54632 = n54626 | n54631 ;
  assign n54633 = n66560 & n54632 ;
  assign n54634 = n53822 & n54231 ;
  assign n82993 = ~n54275 ;
  assign n54277 = n54035 & n82993 ;
  assign n54635 = n53832 | n54035 ;
  assign n82994 = ~n54635 ;
  assign n54636 = n54031 & n82994 ;
  assign n54637 = n54277 | n54636 ;
  assign n54638 = n67021 & n54637 ;
  assign n54639 = n82892 & n54638 ;
  assign n54640 = n54634 | n54639 ;
  assign n54641 = n66505 & n54640 ;
  assign n82995 = ~n54639 ;
  assign n54862 = x81 & n82995 ;
  assign n82996 = ~n54634 ;
  assign n54863 = n82996 & n54862 ;
  assign n54864 = n54641 | n54863 ;
  assign n54642 = n53831 & n54231 ;
  assign n82997 = ~n54026 ;
  assign n54030 = n82997 & n54029 ;
  assign n54643 = n53840 | n54029 ;
  assign n82998 = ~n54643 ;
  assign n54644 = n54271 & n82998 ;
  assign n54645 = n54030 | n54644 ;
  assign n54646 = n67021 & n54645 ;
  assign n54647 = n82892 & n54646 ;
  assign n54648 = n54642 | n54647 ;
  assign n54649 = n66379 & n54648 ;
  assign n54650 = n53839 & n54231 ;
  assign n82999 = ~n54270 ;
  assign n54272 = n54024 & n82999 ;
  assign n54651 = n53849 | n54024 ;
  assign n83000 = ~n54651 ;
  assign n54652 = n54020 & n83000 ;
  assign n54653 = n54272 | n54652 ;
  assign n54654 = n67021 & n54653 ;
  assign n54655 = n82892 & n54654 ;
  assign n54656 = n54650 | n54655 ;
  assign n54657 = n66299 & n54656 ;
  assign n83001 = ~n54655 ;
  assign n54852 = x79 & n83001 ;
  assign n83002 = ~n54650 ;
  assign n54853 = n83002 & n54852 ;
  assign n54854 = n54657 | n54853 ;
  assign n54658 = n53848 & n54231 ;
  assign n83003 = ~n54015 ;
  assign n54019 = n83003 & n54018 ;
  assign n54659 = n53858 | n54018 ;
  assign n83004 = ~n54659 ;
  assign n54660 = n54266 & n83004 ;
  assign n54661 = n54019 | n54660 ;
  assign n54662 = n67021 & n54661 ;
  assign n54663 = n82892 & n54662 ;
  assign n54664 = n54658 | n54663 ;
  assign n54665 = n66244 & n54664 ;
  assign n54666 = n53857 & n54231 ;
  assign n83005 = ~n54265 ;
  assign n54267 = n54013 & n83005 ;
  assign n54667 = n53866 | n54013 ;
  assign n83006 = ~n54667 ;
  assign n54668 = n54009 & n83006 ;
  assign n54669 = n54267 | n54668 ;
  assign n54670 = n67021 & n54669 ;
  assign n54671 = n82892 & n54670 ;
  assign n54672 = n54666 | n54671 ;
  assign n54673 = n66145 & n54672 ;
  assign n83007 = ~n54671 ;
  assign n54840 = x77 & n83007 ;
  assign n83008 = ~n54666 ;
  assign n54841 = n83008 & n54840 ;
  assign n54842 = n54673 | n54841 ;
  assign n54674 = n53865 & n54231 ;
  assign n83009 = ~n54004 ;
  assign n54008 = n83009 & n54007 ;
  assign n54675 = n53875 | n54007 ;
  assign n83010 = ~n54675 ;
  assign n54676 = n54261 & n83010 ;
  assign n54677 = n54008 | n54676 ;
  assign n54678 = n67021 & n54677 ;
  assign n54679 = n82892 & n54678 ;
  assign n54680 = n54674 | n54679 ;
  assign n54681 = n66081 & n54680 ;
  assign n54682 = n53874 & n54231 ;
  assign n83011 = ~n54260 ;
  assign n54262 = n54002 & n83011 ;
  assign n54683 = n53884 | n54002 ;
  assign n83012 = ~n54683 ;
  assign n54684 = n53998 & n83012 ;
  assign n54685 = n54262 | n54684 ;
  assign n54686 = n67021 & n54685 ;
  assign n54687 = n82892 & n54686 ;
  assign n54688 = n54682 | n54687 ;
  assign n54689 = n66043 & n54688 ;
  assign n83013 = ~n54687 ;
  assign n54830 = x75 & n83013 ;
  assign n83014 = ~n54682 ;
  assign n54831 = n83014 & n54830 ;
  assign n54832 = n54689 | n54831 ;
  assign n54690 = n53883 & n54231 ;
  assign n83015 = ~n53993 ;
  assign n53997 = n83015 & n53996 ;
  assign n54691 = n53893 | n53996 ;
  assign n83016 = ~n54691 ;
  assign n54692 = n54256 & n83016 ;
  assign n54693 = n53997 | n54692 ;
  assign n54694 = n67021 & n54693 ;
  assign n54695 = n82892 & n54694 ;
  assign n54696 = n54690 | n54695 ;
  assign n54697 = n65960 & n54696 ;
  assign n54698 = n53892 & n54231 ;
  assign n83017 = ~n54255 ;
  assign n54257 = n53991 & n83017 ;
  assign n54699 = n53902 | n53991 ;
  assign n83018 = ~n54699 ;
  assign n54700 = n53987 & n83018 ;
  assign n54701 = n54257 | n54700 ;
  assign n54702 = n67021 & n54701 ;
  assign n54703 = n82892 & n54702 ;
  assign n54704 = n54698 | n54703 ;
  assign n54705 = n65909 & n54704 ;
  assign n83019 = ~n54703 ;
  assign n54818 = x73 & n83019 ;
  assign n83020 = ~n54698 ;
  assign n54819 = n83020 & n54818 ;
  assign n54820 = n54705 | n54819 ;
  assign n54706 = n53901 & n54231 ;
  assign n83021 = ~n53982 ;
  assign n53986 = n83021 & n53985 ;
  assign n54707 = n53980 | n54250 ;
  assign n54708 = n53911 | n53985 ;
  assign n83022 = ~n54708 ;
  assign n54709 = n54707 & n83022 ;
  assign n54710 = n53986 | n54709 ;
  assign n54711 = n67021 & n54710 ;
  assign n54712 = n82892 & n54711 ;
  assign n54713 = n54706 | n54712 ;
  assign n54714 = n65877 & n54713 ;
  assign n54715 = n53910 & n54231 ;
  assign n83023 = ~n54250 ;
  assign n54252 = n53980 & n83023 ;
  assign n54716 = n53973 | n54247 ;
  assign n54717 = n53920 | n53980 ;
  assign n83024 = ~n54717 ;
  assign n54718 = n54716 & n83024 ;
  assign n54719 = n54252 | n54718 ;
  assign n54720 = n67021 & n54719 ;
  assign n54721 = n82892 & n54720 ;
  assign n54722 = n54715 | n54721 ;
  assign n54723 = n65820 & n54722 ;
  assign n83025 = ~n54721 ;
  assign n54808 = x71 & n83025 ;
  assign n83026 = ~n54715 ;
  assign n54809 = n83026 & n54808 ;
  assign n54810 = n54723 | n54809 ;
  assign n54724 = n53919 & n54231 ;
  assign n83027 = ~n53973 ;
  assign n54248 = n83027 & n54247 ;
  assign n54725 = n53929 | n54247 ;
  assign n83028 = ~n54725 ;
  assign n54726 = n54245 & n83028 ;
  assign n54727 = n54248 | n54726 ;
  assign n54728 = n67021 & n54727 ;
  assign n54729 = n82892 & n54728 ;
  assign n54730 = n54724 | n54729 ;
  assign n54731 = n65791 & n54730 ;
  assign n54732 = n53928 & n54231 ;
  assign n83029 = ~n54243 ;
  assign n54244 = n53971 & n83029 ;
  assign n54733 = n53964 | n54240 ;
  assign n54734 = n53937 | n53971 ;
  assign n83030 = ~n54734 ;
  assign n54735 = n54733 & n83030 ;
  assign n54736 = n54244 | n54735 ;
  assign n54737 = n67021 & n54736 ;
  assign n54738 = n82892 & n54737 ;
  assign n54739 = n54732 | n54738 ;
  assign n54740 = n65772 & n54739 ;
  assign n83031 = ~n54738 ;
  assign n54797 = x69 & n83031 ;
  assign n83032 = ~n54732 ;
  assign n54798 = n83032 & n54797 ;
  assign n54799 = n54740 | n54798 ;
  assign n54741 = n53936 & n54231 ;
  assign n83033 = ~n53964 ;
  assign n54241 = n83033 & n54240 ;
  assign n54742 = n53945 | n54240 ;
  assign n83034 = ~n54742 ;
  assign n54743 = n53963 & n83034 ;
  assign n54744 = n54241 | n54743 ;
  assign n54745 = n67021 & n54744 ;
  assign n54746 = n82892 & n54745 ;
  assign n54747 = n54741 | n54746 ;
  assign n54748 = n65746 & n54747 ;
  assign n54749 = n53944 & n54231 ;
  assign n54750 = n53958 | n53962 ;
  assign n83035 = ~n54750 ;
  assign n54751 = n54236 & n83035 ;
  assign n83036 = ~n54237 ;
  assign n54752 = n53962 & n83036 ;
  assign n54753 = n54751 | n54752 ;
  assign n54754 = n67021 & n54753 ;
  assign n54755 = n82892 & n54754 ;
  assign n54756 = n54749 | n54755 ;
  assign n54757 = n65721 & n54756 ;
  assign n83037 = ~n54755 ;
  assign n54787 = x67 & n83037 ;
  assign n83038 = ~n54749 ;
  assign n54788 = n83038 & n54787 ;
  assign n54789 = n54757 | n54788 ;
  assign n54758 = n54231 & n54233 ;
  assign n54759 = n21731 & n53955 ;
  assign n54760 = n82737 & n54759 ;
  assign n54761 = n65429 | n54760 ;
  assign n83039 = ~n54761 ;
  assign n54762 = n54236 & n83039 ;
  assign n54763 = n82892 & n54762 ;
  assign n54764 = n54758 | n54763 ;
  assign n54765 = n65686 & n54764 ;
  assign n54766 = n22540 & n82892 ;
  assign n83040 = ~n54766 ;
  assign n54767 = x12 & n83040 ;
  assign n54768 = n22550 & n82892 ;
  assign n54769 = n54767 | n54768 ;
  assign n54770 = x65 & n54769 ;
  assign n54362 = n54222 | n54360 ;
  assign n54771 = n82885 & n54362 ;
  assign n54772 = n54227 | n54771 ;
  assign n54773 = n82888 & n54772 ;
  assign n83041 = ~n54773 ;
  assign n54774 = n22540 & n83041 ;
  assign n83042 = ~n54774 ;
  assign n54775 = x12 & n83042 ;
  assign n54776 = x65 | n54768 ;
  assign n54777 = n54775 | n54776 ;
  assign n83043 = ~n54770 ;
  assign n54778 = n83043 & n54777 ;
  assign n54779 = n22557 | n54778 ;
  assign n54780 = n54768 | n54775 ;
  assign n54781 = n65670 & n54780 ;
  assign n83044 = ~n54781 ;
  assign n54782 = n54779 & n83044 ;
  assign n83045 = ~n54763 ;
  assign n54783 = x66 & n83045 ;
  assign n83046 = ~n54758 ;
  assign n54784 = n83046 & n54783 ;
  assign n54785 = n54765 | n54784 ;
  assign n54786 = n54782 | n54785 ;
  assign n83047 = ~n54765 ;
  assign n54790 = n83047 & n54786 ;
  assign n54791 = n54789 | n54790 ;
  assign n83048 = ~n54757 ;
  assign n54792 = n83048 & n54791 ;
  assign n83049 = ~n54746 ;
  assign n54793 = x68 & n83049 ;
  assign n83050 = ~n54741 ;
  assign n54794 = n83050 & n54793 ;
  assign n54795 = n54748 | n54794 ;
  assign n54796 = n54792 | n54795 ;
  assign n83051 = ~n54748 ;
  assign n54800 = n83051 & n54796 ;
  assign n54801 = n54799 | n54800 ;
  assign n83052 = ~n54740 ;
  assign n54802 = n83052 & n54801 ;
  assign n83053 = ~n54729 ;
  assign n54803 = x70 & n83053 ;
  assign n83054 = ~n54724 ;
  assign n54804 = n83054 & n54803 ;
  assign n54805 = n54731 | n54804 ;
  assign n54807 = n54802 | n54805 ;
  assign n83055 = ~n54731 ;
  assign n54811 = n83055 & n54807 ;
  assign n54812 = n54810 | n54811 ;
  assign n83056 = ~n54723 ;
  assign n54813 = n83056 & n54812 ;
  assign n83057 = ~n54712 ;
  assign n54814 = x72 & n83057 ;
  assign n83058 = ~n54706 ;
  assign n54815 = n83058 & n54814 ;
  assign n54816 = n54714 | n54815 ;
  assign n54817 = n54813 | n54816 ;
  assign n83059 = ~n54714 ;
  assign n54822 = n83059 & n54817 ;
  assign n54823 = n54820 | n54822 ;
  assign n83060 = ~n54705 ;
  assign n54824 = n83060 & n54823 ;
  assign n83061 = ~n54695 ;
  assign n54825 = x74 & n83061 ;
  assign n83062 = ~n54690 ;
  assign n54826 = n83062 & n54825 ;
  assign n54827 = n54697 | n54826 ;
  assign n54829 = n54824 | n54827 ;
  assign n83063 = ~n54697 ;
  assign n54833 = n83063 & n54829 ;
  assign n54834 = n54832 | n54833 ;
  assign n83064 = ~n54689 ;
  assign n54835 = n83064 & n54834 ;
  assign n83065 = ~n54679 ;
  assign n54836 = x76 & n83065 ;
  assign n83066 = ~n54674 ;
  assign n54837 = n83066 & n54836 ;
  assign n54838 = n54681 | n54837 ;
  assign n54839 = n54835 | n54838 ;
  assign n83067 = ~n54681 ;
  assign n54844 = n83067 & n54839 ;
  assign n54845 = n54842 | n54844 ;
  assign n83068 = ~n54673 ;
  assign n54846 = n83068 & n54845 ;
  assign n83069 = ~n54663 ;
  assign n54847 = x78 & n83069 ;
  assign n83070 = ~n54658 ;
  assign n54848 = n83070 & n54847 ;
  assign n54849 = n54665 | n54848 ;
  assign n54851 = n54846 | n54849 ;
  assign n83071 = ~n54665 ;
  assign n54855 = n83071 & n54851 ;
  assign n54856 = n54854 | n54855 ;
  assign n83072 = ~n54657 ;
  assign n54857 = n83072 & n54856 ;
  assign n83073 = ~n54647 ;
  assign n54858 = x80 & n83073 ;
  assign n83074 = ~n54642 ;
  assign n54859 = n83074 & n54858 ;
  assign n54860 = n54649 | n54859 ;
  assign n54861 = n54857 | n54860 ;
  assign n83075 = ~n54649 ;
  assign n54866 = n83075 & n54861 ;
  assign n54867 = n54864 | n54866 ;
  assign n83076 = ~n54641 ;
  assign n54868 = n83076 & n54867 ;
  assign n83077 = ~n54631 ;
  assign n54869 = x82 & n83077 ;
  assign n83078 = ~n54626 ;
  assign n54870 = n83078 & n54869 ;
  assign n54871 = n54633 | n54870 ;
  assign n54873 = n54868 | n54871 ;
  assign n83079 = ~n54633 ;
  assign n54877 = n83079 & n54873 ;
  assign n54878 = n54876 | n54877 ;
  assign n83080 = ~n54625 ;
  assign n54879 = n83080 & n54878 ;
  assign n83081 = ~n54615 ;
  assign n54880 = x84 & n83081 ;
  assign n83082 = ~n54610 ;
  assign n54881 = n83082 & n54880 ;
  assign n54882 = n54617 | n54881 ;
  assign n54884 = n54879 | n54882 ;
  assign n83083 = ~n54617 ;
  assign n54888 = n83083 & n54884 ;
  assign n54889 = n54887 | n54888 ;
  assign n83084 = ~n54609 ;
  assign n54890 = n83084 & n54889 ;
  assign n83085 = ~n54599 ;
  assign n54891 = x86 & n83085 ;
  assign n83086 = ~n54594 ;
  assign n54892 = n83086 & n54891 ;
  assign n54893 = n54601 | n54892 ;
  assign n54894 = n54890 | n54893 ;
  assign n83087 = ~n54601 ;
  assign n54898 = n83087 & n54894 ;
  assign n54899 = n54897 | n54898 ;
  assign n83088 = ~n54593 ;
  assign n54900 = n83088 & n54899 ;
  assign n83089 = ~n54583 ;
  assign n54901 = x88 & n83089 ;
  assign n83090 = ~n54578 ;
  assign n54902 = n83090 & n54901 ;
  assign n54903 = n54585 | n54902 ;
  assign n54904 = n54900 | n54903 ;
  assign n83091 = ~n54585 ;
  assign n54908 = n83091 & n54904 ;
  assign n54909 = n54907 | n54908 ;
  assign n83092 = ~n54577 ;
  assign n54910 = n83092 & n54909 ;
  assign n83093 = ~n54567 ;
  assign n54911 = x90 & n83093 ;
  assign n83094 = ~n54562 ;
  assign n54912 = n83094 & n54911 ;
  assign n54913 = n54569 | n54912 ;
  assign n54914 = n54910 | n54913 ;
  assign n83095 = ~n54569 ;
  assign n54918 = n83095 & n54914 ;
  assign n54919 = n54917 | n54918 ;
  assign n83096 = ~n54561 ;
  assign n54920 = n83096 & n54919 ;
  assign n83097 = ~n54551 ;
  assign n54921 = x92 & n83097 ;
  assign n83098 = ~n54546 ;
  assign n54922 = n83098 & n54921 ;
  assign n54923 = n54553 | n54922 ;
  assign n54924 = n54920 | n54923 ;
  assign n83099 = ~n54553 ;
  assign n54929 = n83099 & n54924 ;
  assign n54930 = n54927 | n54929 ;
  assign n83100 = ~n54545 ;
  assign n54931 = n83100 & n54930 ;
  assign n83101 = ~n54535 ;
  assign n54932 = x94 & n83101 ;
  assign n83102 = ~n54530 ;
  assign n54933 = n83102 & n54932 ;
  assign n54934 = n54537 | n54933 ;
  assign n54935 = n54931 | n54934 ;
  assign n83103 = ~n54537 ;
  assign n54939 = n83103 & n54935 ;
  assign n54940 = n54938 | n54939 ;
  assign n83104 = ~n54529 ;
  assign n54941 = n83104 & n54940 ;
  assign n83105 = ~n54519 ;
  assign n54942 = x96 & n83105 ;
  assign n83106 = ~n54514 ;
  assign n54943 = n83106 & n54942 ;
  assign n54944 = n54521 | n54943 ;
  assign n54945 = n54941 | n54944 ;
  assign n83107 = ~n54521 ;
  assign n54949 = n83107 & n54945 ;
  assign n54950 = n54948 | n54949 ;
  assign n83108 = ~n54513 ;
  assign n54951 = n83108 & n54950 ;
  assign n83109 = ~n54503 ;
  assign n54952 = x98 & n83109 ;
  assign n83110 = ~n54498 ;
  assign n54953 = n83110 & n54952 ;
  assign n54954 = n54505 | n54953 ;
  assign n54955 = n54951 | n54954 ;
  assign n83111 = ~n54505 ;
  assign n54959 = n83111 & n54955 ;
  assign n54960 = n54958 | n54959 ;
  assign n83112 = ~n54497 ;
  assign n54961 = n83112 & n54960 ;
  assign n83113 = ~n54487 ;
  assign n54962 = x100 & n83113 ;
  assign n83114 = ~n54482 ;
  assign n54963 = n83114 & n54962 ;
  assign n54964 = n54489 | n54963 ;
  assign n54965 = n54961 | n54964 ;
  assign n83115 = ~n54489 ;
  assign n54970 = n83115 & n54965 ;
  assign n54971 = n54968 | n54970 ;
  assign n83116 = ~n54481 ;
  assign n54972 = n83116 & n54971 ;
  assign n83117 = ~n54471 ;
  assign n54973 = x102 & n83117 ;
  assign n83118 = ~n54466 ;
  assign n54974 = n83118 & n54973 ;
  assign n54975 = n54473 | n54974 ;
  assign n54976 = n54972 | n54975 ;
  assign n83119 = ~n54473 ;
  assign n54981 = n83119 & n54976 ;
  assign n54982 = n54979 | n54981 ;
  assign n83120 = ~n54465 ;
  assign n54983 = n83120 & n54982 ;
  assign n83121 = ~n54455 ;
  assign n54984 = x104 & n83121 ;
  assign n83122 = ~n54450 ;
  assign n54985 = n83122 & n54984 ;
  assign n54986 = n54457 | n54985 ;
  assign n54987 = n54983 | n54986 ;
  assign n83123 = ~n54457 ;
  assign n54991 = n83123 & n54987 ;
  assign n54992 = n54990 | n54991 ;
  assign n83124 = ~n54449 ;
  assign n54993 = n83124 & n54992 ;
  assign n83125 = ~n54439 ;
  assign n54994 = x106 & n83125 ;
  assign n83126 = ~n54434 ;
  assign n54995 = n83126 & n54994 ;
  assign n54996 = n54441 | n54995 ;
  assign n54997 = n54993 | n54996 ;
  assign n83127 = ~n54441 ;
  assign n55002 = n83127 & n54997 ;
  assign n55003 = n55000 | n55002 ;
  assign n83128 = ~n54433 ;
  assign n55004 = n83128 & n55003 ;
  assign n83129 = ~n54423 ;
  assign n55005 = x108 & n83129 ;
  assign n83130 = ~n54418 ;
  assign n55006 = n83130 & n55005 ;
  assign n55007 = n54425 | n55006 ;
  assign n55008 = n55004 | n55007 ;
  assign n83131 = ~n54425 ;
  assign n55012 = n83131 & n55008 ;
  assign n55013 = n55011 | n55012 ;
  assign n83132 = ~n54417 ;
  assign n55014 = n83132 & n55013 ;
  assign n83133 = ~n54407 ;
  assign n55015 = x110 & n83133 ;
  assign n83134 = ~n54402 ;
  assign n55016 = n83134 & n55015 ;
  assign n55017 = n54409 | n55016 ;
  assign n55018 = n55014 | n55017 ;
  assign n83135 = ~n54409 ;
  assign n55022 = n83135 & n55018 ;
  assign n55023 = n55021 | n55022 ;
  assign n83136 = ~n54401 ;
  assign n55024 = n83136 & n55023 ;
  assign n83137 = ~n54391 ;
  assign n55025 = x112 & n83137 ;
  assign n83138 = ~n54386 ;
  assign n55026 = n83138 & n55025 ;
  assign n55027 = n54393 | n55026 ;
  assign n55028 = n55024 | n55027 ;
  assign n83139 = ~n54393 ;
  assign n55032 = n83139 & n55028 ;
  assign n55033 = n55031 | n55032 ;
  assign n83140 = ~n54385 ;
  assign n55034 = n83140 & n55033 ;
  assign n83141 = ~n54375 ;
  assign n55035 = x114 & n83141 ;
  assign n83142 = ~n54370 ;
  assign n55036 = n83142 & n55035 ;
  assign n55037 = n54377 | n55036 ;
  assign n55038 = n55034 | n55037 ;
  assign n83143 = ~n54377 ;
  assign n55042 = n83143 & n55038 ;
  assign n55043 = n55041 | n55042 ;
  assign n83144 = ~n54369 ;
  assign n55044 = n83144 & n55043 ;
  assign n83145 = ~n54224 ;
  assign n54228 = n83145 & n54227 ;
  assign n55045 = n53518 | n54227 ;
  assign n83146 = ~n55045 ;
  assign n55046 = n54362 & n83146 ;
  assign n55047 = n54228 | n55046 ;
  assign n55048 = n54231 | n55047 ;
  assign n83147 = ~n53516 ;
  assign n55049 = n83147 & n54231 ;
  assign n83148 = ~n55049 ;
  assign n55050 = n55048 & n83148 ;
  assign n55051 = n72752 & n55050 ;
  assign n83149 = ~n54231 ;
  assign n55052 = n83149 & n55047 ;
  assign n55053 = n53516 & n54231 ;
  assign n83150 = ~n55053 ;
  assign n55054 = x116 & n83150 ;
  assign n83151 = ~n55052 ;
  assign n55055 = n83151 & n55054 ;
  assign n55056 = n465 | n55055 ;
  assign n55057 = n55051 | n55056 ;
  assign n55058 = n55044 | n55057 ;
  assign n55059 = n67021 & n55050 ;
  assign n83152 = ~n55059 ;
  assign n55060 = n55058 & n83152 ;
  assign n55906 = n54369 | n55055 ;
  assign n55907 = n55051 | n55906 ;
  assign n83153 = ~n55907 ;
  assign n55908 = n55043 & n83153 ;
  assign n55062 = x65 & n54780 ;
  assign n83154 = ~n55062 ;
  assign n55063 = n54777 & n83154 ;
  assign n55064 = n22557 | n55063 ;
  assign n55065 = n83044 & n55064 ;
  assign n55066 = n54785 | n55065 ;
  assign n55067 = n83047 & n55066 ;
  assign n55068 = n54789 | n55067 ;
  assign n55069 = n83048 & n55068 ;
  assign n55070 = n54795 | n55069 ;
  assign n55071 = n83051 & n55070 ;
  assign n55072 = n54799 | n55071 ;
  assign n55073 = n83052 & n55072 ;
  assign n55074 = n54805 | n55073 ;
  assign n55075 = n83055 & n55074 ;
  assign n55076 = n54810 | n55075 ;
  assign n55077 = n83056 & n55076 ;
  assign n55078 = n54816 | n55077 ;
  assign n55079 = n83059 & n55078 ;
  assign n55080 = n54820 | n55079 ;
  assign n55081 = n83060 & n55080 ;
  assign n55082 = n54827 | n55081 ;
  assign n55083 = n83063 & n55082 ;
  assign n55084 = n54832 | n55083 ;
  assign n55085 = n83064 & n55084 ;
  assign n55086 = n54838 | n55085 ;
  assign n55087 = n83067 & n55086 ;
  assign n55088 = n54842 | n55087 ;
  assign n55089 = n83068 & n55088 ;
  assign n55090 = n54849 | n55089 ;
  assign n55091 = n83071 & n55090 ;
  assign n55092 = n54854 | n55091 ;
  assign n55093 = n83072 & n55092 ;
  assign n55094 = n54860 | n55093 ;
  assign n55095 = n83075 & n55094 ;
  assign n55096 = n54864 | n55095 ;
  assign n55097 = n83076 & n55096 ;
  assign n55098 = n54871 | n55097 ;
  assign n55099 = n83079 & n55098 ;
  assign n55100 = n54876 | n55099 ;
  assign n55101 = n83080 & n55100 ;
  assign n55102 = n54882 | n55101 ;
  assign n55103 = n83083 & n55102 ;
  assign n55104 = n54887 | n55103 ;
  assign n55105 = n83084 & n55104 ;
  assign n55106 = n54893 | n55105 ;
  assign n55107 = n83087 & n55106 ;
  assign n55108 = n54897 | n55107 ;
  assign n55109 = n83088 & n55108 ;
  assign n55110 = n54903 | n55109 ;
  assign n55111 = n83091 & n55110 ;
  assign n55112 = n54907 | n55111 ;
  assign n55113 = n83092 & n55112 ;
  assign n55114 = n54913 | n55113 ;
  assign n55115 = n83095 & n55114 ;
  assign n55116 = n54917 | n55115 ;
  assign n55117 = n83096 & n55116 ;
  assign n55118 = n54923 | n55117 ;
  assign n55119 = n83099 & n55118 ;
  assign n55120 = n54927 | n55119 ;
  assign n55121 = n83100 & n55120 ;
  assign n55122 = n54934 | n55121 ;
  assign n55123 = n83103 & n55122 ;
  assign n55124 = n54938 | n55123 ;
  assign n55125 = n83104 & n55124 ;
  assign n55126 = n54944 | n55125 ;
  assign n55127 = n83107 & n55126 ;
  assign n55128 = n54948 | n55127 ;
  assign n55129 = n83108 & n55128 ;
  assign n55130 = n54954 | n55129 ;
  assign n55131 = n83111 & n55130 ;
  assign n55132 = n54958 | n55131 ;
  assign n55133 = n83112 & n55132 ;
  assign n55134 = n54964 | n55133 ;
  assign n55135 = n83115 & n55134 ;
  assign n55136 = n54968 | n55135 ;
  assign n55137 = n83116 & n55136 ;
  assign n55138 = n54975 | n55137 ;
  assign n55139 = n83119 & n55138 ;
  assign n55140 = n54979 | n55139 ;
  assign n55141 = n83120 & n55140 ;
  assign n55142 = n54986 | n55141 ;
  assign n55143 = n83123 & n55142 ;
  assign n55144 = n54990 | n55143 ;
  assign n55145 = n83124 & n55144 ;
  assign n55146 = n54996 | n55145 ;
  assign n55147 = n83127 & n55146 ;
  assign n55148 = n55000 | n55147 ;
  assign n55149 = n83128 & n55148 ;
  assign n55150 = n55007 | n55149 ;
  assign n55151 = n83131 & n55150 ;
  assign n55152 = n55011 | n55151 ;
  assign n55153 = n83132 & n55152 ;
  assign n55154 = n55017 | n55153 ;
  assign n55155 = n83135 & n55154 ;
  assign n55156 = n55021 | n55155 ;
  assign n55157 = n83136 & n55156 ;
  assign n55158 = n55027 | n55157 ;
  assign n55159 = n83139 & n55158 ;
  assign n55160 = n55031 | n55159 ;
  assign n55161 = n83140 & n55160 ;
  assign n55162 = n55037 | n55161 ;
  assign n55163 = n83143 & n55162 ;
  assign n55613 = n55041 | n55163 ;
  assign n55614 = n83144 & n55613 ;
  assign n55909 = n55051 | n55055 ;
  assign n83155 = ~n55614 ;
  assign n55910 = n83155 & n55909 ;
  assign n55911 = n55908 | n55910 ;
  assign n83156 = ~n55060 ;
  assign n55912 = n83156 & n55911 ;
  assign n55913 = n65429 & n53516 ;
  assign n55914 = n55058 & n55913 ;
  assign n55915 = n55912 | n55914 ;
  assign n55921 = n67026 & n55915 ;
  assign n83157 = ~n55042 ;
  assign n55164 = n55041 & n83157 ;
  assign n55165 = n54377 | n55041 ;
  assign n83158 = ~n55165 ;
  assign n55166 = n55162 & n83158 ;
  assign n55167 = n55164 | n55166 ;
  assign n55168 = n83156 & n55167 ;
  assign n55169 = n54368 & n83152 ;
  assign n55170 = n55058 & n55169 ;
  assign n55171 = n55168 | n55170 ;
  assign n55172 = n72752 & n55171 ;
  assign n83159 = ~n55161 ;
  assign n55173 = n55037 & n83159 ;
  assign n55174 = n54385 | n55037 ;
  assign n83160 = ~n55174 ;
  assign n55175 = n55033 & n83160 ;
  assign n55176 = n55173 | n55175 ;
  assign n55177 = n83156 & n55176 ;
  assign n55178 = n54376 & n83152 ;
  assign n55179 = n55058 & n55178 ;
  assign n55180 = n55177 | n55179 ;
  assign n55181 = n72393 & n55180 ;
  assign n83161 = ~n55032 ;
  assign n55182 = n55031 & n83161 ;
  assign n55183 = n54393 | n55031 ;
  assign n83162 = ~n55183 ;
  assign n55184 = n55158 & n83162 ;
  assign n55185 = n55182 | n55184 ;
  assign n55186 = n83156 & n55185 ;
  assign n55187 = n54384 & n83152 ;
  assign n55188 = n55058 & n55187 ;
  assign n55189 = n55186 | n55188 ;
  assign n55190 = n72385 & n55189 ;
  assign n83163 = ~n55157 ;
  assign n55191 = n55027 & n83163 ;
  assign n55192 = n54401 | n55027 ;
  assign n83164 = ~n55192 ;
  assign n55193 = n55023 & n83164 ;
  assign n55194 = n55191 | n55193 ;
  assign n55195 = n83156 & n55194 ;
  assign n55196 = n54392 & n83152 ;
  assign n55197 = n55058 & n55196 ;
  assign n55198 = n55195 | n55197 ;
  assign n55199 = n72025 & n55198 ;
  assign n83165 = ~n55022 ;
  assign n55200 = n55021 & n83165 ;
  assign n55201 = n54409 | n55021 ;
  assign n83166 = ~n55201 ;
  assign n55202 = n55154 & n83166 ;
  assign n55203 = n55200 | n55202 ;
  assign n55204 = n83156 & n55203 ;
  assign n55205 = n54400 & n83152 ;
  assign n55206 = n55058 & n55205 ;
  assign n55207 = n55204 | n55206 ;
  assign n55208 = n71645 & n55207 ;
  assign n83167 = ~n55153 ;
  assign n55209 = n55017 & n83167 ;
  assign n55210 = n54417 | n55017 ;
  assign n83168 = ~n55210 ;
  assign n55211 = n55013 & n83168 ;
  assign n55212 = n55209 | n55211 ;
  assign n55213 = n83156 & n55212 ;
  assign n55214 = n54408 & n83152 ;
  assign n55215 = n55058 & n55214 ;
  assign n55216 = n55213 | n55215 ;
  assign n55217 = n71633 & n55216 ;
  assign n83169 = ~n55012 ;
  assign n55218 = n55011 & n83169 ;
  assign n55219 = n54425 | n55011 ;
  assign n83170 = ~n55219 ;
  assign n55220 = n55150 & n83170 ;
  assign n55221 = n55218 | n55220 ;
  assign n55222 = n83156 & n55221 ;
  assign n55223 = n54416 & n83152 ;
  assign n55224 = n55058 & n55223 ;
  assign n55225 = n55222 | n55224 ;
  assign n55226 = n71253 & n55225 ;
  assign n83171 = ~n55149 ;
  assign n55227 = n55007 & n83171 ;
  assign n55228 = n54433 | n55007 ;
  assign n83172 = ~n55228 ;
  assign n55229 = n55003 & n83172 ;
  assign n55230 = n55227 | n55229 ;
  assign n55231 = n83156 & n55230 ;
  assign n55232 = n54424 & n83152 ;
  assign n55233 = n55058 & n55232 ;
  assign n55234 = n55231 | n55233 ;
  assign n55235 = n70935 & n55234 ;
  assign n83173 = ~n55002 ;
  assign n55236 = n55000 & n83173 ;
  assign n55001 = n54441 | n55000 ;
  assign n83174 = ~n55001 ;
  assign n55237 = n54997 & n83174 ;
  assign n55238 = n55236 | n55237 ;
  assign n55239 = n83156 & n55238 ;
  assign n55240 = n54432 & n83152 ;
  assign n55241 = n55058 & n55240 ;
  assign n55242 = n55239 | n55241 ;
  assign n55243 = n70927 & n55242 ;
  assign n83175 = ~n55145 ;
  assign n55244 = n54996 & n83175 ;
  assign n55245 = n54449 | n54996 ;
  assign n83176 = ~n55245 ;
  assign n55246 = n54992 & n83176 ;
  assign n55247 = n55244 | n55246 ;
  assign n55248 = n83156 & n55247 ;
  assign n55249 = n54440 & n83152 ;
  assign n55250 = n55058 & n55249 ;
  assign n55251 = n55248 | n55250 ;
  assign n55252 = n70609 & n55251 ;
  assign n83177 = ~n54991 ;
  assign n55253 = n54990 & n83177 ;
  assign n55254 = n54457 | n54990 ;
  assign n83178 = ~n55254 ;
  assign n55255 = n55142 & n83178 ;
  assign n55256 = n55253 | n55255 ;
  assign n55257 = n83156 & n55256 ;
  assign n55258 = n54448 & n83152 ;
  assign n55259 = n55058 & n55258 ;
  assign n55260 = n55257 | n55259 ;
  assign n55261 = n70276 & n55260 ;
  assign n83179 = ~n55141 ;
  assign n55262 = n54986 & n83179 ;
  assign n55263 = n54465 | n54986 ;
  assign n83180 = ~n55263 ;
  assign n55264 = n54982 & n83180 ;
  assign n55265 = n55262 | n55264 ;
  assign n55266 = n83156 & n55265 ;
  assign n55267 = n54456 & n83152 ;
  assign n55268 = n55058 & n55267 ;
  assign n55269 = n55266 | n55268 ;
  assign n55270 = n70176 & n55269 ;
  assign n83181 = ~n54981 ;
  assign n55271 = n54979 & n83181 ;
  assign n54980 = n54473 | n54979 ;
  assign n83182 = ~n54980 ;
  assign n55272 = n54976 & n83182 ;
  assign n55273 = n55271 | n55272 ;
  assign n55274 = n83156 & n55273 ;
  assign n55275 = n54464 & n83152 ;
  assign n55276 = n55058 & n55275 ;
  assign n55277 = n55274 | n55276 ;
  assign n55278 = n69857 & n55277 ;
  assign n83183 = ~n55137 ;
  assign n55279 = n54975 & n83183 ;
  assign n55280 = n54481 | n54975 ;
  assign n83184 = ~n55280 ;
  assign n55281 = n54971 & n83184 ;
  assign n55282 = n55279 | n55281 ;
  assign n55283 = n83156 & n55282 ;
  assign n55284 = n54472 & n83152 ;
  assign n55285 = n55058 & n55284 ;
  assign n55286 = n55283 | n55285 ;
  assign n55287 = n69656 & n55286 ;
  assign n83185 = ~n54970 ;
  assign n55288 = n54968 & n83185 ;
  assign n54969 = n54489 | n54968 ;
  assign n83186 = ~n54969 ;
  assign n55289 = n54965 & n83186 ;
  assign n55290 = n55288 | n55289 ;
  assign n55291 = n83156 & n55290 ;
  assign n55292 = n54480 & n83152 ;
  assign n55293 = n55058 & n55292 ;
  assign n55294 = n55291 | n55293 ;
  assign n55295 = n69528 & n55294 ;
  assign n83187 = ~n55133 ;
  assign n55296 = n54964 & n83187 ;
  assign n55297 = n54497 | n54964 ;
  assign n83188 = ~n55297 ;
  assign n55298 = n54960 & n83188 ;
  assign n55299 = n55296 | n55298 ;
  assign n55300 = n83156 & n55299 ;
  assign n55301 = n54488 & n83152 ;
  assign n55302 = n55058 & n55301 ;
  assign n55303 = n55300 | n55302 ;
  assign n55304 = n69261 & n55303 ;
  assign n83189 = ~n54959 ;
  assign n55305 = n54958 & n83189 ;
  assign n55306 = n54505 | n54958 ;
  assign n83190 = ~n55306 ;
  assign n55307 = n55130 & n83190 ;
  assign n55308 = n55305 | n55307 ;
  assign n55309 = n83156 & n55308 ;
  assign n55310 = n54496 & n83152 ;
  assign n55311 = n55058 & n55310 ;
  assign n55312 = n55309 | n55311 ;
  assign n55313 = n69075 & n55312 ;
  assign n83191 = ~n55129 ;
  assign n55314 = n54954 & n83191 ;
  assign n55315 = n54513 | n54954 ;
  assign n83192 = ~n55315 ;
  assign n55316 = n54950 & n83192 ;
  assign n55317 = n55314 | n55316 ;
  assign n55318 = n83156 & n55317 ;
  assign n55319 = n54504 & n83152 ;
  assign n55320 = n55058 & n55319 ;
  assign n55321 = n55318 | n55320 ;
  assign n55322 = n68993 & n55321 ;
  assign n83193 = ~n54949 ;
  assign n55323 = n54948 & n83193 ;
  assign n55324 = n54521 | n54948 ;
  assign n83194 = ~n55324 ;
  assign n55325 = n55126 & n83194 ;
  assign n55326 = n55323 | n55325 ;
  assign n55327 = n83156 & n55326 ;
  assign n55328 = n54512 & n83152 ;
  assign n55329 = n55058 & n55328 ;
  assign n55330 = n55327 | n55329 ;
  assign n55331 = n68716 & n55330 ;
  assign n83195 = ~n55125 ;
  assign n55332 = n54944 & n83195 ;
  assign n55333 = n54529 | n54944 ;
  assign n83196 = ~n55333 ;
  assign n55334 = n54940 & n83196 ;
  assign n55335 = n55332 | n55334 ;
  assign n55336 = n83156 & n55335 ;
  assign n55337 = n54520 & n83152 ;
  assign n55338 = n55058 & n55337 ;
  assign n55339 = n55336 | n55338 ;
  assign n55340 = n68545 & n55339 ;
  assign n83197 = ~n54939 ;
  assign n55341 = n54938 & n83197 ;
  assign n55342 = n54537 | n54938 ;
  assign n83198 = ~n55342 ;
  assign n55343 = n55122 & n83198 ;
  assign n55344 = n55341 | n55343 ;
  assign n55345 = n83156 & n55344 ;
  assign n55346 = n54528 & n83152 ;
  assign n55347 = n55058 & n55346 ;
  assign n55348 = n55345 | n55347 ;
  assign n55349 = n68438 & n55348 ;
  assign n83199 = ~n55121 ;
  assign n55350 = n54934 & n83199 ;
  assign n55351 = n54545 | n54934 ;
  assign n83200 = ~n55351 ;
  assign n55352 = n54930 & n83200 ;
  assign n55353 = n55350 | n55352 ;
  assign n55354 = n83156 & n55353 ;
  assign n55355 = n54536 & n83152 ;
  assign n55356 = n55058 & n55355 ;
  assign n55357 = n55354 | n55356 ;
  assign n55358 = n68214 & n55357 ;
  assign n83201 = ~n54929 ;
  assign n55359 = n54927 & n83201 ;
  assign n54928 = n54553 | n54927 ;
  assign n83202 = ~n54928 ;
  assign n55360 = n54924 & n83202 ;
  assign n55361 = n55359 | n55360 ;
  assign n55362 = n83156 & n55361 ;
  assign n55363 = n54544 & n83152 ;
  assign n55364 = n55058 & n55363 ;
  assign n55365 = n55362 | n55364 ;
  assign n55366 = n68058 & n55365 ;
  assign n83203 = ~n55117 ;
  assign n55367 = n54923 & n83203 ;
  assign n55368 = n54561 | n54923 ;
  assign n83204 = ~n55368 ;
  assign n55369 = n54919 & n83204 ;
  assign n55370 = n55367 | n55369 ;
  assign n55371 = n83156 & n55370 ;
  assign n55372 = n54552 & n83152 ;
  assign n55373 = n55058 & n55372 ;
  assign n55374 = n55371 | n55373 ;
  assign n55375 = n67986 & n55374 ;
  assign n83205 = ~n54918 ;
  assign n55376 = n54917 & n83205 ;
  assign n55377 = n54569 | n54917 ;
  assign n83206 = ~n55377 ;
  assign n55378 = n55114 & n83206 ;
  assign n55379 = n55376 | n55378 ;
  assign n55380 = n83156 & n55379 ;
  assign n55381 = n54560 & n83152 ;
  assign n55382 = n55058 & n55381 ;
  assign n55383 = n55380 | n55382 ;
  assign n55384 = n67763 & n55383 ;
  assign n83207 = ~n55113 ;
  assign n55385 = n54913 & n83207 ;
  assign n55386 = n54577 | n54913 ;
  assign n83208 = ~n55386 ;
  assign n55387 = n54909 & n83208 ;
  assign n55388 = n55385 | n55387 ;
  assign n55389 = n83156 & n55388 ;
  assign n55390 = n54568 & n83152 ;
  assign n55391 = n55058 & n55390 ;
  assign n55392 = n55389 | n55391 ;
  assign n55393 = n67622 & n55392 ;
  assign n83209 = ~n54908 ;
  assign n55394 = n54907 & n83209 ;
  assign n55395 = n54585 | n54907 ;
  assign n83210 = ~n55395 ;
  assign n55396 = n55110 & n83210 ;
  assign n55397 = n55394 | n55396 ;
  assign n55398 = n83156 & n55397 ;
  assign n55399 = n54576 & n83152 ;
  assign n55400 = n55058 & n55399 ;
  assign n55401 = n55398 | n55400 ;
  assign n55402 = n67531 & n55401 ;
  assign n83211 = ~n55109 ;
  assign n55403 = n54903 & n83211 ;
  assign n55404 = n54593 | n54903 ;
  assign n83212 = ~n55404 ;
  assign n55405 = n54899 & n83212 ;
  assign n55406 = n55403 | n55405 ;
  assign n55407 = n83156 & n55406 ;
  assign n55408 = n54584 & n83152 ;
  assign n55409 = n55058 & n55408 ;
  assign n55410 = n55407 | n55409 ;
  assign n55411 = n67348 & n55410 ;
  assign n83213 = ~n54898 ;
  assign n55412 = n54897 & n83213 ;
  assign n55413 = n54601 | n54897 ;
  assign n83214 = ~n55413 ;
  assign n55414 = n55106 & n83214 ;
  assign n55415 = n55412 | n55414 ;
  assign n55416 = n83156 & n55415 ;
  assign n55417 = n54592 & n83152 ;
  assign n55418 = n55058 & n55417 ;
  assign n55419 = n55416 | n55418 ;
  assign n55420 = n67222 & n55419 ;
  assign n83215 = ~n55105 ;
  assign n55421 = n54893 & n83215 ;
  assign n55422 = n54609 | n54893 ;
  assign n83216 = ~n55422 ;
  assign n55423 = n54889 & n83216 ;
  assign n55424 = n55421 | n55423 ;
  assign n55425 = n83156 & n55424 ;
  assign n55426 = n54600 & n83152 ;
  assign n55427 = n55058 & n55426 ;
  assign n55428 = n55425 | n55427 ;
  assign n55429 = n67164 & n55428 ;
  assign n83217 = ~n54888 ;
  assign n55430 = n54887 & n83217 ;
  assign n55431 = n54617 | n54887 ;
  assign n83218 = ~n55431 ;
  assign n55432 = n55102 & n83218 ;
  assign n55433 = n55430 | n55432 ;
  assign n55434 = n83156 & n55433 ;
  assign n55435 = n54608 & n83152 ;
  assign n55436 = n55058 & n55435 ;
  assign n55437 = n55434 | n55436 ;
  assign n55438 = n66979 & n55437 ;
  assign n83219 = ~n55101 ;
  assign n55439 = n54882 & n83219 ;
  assign n54883 = n54625 | n54882 ;
  assign n83220 = ~n54883 ;
  assign n55440 = n83220 & n55100 ;
  assign n55441 = n55439 | n55440 ;
  assign n55442 = n83156 & n55441 ;
  assign n55443 = n54616 & n83152 ;
  assign n55444 = n55058 & n55443 ;
  assign n55445 = n55442 | n55444 ;
  assign n55446 = n66868 & n55445 ;
  assign n83221 = ~n54877 ;
  assign n55447 = n54876 & n83221 ;
  assign n55448 = n54633 | n54876 ;
  assign n83222 = ~n55448 ;
  assign n55449 = n55098 & n83222 ;
  assign n55450 = n55447 | n55449 ;
  assign n55451 = n83156 & n55450 ;
  assign n55452 = n54624 & n83152 ;
  assign n55453 = n55058 & n55452 ;
  assign n55454 = n55451 | n55453 ;
  assign n55455 = n66797 & n55454 ;
  assign n83223 = ~n55097 ;
  assign n55456 = n54871 & n83223 ;
  assign n54872 = n54641 | n54871 ;
  assign n83224 = ~n54872 ;
  assign n55457 = n83224 & n55096 ;
  assign n55458 = n55456 | n55457 ;
  assign n55459 = n83156 & n55458 ;
  assign n55460 = n54632 & n83152 ;
  assign n55461 = n55058 & n55460 ;
  assign n55462 = n55459 | n55461 ;
  assign n55463 = n66654 & n55462 ;
  assign n83225 = ~n54866 ;
  assign n55464 = n54864 & n83225 ;
  assign n54865 = n54649 | n54864 ;
  assign n83226 = ~n54865 ;
  assign n55465 = n54861 & n83226 ;
  assign n55466 = n55464 | n55465 ;
  assign n55467 = n83156 & n55466 ;
  assign n55468 = n54640 & n83152 ;
  assign n55469 = n55058 & n55468 ;
  assign n55470 = n55467 | n55469 ;
  assign n55471 = n66560 & n55470 ;
  assign n83227 = ~n55093 ;
  assign n55472 = n54860 & n83227 ;
  assign n55473 = n54657 | n54860 ;
  assign n83228 = ~n55473 ;
  assign n55474 = n54856 & n83228 ;
  assign n55475 = n55472 | n55474 ;
  assign n55476 = n83156 & n55475 ;
  assign n55477 = n54648 & n83152 ;
  assign n55478 = n55058 & n55477 ;
  assign n55479 = n55476 | n55478 ;
  assign n55480 = n66505 & n55479 ;
  assign n83229 = ~n54855 ;
  assign n55481 = n54854 & n83229 ;
  assign n55482 = n54665 | n54854 ;
  assign n83230 = ~n55482 ;
  assign n55483 = n55090 & n83230 ;
  assign n55484 = n55481 | n55483 ;
  assign n55485 = n83156 & n55484 ;
  assign n55486 = n54656 & n83152 ;
  assign n55487 = n55058 & n55486 ;
  assign n55488 = n55485 | n55487 ;
  assign n55489 = n66379 & n55488 ;
  assign n83231 = ~n55089 ;
  assign n55490 = n54849 & n83231 ;
  assign n54850 = n54673 | n54849 ;
  assign n83232 = ~n54850 ;
  assign n55491 = n83232 & n55088 ;
  assign n55492 = n55490 | n55491 ;
  assign n55493 = n83156 & n55492 ;
  assign n55494 = n54664 & n83152 ;
  assign n55495 = n55058 & n55494 ;
  assign n55496 = n55493 | n55495 ;
  assign n55497 = n66299 & n55496 ;
  assign n83233 = ~n54844 ;
  assign n55498 = n54842 & n83233 ;
  assign n54843 = n54681 | n54842 ;
  assign n83234 = ~n54843 ;
  assign n55499 = n54839 & n83234 ;
  assign n55500 = n55498 | n55499 ;
  assign n55501 = n83156 & n55500 ;
  assign n55502 = n54672 & n83152 ;
  assign n55503 = n55058 & n55502 ;
  assign n55504 = n55501 | n55503 ;
  assign n55505 = n66244 & n55504 ;
  assign n83235 = ~n55085 ;
  assign n55506 = n54838 & n83235 ;
  assign n55507 = n54689 | n54838 ;
  assign n83236 = ~n55507 ;
  assign n55508 = n54834 & n83236 ;
  assign n55509 = n55506 | n55508 ;
  assign n55510 = n83156 & n55509 ;
  assign n55511 = n54680 & n83152 ;
  assign n55512 = n55058 & n55511 ;
  assign n55513 = n55510 | n55512 ;
  assign n55514 = n66145 & n55513 ;
  assign n83237 = ~n54833 ;
  assign n55515 = n54832 & n83237 ;
  assign n55516 = n54697 | n54832 ;
  assign n83238 = ~n55516 ;
  assign n55517 = n55082 & n83238 ;
  assign n55518 = n55515 | n55517 ;
  assign n55519 = n83156 & n55518 ;
  assign n55520 = n54688 & n83152 ;
  assign n55521 = n55058 & n55520 ;
  assign n55522 = n55519 | n55521 ;
  assign n55523 = n66081 & n55522 ;
  assign n83239 = ~n55081 ;
  assign n55524 = n54827 & n83239 ;
  assign n54828 = n54705 | n54827 ;
  assign n83240 = ~n54828 ;
  assign n55525 = n83240 & n55080 ;
  assign n55526 = n55524 | n55525 ;
  assign n55527 = n83156 & n55526 ;
  assign n55528 = n54696 & n83152 ;
  assign n55529 = n55058 & n55528 ;
  assign n55530 = n55527 | n55529 ;
  assign n55531 = n66043 & n55530 ;
  assign n83241 = ~n54822 ;
  assign n55532 = n54820 & n83241 ;
  assign n54821 = n54714 | n54820 ;
  assign n83242 = ~n54821 ;
  assign n55533 = n54817 & n83242 ;
  assign n55534 = n55532 | n55533 ;
  assign n55535 = n83156 & n55534 ;
  assign n55536 = n54704 & n83152 ;
  assign n55537 = n55058 & n55536 ;
  assign n55538 = n55535 | n55537 ;
  assign n55539 = n65960 & n55538 ;
  assign n83243 = ~n55077 ;
  assign n55540 = n54816 & n83243 ;
  assign n55541 = n54723 | n54816 ;
  assign n83244 = ~n55541 ;
  assign n55542 = n54812 & n83244 ;
  assign n55543 = n55540 | n55542 ;
  assign n55544 = n83156 & n55543 ;
  assign n55545 = n54713 & n83152 ;
  assign n55546 = n55058 & n55545 ;
  assign n55547 = n55544 | n55546 ;
  assign n55548 = n65909 & n55547 ;
  assign n83245 = ~n54811 ;
  assign n55549 = n54810 & n83245 ;
  assign n55550 = n54731 | n54810 ;
  assign n83246 = ~n55550 ;
  assign n55551 = n55074 & n83246 ;
  assign n55552 = n55549 | n55551 ;
  assign n55553 = n83156 & n55552 ;
  assign n55554 = n54722 & n83152 ;
  assign n55555 = n55058 & n55554 ;
  assign n55556 = n55553 | n55555 ;
  assign n55557 = n65877 & n55556 ;
  assign n83247 = ~n55073 ;
  assign n55558 = n54805 & n83247 ;
  assign n54806 = n54740 | n54805 ;
  assign n83248 = ~n54806 ;
  assign n55559 = n83248 & n55072 ;
  assign n55560 = n55558 | n55559 ;
  assign n55561 = n83156 & n55560 ;
  assign n55562 = n54730 & n83152 ;
  assign n55563 = n55058 & n55562 ;
  assign n55564 = n55561 | n55563 ;
  assign n55565 = n65820 & n55564 ;
  assign n83249 = ~n54800 ;
  assign n55566 = n54799 & n83249 ;
  assign n55567 = n54748 | n54799 ;
  assign n83250 = ~n55567 ;
  assign n55568 = n55070 & n83250 ;
  assign n55569 = n55566 | n55568 ;
  assign n55570 = n83156 & n55569 ;
  assign n55571 = n54739 & n83152 ;
  assign n55572 = n55058 & n55571 ;
  assign n55573 = n55570 | n55572 ;
  assign n55574 = n65791 & n55573 ;
  assign n83251 = ~n55069 ;
  assign n55576 = n54795 & n83251 ;
  assign n55575 = n54757 | n54795 ;
  assign n83252 = ~n55575 ;
  assign n55577 = n55068 & n83252 ;
  assign n55578 = n55576 | n55577 ;
  assign n55579 = n83156 & n55578 ;
  assign n55580 = n54747 & n83152 ;
  assign n55581 = n55058 & n55580 ;
  assign n55582 = n55579 | n55581 ;
  assign n55583 = n65772 & n55582 ;
  assign n83253 = ~n54790 ;
  assign n55584 = n54789 & n83253 ;
  assign n55585 = n54765 | n54789 ;
  assign n83254 = ~n55585 ;
  assign n55586 = n55066 & n83254 ;
  assign n55587 = n55584 | n55586 ;
  assign n55588 = n83156 & n55587 ;
  assign n55589 = n54756 & n83152 ;
  assign n55590 = n55058 & n55589 ;
  assign n55591 = n55588 | n55590 ;
  assign n55592 = n65746 & n55591 ;
  assign n83255 = ~n55065 ;
  assign n55594 = n54785 & n83255 ;
  assign n55593 = n54781 | n54785 ;
  assign n83256 = ~n55593 ;
  assign n55595 = n55064 & n83256 ;
  assign n55596 = n55594 | n55595 ;
  assign n55597 = n83156 & n55596 ;
  assign n55598 = n54764 & n83152 ;
  assign n55599 = n55058 & n55598 ;
  assign n55600 = n55597 | n55599 ;
  assign n55601 = n65721 & n55600 ;
  assign n55602 = n22557 & n54777 ;
  assign n55603 = n83154 & n55602 ;
  assign n83257 = ~n55603 ;
  assign n55604 = n55064 & n83257 ;
  assign n55605 = n83156 & n55604 ;
  assign n55606 = n54780 & n83152 ;
  assign n55607 = n55058 & n55606 ;
  assign n55608 = n55605 | n55607 ;
  assign n55609 = n65686 & n55608 ;
  assign n55061 = n22557 & n83156 ;
  assign n55610 = x64 & n83156 ;
  assign n83258 = ~n55610 ;
  assign n55611 = x11 & n83258 ;
  assign n55612 = n55061 | n55611 ;
  assign n55624 = n65670 & n55612 ;
  assign n55615 = n55057 | n55614 ;
  assign n55616 = n83152 & n55615 ;
  assign n83259 = ~n55616 ;
  assign n55617 = x64 & n83259 ;
  assign n83260 = ~n55617 ;
  assign n55618 = x11 & n83260 ;
  assign n55619 = n55061 | n55618 ;
  assign n55620 = x65 & n55619 ;
  assign n55621 = x65 | n55061 ;
  assign n55622 = n55618 | n55621 ;
  assign n83261 = ~n55620 ;
  assign n55623 = n83261 & n55622 ;
  assign n55625 = n23402 | n55623 ;
  assign n83262 = ~n55624 ;
  assign n55626 = n83262 & n55625 ;
  assign n83263 = ~n55607 ;
  assign n55627 = x66 & n83263 ;
  assign n83264 = ~n55605 ;
  assign n55628 = n83264 & n55627 ;
  assign n55629 = n55609 | n55628 ;
  assign n55630 = n55626 | n55629 ;
  assign n83265 = ~n55609 ;
  assign n55631 = n83265 & n55630 ;
  assign n83266 = ~n55599 ;
  assign n55632 = x67 & n83266 ;
  assign n83267 = ~n55597 ;
  assign n55633 = n83267 & n55632 ;
  assign n55634 = n55601 | n55633 ;
  assign n55635 = n55631 | n55634 ;
  assign n83268 = ~n55601 ;
  assign n55636 = n83268 & n55635 ;
  assign n83269 = ~n55590 ;
  assign n55637 = x68 & n83269 ;
  assign n83270 = ~n55588 ;
  assign n55638 = n83270 & n55637 ;
  assign n55639 = n55592 | n55638 ;
  assign n55640 = n55636 | n55639 ;
  assign n83271 = ~n55592 ;
  assign n55641 = n83271 & n55640 ;
  assign n83272 = ~n55581 ;
  assign n55642 = x69 & n83272 ;
  assign n83273 = ~n55579 ;
  assign n55643 = n83273 & n55642 ;
  assign n55644 = n55583 | n55643 ;
  assign n55645 = n55641 | n55644 ;
  assign n83274 = ~n55583 ;
  assign n55646 = n83274 & n55645 ;
  assign n83275 = ~n55572 ;
  assign n55647 = x70 & n83275 ;
  assign n83276 = ~n55570 ;
  assign n55648 = n83276 & n55647 ;
  assign n55649 = n55574 | n55648 ;
  assign n55651 = n55646 | n55649 ;
  assign n83277 = ~n55574 ;
  assign n55652 = n83277 & n55651 ;
  assign n83278 = ~n55563 ;
  assign n55653 = x71 & n83278 ;
  assign n83279 = ~n55561 ;
  assign n55654 = n83279 & n55653 ;
  assign n55655 = n55565 | n55654 ;
  assign n55656 = n55652 | n55655 ;
  assign n83280 = ~n55565 ;
  assign n55657 = n83280 & n55656 ;
  assign n83281 = ~n55555 ;
  assign n55658 = x72 & n83281 ;
  assign n83282 = ~n55553 ;
  assign n55659 = n83282 & n55658 ;
  assign n55660 = n55557 | n55659 ;
  assign n55662 = n55657 | n55660 ;
  assign n83283 = ~n55557 ;
  assign n55663 = n83283 & n55662 ;
  assign n83284 = ~n55546 ;
  assign n55664 = x73 & n83284 ;
  assign n83285 = ~n55544 ;
  assign n55665 = n83285 & n55664 ;
  assign n55666 = n55548 | n55665 ;
  assign n55667 = n55663 | n55666 ;
  assign n83286 = ~n55548 ;
  assign n55668 = n83286 & n55667 ;
  assign n83287 = ~n55537 ;
  assign n55669 = x74 & n83287 ;
  assign n83288 = ~n55535 ;
  assign n55670 = n83288 & n55669 ;
  assign n55671 = n55539 | n55670 ;
  assign n55673 = n55668 | n55671 ;
  assign n83289 = ~n55539 ;
  assign n55674 = n83289 & n55673 ;
  assign n83290 = ~n55529 ;
  assign n55675 = x75 & n83290 ;
  assign n83291 = ~n55527 ;
  assign n55676 = n83291 & n55675 ;
  assign n55677 = n55531 | n55676 ;
  assign n55678 = n55674 | n55677 ;
  assign n83292 = ~n55531 ;
  assign n55679 = n83292 & n55678 ;
  assign n83293 = ~n55521 ;
  assign n55680 = x76 & n83293 ;
  assign n83294 = ~n55519 ;
  assign n55681 = n83294 & n55680 ;
  assign n55682 = n55523 | n55681 ;
  assign n55684 = n55679 | n55682 ;
  assign n83295 = ~n55523 ;
  assign n55685 = n83295 & n55684 ;
  assign n83296 = ~n55512 ;
  assign n55686 = x77 & n83296 ;
  assign n83297 = ~n55510 ;
  assign n55687 = n83297 & n55686 ;
  assign n55688 = n55514 | n55687 ;
  assign n55689 = n55685 | n55688 ;
  assign n83298 = ~n55514 ;
  assign n55690 = n83298 & n55689 ;
  assign n83299 = ~n55503 ;
  assign n55691 = x78 & n83299 ;
  assign n83300 = ~n55501 ;
  assign n55692 = n83300 & n55691 ;
  assign n55693 = n55505 | n55692 ;
  assign n55695 = n55690 | n55693 ;
  assign n83301 = ~n55505 ;
  assign n55696 = n83301 & n55695 ;
  assign n83302 = ~n55495 ;
  assign n55697 = x79 & n83302 ;
  assign n83303 = ~n55493 ;
  assign n55698 = n83303 & n55697 ;
  assign n55699 = n55497 | n55698 ;
  assign n55700 = n55696 | n55699 ;
  assign n83304 = ~n55497 ;
  assign n55701 = n83304 & n55700 ;
  assign n83305 = ~n55487 ;
  assign n55702 = x80 & n83305 ;
  assign n83306 = ~n55485 ;
  assign n55703 = n83306 & n55702 ;
  assign n55704 = n55489 | n55703 ;
  assign n55706 = n55701 | n55704 ;
  assign n83307 = ~n55489 ;
  assign n55707 = n83307 & n55706 ;
  assign n83308 = ~n55478 ;
  assign n55708 = x81 & n83308 ;
  assign n83309 = ~n55476 ;
  assign n55709 = n83309 & n55708 ;
  assign n55710 = n55480 | n55709 ;
  assign n55711 = n55707 | n55710 ;
  assign n83310 = ~n55480 ;
  assign n55712 = n83310 & n55711 ;
  assign n83311 = ~n55469 ;
  assign n55713 = x82 & n83311 ;
  assign n83312 = ~n55467 ;
  assign n55714 = n83312 & n55713 ;
  assign n55715 = n55471 | n55714 ;
  assign n55717 = n55712 | n55715 ;
  assign n83313 = ~n55471 ;
  assign n55718 = n83313 & n55717 ;
  assign n83314 = ~n55461 ;
  assign n55719 = x83 & n83314 ;
  assign n83315 = ~n55459 ;
  assign n55720 = n83315 & n55719 ;
  assign n55721 = n55463 | n55720 ;
  assign n55722 = n55718 | n55721 ;
  assign n83316 = ~n55463 ;
  assign n55723 = n83316 & n55722 ;
  assign n83317 = ~n55453 ;
  assign n55724 = x84 & n83317 ;
  assign n83318 = ~n55451 ;
  assign n55725 = n83318 & n55724 ;
  assign n55726 = n55455 | n55725 ;
  assign n55728 = n55723 | n55726 ;
  assign n83319 = ~n55455 ;
  assign n55729 = n83319 & n55728 ;
  assign n83320 = ~n55444 ;
  assign n55730 = x85 & n83320 ;
  assign n83321 = ~n55442 ;
  assign n55731 = n83321 & n55730 ;
  assign n55732 = n55446 | n55731 ;
  assign n55733 = n55729 | n55732 ;
  assign n83322 = ~n55446 ;
  assign n55734 = n83322 & n55733 ;
  assign n83323 = ~n55436 ;
  assign n55735 = x86 & n83323 ;
  assign n83324 = ~n55434 ;
  assign n55736 = n83324 & n55735 ;
  assign n55737 = n55438 | n55736 ;
  assign n55739 = n55734 | n55737 ;
  assign n83325 = ~n55438 ;
  assign n55740 = n83325 & n55739 ;
  assign n83326 = ~n55427 ;
  assign n55741 = x87 & n83326 ;
  assign n83327 = ~n55425 ;
  assign n55742 = n83327 & n55741 ;
  assign n55743 = n55429 | n55742 ;
  assign n55744 = n55740 | n55743 ;
  assign n83328 = ~n55429 ;
  assign n55745 = n83328 & n55744 ;
  assign n83329 = ~n55418 ;
  assign n55746 = x88 & n83329 ;
  assign n83330 = ~n55416 ;
  assign n55747 = n83330 & n55746 ;
  assign n55748 = n55420 | n55747 ;
  assign n55750 = n55745 | n55748 ;
  assign n83331 = ~n55420 ;
  assign n55751 = n83331 & n55750 ;
  assign n83332 = ~n55409 ;
  assign n55752 = x89 & n83332 ;
  assign n83333 = ~n55407 ;
  assign n55753 = n83333 & n55752 ;
  assign n55754 = n55411 | n55753 ;
  assign n55755 = n55751 | n55754 ;
  assign n83334 = ~n55411 ;
  assign n55756 = n83334 & n55755 ;
  assign n83335 = ~n55400 ;
  assign n55757 = x90 & n83335 ;
  assign n83336 = ~n55398 ;
  assign n55758 = n83336 & n55757 ;
  assign n55759 = n55402 | n55758 ;
  assign n55761 = n55756 | n55759 ;
  assign n83337 = ~n55402 ;
  assign n55762 = n83337 & n55761 ;
  assign n83338 = ~n55391 ;
  assign n55763 = x91 & n83338 ;
  assign n83339 = ~n55389 ;
  assign n55764 = n83339 & n55763 ;
  assign n55765 = n55393 | n55764 ;
  assign n55766 = n55762 | n55765 ;
  assign n83340 = ~n55393 ;
  assign n55767 = n83340 & n55766 ;
  assign n83341 = ~n55382 ;
  assign n55768 = x92 & n83341 ;
  assign n83342 = ~n55380 ;
  assign n55769 = n83342 & n55768 ;
  assign n55770 = n55384 | n55769 ;
  assign n55772 = n55767 | n55770 ;
  assign n83343 = ~n55384 ;
  assign n55773 = n83343 & n55772 ;
  assign n83344 = ~n55373 ;
  assign n55774 = x93 & n83344 ;
  assign n83345 = ~n55371 ;
  assign n55775 = n83345 & n55774 ;
  assign n55776 = n55375 | n55775 ;
  assign n55777 = n55773 | n55776 ;
  assign n83346 = ~n55375 ;
  assign n55778 = n83346 & n55777 ;
  assign n83347 = ~n55364 ;
  assign n55779 = x94 & n83347 ;
  assign n83348 = ~n55362 ;
  assign n55780 = n83348 & n55779 ;
  assign n55781 = n55366 | n55780 ;
  assign n55783 = n55778 | n55781 ;
  assign n83349 = ~n55366 ;
  assign n55784 = n83349 & n55783 ;
  assign n83350 = ~n55356 ;
  assign n55785 = x95 & n83350 ;
  assign n83351 = ~n55354 ;
  assign n55786 = n83351 & n55785 ;
  assign n55787 = n55358 | n55786 ;
  assign n55788 = n55784 | n55787 ;
  assign n83352 = ~n55358 ;
  assign n55789 = n83352 & n55788 ;
  assign n83353 = ~n55347 ;
  assign n55790 = x96 & n83353 ;
  assign n83354 = ~n55345 ;
  assign n55791 = n83354 & n55790 ;
  assign n55792 = n55349 | n55791 ;
  assign n55794 = n55789 | n55792 ;
  assign n83355 = ~n55349 ;
  assign n55795 = n83355 & n55794 ;
  assign n83356 = ~n55338 ;
  assign n55796 = x97 & n83356 ;
  assign n83357 = ~n55336 ;
  assign n55797 = n83357 & n55796 ;
  assign n55798 = n55340 | n55797 ;
  assign n55799 = n55795 | n55798 ;
  assign n83358 = ~n55340 ;
  assign n55800 = n83358 & n55799 ;
  assign n83359 = ~n55329 ;
  assign n55801 = x98 & n83359 ;
  assign n83360 = ~n55327 ;
  assign n55802 = n83360 & n55801 ;
  assign n55803 = n55331 | n55802 ;
  assign n55805 = n55800 | n55803 ;
  assign n83361 = ~n55331 ;
  assign n55806 = n83361 & n55805 ;
  assign n83362 = ~n55320 ;
  assign n55807 = x99 & n83362 ;
  assign n83363 = ~n55318 ;
  assign n55808 = n83363 & n55807 ;
  assign n55809 = n55322 | n55808 ;
  assign n55810 = n55806 | n55809 ;
  assign n83364 = ~n55322 ;
  assign n55811 = n83364 & n55810 ;
  assign n83365 = ~n55311 ;
  assign n55812 = x100 & n83365 ;
  assign n83366 = ~n55309 ;
  assign n55813 = n83366 & n55812 ;
  assign n55814 = n55313 | n55813 ;
  assign n55816 = n55811 | n55814 ;
  assign n83367 = ~n55313 ;
  assign n55817 = n83367 & n55816 ;
  assign n83368 = ~n55302 ;
  assign n55818 = x101 & n83368 ;
  assign n83369 = ~n55300 ;
  assign n55819 = n83369 & n55818 ;
  assign n55820 = n55304 | n55819 ;
  assign n55821 = n55817 | n55820 ;
  assign n83370 = ~n55304 ;
  assign n55822 = n83370 & n55821 ;
  assign n83371 = ~n55293 ;
  assign n55823 = x102 & n83371 ;
  assign n83372 = ~n55291 ;
  assign n55824 = n83372 & n55823 ;
  assign n55825 = n55295 | n55824 ;
  assign n55827 = n55822 | n55825 ;
  assign n83373 = ~n55295 ;
  assign n55828 = n83373 & n55827 ;
  assign n83374 = ~n55285 ;
  assign n55829 = x103 & n83374 ;
  assign n83375 = ~n55283 ;
  assign n55830 = n83375 & n55829 ;
  assign n55831 = n55287 | n55830 ;
  assign n55832 = n55828 | n55831 ;
  assign n83376 = ~n55287 ;
  assign n55833 = n83376 & n55832 ;
  assign n83377 = ~n55276 ;
  assign n55834 = x104 & n83377 ;
  assign n83378 = ~n55274 ;
  assign n55835 = n83378 & n55834 ;
  assign n55836 = n55278 | n55835 ;
  assign n55838 = n55833 | n55836 ;
  assign n83379 = ~n55278 ;
  assign n55839 = n83379 & n55838 ;
  assign n83380 = ~n55268 ;
  assign n55840 = x105 & n83380 ;
  assign n83381 = ~n55266 ;
  assign n55841 = n83381 & n55840 ;
  assign n55842 = n55270 | n55841 ;
  assign n55843 = n55839 | n55842 ;
  assign n83382 = ~n55270 ;
  assign n55844 = n83382 & n55843 ;
  assign n83383 = ~n55259 ;
  assign n55845 = x106 & n83383 ;
  assign n83384 = ~n55257 ;
  assign n55846 = n83384 & n55845 ;
  assign n55847 = n55261 | n55846 ;
  assign n55849 = n55844 | n55847 ;
  assign n83385 = ~n55261 ;
  assign n55850 = n83385 & n55849 ;
  assign n83386 = ~n55250 ;
  assign n55851 = x107 & n83386 ;
  assign n83387 = ~n55248 ;
  assign n55852 = n83387 & n55851 ;
  assign n55853 = n55252 | n55852 ;
  assign n55854 = n55850 | n55853 ;
  assign n83388 = ~n55252 ;
  assign n55855 = n83388 & n55854 ;
  assign n83389 = ~n55241 ;
  assign n55856 = x108 & n83389 ;
  assign n83390 = ~n55239 ;
  assign n55857 = n83390 & n55856 ;
  assign n55858 = n55243 | n55857 ;
  assign n55860 = n55855 | n55858 ;
  assign n83391 = ~n55243 ;
  assign n55861 = n83391 & n55860 ;
  assign n83392 = ~n55233 ;
  assign n55862 = x109 & n83392 ;
  assign n83393 = ~n55231 ;
  assign n55863 = n83393 & n55862 ;
  assign n55864 = n55235 | n55863 ;
  assign n55865 = n55861 | n55864 ;
  assign n83394 = ~n55235 ;
  assign n55866 = n83394 & n55865 ;
  assign n83395 = ~n55224 ;
  assign n55867 = x110 & n83395 ;
  assign n83396 = ~n55222 ;
  assign n55868 = n83396 & n55867 ;
  assign n55869 = n55226 | n55868 ;
  assign n55871 = n55866 | n55869 ;
  assign n83397 = ~n55226 ;
  assign n55872 = n83397 & n55871 ;
  assign n83398 = ~n55215 ;
  assign n55873 = x111 & n83398 ;
  assign n83399 = ~n55213 ;
  assign n55874 = n83399 & n55873 ;
  assign n55875 = n55217 | n55874 ;
  assign n55876 = n55872 | n55875 ;
  assign n83400 = ~n55217 ;
  assign n55877 = n83400 & n55876 ;
  assign n83401 = ~n55206 ;
  assign n55878 = x112 & n83401 ;
  assign n83402 = ~n55204 ;
  assign n55879 = n83402 & n55878 ;
  assign n55880 = n55208 | n55879 ;
  assign n55882 = n55877 | n55880 ;
  assign n83403 = ~n55208 ;
  assign n55883 = n83403 & n55882 ;
  assign n83404 = ~n55197 ;
  assign n55884 = x113 & n83404 ;
  assign n83405 = ~n55195 ;
  assign n55885 = n83405 & n55884 ;
  assign n55886 = n55199 | n55885 ;
  assign n55887 = n55883 | n55886 ;
  assign n83406 = ~n55199 ;
  assign n55888 = n83406 & n55887 ;
  assign n83407 = ~n55188 ;
  assign n55889 = x114 & n83407 ;
  assign n83408 = ~n55186 ;
  assign n55890 = n83408 & n55889 ;
  assign n55891 = n55190 | n55890 ;
  assign n55893 = n55888 | n55891 ;
  assign n83409 = ~n55190 ;
  assign n55894 = n83409 & n55893 ;
  assign n83410 = ~n55179 ;
  assign n55895 = x115 & n83410 ;
  assign n83411 = ~n55177 ;
  assign n55896 = n83411 & n55895 ;
  assign n55897 = n55181 | n55896 ;
  assign n55898 = n55894 | n55897 ;
  assign n83412 = ~n55181 ;
  assign n55899 = n83412 & n55898 ;
  assign n83413 = ~n55170 ;
  assign n55900 = x116 & n83413 ;
  assign n83414 = ~n55168 ;
  assign n55901 = n83414 & n55900 ;
  assign n55902 = n55172 | n55901 ;
  assign n55904 = n55899 | n55902 ;
  assign n83415 = ~n55172 ;
  assign n55905 = n83415 & n55904 ;
  assign n55916 = n73177 & n55915 ;
  assign n83416 = ~n55914 ;
  assign n55917 = x117 & n83416 ;
  assign n83417 = ~n55912 ;
  assign n55918 = n83417 & n55917 ;
  assign n55919 = n23684 | n55918 ;
  assign n55920 = n55916 | n55919 ;
  assign n55922 = n55905 | n55920 ;
  assign n83418 = ~n55921 ;
  assign n55923 = n83418 & n55922 ;
  assign n56066 = n55172 | n55918 ;
  assign n56067 = n55916 | n56066 ;
  assign n83419 = ~n56067 ;
  assign n56068 = n55904 & n83419 ;
  assign n55926 = x65 & n55612 ;
  assign n83420 = ~n55926 ;
  assign n55927 = n55622 & n83420 ;
  assign n55928 = n23402 | n55927 ;
  assign n55929 = n83262 & n55928 ;
  assign n55930 = n55629 | n55929 ;
  assign n55931 = n83265 & n55930 ;
  assign n55933 = n55634 | n55931 ;
  assign n55934 = n83268 & n55933 ;
  assign n55936 = n55639 | n55934 ;
  assign n55937 = n83271 & n55936 ;
  assign n55938 = n55644 | n55937 ;
  assign n55940 = n83274 & n55938 ;
  assign n55941 = n55649 | n55940 ;
  assign n55942 = n83277 & n55941 ;
  assign n55943 = n55655 | n55942 ;
  assign n55945 = n83280 & n55943 ;
  assign n55946 = n55660 | n55945 ;
  assign n55947 = n83283 & n55946 ;
  assign n55948 = n55666 | n55947 ;
  assign n55950 = n83286 & n55948 ;
  assign n55951 = n55671 | n55950 ;
  assign n55952 = n83289 & n55951 ;
  assign n55953 = n55677 | n55952 ;
  assign n55955 = n83292 & n55953 ;
  assign n55956 = n55682 | n55955 ;
  assign n55957 = n83295 & n55956 ;
  assign n55958 = n55688 | n55957 ;
  assign n55960 = n83298 & n55958 ;
  assign n55961 = n55693 | n55960 ;
  assign n55962 = n83301 & n55961 ;
  assign n55963 = n55699 | n55962 ;
  assign n55965 = n83304 & n55963 ;
  assign n55966 = n55704 | n55965 ;
  assign n55967 = n83307 & n55966 ;
  assign n55968 = n55710 | n55967 ;
  assign n55970 = n83310 & n55968 ;
  assign n55971 = n55715 | n55970 ;
  assign n55972 = n83313 & n55971 ;
  assign n55973 = n55721 | n55972 ;
  assign n55975 = n83316 & n55973 ;
  assign n55976 = n55726 | n55975 ;
  assign n55977 = n83319 & n55976 ;
  assign n55978 = n55732 | n55977 ;
  assign n55980 = n83322 & n55978 ;
  assign n55981 = n55737 | n55980 ;
  assign n55982 = n83325 & n55981 ;
  assign n55983 = n55743 | n55982 ;
  assign n55985 = n83328 & n55983 ;
  assign n55986 = n55748 | n55985 ;
  assign n55987 = n83331 & n55986 ;
  assign n55988 = n55754 | n55987 ;
  assign n55990 = n83334 & n55988 ;
  assign n55991 = n55759 | n55990 ;
  assign n55992 = n83337 & n55991 ;
  assign n55993 = n55765 | n55992 ;
  assign n55995 = n83340 & n55993 ;
  assign n55996 = n55770 | n55995 ;
  assign n55997 = n83343 & n55996 ;
  assign n55998 = n55776 | n55997 ;
  assign n56000 = n83346 & n55998 ;
  assign n56001 = n55781 | n56000 ;
  assign n56002 = n83349 & n56001 ;
  assign n56003 = n55787 | n56002 ;
  assign n56005 = n83352 & n56003 ;
  assign n56006 = n55792 | n56005 ;
  assign n56007 = n83355 & n56006 ;
  assign n56008 = n55798 | n56007 ;
  assign n56010 = n83358 & n56008 ;
  assign n56011 = n55803 | n56010 ;
  assign n56012 = n83361 & n56011 ;
  assign n56013 = n55809 | n56012 ;
  assign n56015 = n83364 & n56013 ;
  assign n56016 = n55814 | n56015 ;
  assign n56017 = n83367 & n56016 ;
  assign n56018 = n55820 | n56017 ;
  assign n56020 = n83370 & n56018 ;
  assign n56021 = n55825 | n56020 ;
  assign n56022 = n83373 & n56021 ;
  assign n56023 = n55831 | n56022 ;
  assign n56025 = n83376 & n56023 ;
  assign n56026 = n55836 | n56025 ;
  assign n56027 = n83379 & n56026 ;
  assign n56028 = n55842 | n56027 ;
  assign n56030 = n83382 & n56028 ;
  assign n56031 = n55847 | n56030 ;
  assign n56032 = n83385 & n56031 ;
  assign n56033 = n55853 | n56032 ;
  assign n56035 = n83388 & n56033 ;
  assign n56036 = n55858 | n56035 ;
  assign n56037 = n83391 & n56036 ;
  assign n56038 = n55864 | n56037 ;
  assign n56040 = n83394 & n56038 ;
  assign n56041 = n55869 | n56040 ;
  assign n56042 = n83397 & n56041 ;
  assign n56043 = n55875 | n56042 ;
  assign n56045 = n83400 & n56043 ;
  assign n56046 = n55880 | n56045 ;
  assign n56047 = n83403 & n56046 ;
  assign n56048 = n55886 | n56047 ;
  assign n56050 = n83406 & n56048 ;
  assign n56051 = n55891 | n56050 ;
  assign n56052 = n83409 & n56051 ;
  assign n56054 = n55897 | n56052 ;
  assign n56059 = n83412 & n56054 ;
  assign n56060 = n55902 | n56059 ;
  assign n56061 = n83415 & n56060 ;
  assign n56069 = n55916 | n55918 ;
  assign n83421 = ~n56061 ;
  assign n56070 = n83421 & n56069 ;
  assign n56071 = n56068 | n56070 ;
  assign n83422 = ~n55923 ;
  assign n56072 = n83422 & n56071 ;
  assign n56062 = n55920 | n56061 ;
  assign n56073 = n465 & n55915 ;
  assign n56074 = n56062 & n56073 ;
  assign n56075 = n56072 | n56074 ;
  assign n56076 = n73188 & n56075 ;
  assign n83423 = ~n56074 ;
  assign n56807 = x118 & n83423 ;
  assign n83424 = ~n56072 ;
  assign n56808 = n83424 & n56807 ;
  assign n56809 = n56076 | n56808 ;
  assign n83425 = ~n55899 ;
  assign n55903 = n83425 & n55902 ;
  assign n56055 = n55181 | n55902 ;
  assign n83426 = ~n56055 ;
  assign n56056 = n56054 & n83426 ;
  assign n56057 = n55903 | n56056 ;
  assign n56058 = n83422 & n56057 ;
  assign n56063 = n55171 & n83418 ;
  assign n56064 = n56062 & n56063 ;
  assign n56065 = n56058 | n56064 ;
  assign n56077 = n73177 & n56065 ;
  assign n83427 = ~n56052 ;
  assign n56053 = n55897 & n83427 ;
  assign n56078 = n55190 | n55897 ;
  assign n83428 = ~n56078 ;
  assign n56079 = n55893 & n83428 ;
  assign n56080 = n56053 | n56079 ;
  assign n56081 = n83422 & n56080 ;
  assign n56082 = n55180 & n83418 ;
  assign n56083 = n56062 & n56082 ;
  assign n56084 = n56081 | n56083 ;
  assign n56085 = n72752 & n56084 ;
  assign n83429 = ~n56083 ;
  assign n56795 = x116 & n83429 ;
  assign n83430 = ~n56081 ;
  assign n56796 = n83430 & n56795 ;
  assign n56797 = n56085 | n56796 ;
  assign n83431 = ~n55888 ;
  assign n55892 = n83431 & n55891 ;
  assign n56086 = n55199 | n55891 ;
  assign n83432 = ~n56086 ;
  assign n56087 = n56048 & n83432 ;
  assign n56088 = n55892 | n56087 ;
  assign n56089 = n83422 & n56088 ;
  assign n56090 = n55189 & n83418 ;
  assign n56091 = n56062 & n56090 ;
  assign n56092 = n56089 | n56091 ;
  assign n56093 = n72393 & n56092 ;
  assign n83433 = ~n56047 ;
  assign n56049 = n55886 & n83433 ;
  assign n56094 = n55208 | n55886 ;
  assign n83434 = ~n56094 ;
  assign n56095 = n55882 & n83434 ;
  assign n56096 = n56049 | n56095 ;
  assign n56097 = n83422 & n56096 ;
  assign n56098 = n55198 & n83418 ;
  assign n56099 = n56062 & n56098 ;
  assign n56100 = n56097 | n56099 ;
  assign n56101 = n72385 & n56100 ;
  assign n83435 = ~n56099 ;
  assign n56783 = x114 & n83435 ;
  assign n83436 = ~n56097 ;
  assign n56784 = n83436 & n56783 ;
  assign n56785 = n56101 | n56784 ;
  assign n83437 = ~n55877 ;
  assign n55881 = n83437 & n55880 ;
  assign n56102 = n55217 | n55880 ;
  assign n83438 = ~n56102 ;
  assign n56103 = n56043 & n83438 ;
  assign n56104 = n55881 | n56103 ;
  assign n56105 = n83422 & n56104 ;
  assign n56106 = n55207 & n83418 ;
  assign n56107 = n56062 & n56106 ;
  assign n56108 = n56105 | n56107 ;
  assign n56109 = n72025 & n56108 ;
  assign n83439 = ~n56042 ;
  assign n56044 = n55875 & n83439 ;
  assign n56110 = n55226 | n55875 ;
  assign n83440 = ~n56110 ;
  assign n56111 = n55871 & n83440 ;
  assign n56112 = n56044 | n56111 ;
  assign n56113 = n83422 & n56112 ;
  assign n56114 = n55216 & n83418 ;
  assign n56115 = n56062 & n56114 ;
  assign n56116 = n56113 | n56115 ;
  assign n56117 = n71645 & n56116 ;
  assign n83441 = ~n56115 ;
  assign n56771 = x112 & n83441 ;
  assign n83442 = ~n56113 ;
  assign n56772 = n83442 & n56771 ;
  assign n56773 = n56117 | n56772 ;
  assign n83443 = ~n55866 ;
  assign n55870 = n83443 & n55869 ;
  assign n56118 = n55235 | n55869 ;
  assign n83444 = ~n56118 ;
  assign n56119 = n56038 & n83444 ;
  assign n56120 = n55870 | n56119 ;
  assign n56121 = n83422 & n56120 ;
  assign n56122 = n55225 & n83418 ;
  assign n56123 = n56062 & n56122 ;
  assign n56124 = n56121 | n56123 ;
  assign n56125 = n71633 & n56124 ;
  assign n83445 = ~n56037 ;
  assign n56039 = n55864 & n83445 ;
  assign n56126 = n55243 | n55864 ;
  assign n83446 = ~n56126 ;
  assign n56127 = n55860 & n83446 ;
  assign n56128 = n56039 | n56127 ;
  assign n56129 = n83422 & n56128 ;
  assign n56130 = n55234 & n83418 ;
  assign n56131 = n56062 & n56130 ;
  assign n56132 = n56129 | n56131 ;
  assign n56133 = n71253 & n56132 ;
  assign n83447 = ~n56131 ;
  assign n56759 = x110 & n83447 ;
  assign n83448 = ~n56129 ;
  assign n56760 = n83448 & n56759 ;
  assign n56761 = n56133 | n56760 ;
  assign n83449 = ~n55855 ;
  assign n55859 = n83449 & n55858 ;
  assign n56134 = n55252 | n55858 ;
  assign n83450 = ~n56134 ;
  assign n56135 = n56033 & n83450 ;
  assign n56136 = n55859 | n56135 ;
  assign n56137 = n83422 & n56136 ;
  assign n56138 = n55242 & n83418 ;
  assign n56139 = n56062 & n56138 ;
  assign n56140 = n56137 | n56139 ;
  assign n56141 = n70935 & n56140 ;
  assign n83451 = ~n56032 ;
  assign n56034 = n55853 & n83451 ;
  assign n56142 = n55261 | n55853 ;
  assign n83452 = ~n56142 ;
  assign n56143 = n55849 & n83452 ;
  assign n56144 = n56034 | n56143 ;
  assign n56145 = n83422 & n56144 ;
  assign n56146 = n55251 & n83418 ;
  assign n56147 = n56062 & n56146 ;
  assign n56148 = n56145 | n56147 ;
  assign n56149 = n70927 & n56148 ;
  assign n83453 = ~n56147 ;
  assign n56747 = x108 & n83453 ;
  assign n83454 = ~n56145 ;
  assign n56748 = n83454 & n56747 ;
  assign n56749 = n56149 | n56748 ;
  assign n83455 = ~n55844 ;
  assign n55848 = n83455 & n55847 ;
  assign n56150 = n55270 | n55847 ;
  assign n83456 = ~n56150 ;
  assign n56151 = n56028 & n83456 ;
  assign n56152 = n55848 | n56151 ;
  assign n56153 = n83422 & n56152 ;
  assign n56154 = n55260 & n83418 ;
  assign n56155 = n56062 & n56154 ;
  assign n56156 = n56153 | n56155 ;
  assign n56157 = n70609 & n56156 ;
  assign n83457 = ~n56027 ;
  assign n56029 = n55842 & n83457 ;
  assign n56158 = n55278 | n55842 ;
  assign n83458 = ~n56158 ;
  assign n56159 = n55838 & n83458 ;
  assign n56160 = n56029 | n56159 ;
  assign n56161 = n83422 & n56160 ;
  assign n56162 = n55269 & n83418 ;
  assign n56163 = n56062 & n56162 ;
  assign n56164 = n56161 | n56163 ;
  assign n56165 = n70276 & n56164 ;
  assign n83459 = ~n56163 ;
  assign n56735 = x106 & n83459 ;
  assign n83460 = ~n56161 ;
  assign n56736 = n83460 & n56735 ;
  assign n56737 = n56165 | n56736 ;
  assign n83461 = ~n55833 ;
  assign n55837 = n83461 & n55836 ;
  assign n56166 = n55287 | n55836 ;
  assign n83462 = ~n56166 ;
  assign n56167 = n56023 & n83462 ;
  assign n56168 = n55837 | n56167 ;
  assign n56169 = n83422 & n56168 ;
  assign n56170 = n55277 & n83418 ;
  assign n56171 = n56062 & n56170 ;
  assign n56172 = n56169 | n56171 ;
  assign n56173 = n70176 & n56172 ;
  assign n83463 = ~n56022 ;
  assign n56024 = n55831 & n83463 ;
  assign n56174 = n55295 | n55831 ;
  assign n83464 = ~n56174 ;
  assign n56175 = n55827 & n83464 ;
  assign n56176 = n56024 | n56175 ;
  assign n56177 = n83422 & n56176 ;
  assign n56178 = n55286 & n83418 ;
  assign n56179 = n56062 & n56178 ;
  assign n56180 = n56177 | n56179 ;
  assign n56181 = n69857 & n56180 ;
  assign n83465 = ~n56179 ;
  assign n56723 = x104 & n83465 ;
  assign n83466 = ~n56177 ;
  assign n56724 = n83466 & n56723 ;
  assign n56725 = n56181 | n56724 ;
  assign n83467 = ~n55822 ;
  assign n55826 = n83467 & n55825 ;
  assign n56182 = n55304 | n55825 ;
  assign n83468 = ~n56182 ;
  assign n56183 = n56018 & n83468 ;
  assign n56184 = n55826 | n56183 ;
  assign n56185 = n83422 & n56184 ;
  assign n56186 = n55294 & n83418 ;
  assign n56187 = n56062 & n56186 ;
  assign n56188 = n56185 | n56187 ;
  assign n56189 = n69656 & n56188 ;
  assign n83469 = ~n56017 ;
  assign n56019 = n55820 & n83469 ;
  assign n56190 = n55313 | n55820 ;
  assign n83470 = ~n56190 ;
  assign n56191 = n55816 & n83470 ;
  assign n56192 = n56019 | n56191 ;
  assign n56193 = n83422 & n56192 ;
  assign n56194 = n55303 & n83418 ;
  assign n56195 = n56062 & n56194 ;
  assign n56196 = n56193 | n56195 ;
  assign n56197 = n69528 & n56196 ;
  assign n83471 = ~n56195 ;
  assign n56711 = x102 & n83471 ;
  assign n83472 = ~n56193 ;
  assign n56712 = n83472 & n56711 ;
  assign n56713 = n56197 | n56712 ;
  assign n83473 = ~n55811 ;
  assign n55815 = n83473 & n55814 ;
  assign n56198 = n55322 | n55814 ;
  assign n83474 = ~n56198 ;
  assign n56199 = n56013 & n83474 ;
  assign n56200 = n55815 | n56199 ;
  assign n56201 = n83422 & n56200 ;
  assign n56202 = n55312 & n83418 ;
  assign n56203 = n56062 & n56202 ;
  assign n56204 = n56201 | n56203 ;
  assign n56205 = n69261 & n56204 ;
  assign n83475 = ~n56012 ;
  assign n56014 = n55809 & n83475 ;
  assign n56206 = n55331 | n55809 ;
  assign n83476 = ~n56206 ;
  assign n56207 = n55805 & n83476 ;
  assign n56208 = n56014 | n56207 ;
  assign n56209 = n83422 & n56208 ;
  assign n56210 = n55321 & n83418 ;
  assign n56211 = n56062 & n56210 ;
  assign n56212 = n56209 | n56211 ;
  assign n56213 = n69075 & n56212 ;
  assign n83477 = ~n56211 ;
  assign n56699 = x100 & n83477 ;
  assign n83478 = ~n56209 ;
  assign n56700 = n83478 & n56699 ;
  assign n56701 = n56213 | n56700 ;
  assign n83479 = ~n55800 ;
  assign n55804 = n83479 & n55803 ;
  assign n56214 = n55340 | n55803 ;
  assign n83480 = ~n56214 ;
  assign n56215 = n56008 & n83480 ;
  assign n56216 = n55804 | n56215 ;
  assign n56217 = n83422 & n56216 ;
  assign n56218 = n55330 & n83418 ;
  assign n56219 = n56062 & n56218 ;
  assign n56220 = n56217 | n56219 ;
  assign n56221 = n68993 & n56220 ;
  assign n83481 = ~n56007 ;
  assign n56009 = n55798 & n83481 ;
  assign n56222 = n55349 | n55798 ;
  assign n83482 = ~n56222 ;
  assign n56223 = n55794 & n83482 ;
  assign n56224 = n56009 | n56223 ;
  assign n56225 = n83422 & n56224 ;
  assign n56226 = n55339 & n83418 ;
  assign n56227 = n56062 & n56226 ;
  assign n56228 = n56225 | n56227 ;
  assign n56229 = n68716 & n56228 ;
  assign n83483 = ~n56227 ;
  assign n56687 = x98 & n83483 ;
  assign n83484 = ~n56225 ;
  assign n56688 = n83484 & n56687 ;
  assign n56689 = n56229 | n56688 ;
  assign n83485 = ~n55789 ;
  assign n55793 = n83485 & n55792 ;
  assign n56230 = n55358 | n55792 ;
  assign n83486 = ~n56230 ;
  assign n56231 = n56003 & n83486 ;
  assign n56232 = n55793 | n56231 ;
  assign n56233 = n83422 & n56232 ;
  assign n56234 = n55348 & n83418 ;
  assign n56235 = n56062 & n56234 ;
  assign n56236 = n56233 | n56235 ;
  assign n56237 = n68545 & n56236 ;
  assign n83487 = ~n56002 ;
  assign n56004 = n55787 & n83487 ;
  assign n56238 = n55366 | n55787 ;
  assign n83488 = ~n56238 ;
  assign n56239 = n55783 & n83488 ;
  assign n56240 = n56004 | n56239 ;
  assign n56241 = n83422 & n56240 ;
  assign n56242 = n55357 & n83418 ;
  assign n56243 = n56062 & n56242 ;
  assign n56244 = n56241 | n56243 ;
  assign n56245 = n68438 & n56244 ;
  assign n83489 = ~n56243 ;
  assign n56675 = x96 & n83489 ;
  assign n83490 = ~n56241 ;
  assign n56676 = n83490 & n56675 ;
  assign n56677 = n56245 | n56676 ;
  assign n83491 = ~n55778 ;
  assign n55782 = n83491 & n55781 ;
  assign n56246 = n55375 | n55781 ;
  assign n83492 = ~n56246 ;
  assign n56247 = n55998 & n83492 ;
  assign n56248 = n55782 | n56247 ;
  assign n56249 = n83422 & n56248 ;
  assign n56250 = n55365 & n83418 ;
  assign n56251 = n56062 & n56250 ;
  assign n56252 = n56249 | n56251 ;
  assign n56253 = n68214 & n56252 ;
  assign n83493 = ~n55997 ;
  assign n55999 = n55776 & n83493 ;
  assign n56254 = n55384 | n55776 ;
  assign n83494 = ~n56254 ;
  assign n56255 = n55772 & n83494 ;
  assign n56256 = n55999 | n56255 ;
  assign n56257 = n83422 & n56256 ;
  assign n56258 = n55374 & n83418 ;
  assign n56259 = n56062 & n56258 ;
  assign n56260 = n56257 | n56259 ;
  assign n56261 = n68058 & n56260 ;
  assign n83495 = ~n56259 ;
  assign n56663 = x94 & n83495 ;
  assign n83496 = ~n56257 ;
  assign n56664 = n83496 & n56663 ;
  assign n56665 = n56261 | n56664 ;
  assign n83497 = ~n55767 ;
  assign n55771 = n83497 & n55770 ;
  assign n56262 = n55393 | n55770 ;
  assign n83498 = ~n56262 ;
  assign n56263 = n55993 & n83498 ;
  assign n56264 = n55771 | n56263 ;
  assign n56265 = n83422 & n56264 ;
  assign n56266 = n55383 & n83418 ;
  assign n56267 = n56062 & n56266 ;
  assign n56268 = n56265 | n56267 ;
  assign n56269 = n67986 & n56268 ;
  assign n83499 = ~n55992 ;
  assign n55994 = n55765 & n83499 ;
  assign n56270 = n55402 | n55765 ;
  assign n83500 = ~n56270 ;
  assign n56271 = n55761 & n83500 ;
  assign n56272 = n55994 | n56271 ;
  assign n56273 = n83422 & n56272 ;
  assign n56274 = n55392 & n83418 ;
  assign n56275 = n56062 & n56274 ;
  assign n56276 = n56273 | n56275 ;
  assign n56277 = n67763 & n56276 ;
  assign n83501 = ~n56275 ;
  assign n56651 = x92 & n83501 ;
  assign n83502 = ~n56273 ;
  assign n56652 = n83502 & n56651 ;
  assign n56653 = n56277 | n56652 ;
  assign n83503 = ~n55756 ;
  assign n55760 = n83503 & n55759 ;
  assign n56278 = n55411 | n55759 ;
  assign n83504 = ~n56278 ;
  assign n56279 = n55988 & n83504 ;
  assign n56280 = n55760 | n56279 ;
  assign n56281 = n83422 & n56280 ;
  assign n56282 = n55401 & n83418 ;
  assign n56283 = n56062 & n56282 ;
  assign n56284 = n56281 | n56283 ;
  assign n56285 = n67622 & n56284 ;
  assign n83505 = ~n55987 ;
  assign n55989 = n55754 & n83505 ;
  assign n56286 = n55420 | n55754 ;
  assign n83506 = ~n56286 ;
  assign n56287 = n55750 & n83506 ;
  assign n56288 = n55989 | n56287 ;
  assign n56289 = n83422 & n56288 ;
  assign n56290 = n55410 & n83418 ;
  assign n56291 = n56062 & n56290 ;
  assign n56292 = n56289 | n56291 ;
  assign n56293 = n67531 & n56292 ;
  assign n83507 = ~n56291 ;
  assign n56639 = x90 & n83507 ;
  assign n83508 = ~n56289 ;
  assign n56640 = n83508 & n56639 ;
  assign n56641 = n56293 | n56640 ;
  assign n83509 = ~n55745 ;
  assign n55749 = n83509 & n55748 ;
  assign n56294 = n55429 | n55748 ;
  assign n83510 = ~n56294 ;
  assign n56295 = n55983 & n83510 ;
  assign n56296 = n55749 | n56295 ;
  assign n56297 = n83422 & n56296 ;
  assign n56298 = n55419 & n83418 ;
  assign n56299 = n56062 & n56298 ;
  assign n56300 = n56297 | n56299 ;
  assign n56301 = n67348 & n56300 ;
  assign n83511 = ~n55982 ;
  assign n55984 = n55743 & n83511 ;
  assign n56302 = n55438 | n55743 ;
  assign n83512 = ~n56302 ;
  assign n56303 = n55739 & n83512 ;
  assign n56304 = n55984 | n56303 ;
  assign n56305 = n83422 & n56304 ;
  assign n56306 = n55428 & n83418 ;
  assign n56307 = n56062 & n56306 ;
  assign n56308 = n56305 | n56307 ;
  assign n56309 = n67222 & n56308 ;
  assign n83513 = ~n56307 ;
  assign n56627 = x88 & n83513 ;
  assign n83514 = ~n56305 ;
  assign n56628 = n83514 & n56627 ;
  assign n56629 = n56309 | n56628 ;
  assign n83515 = ~n55734 ;
  assign n55738 = n83515 & n55737 ;
  assign n56310 = n55446 | n55737 ;
  assign n83516 = ~n56310 ;
  assign n56311 = n55978 & n83516 ;
  assign n56312 = n55738 | n56311 ;
  assign n56313 = n83422 & n56312 ;
  assign n56314 = n55437 & n83418 ;
  assign n56315 = n56062 & n56314 ;
  assign n56316 = n56313 | n56315 ;
  assign n56317 = n67164 & n56316 ;
  assign n83517 = ~n55977 ;
  assign n55979 = n55732 & n83517 ;
  assign n56318 = n55455 | n55732 ;
  assign n83518 = ~n56318 ;
  assign n56319 = n55728 & n83518 ;
  assign n56320 = n55979 | n56319 ;
  assign n56321 = n83422 & n56320 ;
  assign n56322 = n55445 & n83418 ;
  assign n56323 = n56062 & n56322 ;
  assign n56324 = n56321 | n56323 ;
  assign n56325 = n66979 & n56324 ;
  assign n83519 = ~n56323 ;
  assign n56615 = x86 & n83519 ;
  assign n83520 = ~n56321 ;
  assign n56616 = n83520 & n56615 ;
  assign n56617 = n56325 | n56616 ;
  assign n83521 = ~n55723 ;
  assign n55727 = n83521 & n55726 ;
  assign n56326 = n55463 | n55726 ;
  assign n83522 = ~n56326 ;
  assign n56327 = n55973 & n83522 ;
  assign n56328 = n55727 | n56327 ;
  assign n56329 = n83422 & n56328 ;
  assign n56330 = n55454 & n83418 ;
  assign n56331 = n56062 & n56330 ;
  assign n56332 = n56329 | n56331 ;
  assign n56333 = n66868 & n56332 ;
  assign n83523 = ~n55972 ;
  assign n55974 = n55721 & n83523 ;
  assign n56334 = n55471 | n55721 ;
  assign n83524 = ~n56334 ;
  assign n56335 = n55717 & n83524 ;
  assign n56336 = n55974 | n56335 ;
  assign n56337 = n83422 & n56336 ;
  assign n56338 = n55462 & n83418 ;
  assign n56339 = n56062 & n56338 ;
  assign n56340 = n56337 | n56339 ;
  assign n56341 = n66797 & n56340 ;
  assign n83525 = ~n56339 ;
  assign n56603 = x84 & n83525 ;
  assign n83526 = ~n56337 ;
  assign n56604 = n83526 & n56603 ;
  assign n56605 = n56341 | n56604 ;
  assign n83527 = ~n55712 ;
  assign n55716 = n83527 & n55715 ;
  assign n56342 = n55480 | n55715 ;
  assign n83528 = ~n56342 ;
  assign n56343 = n55968 & n83528 ;
  assign n56344 = n55716 | n56343 ;
  assign n56345 = n83422 & n56344 ;
  assign n56346 = n55470 & n83418 ;
  assign n56347 = n56062 & n56346 ;
  assign n56348 = n56345 | n56347 ;
  assign n56349 = n66654 & n56348 ;
  assign n83529 = ~n55967 ;
  assign n55969 = n55710 & n83529 ;
  assign n56350 = n55489 | n55710 ;
  assign n83530 = ~n56350 ;
  assign n56351 = n55706 & n83530 ;
  assign n56352 = n55969 | n56351 ;
  assign n56353 = n83422 & n56352 ;
  assign n56354 = n55479 & n83418 ;
  assign n56355 = n56062 & n56354 ;
  assign n56356 = n56353 | n56355 ;
  assign n56357 = n66560 & n56356 ;
  assign n83531 = ~n56355 ;
  assign n56591 = x82 & n83531 ;
  assign n83532 = ~n56353 ;
  assign n56592 = n83532 & n56591 ;
  assign n56593 = n56357 | n56592 ;
  assign n83533 = ~n55701 ;
  assign n55705 = n83533 & n55704 ;
  assign n56358 = n55497 | n55704 ;
  assign n83534 = ~n56358 ;
  assign n56359 = n55963 & n83534 ;
  assign n56360 = n55705 | n56359 ;
  assign n56361 = n83422 & n56360 ;
  assign n56362 = n55488 & n83418 ;
  assign n56363 = n56062 & n56362 ;
  assign n56364 = n56361 | n56363 ;
  assign n56365 = n66505 & n56364 ;
  assign n83535 = ~n55962 ;
  assign n55964 = n55699 & n83535 ;
  assign n56366 = n55505 | n55699 ;
  assign n83536 = ~n56366 ;
  assign n56367 = n55695 & n83536 ;
  assign n56368 = n55964 | n56367 ;
  assign n56369 = n83422 & n56368 ;
  assign n56370 = n55496 & n83418 ;
  assign n56371 = n56062 & n56370 ;
  assign n56372 = n56369 | n56371 ;
  assign n56373 = n66379 & n56372 ;
  assign n83537 = ~n56371 ;
  assign n56579 = x80 & n83537 ;
  assign n83538 = ~n56369 ;
  assign n56580 = n83538 & n56579 ;
  assign n56581 = n56373 | n56580 ;
  assign n83539 = ~n55690 ;
  assign n55694 = n83539 & n55693 ;
  assign n56374 = n55514 | n55693 ;
  assign n83540 = ~n56374 ;
  assign n56375 = n55958 & n83540 ;
  assign n56376 = n55694 | n56375 ;
  assign n56377 = n83422 & n56376 ;
  assign n56378 = n55504 & n83418 ;
  assign n56379 = n56062 & n56378 ;
  assign n56380 = n56377 | n56379 ;
  assign n56381 = n66299 & n56380 ;
  assign n83541 = ~n55957 ;
  assign n55959 = n55688 & n83541 ;
  assign n56382 = n55523 | n55688 ;
  assign n83542 = ~n56382 ;
  assign n56383 = n55684 & n83542 ;
  assign n56384 = n55959 | n56383 ;
  assign n56385 = n83422 & n56384 ;
  assign n56386 = n55513 & n83418 ;
  assign n56387 = n56062 & n56386 ;
  assign n56388 = n56385 | n56387 ;
  assign n56389 = n66244 & n56388 ;
  assign n83543 = ~n56387 ;
  assign n56567 = x78 & n83543 ;
  assign n83544 = ~n56385 ;
  assign n56568 = n83544 & n56567 ;
  assign n56569 = n56389 | n56568 ;
  assign n83545 = ~n55679 ;
  assign n55683 = n83545 & n55682 ;
  assign n56390 = n55531 | n55682 ;
  assign n83546 = ~n56390 ;
  assign n56391 = n55953 & n83546 ;
  assign n56392 = n55683 | n56391 ;
  assign n56393 = n83422 & n56392 ;
  assign n56394 = n55522 & n83418 ;
  assign n56395 = n56062 & n56394 ;
  assign n56396 = n56393 | n56395 ;
  assign n56397 = n66145 & n56396 ;
  assign n83547 = ~n55952 ;
  assign n55954 = n55677 & n83547 ;
  assign n56398 = n55539 | n55677 ;
  assign n83548 = ~n56398 ;
  assign n56399 = n55673 & n83548 ;
  assign n56400 = n55954 | n56399 ;
  assign n56401 = n83422 & n56400 ;
  assign n56402 = n55530 & n83418 ;
  assign n56403 = n56062 & n56402 ;
  assign n56404 = n56401 | n56403 ;
  assign n56405 = n66081 & n56404 ;
  assign n83549 = ~n56403 ;
  assign n56555 = x76 & n83549 ;
  assign n83550 = ~n56401 ;
  assign n56556 = n83550 & n56555 ;
  assign n56557 = n56405 | n56556 ;
  assign n83551 = ~n55668 ;
  assign n55672 = n83551 & n55671 ;
  assign n56406 = n55548 | n55671 ;
  assign n83552 = ~n56406 ;
  assign n56407 = n55948 & n83552 ;
  assign n56408 = n55672 | n56407 ;
  assign n56409 = n83422 & n56408 ;
  assign n56410 = n55538 & n83418 ;
  assign n56411 = n56062 & n56410 ;
  assign n56412 = n56409 | n56411 ;
  assign n56413 = n66043 & n56412 ;
  assign n83553 = ~n55947 ;
  assign n55949 = n55666 & n83553 ;
  assign n56414 = n55557 | n55666 ;
  assign n83554 = ~n56414 ;
  assign n56415 = n55662 & n83554 ;
  assign n56416 = n55949 | n56415 ;
  assign n56417 = n83422 & n56416 ;
  assign n56418 = n55547 & n83418 ;
  assign n56419 = n56062 & n56418 ;
  assign n56420 = n56417 | n56419 ;
  assign n56421 = n65960 & n56420 ;
  assign n83555 = ~n56419 ;
  assign n56543 = x74 & n83555 ;
  assign n83556 = ~n56417 ;
  assign n56544 = n83556 & n56543 ;
  assign n56545 = n56421 | n56544 ;
  assign n83557 = ~n55657 ;
  assign n55661 = n83557 & n55660 ;
  assign n56422 = n55565 | n55660 ;
  assign n83558 = ~n56422 ;
  assign n56423 = n55943 & n83558 ;
  assign n56424 = n55661 | n56423 ;
  assign n56425 = n83422 & n56424 ;
  assign n56426 = n55556 & n83418 ;
  assign n56427 = n56062 & n56426 ;
  assign n56428 = n56425 | n56427 ;
  assign n56429 = n65909 & n56428 ;
  assign n83559 = ~n55942 ;
  assign n55944 = n55655 & n83559 ;
  assign n56430 = n55574 | n55655 ;
  assign n83560 = ~n56430 ;
  assign n56431 = n55651 & n83560 ;
  assign n56432 = n55944 | n56431 ;
  assign n56433 = n83422 & n56432 ;
  assign n56434 = n55564 & n83418 ;
  assign n56435 = n56062 & n56434 ;
  assign n56436 = n56433 | n56435 ;
  assign n56437 = n65877 & n56436 ;
  assign n83561 = ~n56435 ;
  assign n56531 = x72 & n83561 ;
  assign n83562 = ~n56433 ;
  assign n56532 = n83562 & n56531 ;
  assign n56533 = n56437 | n56532 ;
  assign n83563 = ~n55646 ;
  assign n55650 = n83563 & n55649 ;
  assign n56438 = n55583 | n55649 ;
  assign n83564 = ~n56438 ;
  assign n56439 = n55938 & n83564 ;
  assign n56440 = n55650 | n56439 ;
  assign n56441 = n83422 & n56440 ;
  assign n56442 = n55573 & n83418 ;
  assign n56443 = n56062 & n56442 ;
  assign n56444 = n56441 | n56443 ;
  assign n56445 = n65820 & n56444 ;
  assign n83565 = ~n55937 ;
  assign n55939 = n55644 & n83565 ;
  assign n56446 = n55592 | n55644 ;
  assign n83566 = ~n56446 ;
  assign n56447 = n55640 & n83566 ;
  assign n56448 = n55939 | n56447 ;
  assign n56449 = n83422 & n56448 ;
  assign n56450 = n55582 & n83418 ;
  assign n56451 = n56062 & n56450 ;
  assign n56452 = n56449 | n56451 ;
  assign n56453 = n65791 & n56452 ;
  assign n83567 = ~n56451 ;
  assign n56519 = x70 & n83567 ;
  assign n83568 = ~n56449 ;
  assign n56520 = n83568 & n56519 ;
  assign n56521 = n56453 | n56520 ;
  assign n83569 = ~n55636 ;
  assign n55935 = n83569 & n55639 ;
  assign n56454 = n55601 | n55639 ;
  assign n83570 = ~n56454 ;
  assign n56455 = n55933 & n83570 ;
  assign n56456 = n55935 | n56455 ;
  assign n56457 = n83422 & n56456 ;
  assign n56458 = n55591 & n83418 ;
  assign n56459 = n56062 & n56458 ;
  assign n56460 = n56457 | n56459 ;
  assign n56461 = n65772 & n56460 ;
  assign n83571 = ~n55931 ;
  assign n55932 = n55634 & n83571 ;
  assign n56462 = n55609 | n55634 ;
  assign n83572 = ~n56462 ;
  assign n56463 = n55930 & n83572 ;
  assign n56464 = n55932 | n56463 ;
  assign n56465 = n83422 & n56464 ;
  assign n56466 = n55600 & n83418 ;
  assign n56467 = n56062 & n56466 ;
  assign n56468 = n56465 | n56467 ;
  assign n56469 = n65746 & n56468 ;
  assign n83573 = ~n56467 ;
  assign n56508 = x68 & n83573 ;
  assign n83574 = ~n56465 ;
  assign n56509 = n83574 & n56508 ;
  assign n56510 = n56469 | n56509 ;
  assign n83575 = ~n55929 ;
  assign n56471 = n55629 & n83575 ;
  assign n56470 = n55624 | n55629 ;
  assign n83576 = ~n56470 ;
  assign n56472 = n55625 & n83576 ;
  assign n56473 = n56471 | n56472 ;
  assign n56474 = n83422 & n56473 ;
  assign n56475 = n55608 & n83418 ;
  assign n56476 = n56062 & n56475 ;
  assign n56477 = n56474 | n56476 ;
  assign n56478 = n65721 & n56477 ;
  assign n56479 = n23402 & n55622 ;
  assign n56480 = n83420 & n56479 ;
  assign n83577 = ~n56480 ;
  assign n56481 = n55625 & n83577 ;
  assign n56482 = n83422 & n56481 ;
  assign n56483 = n55612 & n83418 ;
  assign n56484 = n56062 & n56483 ;
  assign n56485 = n56482 | n56484 ;
  assign n56486 = n65686 & n56485 ;
  assign n83578 = ~n56484 ;
  assign n56498 = x66 & n83578 ;
  assign n83579 = ~n56482 ;
  assign n56499 = n83579 & n56498 ;
  assign n56500 = n56486 | n56499 ;
  assign n55924 = n23402 & n83422 ;
  assign n55925 = x64 & n83422 ;
  assign n83580 = ~n55925 ;
  assign n56487 = x10 & n83580 ;
  assign n56488 = n55924 | n56487 ;
  assign n56489 = x65 & n56488 ;
  assign n56490 = n83418 & n56062 ;
  assign n83581 = ~n56490 ;
  assign n56491 = n23402 & n83581 ;
  assign n56492 = x65 | n56491 ;
  assign n56493 = n56487 | n56492 ;
  assign n83582 = ~n56489 ;
  assign n56494 = n83582 & n56493 ;
  assign n56496 = n24281 | n56494 ;
  assign n56497 = n65670 & n56488 ;
  assign n83583 = ~n56497 ;
  assign n56501 = n56496 & n83583 ;
  assign n56502 = n56500 | n56501 ;
  assign n83584 = ~n56486 ;
  assign n56503 = n83584 & n56502 ;
  assign n83585 = ~n56476 ;
  assign n56504 = x67 & n83585 ;
  assign n83586 = ~n56474 ;
  assign n56505 = n83586 & n56504 ;
  assign n56506 = n56478 | n56505 ;
  assign n56507 = n56503 | n56506 ;
  assign n83587 = ~n56478 ;
  assign n56511 = n83587 & n56507 ;
  assign n56512 = n56510 | n56511 ;
  assign n83588 = ~n56469 ;
  assign n56513 = n83588 & n56512 ;
  assign n83589 = ~n56459 ;
  assign n56514 = x69 & n83589 ;
  assign n83590 = ~n56457 ;
  assign n56515 = n83590 & n56514 ;
  assign n56516 = n56461 | n56515 ;
  assign n56518 = n56513 | n56516 ;
  assign n83591 = ~n56461 ;
  assign n56523 = n83591 & n56518 ;
  assign n56524 = n56521 | n56523 ;
  assign n83592 = ~n56453 ;
  assign n56525 = n83592 & n56524 ;
  assign n83593 = ~n56443 ;
  assign n56526 = x71 & n83593 ;
  assign n83594 = ~n56441 ;
  assign n56527 = n83594 & n56526 ;
  assign n56528 = n56445 | n56527 ;
  assign n56530 = n56525 | n56528 ;
  assign n83595 = ~n56445 ;
  assign n56535 = n83595 & n56530 ;
  assign n56536 = n56533 | n56535 ;
  assign n83596 = ~n56437 ;
  assign n56537 = n83596 & n56536 ;
  assign n83597 = ~n56427 ;
  assign n56538 = x73 & n83597 ;
  assign n83598 = ~n56425 ;
  assign n56539 = n83598 & n56538 ;
  assign n56540 = n56429 | n56539 ;
  assign n56542 = n56537 | n56540 ;
  assign n83599 = ~n56429 ;
  assign n56547 = n83599 & n56542 ;
  assign n56548 = n56545 | n56547 ;
  assign n83600 = ~n56421 ;
  assign n56549 = n83600 & n56548 ;
  assign n83601 = ~n56411 ;
  assign n56550 = x75 & n83601 ;
  assign n83602 = ~n56409 ;
  assign n56551 = n83602 & n56550 ;
  assign n56552 = n56413 | n56551 ;
  assign n56554 = n56549 | n56552 ;
  assign n83603 = ~n56413 ;
  assign n56559 = n83603 & n56554 ;
  assign n56560 = n56557 | n56559 ;
  assign n83604 = ~n56405 ;
  assign n56561 = n83604 & n56560 ;
  assign n83605 = ~n56395 ;
  assign n56562 = x77 & n83605 ;
  assign n83606 = ~n56393 ;
  assign n56563 = n83606 & n56562 ;
  assign n56564 = n56397 | n56563 ;
  assign n56566 = n56561 | n56564 ;
  assign n83607 = ~n56397 ;
  assign n56571 = n83607 & n56566 ;
  assign n56572 = n56569 | n56571 ;
  assign n83608 = ~n56389 ;
  assign n56573 = n83608 & n56572 ;
  assign n83609 = ~n56379 ;
  assign n56574 = x79 & n83609 ;
  assign n83610 = ~n56377 ;
  assign n56575 = n83610 & n56574 ;
  assign n56576 = n56381 | n56575 ;
  assign n56578 = n56573 | n56576 ;
  assign n83611 = ~n56381 ;
  assign n56583 = n83611 & n56578 ;
  assign n56584 = n56581 | n56583 ;
  assign n83612 = ~n56373 ;
  assign n56585 = n83612 & n56584 ;
  assign n83613 = ~n56363 ;
  assign n56586 = x81 & n83613 ;
  assign n83614 = ~n56361 ;
  assign n56587 = n83614 & n56586 ;
  assign n56588 = n56365 | n56587 ;
  assign n56590 = n56585 | n56588 ;
  assign n83615 = ~n56365 ;
  assign n56595 = n83615 & n56590 ;
  assign n56596 = n56593 | n56595 ;
  assign n83616 = ~n56357 ;
  assign n56597 = n83616 & n56596 ;
  assign n83617 = ~n56347 ;
  assign n56598 = x83 & n83617 ;
  assign n83618 = ~n56345 ;
  assign n56599 = n83618 & n56598 ;
  assign n56600 = n56349 | n56599 ;
  assign n56602 = n56597 | n56600 ;
  assign n83619 = ~n56349 ;
  assign n56607 = n83619 & n56602 ;
  assign n56608 = n56605 | n56607 ;
  assign n83620 = ~n56341 ;
  assign n56609 = n83620 & n56608 ;
  assign n83621 = ~n56331 ;
  assign n56610 = x85 & n83621 ;
  assign n83622 = ~n56329 ;
  assign n56611 = n83622 & n56610 ;
  assign n56612 = n56333 | n56611 ;
  assign n56614 = n56609 | n56612 ;
  assign n83623 = ~n56333 ;
  assign n56619 = n83623 & n56614 ;
  assign n56620 = n56617 | n56619 ;
  assign n83624 = ~n56325 ;
  assign n56621 = n83624 & n56620 ;
  assign n83625 = ~n56315 ;
  assign n56622 = x87 & n83625 ;
  assign n83626 = ~n56313 ;
  assign n56623 = n83626 & n56622 ;
  assign n56624 = n56317 | n56623 ;
  assign n56626 = n56621 | n56624 ;
  assign n83627 = ~n56317 ;
  assign n56631 = n83627 & n56626 ;
  assign n56632 = n56629 | n56631 ;
  assign n83628 = ~n56309 ;
  assign n56633 = n83628 & n56632 ;
  assign n83629 = ~n56299 ;
  assign n56634 = x89 & n83629 ;
  assign n83630 = ~n56297 ;
  assign n56635 = n83630 & n56634 ;
  assign n56636 = n56301 | n56635 ;
  assign n56638 = n56633 | n56636 ;
  assign n83631 = ~n56301 ;
  assign n56643 = n83631 & n56638 ;
  assign n56644 = n56641 | n56643 ;
  assign n83632 = ~n56293 ;
  assign n56645 = n83632 & n56644 ;
  assign n83633 = ~n56283 ;
  assign n56646 = x91 & n83633 ;
  assign n83634 = ~n56281 ;
  assign n56647 = n83634 & n56646 ;
  assign n56648 = n56285 | n56647 ;
  assign n56650 = n56645 | n56648 ;
  assign n83635 = ~n56285 ;
  assign n56655 = n83635 & n56650 ;
  assign n56656 = n56653 | n56655 ;
  assign n83636 = ~n56277 ;
  assign n56657 = n83636 & n56656 ;
  assign n83637 = ~n56267 ;
  assign n56658 = x93 & n83637 ;
  assign n83638 = ~n56265 ;
  assign n56659 = n83638 & n56658 ;
  assign n56660 = n56269 | n56659 ;
  assign n56662 = n56657 | n56660 ;
  assign n83639 = ~n56269 ;
  assign n56667 = n83639 & n56662 ;
  assign n56668 = n56665 | n56667 ;
  assign n83640 = ~n56261 ;
  assign n56669 = n83640 & n56668 ;
  assign n83641 = ~n56251 ;
  assign n56670 = x95 & n83641 ;
  assign n83642 = ~n56249 ;
  assign n56671 = n83642 & n56670 ;
  assign n56672 = n56253 | n56671 ;
  assign n56674 = n56669 | n56672 ;
  assign n83643 = ~n56253 ;
  assign n56679 = n83643 & n56674 ;
  assign n56680 = n56677 | n56679 ;
  assign n83644 = ~n56245 ;
  assign n56681 = n83644 & n56680 ;
  assign n83645 = ~n56235 ;
  assign n56682 = x97 & n83645 ;
  assign n83646 = ~n56233 ;
  assign n56683 = n83646 & n56682 ;
  assign n56684 = n56237 | n56683 ;
  assign n56686 = n56681 | n56684 ;
  assign n83647 = ~n56237 ;
  assign n56691 = n83647 & n56686 ;
  assign n56692 = n56689 | n56691 ;
  assign n83648 = ~n56229 ;
  assign n56693 = n83648 & n56692 ;
  assign n83649 = ~n56219 ;
  assign n56694 = x99 & n83649 ;
  assign n83650 = ~n56217 ;
  assign n56695 = n83650 & n56694 ;
  assign n56696 = n56221 | n56695 ;
  assign n56698 = n56693 | n56696 ;
  assign n83651 = ~n56221 ;
  assign n56703 = n83651 & n56698 ;
  assign n56704 = n56701 | n56703 ;
  assign n83652 = ~n56213 ;
  assign n56705 = n83652 & n56704 ;
  assign n83653 = ~n56203 ;
  assign n56706 = x101 & n83653 ;
  assign n83654 = ~n56201 ;
  assign n56707 = n83654 & n56706 ;
  assign n56708 = n56205 | n56707 ;
  assign n56710 = n56705 | n56708 ;
  assign n83655 = ~n56205 ;
  assign n56715 = n83655 & n56710 ;
  assign n56716 = n56713 | n56715 ;
  assign n83656 = ~n56197 ;
  assign n56717 = n83656 & n56716 ;
  assign n83657 = ~n56187 ;
  assign n56718 = x103 & n83657 ;
  assign n83658 = ~n56185 ;
  assign n56719 = n83658 & n56718 ;
  assign n56720 = n56189 | n56719 ;
  assign n56722 = n56717 | n56720 ;
  assign n83659 = ~n56189 ;
  assign n56727 = n83659 & n56722 ;
  assign n56728 = n56725 | n56727 ;
  assign n83660 = ~n56181 ;
  assign n56729 = n83660 & n56728 ;
  assign n83661 = ~n56171 ;
  assign n56730 = x105 & n83661 ;
  assign n83662 = ~n56169 ;
  assign n56731 = n83662 & n56730 ;
  assign n56732 = n56173 | n56731 ;
  assign n56734 = n56729 | n56732 ;
  assign n83663 = ~n56173 ;
  assign n56739 = n83663 & n56734 ;
  assign n56740 = n56737 | n56739 ;
  assign n83664 = ~n56165 ;
  assign n56741 = n83664 & n56740 ;
  assign n83665 = ~n56155 ;
  assign n56742 = x107 & n83665 ;
  assign n83666 = ~n56153 ;
  assign n56743 = n83666 & n56742 ;
  assign n56744 = n56157 | n56743 ;
  assign n56746 = n56741 | n56744 ;
  assign n83667 = ~n56157 ;
  assign n56751 = n83667 & n56746 ;
  assign n56752 = n56749 | n56751 ;
  assign n83668 = ~n56149 ;
  assign n56753 = n83668 & n56752 ;
  assign n83669 = ~n56139 ;
  assign n56754 = x109 & n83669 ;
  assign n83670 = ~n56137 ;
  assign n56755 = n83670 & n56754 ;
  assign n56756 = n56141 | n56755 ;
  assign n56758 = n56753 | n56756 ;
  assign n83671 = ~n56141 ;
  assign n56763 = n83671 & n56758 ;
  assign n56764 = n56761 | n56763 ;
  assign n83672 = ~n56133 ;
  assign n56765 = n83672 & n56764 ;
  assign n83673 = ~n56123 ;
  assign n56766 = x111 & n83673 ;
  assign n83674 = ~n56121 ;
  assign n56767 = n83674 & n56766 ;
  assign n56768 = n56125 | n56767 ;
  assign n56770 = n56765 | n56768 ;
  assign n83675 = ~n56125 ;
  assign n56775 = n83675 & n56770 ;
  assign n56776 = n56773 | n56775 ;
  assign n83676 = ~n56117 ;
  assign n56777 = n83676 & n56776 ;
  assign n83677 = ~n56107 ;
  assign n56778 = x113 & n83677 ;
  assign n83678 = ~n56105 ;
  assign n56779 = n83678 & n56778 ;
  assign n56780 = n56109 | n56779 ;
  assign n56782 = n56777 | n56780 ;
  assign n83679 = ~n56109 ;
  assign n56787 = n83679 & n56782 ;
  assign n56788 = n56785 | n56787 ;
  assign n83680 = ~n56101 ;
  assign n56789 = n83680 & n56788 ;
  assign n83681 = ~n56091 ;
  assign n56790 = x115 & n83681 ;
  assign n83682 = ~n56089 ;
  assign n56791 = n83682 & n56790 ;
  assign n56792 = n56093 | n56791 ;
  assign n56794 = n56789 | n56792 ;
  assign n83683 = ~n56093 ;
  assign n56799 = n83683 & n56794 ;
  assign n56800 = n56797 | n56799 ;
  assign n83684 = ~n56085 ;
  assign n56801 = n83684 & n56800 ;
  assign n83685 = ~n56064 ;
  assign n56802 = x117 & n83685 ;
  assign n83686 = ~n56058 ;
  assign n56803 = n83686 & n56802 ;
  assign n56804 = n56077 | n56803 ;
  assign n56806 = n56801 | n56804 ;
  assign n83687 = ~n56077 ;
  assign n56810 = n83687 & n56806 ;
  assign n56811 = n56809 | n56810 ;
  assign n83688 = ~n56076 ;
  assign n56812 = n83688 & n56811 ;
  assign n56813 = n24576 | n56812 ;
  assign n83689 = ~n56075 ;
  assign n56814 = n83689 & n56813 ;
  assign n83690 = ~n56810 ;
  assign n57657 = n56809 & n83690 ;
  assign n56817 = x64 & n83581 ;
  assign n83691 = ~n56817 ;
  assign n56818 = x10 & n83691 ;
  assign n56819 = n55924 | n56818 ;
  assign n56820 = x65 & n56819 ;
  assign n83692 = ~n56820 ;
  assign n56821 = n56493 & n83692 ;
  assign n56822 = n24281 | n56821 ;
  assign n56823 = n83583 & n56822 ;
  assign n56825 = n56500 | n56823 ;
  assign n56826 = n83584 & n56825 ;
  assign n56827 = n56506 | n56826 ;
  assign n56828 = n83587 & n56827 ;
  assign n56829 = n56510 | n56828 ;
  assign n56830 = n83588 & n56829 ;
  assign n56831 = n56516 | n56830 ;
  assign n56832 = n83591 & n56831 ;
  assign n56833 = n56521 | n56832 ;
  assign n56834 = n83592 & n56833 ;
  assign n56835 = n56528 | n56834 ;
  assign n56836 = n83595 & n56835 ;
  assign n56837 = n56533 | n56836 ;
  assign n56838 = n83596 & n56837 ;
  assign n56839 = n56540 | n56838 ;
  assign n56840 = n83599 & n56839 ;
  assign n56841 = n56545 | n56840 ;
  assign n56842 = n83600 & n56841 ;
  assign n56843 = n56552 | n56842 ;
  assign n56844 = n83603 & n56843 ;
  assign n56845 = n56557 | n56844 ;
  assign n56846 = n83604 & n56845 ;
  assign n56847 = n56564 | n56846 ;
  assign n56848 = n83607 & n56847 ;
  assign n56849 = n56569 | n56848 ;
  assign n56850 = n83608 & n56849 ;
  assign n56851 = n56576 | n56850 ;
  assign n56852 = n83611 & n56851 ;
  assign n56853 = n56581 | n56852 ;
  assign n56854 = n83612 & n56853 ;
  assign n56855 = n56588 | n56854 ;
  assign n56856 = n83615 & n56855 ;
  assign n56857 = n56593 | n56856 ;
  assign n56858 = n83616 & n56857 ;
  assign n56859 = n56600 | n56858 ;
  assign n56860 = n83619 & n56859 ;
  assign n56861 = n56605 | n56860 ;
  assign n56862 = n83620 & n56861 ;
  assign n56863 = n56612 | n56862 ;
  assign n56864 = n83623 & n56863 ;
  assign n56865 = n56617 | n56864 ;
  assign n56866 = n83624 & n56865 ;
  assign n56867 = n56624 | n56866 ;
  assign n56868 = n83627 & n56867 ;
  assign n56869 = n56629 | n56868 ;
  assign n56870 = n83628 & n56869 ;
  assign n56871 = n56636 | n56870 ;
  assign n56872 = n83631 & n56871 ;
  assign n56873 = n56641 | n56872 ;
  assign n56874 = n83632 & n56873 ;
  assign n56875 = n56648 | n56874 ;
  assign n56876 = n83635 & n56875 ;
  assign n56877 = n56653 | n56876 ;
  assign n56878 = n83636 & n56877 ;
  assign n56879 = n56660 | n56878 ;
  assign n56880 = n83639 & n56879 ;
  assign n56881 = n56665 | n56880 ;
  assign n56882 = n83640 & n56881 ;
  assign n56883 = n56672 | n56882 ;
  assign n56884 = n83643 & n56883 ;
  assign n56885 = n56677 | n56884 ;
  assign n56886 = n83644 & n56885 ;
  assign n56887 = n56684 | n56886 ;
  assign n56888 = n83647 & n56887 ;
  assign n56889 = n56689 | n56888 ;
  assign n56890 = n83648 & n56889 ;
  assign n56891 = n56696 | n56890 ;
  assign n56892 = n83651 & n56891 ;
  assign n56893 = n56701 | n56892 ;
  assign n56894 = n83652 & n56893 ;
  assign n56895 = n56708 | n56894 ;
  assign n56896 = n83655 & n56895 ;
  assign n56897 = n56713 | n56896 ;
  assign n56898 = n83656 & n56897 ;
  assign n56899 = n56720 | n56898 ;
  assign n56900 = n83659 & n56899 ;
  assign n56901 = n56725 | n56900 ;
  assign n56902 = n83660 & n56901 ;
  assign n56903 = n56732 | n56902 ;
  assign n56904 = n83663 & n56903 ;
  assign n56905 = n56737 | n56904 ;
  assign n56906 = n83664 & n56905 ;
  assign n56907 = n56744 | n56906 ;
  assign n56908 = n83667 & n56907 ;
  assign n56909 = n56749 | n56908 ;
  assign n56910 = n83668 & n56909 ;
  assign n56911 = n56756 | n56910 ;
  assign n56912 = n83671 & n56911 ;
  assign n56913 = n56761 | n56912 ;
  assign n56914 = n83672 & n56913 ;
  assign n56915 = n56768 | n56914 ;
  assign n56916 = n83675 & n56915 ;
  assign n56917 = n56773 | n56916 ;
  assign n56918 = n83676 & n56917 ;
  assign n56919 = n56780 | n56918 ;
  assign n56920 = n83679 & n56919 ;
  assign n56921 = n56785 | n56920 ;
  assign n56922 = n83680 & n56921 ;
  assign n56923 = n56792 | n56922 ;
  assign n56924 = n83683 & n56923 ;
  assign n56925 = n56797 | n56924 ;
  assign n56927 = n83684 & n56925 ;
  assign n57351 = n56804 | n56927 ;
  assign n57658 = n56077 | n56809 ;
  assign n83693 = ~n57658 ;
  assign n57659 = n57351 & n83693 ;
  assign n57660 = n57657 | n57659 ;
  assign n57661 = n56813 | n57660 ;
  assign n83694 = ~n56814 ;
  assign n57662 = n83694 & n57661 ;
  assign n57670 = n73458 & n57662 ;
  assign n56816 = n56065 & n56813 ;
  assign n56805 = n56085 | n56804 ;
  assign n83695 = ~n56805 ;
  assign n56926 = n83695 & n56925 ;
  assign n83696 = ~n56927 ;
  assign n56928 = n56804 & n83696 ;
  assign n56929 = n56926 | n56928 ;
  assign n56930 = n73458 & n56929 ;
  assign n83697 = ~n56812 ;
  assign n56931 = n83697 & n56930 ;
  assign n56932 = n56816 | n56931 ;
  assign n56933 = n73188 & n56932 ;
  assign n56934 = n56084 & n56813 ;
  assign n56798 = n56093 | n56797 ;
  assign n83698 = ~n56798 ;
  assign n56935 = n56794 & n83698 ;
  assign n83699 = ~n56799 ;
  assign n56936 = n56797 & n83699 ;
  assign n56937 = n56935 | n56936 ;
  assign n56938 = n73458 & n56937 ;
  assign n56939 = n83697 & n56938 ;
  assign n56940 = n56934 | n56939 ;
  assign n56941 = n73177 & n56940 ;
  assign n56942 = n56092 & n56813 ;
  assign n56793 = n56101 | n56792 ;
  assign n83700 = ~n56793 ;
  assign n56943 = n83700 & n56921 ;
  assign n83701 = ~n56922 ;
  assign n56944 = n56792 & n83701 ;
  assign n56945 = n56943 | n56944 ;
  assign n56946 = n73458 & n56945 ;
  assign n56947 = n83697 & n56946 ;
  assign n56948 = n56942 | n56947 ;
  assign n56949 = n72752 & n56948 ;
  assign n56950 = n56100 & n56813 ;
  assign n56786 = n56109 | n56785 ;
  assign n83702 = ~n56786 ;
  assign n56951 = n56782 & n83702 ;
  assign n83703 = ~n56787 ;
  assign n56952 = n56785 & n83703 ;
  assign n56953 = n56951 | n56952 ;
  assign n56954 = n73458 & n56953 ;
  assign n56955 = n83697 & n56954 ;
  assign n56956 = n56950 | n56955 ;
  assign n56957 = n72393 & n56956 ;
  assign n56958 = n56108 & n56813 ;
  assign n56781 = n56117 | n56780 ;
  assign n83704 = ~n56781 ;
  assign n56959 = n83704 & n56917 ;
  assign n83705 = ~n56918 ;
  assign n56960 = n56780 & n83705 ;
  assign n56961 = n56959 | n56960 ;
  assign n56962 = n73458 & n56961 ;
  assign n56963 = n83697 & n56962 ;
  assign n56964 = n56958 | n56963 ;
  assign n56965 = n72385 & n56964 ;
  assign n56966 = n56116 & n56813 ;
  assign n56774 = n56125 | n56773 ;
  assign n83706 = ~n56774 ;
  assign n56967 = n56770 & n83706 ;
  assign n83707 = ~n56775 ;
  assign n56968 = n56773 & n83707 ;
  assign n56969 = n56967 | n56968 ;
  assign n56970 = n73458 & n56969 ;
  assign n56971 = n83697 & n56970 ;
  assign n56972 = n56966 | n56971 ;
  assign n56973 = n72025 & n56972 ;
  assign n56974 = n56124 & n56813 ;
  assign n56769 = n56133 | n56768 ;
  assign n83708 = ~n56769 ;
  assign n56975 = n83708 & n56913 ;
  assign n83709 = ~n56914 ;
  assign n56976 = n56768 & n83709 ;
  assign n56977 = n56975 | n56976 ;
  assign n56978 = n73458 & n56977 ;
  assign n56979 = n83697 & n56978 ;
  assign n56980 = n56974 | n56979 ;
  assign n56981 = n71645 & n56980 ;
  assign n56982 = n56132 & n56813 ;
  assign n56762 = n56141 | n56761 ;
  assign n83710 = ~n56762 ;
  assign n56983 = n56758 & n83710 ;
  assign n83711 = ~n56763 ;
  assign n56984 = n56761 & n83711 ;
  assign n56985 = n56983 | n56984 ;
  assign n56986 = n73458 & n56985 ;
  assign n56987 = n83697 & n56986 ;
  assign n56988 = n56982 | n56987 ;
  assign n56989 = n71633 & n56988 ;
  assign n56990 = n56140 & n56813 ;
  assign n56757 = n56149 | n56756 ;
  assign n83712 = ~n56757 ;
  assign n56991 = n83712 & n56909 ;
  assign n83713 = ~n56910 ;
  assign n56992 = n56756 & n83713 ;
  assign n56993 = n56991 | n56992 ;
  assign n56994 = n73458 & n56993 ;
  assign n56995 = n83697 & n56994 ;
  assign n56996 = n56990 | n56995 ;
  assign n56997 = n71253 & n56996 ;
  assign n56998 = n56148 & n56813 ;
  assign n56750 = n56157 | n56749 ;
  assign n83714 = ~n56750 ;
  assign n56999 = n56746 & n83714 ;
  assign n83715 = ~n56751 ;
  assign n57000 = n56749 & n83715 ;
  assign n57001 = n56999 | n57000 ;
  assign n57002 = n73458 & n57001 ;
  assign n57003 = n83697 & n57002 ;
  assign n57004 = n56998 | n57003 ;
  assign n57005 = n70935 & n57004 ;
  assign n57006 = n56156 & n56813 ;
  assign n56745 = n56165 | n56744 ;
  assign n83716 = ~n56745 ;
  assign n57007 = n83716 & n56905 ;
  assign n83717 = ~n56906 ;
  assign n57008 = n56744 & n83717 ;
  assign n57009 = n57007 | n57008 ;
  assign n57010 = n73458 & n57009 ;
  assign n57011 = n83697 & n57010 ;
  assign n57012 = n57006 | n57011 ;
  assign n57013 = n70927 & n57012 ;
  assign n57014 = n56164 & n56813 ;
  assign n56738 = n56173 | n56737 ;
  assign n83718 = ~n56738 ;
  assign n57015 = n56734 & n83718 ;
  assign n83719 = ~n56739 ;
  assign n57016 = n56737 & n83719 ;
  assign n57017 = n57015 | n57016 ;
  assign n57018 = n73458 & n57017 ;
  assign n57019 = n83697 & n57018 ;
  assign n57020 = n57014 | n57019 ;
  assign n57021 = n70609 & n57020 ;
  assign n57022 = n56172 & n56813 ;
  assign n56733 = n56181 | n56732 ;
  assign n83720 = ~n56733 ;
  assign n57023 = n83720 & n56901 ;
  assign n83721 = ~n56902 ;
  assign n57024 = n56732 & n83721 ;
  assign n57025 = n57023 | n57024 ;
  assign n57026 = n73458 & n57025 ;
  assign n57027 = n83697 & n57026 ;
  assign n57028 = n57022 | n57027 ;
  assign n57029 = n70276 & n57028 ;
  assign n57030 = n56180 & n56813 ;
  assign n56726 = n56189 | n56725 ;
  assign n83722 = ~n56726 ;
  assign n57031 = n56722 & n83722 ;
  assign n83723 = ~n56727 ;
  assign n57032 = n56725 & n83723 ;
  assign n57033 = n57031 | n57032 ;
  assign n57034 = n73458 & n57033 ;
  assign n57035 = n83697 & n57034 ;
  assign n57036 = n57030 | n57035 ;
  assign n57037 = n70176 & n57036 ;
  assign n57038 = n56188 & n56813 ;
  assign n56721 = n56197 | n56720 ;
  assign n83724 = ~n56721 ;
  assign n57039 = n83724 & n56897 ;
  assign n83725 = ~n56898 ;
  assign n57040 = n56720 & n83725 ;
  assign n57041 = n57039 | n57040 ;
  assign n57042 = n73458 & n57041 ;
  assign n57043 = n83697 & n57042 ;
  assign n57044 = n57038 | n57043 ;
  assign n57045 = n69857 & n57044 ;
  assign n57046 = n56196 & n56813 ;
  assign n56714 = n56205 | n56713 ;
  assign n83726 = ~n56714 ;
  assign n57047 = n56710 & n83726 ;
  assign n83727 = ~n56715 ;
  assign n57048 = n56713 & n83727 ;
  assign n57049 = n57047 | n57048 ;
  assign n57050 = n73458 & n57049 ;
  assign n57051 = n83697 & n57050 ;
  assign n57052 = n57046 | n57051 ;
  assign n57053 = n69656 & n57052 ;
  assign n57054 = n56204 & n56813 ;
  assign n56709 = n56213 | n56708 ;
  assign n83728 = ~n56709 ;
  assign n57055 = n83728 & n56893 ;
  assign n83729 = ~n56894 ;
  assign n57056 = n56708 & n83729 ;
  assign n57057 = n57055 | n57056 ;
  assign n57058 = n73458 & n57057 ;
  assign n57059 = n83697 & n57058 ;
  assign n57060 = n57054 | n57059 ;
  assign n57061 = n69528 & n57060 ;
  assign n57062 = n56212 & n56813 ;
  assign n56702 = n56221 | n56701 ;
  assign n83730 = ~n56702 ;
  assign n57063 = n56698 & n83730 ;
  assign n83731 = ~n56703 ;
  assign n57064 = n56701 & n83731 ;
  assign n57065 = n57063 | n57064 ;
  assign n57066 = n73458 & n57065 ;
  assign n57067 = n83697 & n57066 ;
  assign n57068 = n57062 | n57067 ;
  assign n57069 = n69261 & n57068 ;
  assign n57070 = n56220 & n56813 ;
  assign n56697 = n56229 | n56696 ;
  assign n83732 = ~n56697 ;
  assign n57071 = n83732 & n56889 ;
  assign n83733 = ~n56890 ;
  assign n57072 = n56696 & n83733 ;
  assign n57073 = n57071 | n57072 ;
  assign n57074 = n73458 & n57073 ;
  assign n57075 = n83697 & n57074 ;
  assign n57076 = n57070 | n57075 ;
  assign n57077 = n69075 & n57076 ;
  assign n57078 = n56228 & n56813 ;
  assign n56690 = n56237 | n56689 ;
  assign n83734 = ~n56690 ;
  assign n57079 = n56686 & n83734 ;
  assign n83735 = ~n56691 ;
  assign n57080 = n56689 & n83735 ;
  assign n57081 = n57079 | n57080 ;
  assign n57082 = n73458 & n57081 ;
  assign n57083 = n83697 & n57082 ;
  assign n57084 = n57078 | n57083 ;
  assign n57085 = n68993 & n57084 ;
  assign n57086 = n56236 & n56813 ;
  assign n56685 = n56245 | n56684 ;
  assign n83736 = ~n56685 ;
  assign n57087 = n83736 & n56885 ;
  assign n83737 = ~n56886 ;
  assign n57088 = n56684 & n83737 ;
  assign n57089 = n57087 | n57088 ;
  assign n57090 = n73458 & n57089 ;
  assign n57091 = n83697 & n57090 ;
  assign n57092 = n57086 | n57091 ;
  assign n57093 = n68716 & n57092 ;
  assign n57094 = n56244 & n56813 ;
  assign n56678 = n56253 | n56677 ;
  assign n83738 = ~n56678 ;
  assign n57095 = n56674 & n83738 ;
  assign n83739 = ~n56679 ;
  assign n57096 = n56677 & n83739 ;
  assign n57097 = n57095 | n57096 ;
  assign n57098 = n73458 & n57097 ;
  assign n57099 = n83697 & n57098 ;
  assign n57100 = n57094 | n57099 ;
  assign n57101 = n68545 & n57100 ;
  assign n57102 = n56252 & n56813 ;
  assign n56673 = n56261 | n56672 ;
  assign n83740 = ~n56673 ;
  assign n57103 = n83740 & n56881 ;
  assign n83741 = ~n56882 ;
  assign n57104 = n56672 & n83741 ;
  assign n57105 = n57103 | n57104 ;
  assign n57106 = n73458 & n57105 ;
  assign n57107 = n83697 & n57106 ;
  assign n57108 = n57102 | n57107 ;
  assign n57109 = n68438 & n57108 ;
  assign n57110 = n56260 & n56813 ;
  assign n56666 = n56269 | n56665 ;
  assign n83742 = ~n56666 ;
  assign n57111 = n56662 & n83742 ;
  assign n83743 = ~n56667 ;
  assign n57112 = n56665 & n83743 ;
  assign n57113 = n57111 | n57112 ;
  assign n57114 = n73458 & n57113 ;
  assign n57115 = n83697 & n57114 ;
  assign n57116 = n57110 | n57115 ;
  assign n57117 = n68214 & n57116 ;
  assign n57118 = n56268 & n56813 ;
  assign n56661 = n56277 | n56660 ;
  assign n83744 = ~n56661 ;
  assign n57119 = n83744 & n56877 ;
  assign n83745 = ~n56878 ;
  assign n57120 = n56660 & n83745 ;
  assign n57121 = n57119 | n57120 ;
  assign n57122 = n73458 & n57121 ;
  assign n57123 = n83697 & n57122 ;
  assign n57124 = n57118 | n57123 ;
  assign n57125 = n68058 & n57124 ;
  assign n57126 = n56276 & n56813 ;
  assign n56654 = n56285 | n56653 ;
  assign n83746 = ~n56654 ;
  assign n57127 = n56650 & n83746 ;
  assign n83747 = ~n56655 ;
  assign n57128 = n56653 & n83747 ;
  assign n57129 = n57127 | n57128 ;
  assign n57130 = n73458 & n57129 ;
  assign n57131 = n83697 & n57130 ;
  assign n57132 = n57126 | n57131 ;
  assign n57133 = n67986 & n57132 ;
  assign n57134 = n56284 & n56813 ;
  assign n56649 = n56293 | n56648 ;
  assign n83748 = ~n56649 ;
  assign n57135 = n83748 & n56873 ;
  assign n83749 = ~n56874 ;
  assign n57136 = n56648 & n83749 ;
  assign n57137 = n57135 | n57136 ;
  assign n57138 = n73458 & n57137 ;
  assign n57139 = n83697 & n57138 ;
  assign n57140 = n57134 | n57139 ;
  assign n57141 = n67763 & n57140 ;
  assign n57142 = n56292 & n56813 ;
  assign n56642 = n56301 | n56641 ;
  assign n83750 = ~n56642 ;
  assign n57143 = n56638 & n83750 ;
  assign n83751 = ~n56643 ;
  assign n57144 = n56641 & n83751 ;
  assign n57145 = n57143 | n57144 ;
  assign n57146 = n73458 & n57145 ;
  assign n57147 = n83697 & n57146 ;
  assign n57148 = n57142 | n57147 ;
  assign n57149 = n67622 & n57148 ;
  assign n57150 = n56300 & n56813 ;
  assign n56637 = n56309 | n56636 ;
  assign n83752 = ~n56637 ;
  assign n57151 = n83752 & n56869 ;
  assign n83753 = ~n56870 ;
  assign n57152 = n56636 & n83753 ;
  assign n57153 = n57151 | n57152 ;
  assign n57154 = n73458 & n57153 ;
  assign n57155 = n83697 & n57154 ;
  assign n57156 = n57150 | n57155 ;
  assign n57157 = n67531 & n57156 ;
  assign n57158 = n56308 & n56813 ;
  assign n56630 = n56317 | n56629 ;
  assign n83754 = ~n56630 ;
  assign n57159 = n56626 & n83754 ;
  assign n83755 = ~n56631 ;
  assign n57160 = n56629 & n83755 ;
  assign n57161 = n57159 | n57160 ;
  assign n57162 = n73458 & n57161 ;
  assign n57163 = n83697 & n57162 ;
  assign n57164 = n57158 | n57163 ;
  assign n57165 = n67348 & n57164 ;
  assign n57166 = n56316 & n56813 ;
  assign n56625 = n56325 | n56624 ;
  assign n83756 = ~n56625 ;
  assign n57167 = n83756 & n56865 ;
  assign n83757 = ~n56866 ;
  assign n57168 = n56624 & n83757 ;
  assign n57169 = n57167 | n57168 ;
  assign n57170 = n73458 & n57169 ;
  assign n57171 = n83697 & n57170 ;
  assign n57172 = n57166 | n57171 ;
  assign n57173 = n67222 & n57172 ;
  assign n57174 = n56324 & n56813 ;
  assign n56618 = n56333 | n56617 ;
  assign n83758 = ~n56618 ;
  assign n57175 = n56614 & n83758 ;
  assign n83759 = ~n56619 ;
  assign n57176 = n56617 & n83759 ;
  assign n57177 = n57175 | n57176 ;
  assign n57178 = n73458 & n57177 ;
  assign n57179 = n83697 & n57178 ;
  assign n57180 = n57174 | n57179 ;
  assign n57181 = n67164 & n57180 ;
  assign n57182 = n56332 & n56813 ;
  assign n56613 = n56341 | n56612 ;
  assign n83760 = ~n56613 ;
  assign n57183 = n83760 & n56861 ;
  assign n83761 = ~n56862 ;
  assign n57184 = n56612 & n83761 ;
  assign n57185 = n57183 | n57184 ;
  assign n57186 = n73458 & n57185 ;
  assign n57187 = n83697 & n57186 ;
  assign n57188 = n57182 | n57187 ;
  assign n57189 = n66979 & n57188 ;
  assign n57190 = n56340 & n56813 ;
  assign n56606 = n56349 | n56605 ;
  assign n83762 = ~n56606 ;
  assign n57191 = n56602 & n83762 ;
  assign n83763 = ~n56607 ;
  assign n57192 = n56605 & n83763 ;
  assign n57193 = n57191 | n57192 ;
  assign n57194 = n73458 & n57193 ;
  assign n57195 = n83697 & n57194 ;
  assign n57196 = n57190 | n57195 ;
  assign n57197 = n66868 & n57196 ;
  assign n57198 = n56348 & n56813 ;
  assign n56601 = n56357 | n56600 ;
  assign n83764 = ~n56601 ;
  assign n57199 = n83764 & n56857 ;
  assign n83765 = ~n56858 ;
  assign n57200 = n56600 & n83765 ;
  assign n57201 = n57199 | n57200 ;
  assign n57202 = n73458 & n57201 ;
  assign n57203 = n83697 & n57202 ;
  assign n57204 = n57198 | n57203 ;
  assign n57205 = n66797 & n57204 ;
  assign n57206 = n56356 & n56813 ;
  assign n56594 = n56365 | n56593 ;
  assign n83766 = ~n56594 ;
  assign n57207 = n56590 & n83766 ;
  assign n83767 = ~n56595 ;
  assign n57208 = n56593 & n83767 ;
  assign n57209 = n57207 | n57208 ;
  assign n57210 = n73458 & n57209 ;
  assign n57211 = n83697 & n57210 ;
  assign n57212 = n57206 | n57211 ;
  assign n57213 = n66654 & n57212 ;
  assign n57214 = n56364 & n56813 ;
  assign n56589 = n56373 | n56588 ;
  assign n83768 = ~n56589 ;
  assign n57215 = n83768 & n56853 ;
  assign n83769 = ~n56854 ;
  assign n57216 = n56588 & n83769 ;
  assign n57217 = n57215 | n57216 ;
  assign n57218 = n73458 & n57217 ;
  assign n57219 = n83697 & n57218 ;
  assign n57220 = n57214 | n57219 ;
  assign n57221 = n66560 & n57220 ;
  assign n57222 = n56372 & n56813 ;
  assign n56582 = n56381 | n56581 ;
  assign n83770 = ~n56582 ;
  assign n57223 = n56578 & n83770 ;
  assign n83771 = ~n56583 ;
  assign n57224 = n56581 & n83771 ;
  assign n57225 = n57223 | n57224 ;
  assign n57226 = n73458 & n57225 ;
  assign n57227 = n83697 & n57226 ;
  assign n57228 = n57222 | n57227 ;
  assign n57229 = n66505 & n57228 ;
  assign n57230 = n56380 & n56813 ;
  assign n56577 = n56389 | n56576 ;
  assign n83772 = ~n56577 ;
  assign n57231 = n83772 & n56849 ;
  assign n83773 = ~n56850 ;
  assign n57232 = n56576 & n83773 ;
  assign n57233 = n57231 | n57232 ;
  assign n57234 = n73458 & n57233 ;
  assign n57235 = n83697 & n57234 ;
  assign n57236 = n57230 | n57235 ;
  assign n57237 = n66379 & n57236 ;
  assign n57238 = n56388 & n56813 ;
  assign n56570 = n56397 | n56569 ;
  assign n83774 = ~n56570 ;
  assign n57239 = n56566 & n83774 ;
  assign n83775 = ~n56571 ;
  assign n57240 = n56569 & n83775 ;
  assign n57241 = n57239 | n57240 ;
  assign n57242 = n73458 & n57241 ;
  assign n57243 = n83697 & n57242 ;
  assign n57244 = n57238 | n57243 ;
  assign n57245 = n66299 & n57244 ;
  assign n57246 = n56396 & n56813 ;
  assign n56565 = n56405 | n56564 ;
  assign n83776 = ~n56565 ;
  assign n57247 = n83776 & n56845 ;
  assign n83777 = ~n56846 ;
  assign n57248 = n56564 & n83777 ;
  assign n57249 = n57247 | n57248 ;
  assign n57250 = n73458 & n57249 ;
  assign n57251 = n83697 & n57250 ;
  assign n57252 = n57246 | n57251 ;
  assign n57253 = n66244 & n57252 ;
  assign n57254 = n56404 & n56813 ;
  assign n56558 = n56413 | n56557 ;
  assign n83778 = ~n56558 ;
  assign n57255 = n56554 & n83778 ;
  assign n83779 = ~n56559 ;
  assign n57256 = n56557 & n83779 ;
  assign n57257 = n57255 | n57256 ;
  assign n57258 = n73458 & n57257 ;
  assign n57259 = n83697 & n57258 ;
  assign n57260 = n57254 | n57259 ;
  assign n57261 = n66145 & n57260 ;
  assign n57262 = n56412 & n56813 ;
  assign n56553 = n56421 | n56552 ;
  assign n83780 = ~n56553 ;
  assign n57263 = n83780 & n56841 ;
  assign n83781 = ~n56842 ;
  assign n57264 = n56552 & n83781 ;
  assign n57265 = n57263 | n57264 ;
  assign n57266 = n73458 & n57265 ;
  assign n57267 = n83697 & n57266 ;
  assign n57268 = n57262 | n57267 ;
  assign n57269 = n66081 & n57268 ;
  assign n57270 = n56420 & n56813 ;
  assign n56546 = n56429 | n56545 ;
  assign n83782 = ~n56546 ;
  assign n57271 = n56542 & n83782 ;
  assign n83783 = ~n56547 ;
  assign n57272 = n56545 & n83783 ;
  assign n57273 = n57271 | n57272 ;
  assign n57274 = n73458 & n57273 ;
  assign n57275 = n83697 & n57274 ;
  assign n57276 = n57270 | n57275 ;
  assign n57277 = n66043 & n57276 ;
  assign n57278 = n56428 & n56813 ;
  assign n56541 = n56437 | n56540 ;
  assign n83784 = ~n56541 ;
  assign n57279 = n83784 & n56837 ;
  assign n83785 = ~n56838 ;
  assign n57280 = n56540 & n83785 ;
  assign n57281 = n57279 | n57280 ;
  assign n57282 = n73458 & n57281 ;
  assign n57283 = n83697 & n57282 ;
  assign n57284 = n57278 | n57283 ;
  assign n57285 = n65960 & n57284 ;
  assign n57286 = n56436 & n56813 ;
  assign n56534 = n56445 | n56533 ;
  assign n83786 = ~n56534 ;
  assign n57287 = n56530 & n83786 ;
  assign n83787 = ~n56535 ;
  assign n57288 = n56533 & n83787 ;
  assign n57289 = n57287 | n57288 ;
  assign n57290 = n73458 & n57289 ;
  assign n57291 = n83697 & n57290 ;
  assign n57292 = n57286 | n57291 ;
  assign n57293 = n65909 & n57292 ;
  assign n57294 = n56444 & n56813 ;
  assign n56529 = n56453 | n56528 ;
  assign n83788 = ~n56529 ;
  assign n57295 = n83788 & n56833 ;
  assign n83789 = ~n56834 ;
  assign n57296 = n56528 & n83789 ;
  assign n57297 = n57295 | n57296 ;
  assign n57298 = n73458 & n57297 ;
  assign n57299 = n83697 & n57298 ;
  assign n57300 = n57294 | n57299 ;
  assign n57301 = n65877 & n57300 ;
  assign n57302 = n56452 & n56813 ;
  assign n56522 = n56461 | n56521 ;
  assign n83790 = ~n56522 ;
  assign n57303 = n56518 & n83790 ;
  assign n83791 = ~n56523 ;
  assign n57304 = n56521 & n83791 ;
  assign n57305 = n57303 | n57304 ;
  assign n57306 = n73458 & n57305 ;
  assign n57307 = n83697 & n57306 ;
  assign n57308 = n57302 | n57307 ;
  assign n57309 = n65820 & n57308 ;
  assign n57310 = n56460 & n56813 ;
  assign n56517 = n56469 | n56516 ;
  assign n83792 = ~n56517 ;
  assign n57311 = n83792 & n56829 ;
  assign n83793 = ~n56830 ;
  assign n57312 = n56516 & n83793 ;
  assign n57313 = n57311 | n57312 ;
  assign n57314 = n73458 & n57313 ;
  assign n57315 = n83697 & n57314 ;
  assign n57316 = n57310 | n57315 ;
  assign n57317 = n65791 & n57316 ;
  assign n57318 = n56468 & n56813 ;
  assign n57319 = n56478 | n56510 ;
  assign n83794 = ~n57319 ;
  assign n57320 = n56507 & n83794 ;
  assign n83795 = ~n56511 ;
  assign n57321 = n56510 & n83795 ;
  assign n57322 = n57320 | n57321 ;
  assign n57323 = n73458 & n57322 ;
  assign n57324 = n83697 & n57323 ;
  assign n57325 = n57318 | n57324 ;
  assign n57326 = n65772 & n57325 ;
  assign n57327 = n56477 & n56813 ;
  assign n57328 = n56486 | n56506 ;
  assign n83796 = ~n57328 ;
  assign n57329 = n56502 & n83796 ;
  assign n83797 = ~n56826 ;
  assign n57330 = n56506 & n83797 ;
  assign n57331 = n57329 | n57330 ;
  assign n57332 = n73458 & n57331 ;
  assign n57333 = n83697 & n57332 ;
  assign n57334 = n57327 | n57333 ;
  assign n57335 = n65746 & n57334 ;
  assign n57336 = n56485 & n56813 ;
  assign n56824 = n56497 | n56500 ;
  assign n83798 = ~n56824 ;
  assign n57337 = n56822 & n83798 ;
  assign n83799 = ~n56501 ;
  assign n57338 = n56500 & n83799 ;
  assign n57339 = n57337 | n57338 ;
  assign n57340 = n73458 & n57339 ;
  assign n57341 = n83697 & n57340 ;
  assign n57342 = n57336 | n57341 ;
  assign n57343 = n65721 & n57342 ;
  assign n56815 = n56488 & n56813 ;
  assign n56495 = n24281 & n56493 ;
  assign n57344 = n56495 & n83692 ;
  assign n57345 = n24576 | n57344 ;
  assign n83800 = ~n57345 ;
  assign n57346 = n56822 & n83800 ;
  assign n57347 = n83697 & n57346 ;
  assign n57348 = n56815 | n57347 ;
  assign n57349 = n65686 & n57348 ;
  assign n57350 = n25150 & n83697 ;
  assign n57352 = n83687 & n57351 ;
  assign n57353 = n56809 | n57352 ;
  assign n57354 = n83688 & n57353 ;
  assign n83801 = ~n57354 ;
  assign n57355 = n25145 & n83801 ;
  assign n83802 = ~n57355 ;
  assign n57356 = x9 & n83802 ;
  assign n57357 = n57350 | n57356 ;
  assign n57365 = n65670 & n57357 ;
  assign n57358 = n25145 & n83697 ;
  assign n83803 = ~n57358 ;
  assign n57359 = x9 & n83803 ;
  assign n57360 = n57350 | n57359 ;
  assign n57361 = x65 & n57360 ;
  assign n57362 = x65 | n57350 ;
  assign n57363 = n57359 | n57362 ;
  assign n83804 = ~n57361 ;
  assign n57364 = n83804 & n57363 ;
  assign n57366 = n25157 | n57364 ;
  assign n83805 = ~n57365 ;
  assign n57367 = n83805 & n57366 ;
  assign n83806 = ~n57347 ;
  assign n57368 = x66 & n83806 ;
  assign n83807 = ~n56815 ;
  assign n57369 = n83807 & n57368 ;
  assign n57370 = n57367 | n57369 ;
  assign n83808 = ~n57349 ;
  assign n57371 = n83808 & n57370 ;
  assign n83809 = ~n57341 ;
  assign n57372 = x67 & n83809 ;
  assign n83810 = ~n57336 ;
  assign n57373 = n83810 & n57372 ;
  assign n57374 = n57343 | n57373 ;
  assign n57375 = n57371 | n57374 ;
  assign n83811 = ~n57343 ;
  assign n57376 = n83811 & n57375 ;
  assign n83812 = ~n57333 ;
  assign n57377 = x68 & n83812 ;
  assign n83813 = ~n57327 ;
  assign n57378 = n83813 & n57377 ;
  assign n57379 = n57335 | n57378 ;
  assign n57380 = n57376 | n57379 ;
  assign n83814 = ~n57335 ;
  assign n57381 = n83814 & n57380 ;
  assign n83815 = ~n57324 ;
  assign n57382 = x69 & n83815 ;
  assign n83816 = ~n57318 ;
  assign n57383 = n83816 & n57382 ;
  assign n57384 = n57326 | n57383 ;
  assign n57385 = n57381 | n57384 ;
  assign n83817 = ~n57326 ;
  assign n57386 = n83817 & n57385 ;
  assign n83818 = ~n57315 ;
  assign n57387 = x70 & n83818 ;
  assign n83819 = ~n57310 ;
  assign n57388 = n83819 & n57387 ;
  assign n57389 = n57317 | n57388 ;
  assign n57391 = n57386 | n57389 ;
  assign n83820 = ~n57317 ;
  assign n57392 = n83820 & n57391 ;
  assign n83821 = ~n57307 ;
  assign n57393 = x71 & n83821 ;
  assign n83822 = ~n57302 ;
  assign n57394 = n83822 & n57393 ;
  assign n57395 = n57309 | n57394 ;
  assign n57396 = n57392 | n57395 ;
  assign n83823 = ~n57309 ;
  assign n57397 = n83823 & n57396 ;
  assign n83824 = ~n57299 ;
  assign n57398 = x72 & n83824 ;
  assign n83825 = ~n57294 ;
  assign n57399 = n83825 & n57398 ;
  assign n57400 = n57301 | n57399 ;
  assign n57402 = n57397 | n57400 ;
  assign n83826 = ~n57301 ;
  assign n57403 = n83826 & n57402 ;
  assign n83827 = ~n57291 ;
  assign n57404 = x73 & n83827 ;
  assign n83828 = ~n57286 ;
  assign n57405 = n83828 & n57404 ;
  assign n57406 = n57293 | n57405 ;
  assign n57407 = n57403 | n57406 ;
  assign n83829 = ~n57293 ;
  assign n57408 = n83829 & n57407 ;
  assign n83830 = ~n57283 ;
  assign n57409 = x74 & n83830 ;
  assign n83831 = ~n57278 ;
  assign n57410 = n83831 & n57409 ;
  assign n57411 = n57285 | n57410 ;
  assign n57413 = n57408 | n57411 ;
  assign n83832 = ~n57285 ;
  assign n57414 = n83832 & n57413 ;
  assign n83833 = ~n57275 ;
  assign n57415 = x75 & n83833 ;
  assign n83834 = ~n57270 ;
  assign n57416 = n83834 & n57415 ;
  assign n57417 = n57277 | n57416 ;
  assign n57418 = n57414 | n57417 ;
  assign n83835 = ~n57277 ;
  assign n57419 = n83835 & n57418 ;
  assign n83836 = ~n57267 ;
  assign n57420 = x76 & n83836 ;
  assign n83837 = ~n57262 ;
  assign n57421 = n83837 & n57420 ;
  assign n57422 = n57269 | n57421 ;
  assign n57424 = n57419 | n57422 ;
  assign n83838 = ~n57269 ;
  assign n57425 = n83838 & n57424 ;
  assign n83839 = ~n57259 ;
  assign n57426 = x77 & n83839 ;
  assign n83840 = ~n57254 ;
  assign n57427 = n83840 & n57426 ;
  assign n57428 = n57261 | n57427 ;
  assign n57429 = n57425 | n57428 ;
  assign n83841 = ~n57261 ;
  assign n57430 = n83841 & n57429 ;
  assign n83842 = ~n57251 ;
  assign n57431 = x78 & n83842 ;
  assign n83843 = ~n57246 ;
  assign n57432 = n83843 & n57431 ;
  assign n57433 = n57253 | n57432 ;
  assign n57435 = n57430 | n57433 ;
  assign n83844 = ~n57253 ;
  assign n57436 = n83844 & n57435 ;
  assign n83845 = ~n57243 ;
  assign n57437 = x79 & n83845 ;
  assign n83846 = ~n57238 ;
  assign n57438 = n83846 & n57437 ;
  assign n57439 = n57245 | n57438 ;
  assign n57440 = n57436 | n57439 ;
  assign n83847 = ~n57245 ;
  assign n57441 = n83847 & n57440 ;
  assign n83848 = ~n57235 ;
  assign n57442 = x80 & n83848 ;
  assign n83849 = ~n57230 ;
  assign n57443 = n83849 & n57442 ;
  assign n57444 = n57237 | n57443 ;
  assign n57446 = n57441 | n57444 ;
  assign n83850 = ~n57237 ;
  assign n57447 = n83850 & n57446 ;
  assign n83851 = ~n57227 ;
  assign n57448 = x81 & n83851 ;
  assign n83852 = ~n57222 ;
  assign n57449 = n83852 & n57448 ;
  assign n57450 = n57229 | n57449 ;
  assign n57451 = n57447 | n57450 ;
  assign n83853 = ~n57229 ;
  assign n57452 = n83853 & n57451 ;
  assign n83854 = ~n57219 ;
  assign n57453 = x82 & n83854 ;
  assign n83855 = ~n57214 ;
  assign n57454 = n83855 & n57453 ;
  assign n57455 = n57221 | n57454 ;
  assign n57457 = n57452 | n57455 ;
  assign n83856 = ~n57221 ;
  assign n57458 = n83856 & n57457 ;
  assign n83857 = ~n57211 ;
  assign n57459 = x83 & n83857 ;
  assign n83858 = ~n57206 ;
  assign n57460 = n83858 & n57459 ;
  assign n57461 = n57213 | n57460 ;
  assign n57462 = n57458 | n57461 ;
  assign n83859 = ~n57213 ;
  assign n57463 = n83859 & n57462 ;
  assign n83860 = ~n57203 ;
  assign n57464 = x84 & n83860 ;
  assign n83861 = ~n57198 ;
  assign n57465 = n83861 & n57464 ;
  assign n57466 = n57205 | n57465 ;
  assign n57468 = n57463 | n57466 ;
  assign n83862 = ~n57205 ;
  assign n57469 = n83862 & n57468 ;
  assign n83863 = ~n57195 ;
  assign n57470 = x85 & n83863 ;
  assign n83864 = ~n57190 ;
  assign n57471 = n83864 & n57470 ;
  assign n57472 = n57197 | n57471 ;
  assign n57473 = n57469 | n57472 ;
  assign n83865 = ~n57197 ;
  assign n57474 = n83865 & n57473 ;
  assign n83866 = ~n57187 ;
  assign n57475 = x86 & n83866 ;
  assign n83867 = ~n57182 ;
  assign n57476 = n83867 & n57475 ;
  assign n57477 = n57189 | n57476 ;
  assign n57479 = n57474 | n57477 ;
  assign n83868 = ~n57189 ;
  assign n57480 = n83868 & n57479 ;
  assign n83869 = ~n57179 ;
  assign n57481 = x87 & n83869 ;
  assign n83870 = ~n57174 ;
  assign n57482 = n83870 & n57481 ;
  assign n57483 = n57181 | n57482 ;
  assign n57484 = n57480 | n57483 ;
  assign n83871 = ~n57181 ;
  assign n57485 = n83871 & n57484 ;
  assign n83872 = ~n57171 ;
  assign n57486 = x88 & n83872 ;
  assign n83873 = ~n57166 ;
  assign n57487 = n83873 & n57486 ;
  assign n57488 = n57173 | n57487 ;
  assign n57490 = n57485 | n57488 ;
  assign n83874 = ~n57173 ;
  assign n57491 = n83874 & n57490 ;
  assign n83875 = ~n57163 ;
  assign n57492 = x89 & n83875 ;
  assign n83876 = ~n57158 ;
  assign n57493 = n83876 & n57492 ;
  assign n57494 = n57165 | n57493 ;
  assign n57495 = n57491 | n57494 ;
  assign n83877 = ~n57165 ;
  assign n57496 = n83877 & n57495 ;
  assign n83878 = ~n57155 ;
  assign n57497 = x90 & n83878 ;
  assign n83879 = ~n57150 ;
  assign n57498 = n83879 & n57497 ;
  assign n57499 = n57157 | n57498 ;
  assign n57501 = n57496 | n57499 ;
  assign n83880 = ~n57157 ;
  assign n57502 = n83880 & n57501 ;
  assign n83881 = ~n57147 ;
  assign n57503 = x91 & n83881 ;
  assign n83882 = ~n57142 ;
  assign n57504 = n83882 & n57503 ;
  assign n57505 = n57149 | n57504 ;
  assign n57506 = n57502 | n57505 ;
  assign n83883 = ~n57149 ;
  assign n57507 = n83883 & n57506 ;
  assign n83884 = ~n57139 ;
  assign n57508 = x92 & n83884 ;
  assign n83885 = ~n57134 ;
  assign n57509 = n83885 & n57508 ;
  assign n57510 = n57141 | n57509 ;
  assign n57512 = n57507 | n57510 ;
  assign n83886 = ~n57141 ;
  assign n57513 = n83886 & n57512 ;
  assign n83887 = ~n57131 ;
  assign n57514 = x93 & n83887 ;
  assign n83888 = ~n57126 ;
  assign n57515 = n83888 & n57514 ;
  assign n57516 = n57133 | n57515 ;
  assign n57517 = n57513 | n57516 ;
  assign n83889 = ~n57133 ;
  assign n57518 = n83889 & n57517 ;
  assign n83890 = ~n57123 ;
  assign n57519 = x94 & n83890 ;
  assign n83891 = ~n57118 ;
  assign n57520 = n83891 & n57519 ;
  assign n57521 = n57125 | n57520 ;
  assign n57523 = n57518 | n57521 ;
  assign n83892 = ~n57125 ;
  assign n57524 = n83892 & n57523 ;
  assign n83893 = ~n57115 ;
  assign n57525 = x95 & n83893 ;
  assign n83894 = ~n57110 ;
  assign n57526 = n83894 & n57525 ;
  assign n57527 = n57117 | n57526 ;
  assign n57528 = n57524 | n57527 ;
  assign n83895 = ~n57117 ;
  assign n57529 = n83895 & n57528 ;
  assign n83896 = ~n57107 ;
  assign n57530 = x96 & n83896 ;
  assign n83897 = ~n57102 ;
  assign n57531 = n83897 & n57530 ;
  assign n57532 = n57109 | n57531 ;
  assign n57534 = n57529 | n57532 ;
  assign n83898 = ~n57109 ;
  assign n57535 = n83898 & n57534 ;
  assign n83899 = ~n57099 ;
  assign n57536 = x97 & n83899 ;
  assign n83900 = ~n57094 ;
  assign n57537 = n83900 & n57536 ;
  assign n57538 = n57101 | n57537 ;
  assign n57539 = n57535 | n57538 ;
  assign n83901 = ~n57101 ;
  assign n57540 = n83901 & n57539 ;
  assign n83902 = ~n57091 ;
  assign n57541 = x98 & n83902 ;
  assign n83903 = ~n57086 ;
  assign n57542 = n83903 & n57541 ;
  assign n57543 = n57093 | n57542 ;
  assign n57545 = n57540 | n57543 ;
  assign n83904 = ~n57093 ;
  assign n57546 = n83904 & n57545 ;
  assign n83905 = ~n57083 ;
  assign n57547 = x99 & n83905 ;
  assign n83906 = ~n57078 ;
  assign n57548 = n83906 & n57547 ;
  assign n57549 = n57085 | n57548 ;
  assign n57550 = n57546 | n57549 ;
  assign n83907 = ~n57085 ;
  assign n57551 = n83907 & n57550 ;
  assign n83908 = ~n57075 ;
  assign n57552 = x100 & n83908 ;
  assign n83909 = ~n57070 ;
  assign n57553 = n83909 & n57552 ;
  assign n57554 = n57077 | n57553 ;
  assign n57556 = n57551 | n57554 ;
  assign n83910 = ~n57077 ;
  assign n57557 = n83910 & n57556 ;
  assign n83911 = ~n57067 ;
  assign n57558 = x101 & n83911 ;
  assign n83912 = ~n57062 ;
  assign n57559 = n83912 & n57558 ;
  assign n57560 = n57069 | n57559 ;
  assign n57561 = n57557 | n57560 ;
  assign n83913 = ~n57069 ;
  assign n57562 = n83913 & n57561 ;
  assign n83914 = ~n57059 ;
  assign n57563 = x102 & n83914 ;
  assign n83915 = ~n57054 ;
  assign n57564 = n83915 & n57563 ;
  assign n57565 = n57061 | n57564 ;
  assign n57567 = n57562 | n57565 ;
  assign n83916 = ~n57061 ;
  assign n57568 = n83916 & n57567 ;
  assign n83917 = ~n57051 ;
  assign n57569 = x103 & n83917 ;
  assign n83918 = ~n57046 ;
  assign n57570 = n83918 & n57569 ;
  assign n57571 = n57053 | n57570 ;
  assign n57572 = n57568 | n57571 ;
  assign n83919 = ~n57053 ;
  assign n57573 = n83919 & n57572 ;
  assign n83920 = ~n57043 ;
  assign n57574 = x104 & n83920 ;
  assign n83921 = ~n57038 ;
  assign n57575 = n83921 & n57574 ;
  assign n57576 = n57045 | n57575 ;
  assign n57578 = n57573 | n57576 ;
  assign n83922 = ~n57045 ;
  assign n57579 = n83922 & n57578 ;
  assign n83923 = ~n57035 ;
  assign n57580 = x105 & n83923 ;
  assign n83924 = ~n57030 ;
  assign n57581 = n83924 & n57580 ;
  assign n57582 = n57037 | n57581 ;
  assign n57583 = n57579 | n57582 ;
  assign n83925 = ~n57037 ;
  assign n57584 = n83925 & n57583 ;
  assign n83926 = ~n57027 ;
  assign n57585 = x106 & n83926 ;
  assign n83927 = ~n57022 ;
  assign n57586 = n83927 & n57585 ;
  assign n57587 = n57029 | n57586 ;
  assign n57589 = n57584 | n57587 ;
  assign n83928 = ~n57029 ;
  assign n57590 = n83928 & n57589 ;
  assign n83929 = ~n57019 ;
  assign n57591 = x107 & n83929 ;
  assign n83930 = ~n57014 ;
  assign n57592 = n83930 & n57591 ;
  assign n57593 = n57021 | n57592 ;
  assign n57594 = n57590 | n57593 ;
  assign n83931 = ~n57021 ;
  assign n57595 = n83931 & n57594 ;
  assign n83932 = ~n57011 ;
  assign n57596 = x108 & n83932 ;
  assign n83933 = ~n57006 ;
  assign n57597 = n83933 & n57596 ;
  assign n57598 = n57013 | n57597 ;
  assign n57600 = n57595 | n57598 ;
  assign n83934 = ~n57013 ;
  assign n57601 = n83934 & n57600 ;
  assign n83935 = ~n57003 ;
  assign n57602 = x109 & n83935 ;
  assign n83936 = ~n56998 ;
  assign n57603 = n83936 & n57602 ;
  assign n57604 = n57005 | n57603 ;
  assign n57605 = n57601 | n57604 ;
  assign n83937 = ~n57005 ;
  assign n57606 = n83937 & n57605 ;
  assign n83938 = ~n56995 ;
  assign n57607 = x110 & n83938 ;
  assign n83939 = ~n56990 ;
  assign n57608 = n83939 & n57607 ;
  assign n57609 = n56997 | n57608 ;
  assign n57611 = n57606 | n57609 ;
  assign n83940 = ~n56997 ;
  assign n57612 = n83940 & n57611 ;
  assign n83941 = ~n56987 ;
  assign n57613 = x111 & n83941 ;
  assign n83942 = ~n56982 ;
  assign n57614 = n83942 & n57613 ;
  assign n57615 = n56989 | n57614 ;
  assign n57616 = n57612 | n57615 ;
  assign n83943 = ~n56989 ;
  assign n57617 = n83943 & n57616 ;
  assign n83944 = ~n56979 ;
  assign n57618 = x112 & n83944 ;
  assign n83945 = ~n56974 ;
  assign n57619 = n83945 & n57618 ;
  assign n57620 = n56981 | n57619 ;
  assign n57622 = n57617 | n57620 ;
  assign n83946 = ~n56981 ;
  assign n57623 = n83946 & n57622 ;
  assign n83947 = ~n56971 ;
  assign n57624 = x113 & n83947 ;
  assign n83948 = ~n56966 ;
  assign n57625 = n83948 & n57624 ;
  assign n57626 = n56973 | n57625 ;
  assign n57627 = n57623 | n57626 ;
  assign n83949 = ~n56973 ;
  assign n57628 = n83949 & n57627 ;
  assign n83950 = ~n56963 ;
  assign n57629 = x114 & n83950 ;
  assign n83951 = ~n56958 ;
  assign n57630 = n83951 & n57629 ;
  assign n57631 = n56965 | n57630 ;
  assign n57633 = n57628 | n57631 ;
  assign n83952 = ~n56965 ;
  assign n57634 = n83952 & n57633 ;
  assign n83953 = ~n56955 ;
  assign n57635 = x115 & n83953 ;
  assign n83954 = ~n56950 ;
  assign n57636 = n83954 & n57635 ;
  assign n57637 = n56957 | n57636 ;
  assign n57638 = n57634 | n57637 ;
  assign n83955 = ~n56957 ;
  assign n57639 = n83955 & n57638 ;
  assign n83956 = ~n56947 ;
  assign n57640 = x116 & n83956 ;
  assign n83957 = ~n56942 ;
  assign n57641 = n83957 & n57640 ;
  assign n57642 = n56949 | n57641 ;
  assign n57644 = n57639 | n57642 ;
  assign n83958 = ~n56949 ;
  assign n57645 = n83958 & n57644 ;
  assign n83959 = ~n56939 ;
  assign n57646 = x117 & n83959 ;
  assign n83960 = ~n56934 ;
  assign n57647 = n83960 & n57646 ;
  assign n57648 = n56941 | n57647 ;
  assign n57649 = n57645 | n57648 ;
  assign n83961 = ~n56941 ;
  assign n57650 = n83961 & n57649 ;
  assign n83962 = ~n56931 ;
  assign n57651 = x118 & n83962 ;
  assign n83963 = ~n56816 ;
  assign n57652 = n83963 & n57651 ;
  assign n57653 = n56933 | n57652 ;
  assign n57655 = n57650 | n57653 ;
  assign n83964 = ~n56933 ;
  assign n57656 = n83964 & n57655 ;
  assign n57663 = n73617 & n57662 ;
  assign n83965 = ~n56813 ;
  assign n57664 = n83965 & n57660 ;
  assign n57665 = n56075 & n56813 ;
  assign n83966 = ~n57665 ;
  assign n57666 = x119 & n83966 ;
  assign n83967 = ~n57664 ;
  assign n57667 = n83967 & n57666 ;
  assign n57668 = n66655 | n57667 ;
  assign n57669 = n57663 | n57668 ;
  assign n57671 = n57656 | n57669 ;
  assign n83968 = ~n57670 ;
  assign n57672 = n83968 & n57671 ;
  assign n83969 = ~n57650 ;
  assign n57654 = n83969 & n57653 ;
  assign n57675 = x65 & n57357 ;
  assign n83970 = ~n57675 ;
  assign n57676 = n57363 & n83970 ;
  assign n57677 = n25157 | n57676 ;
  assign n57678 = n83805 & n57677 ;
  assign n57679 = n57349 | n57369 ;
  assign n57681 = n57678 | n57679 ;
  assign n57682 = n83808 & n57681 ;
  assign n57683 = n57373 | n57682 ;
  assign n57685 = n83811 & n57683 ;
  assign n57687 = n57379 | n57685 ;
  assign n57688 = n83814 & n57687 ;
  assign n57690 = n57384 | n57688 ;
  assign n57691 = n83817 & n57690 ;
  assign n57692 = n57389 | n57691 ;
  assign n57693 = n83820 & n57692 ;
  assign n57694 = n57395 | n57693 ;
  assign n57696 = n83823 & n57694 ;
  assign n57697 = n57400 | n57696 ;
  assign n57698 = n83826 & n57697 ;
  assign n57699 = n57406 | n57698 ;
  assign n57701 = n83829 & n57699 ;
  assign n57702 = n57411 | n57701 ;
  assign n57703 = n83832 & n57702 ;
  assign n57704 = n57417 | n57703 ;
  assign n57706 = n83835 & n57704 ;
  assign n57707 = n57422 | n57706 ;
  assign n57708 = n83838 & n57707 ;
  assign n57709 = n57428 | n57708 ;
  assign n57711 = n83841 & n57709 ;
  assign n57712 = n57433 | n57711 ;
  assign n57713 = n83844 & n57712 ;
  assign n57714 = n57439 | n57713 ;
  assign n57716 = n83847 & n57714 ;
  assign n57717 = n57444 | n57716 ;
  assign n57718 = n83850 & n57717 ;
  assign n57719 = n57450 | n57718 ;
  assign n57721 = n83853 & n57719 ;
  assign n57722 = n57455 | n57721 ;
  assign n57723 = n83856 & n57722 ;
  assign n57724 = n57461 | n57723 ;
  assign n57726 = n83859 & n57724 ;
  assign n57727 = n57466 | n57726 ;
  assign n57728 = n83862 & n57727 ;
  assign n57729 = n57472 | n57728 ;
  assign n57731 = n83865 & n57729 ;
  assign n57732 = n57477 | n57731 ;
  assign n57733 = n83868 & n57732 ;
  assign n57734 = n57483 | n57733 ;
  assign n57736 = n83871 & n57734 ;
  assign n57737 = n57488 | n57736 ;
  assign n57738 = n83874 & n57737 ;
  assign n57739 = n57494 | n57738 ;
  assign n57741 = n83877 & n57739 ;
  assign n57742 = n57499 | n57741 ;
  assign n57743 = n83880 & n57742 ;
  assign n57744 = n57505 | n57743 ;
  assign n57746 = n83883 & n57744 ;
  assign n57747 = n57510 | n57746 ;
  assign n57748 = n83886 & n57747 ;
  assign n57749 = n57516 | n57748 ;
  assign n57751 = n83889 & n57749 ;
  assign n57752 = n57521 | n57751 ;
  assign n57753 = n83892 & n57752 ;
  assign n57754 = n57527 | n57753 ;
  assign n57756 = n83895 & n57754 ;
  assign n57757 = n57532 | n57756 ;
  assign n57758 = n83898 & n57757 ;
  assign n57759 = n57538 | n57758 ;
  assign n57761 = n83901 & n57759 ;
  assign n57762 = n57543 | n57761 ;
  assign n57763 = n83904 & n57762 ;
  assign n57764 = n57549 | n57763 ;
  assign n57766 = n83907 & n57764 ;
  assign n57767 = n57554 | n57766 ;
  assign n57768 = n83910 & n57767 ;
  assign n57769 = n57560 | n57768 ;
  assign n57771 = n83913 & n57769 ;
  assign n57772 = n57565 | n57771 ;
  assign n57773 = n83916 & n57772 ;
  assign n57774 = n57571 | n57773 ;
  assign n57776 = n83919 & n57774 ;
  assign n57777 = n57576 | n57776 ;
  assign n57778 = n83922 & n57777 ;
  assign n57779 = n57582 | n57778 ;
  assign n57781 = n83925 & n57779 ;
  assign n57782 = n57587 | n57781 ;
  assign n57783 = n83928 & n57782 ;
  assign n57784 = n57593 | n57783 ;
  assign n57786 = n83931 & n57784 ;
  assign n57787 = n57598 | n57786 ;
  assign n57788 = n83934 & n57787 ;
  assign n57789 = n57604 | n57788 ;
  assign n57791 = n83937 & n57789 ;
  assign n57792 = n57609 | n57791 ;
  assign n57793 = n83940 & n57792 ;
  assign n57794 = n57615 | n57793 ;
  assign n57796 = n83943 & n57794 ;
  assign n57797 = n57620 | n57796 ;
  assign n57798 = n83946 & n57797 ;
  assign n57799 = n57626 | n57798 ;
  assign n57801 = n83949 & n57799 ;
  assign n57802 = n57631 | n57801 ;
  assign n57803 = n83952 & n57802 ;
  assign n57804 = n57637 | n57803 ;
  assign n57806 = n83955 & n57804 ;
  assign n57807 = n57642 | n57806 ;
  assign n57808 = n83958 & n57807 ;
  assign n57810 = n57648 | n57808 ;
  assign n57811 = n56941 | n57653 ;
  assign n83971 = ~n57811 ;
  assign n57812 = n57810 & n83971 ;
  assign n57813 = n57654 | n57812 ;
  assign n83972 = ~n57672 ;
  assign n57814 = n83972 & n57813 ;
  assign n57815 = n83961 & n57810 ;
  assign n57816 = n57653 | n57815 ;
  assign n57817 = n83964 & n57816 ;
  assign n57818 = n57669 | n57817 ;
  assign n57819 = n56932 & n83968 ;
  assign n57820 = n57818 & n57819 ;
  assign n57821 = n57814 | n57820 ;
  assign n57822 = n73617 & n57821 ;
  assign n83973 = ~n57820 ;
  assign n58531 = x119 & n83973 ;
  assign n83974 = ~n57814 ;
  assign n58532 = n83974 & n58531 ;
  assign n58533 = n57822 | n58532 ;
  assign n83975 = ~n57808 ;
  assign n57809 = n57648 & n83975 ;
  assign n57823 = n56949 | n57648 ;
  assign n83976 = ~n57823 ;
  assign n57824 = n57644 & n83976 ;
  assign n57825 = n57809 | n57824 ;
  assign n57826 = n83972 & n57825 ;
  assign n57827 = n56940 & n83968 ;
  assign n57828 = n57818 & n57827 ;
  assign n57829 = n57826 | n57828 ;
  assign n57830 = n73188 & n57829 ;
  assign n83977 = ~n57639 ;
  assign n57643 = n83977 & n57642 ;
  assign n57831 = n56957 | n57642 ;
  assign n83978 = ~n57831 ;
  assign n57832 = n57804 & n83978 ;
  assign n57833 = n57643 | n57832 ;
  assign n57834 = n83972 & n57833 ;
  assign n57835 = n56948 & n83968 ;
  assign n57836 = n57818 & n57835 ;
  assign n57837 = n57834 | n57836 ;
  assign n57838 = n73177 & n57837 ;
  assign n83979 = ~n57836 ;
  assign n58521 = x117 & n83979 ;
  assign n83980 = ~n57834 ;
  assign n58522 = n83980 & n58521 ;
  assign n58523 = n57838 | n58522 ;
  assign n83981 = ~n57803 ;
  assign n57805 = n57637 & n83981 ;
  assign n57839 = n56965 | n57637 ;
  assign n83982 = ~n57839 ;
  assign n57840 = n57633 & n83982 ;
  assign n57841 = n57805 | n57840 ;
  assign n57842 = n83972 & n57841 ;
  assign n57843 = n56956 & n83968 ;
  assign n57844 = n57818 & n57843 ;
  assign n57845 = n57842 | n57844 ;
  assign n57846 = n72752 & n57845 ;
  assign n83983 = ~n57628 ;
  assign n57632 = n83983 & n57631 ;
  assign n57847 = n56973 | n57631 ;
  assign n83984 = ~n57847 ;
  assign n57848 = n57799 & n83984 ;
  assign n57849 = n57632 | n57848 ;
  assign n57850 = n83972 & n57849 ;
  assign n57851 = n56964 & n83968 ;
  assign n57852 = n57818 & n57851 ;
  assign n57853 = n57850 | n57852 ;
  assign n57854 = n72393 & n57853 ;
  assign n83985 = ~n57852 ;
  assign n58511 = x115 & n83985 ;
  assign n83986 = ~n57850 ;
  assign n58512 = n83986 & n58511 ;
  assign n58513 = n57854 | n58512 ;
  assign n83987 = ~n57798 ;
  assign n57800 = n57626 & n83987 ;
  assign n57855 = n56981 | n57626 ;
  assign n83988 = ~n57855 ;
  assign n57856 = n57622 & n83988 ;
  assign n57857 = n57800 | n57856 ;
  assign n57858 = n83972 & n57857 ;
  assign n57859 = n56972 & n83968 ;
  assign n57860 = n57818 & n57859 ;
  assign n57861 = n57858 | n57860 ;
  assign n57862 = n72385 & n57861 ;
  assign n83989 = ~n57617 ;
  assign n57621 = n83989 & n57620 ;
  assign n57863 = n56989 | n57620 ;
  assign n83990 = ~n57863 ;
  assign n57864 = n57794 & n83990 ;
  assign n57865 = n57621 | n57864 ;
  assign n57866 = n83972 & n57865 ;
  assign n57867 = n56980 & n83968 ;
  assign n57868 = n57818 & n57867 ;
  assign n57869 = n57866 | n57868 ;
  assign n57870 = n72025 & n57869 ;
  assign n83991 = ~n57868 ;
  assign n58501 = x113 & n83991 ;
  assign n83992 = ~n57866 ;
  assign n58502 = n83992 & n58501 ;
  assign n58503 = n57870 | n58502 ;
  assign n83993 = ~n57793 ;
  assign n57795 = n57615 & n83993 ;
  assign n57871 = n56997 | n57615 ;
  assign n83994 = ~n57871 ;
  assign n57872 = n57611 & n83994 ;
  assign n57873 = n57795 | n57872 ;
  assign n57874 = n83972 & n57873 ;
  assign n57875 = n56988 & n83968 ;
  assign n57876 = n57818 & n57875 ;
  assign n57877 = n57874 | n57876 ;
  assign n57878 = n71645 & n57877 ;
  assign n83995 = ~n57606 ;
  assign n57610 = n83995 & n57609 ;
  assign n57879 = n57005 | n57609 ;
  assign n83996 = ~n57879 ;
  assign n57880 = n57789 & n83996 ;
  assign n57881 = n57610 | n57880 ;
  assign n57882 = n83972 & n57881 ;
  assign n57883 = n56996 & n83968 ;
  assign n57884 = n57818 & n57883 ;
  assign n57885 = n57882 | n57884 ;
  assign n57886 = n71633 & n57885 ;
  assign n83997 = ~n57884 ;
  assign n58491 = x111 & n83997 ;
  assign n83998 = ~n57882 ;
  assign n58492 = n83998 & n58491 ;
  assign n58493 = n57886 | n58492 ;
  assign n83999 = ~n57788 ;
  assign n57790 = n57604 & n83999 ;
  assign n57887 = n57013 | n57604 ;
  assign n84000 = ~n57887 ;
  assign n57888 = n57600 & n84000 ;
  assign n57889 = n57790 | n57888 ;
  assign n57890 = n83972 & n57889 ;
  assign n57891 = n57004 & n83968 ;
  assign n57892 = n57818 & n57891 ;
  assign n57893 = n57890 | n57892 ;
  assign n57894 = n71253 & n57893 ;
  assign n84001 = ~n57595 ;
  assign n57599 = n84001 & n57598 ;
  assign n57895 = n57021 | n57598 ;
  assign n84002 = ~n57895 ;
  assign n57896 = n57784 & n84002 ;
  assign n57897 = n57599 | n57896 ;
  assign n57898 = n83972 & n57897 ;
  assign n57899 = n57012 & n83968 ;
  assign n57900 = n57818 & n57899 ;
  assign n57901 = n57898 | n57900 ;
  assign n57902 = n70935 & n57901 ;
  assign n84003 = ~n57900 ;
  assign n58481 = x109 & n84003 ;
  assign n84004 = ~n57898 ;
  assign n58482 = n84004 & n58481 ;
  assign n58483 = n57902 | n58482 ;
  assign n84005 = ~n57783 ;
  assign n57785 = n57593 & n84005 ;
  assign n57903 = n57029 | n57593 ;
  assign n84006 = ~n57903 ;
  assign n57904 = n57589 & n84006 ;
  assign n57905 = n57785 | n57904 ;
  assign n57906 = n83972 & n57905 ;
  assign n57907 = n57020 & n83968 ;
  assign n57908 = n57818 & n57907 ;
  assign n57909 = n57906 | n57908 ;
  assign n57910 = n70927 & n57909 ;
  assign n84007 = ~n57584 ;
  assign n57588 = n84007 & n57587 ;
  assign n57911 = n57037 | n57587 ;
  assign n84008 = ~n57911 ;
  assign n57912 = n57779 & n84008 ;
  assign n57913 = n57588 | n57912 ;
  assign n57914 = n83972 & n57913 ;
  assign n57915 = n57028 & n83968 ;
  assign n57916 = n57818 & n57915 ;
  assign n57917 = n57914 | n57916 ;
  assign n57918 = n70609 & n57917 ;
  assign n84009 = ~n57916 ;
  assign n58471 = x107 & n84009 ;
  assign n84010 = ~n57914 ;
  assign n58472 = n84010 & n58471 ;
  assign n58473 = n57918 | n58472 ;
  assign n84011 = ~n57778 ;
  assign n57780 = n57582 & n84011 ;
  assign n57919 = n57045 | n57582 ;
  assign n84012 = ~n57919 ;
  assign n57920 = n57578 & n84012 ;
  assign n57921 = n57780 | n57920 ;
  assign n57922 = n83972 & n57921 ;
  assign n57923 = n57036 & n83968 ;
  assign n57924 = n57818 & n57923 ;
  assign n57925 = n57922 | n57924 ;
  assign n57926 = n70276 & n57925 ;
  assign n84013 = ~n57573 ;
  assign n57577 = n84013 & n57576 ;
  assign n57927 = n57053 | n57576 ;
  assign n84014 = ~n57927 ;
  assign n57928 = n57774 & n84014 ;
  assign n57929 = n57577 | n57928 ;
  assign n57930 = n83972 & n57929 ;
  assign n57931 = n57044 & n83968 ;
  assign n57932 = n57818 & n57931 ;
  assign n57933 = n57930 | n57932 ;
  assign n57934 = n70176 & n57933 ;
  assign n84015 = ~n57932 ;
  assign n58460 = x105 & n84015 ;
  assign n84016 = ~n57930 ;
  assign n58461 = n84016 & n58460 ;
  assign n58462 = n57934 | n58461 ;
  assign n84017 = ~n57773 ;
  assign n57775 = n57571 & n84017 ;
  assign n57935 = n57061 | n57571 ;
  assign n84018 = ~n57935 ;
  assign n57936 = n57567 & n84018 ;
  assign n57937 = n57775 | n57936 ;
  assign n57938 = n83972 & n57937 ;
  assign n57939 = n57052 & n83968 ;
  assign n57940 = n57818 & n57939 ;
  assign n57941 = n57938 | n57940 ;
  assign n57942 = n69857 & n57941 ;
  assign n84019 = ~n57562 ;
  assign n57566 = n84019 & n57565 ;
  assign n57943 = n57069 | n57565 ;
  assign n84020 = ~n57943 ;
  assign n57944 = n57769 & n84020 ;
  assign n57945 = n57566 | n57944 ;
  assign n57946 = n83972 & n57945 ;
  assign n57947 = n57060 & n83968 ;
  assign n57948 = n57818 & n57947 ;
  assign n57949 = n57946 | n57948 ;
  assign n57950 = n69656 & n57949 ;
  assign n84021 = ~n57948 ;
  assign n58450 = x103 & n84021 ;
  assign n84022 = ~n57946 ;
  assign n58451 = n84022 & n58450 ;
  assign n58452 = n57950 | n58451 ;
  assign n84023 = ~n57768 ;
  assign n57770 = n57560 & n84023 ;
  assign n57951 = n57077 | n57560 ;
  assign n84024 = ~n57951 ;
  assign n57952 = n57556 & n84024 ;
  assign n57953 = n57770 | n57952 ;
  assign n57954 = n83972 & n57953 ;
  assign n57955 = n57068 & n83968 ;
  assign n57956 = n57818 & n57955 ;
  assign n57957 = n57954 | n57956 ;
  assign n57958 = n69528 & n57957 ;
  assign n84025 = ~n57551 ;
  assign n57555 = n84025 & n57554 ;
  assign n57959 = n57085 | n57554 ;
  assign n84026 = ~n57959 ;
  assign n57960 = n57764 & n84026 ;
  assign n57961 = n57555 | n57960 ;
  assign n57962 = n83972 & n57961 ;
  assign n57963 = n57076 & n83968 ;
  assign n57964 = n57818 & n57963 ;
  assign n57965 = n57962 | n57964 ;
  assign n57966 = n69261 & n57965 ;
  assign n84027 = ~n57964 ;
  assign n58440 = x101 & n84027 ;
  assign n84028 = ~n57962 ;
  assign n58441 = n84028 & n58440 ;
  assign n58442 = n57966 | n58441 ;
  assign n84029 = ~n57763 ;
  assign n57765 = n57549 & n84029 ;
  assign n57967 = n57093 | n57549 ;
  assign n84030 = ~n57967 ;
  assign n57968 = n57545 & n84030 ;
  assign n57969 = n57765 | n57968 ;
  assign n57970 = n83972 & n57969 ;
  assign n57971 = n57084 & n83968 ;
  assign n57972 = n57818 & n57971 ;
  assign n57973 = n57970 | n57972 ;
  assign n57974 = n69075 & n57973 ;
  assign n84031 = ~n57540 ;
  assign n57544 = n84031 & n57543 ;
  assign n57975 = n57101 | n57543 ;
  assign n84032 = ~n57975 ;
  assign n57976 = n57759 & n84032 ;
  assign n57977 = n57544 | n57976 ;
  assign n57978 = n83972 & n57977 ;
  assign n57979 = n57092 & n83968 ;
  assign n57980 = n57818 & n57979 ;
  assign n57981 = n57978 | n57980 ;
  assign n57982 = n68993 & n57981 ;
  assign n84033 = ~n57980 ;
  assign n58429 = x99 & n84033 ;
  assign n84034 = ~n57978 ;
  assign n58430 = n84034 & n58429 ;
  assign n58431 = n57982 | n58430 ;
  assign n84035 = ~n57758 ;
  assign n57760 = n57538 & n84035 ;
  assign n57983 = n57109 | n57538 ;
  assign n84036 = ~n57983 ;
  assign n57984 = n57534 & n84036 ;
  assign n57985 = n57760 | n57984 ;
  assign n57986 = n83972 & n57985 ;
  assign n57987 = n57100 & n83968 ;
  assign n57988 = n57818 & n57987 ;
  assign n57989 = n57986 | n57988 ;
  assign n57990 = n68716 & n57989 ;
  assign n84037 = ~n57529 ;
  assign n57533 = n84037 & n57532 ;
  assign n57991 = n57117 | n57532 ;
  assign n84038 = ~n57991 ;
  assign n57992 = n57754 & n84038 ;
  assign n57993 = n57533 | n57992 ;
  assign n57994 = n83972 & n57993 ;
  assign n57995 = n57108 & n83968 ;
  assign n57996 = n57818 & n57995 ;
  assign n57997 = n57994 | n57996 ;
  assign n57998 = n68545 & n57997 ;
  assign n84039 = ~n57996 ;
  assign n58419 = x97 & n84039 ;
  assign n84040 = ~n57994 ;
  assign n58420 = n84040 & n58419 ;
  assign n58421 = n57998 | n58420 ;
  assign n84041 = ~n57753 ;
  assign n57755 = n57527 & n84041 ;
  assign n57999 = n57125 | n57527 ;
  assign n84042 = ~n57999 ;
  assign n58000 = n57523 & n84042 ;
  assign n58001 = n57755 | n58000 ;
  assign n58002 = n83972 & n58001 ;
  assign n58003 = n57116 & n83968 ;
  assign n58004 = n57818 & n58003 ;
  assign n58005 = n58002 | n58004 ;
  assign n58006 = n68438 & n58005 ;
  assign n84043 = ~n57518 ;
  assign n57522 = n84043 & n57521 ;
  assign n58007 = n57133 | n57521 ;
  assign n84044 = ~n58007 ;
  assign n58008 = n57749 & n84044 ;
  assign n58009 = n57522 | n58008 ;
  assign n58010 = n83972 & n58009 ;
  assign n58011 = n57124 & n83968 ;
  assign n58012 = n57818 & n58011 ;
  assign n58013 = n58010 | n58012 ;
  assign n58014 = n68214 & n58013 ;
  assign n84045 = ~n58012 ;
  assign n58409 = x95 & n84045 ;
  assign n84046 = ~n58010 ;
  assign n58410 = n84046 & n58409 ;
  assign n58411 = n58014 | n58410 ;
  assign n84047 = ~n57748 ;
  assign n57750 = n57516 & n84047 ;
  assign n58015 = n57141 | n57516 ;
  assign n84048 = ~n58015 ;
  assign n58016 = n57512 & n84048 ;
  assign n58017 = n57750 | n58016 ;
  assign n58018 = n83972 & n58017 ;
  assign n58019 = n57132 & n83968 ;
  assign n58020 = n57818 & n58019 ;
  assign n58021 = n58018 | n58020 ;
  assign n58022 = n68058 & n58021 ;
  assign n84049 = ~n57507 ;
  assign n57511 = n84049 & n57510 ;
  assign n58023 = n57149 | n57510 ;
  assign n84050 = ~n58023 ;
  assign n58024 = n57744 & n84050 ;
  assign n58025 = n57511 | n58024 ;
  assign n58026 = n83972 & n58025 ;
  assign n58027 = n57140 & n83968 ;
  assign n58028 = n57818 & n58027 ;
  assign n58029 = n58026 | n58028 ;
  assign n58030 = n67986 & n58029 ;
  assign n84051 = ~n58028 ;
  assign n58398 = x93 & n84051 ;
  assign n84052 = ~n58026 ;
  assign n58399 = n84052 & n58398 ;
  assign n58400 = n58030 | n58399 ;
  assign n84053 = ~n57743 ;
  assign n57745 = n57505 & n84053 ;
  assign n58031 = n57157 | n57505 ;
  assign n84054 = ~n58031 ;
  assign n58032 = n57501 & n84054 ;
  assign n58033 = n57745 | n58032 ;
  assign n58034 = n83972 & n58033 ;
  assign n58035 = n57148 & n83968 ;
  assign n58036 = n57818 & n58035 ;
  assign n58037 = n58034 | n58036 ;
  assign n58038 = n67763 & n58037 ;
  assign n84055 = ~n57496 ;
  assign n57500 = n84055 & n57499 ;
  assign n58039 = n57165 | n57499 ;
  assign n84056 = ~n58039 ;
  assign n58040 = n57739 & n84056 ;
  assign n58041 = n57500 | n58040 ;
  assign n58042 = n83972 & n58041 ;
  assign n58043 = n57156 & n83968 ;
  assign n58044 = n57818 & n58043 ;
  assign n58045 = n58042 | n58044 ;
  assign n58046 = n67622 & n58045 ;
  assign n84057 = ~n58044 ;
  assign n58388 = x91 & n84057 ;
  assign n84058 = ~n58042 ;
  assign n58389 = n84058 & n58388 ;
  assign n58390 = n58046 | n58389 ;
  assign n84059 = ~n57738 ;
  assign n57740 = n57494 & n84059 ;
  assign n58047 = n57173 | n57494 ;
  assign n84060 = ~n58047 ;
  assign n58048 = n57490 & n84060 ;
  assign n58049 = n57740 | n58048 ;
  assign n58050 = n83972 & n58049 ;
  assign n58051 = n57164 & n83968 ;
  assign n58052 = n57818 & n58051 ;
  assign n58053 = n58050 | n58052 ;
  assign n58054 = n67531 & n58053 ;
  assign n84061 = ~n57485 ;
  assign n57489 = n84061 & n57488 ;
  assign n58055 = n57181 | n57488 ;
  assign n84062 = ~n58055 ;
  assign n58056 = n57734 & n84062 ;
  assign n58057 = n57489 | n58056 ;
  assign n58058 = n83972 & n58057 ;
  assign n58059 = n57172 & n83968 ;
  assign n58060 = n57818 & n58059 ;
  assign n58061 = n58058 | n58060 ;
  assign n58062 = n67348 & n58061 ;
  assign n84063 = ~n58060 ;
  assign n58377 = x89 & n84063 ;
  assign n84064 = ~n58058 ;
  assign n58378 = n84064 & n58377 ;
  assign n58379 = n58062 | n58378 ;
  assign n84065 = ~n57733 ;
  assign n57735 = n57483 & n84065 ;
  assign n58063 = n57189 | n57483 ;
  assign n84066 = ~n58063 ;
  assign n58064 = n57479 & n84066 ;
  assign n58065 = n57735 | n58064 ;
  assign n58066 = n83972 & n58065 ;
  assign n58067 = n57180 & n83968 ;
  assign n58068 = n57818 & n58067 ;
  assign n58069 = n58066 | n58068 ;
  assign n58070 = n67222 & n58069 ;
  assign n84067 = ~n57474 ;
  assign n57478 = n84067 & n57477 ;
  assign n58071 = n57197 | n57477 ;
  assign n84068 = ~n58071 ;
  assign n58072 = n57729 & n84068 ;
  assign n58073 = n57478 | n58072 ;
  assign n58074 = n83972 & n58073 ;
  assign n58075 = n57188 & n83968 ;
  assign n58076 = n57818 & n58075 ;
  assign n58077 = n58074 | n58076 ;
  assign n58078 = n67164 & n58077 ;
  assign n84069 = ~n58076 ;
  assign n58367 = x87 & n84069 ;
  assign n84070 = ~n58074 ;
  assign n58368 = n84070 & n58367 ;
  assign n58369 = n58078 | n58368 ;
  assign n84071 = ~n57728 ;
  assign n57730 = n57472 & n84071 ;
  assign n58079 = n57205 | n57472 ;
  assign n84072 = ~n58079 ;
  assign n58080 = n57468 & n84072 ;
  assign n58081 = n57730 | n58080 ;
  assign n58082 = n83972 & n58081 ;
  assign n58083 = n57196 & n83968 ;
  assign n58084 = n57818 & n58083 ;
  assign n58085 = n58082 | n58084 ;
  assign n58086 = n66979 & n58085 ;
  assign n84073 = ~n57463 ;
  assign n57467 = n84073 & n57466 ;
  assign n58087 = n57213 | n57466 ;
  assign n84074 = ~n58087 ;
  assign n58088 = n57724 & n84074 ;
  assign n58089 = n57467 | n58088 ;
  assign n58090 = n83972 & n58089 ;
  assign n58091 = n57204 & n83968 ;
  assign n58092 = n57818 & n58091 ;
  assign n58093 = n58090 | n58092 ;
  assign n58094 = n66868 & n58093 ;
  assign n84075 = ~n58092 ;
  assign n58357 = x85 & n84075 ;
  assign n84076 = ~n58090 ;
  assign n58358 = n84076 & n58357 ;
  assign n58359 = n58094 | n58358 ;
  assign n84077 = ~n57723 ;
  assign n57725 = n57461 & n84077 ;
  assign n58095 = n57221 | n57461 ;
  assign n84078 = ~n58095 ;
  assign n58096 = n57457 & n84078 ;
  assign n58097 = n57725 | n58096 ;
  assign n58098 = n83972 & n58097 ;
  assign n58099 = n57212 & n83968 ;
  assign n58100 = n57818 & n58099 ;
  assign n58101 = n58098 | n58100 ;
  assign n58102 = n66797 & n58101 ;
  assign n84079 = ~n57452 ;
  assign n57456 = n84079 & n57455 ;
  assign n58103 = n57229 | n57455 ;
  assign n84080 = ~n58103 ;
  assign n58104 = n57719 & n84080 ;
  assign n58105 = n57456 | n58104 ;
  assign n58106 = n83972 & n58105 ;
  assign n58107 = n57220 & n83968 ;
  assign n58108 = n57818 & n58107 ;
  assign n58109 = n58106 | n58108 ;
  assign n58110 = n66654 & n58109 ;
  assign n84081 = ~n58108 ;
  assign n58347 = x83 & n84081 ;
  assign n84082 = ~n58106 ;
  assign n58348 = n84082 & n58347 ;
  assign n58349 = n58110 | n58348 ;
  assign n84083 = ~n57718 ;
  assign n57720 = n57450 & n84083 ;
  assign n58111 = n57237 | n57450 ;
  assign n84084 = ~n58111 ;
  assign n58112 = n57446 & n84084 ;
  assign n58113 = n57720 | n58112 ;
  assign n58114 = n83972 & n58113 ;
  assign n58115 = n57228 & n83968 ;
  assign n58116 = n57818 & n58115 ;
  assign n58117 = n58114 | n58116 ;
  assign n58118 = n66560 & n58117 ;
  assign n84085 = ~n57441 ;
  assign n57445 = n84085 & n57444 ;
  assign n58119 = n57245 | n57444 ;
  assign n84086 = ~n58119 ;
  assign n58120 = n57714 & n84086 ;
  assign n58121 = n57445 | n58120 ;
  assign n58122 = n83972 & n58121 ;
  assign n58123 = n57236 & n83968 ;
  assign n58124 = n57818 & n58123 ;
  assign n58125 = n58122 | n58124 ;
  assign n58126 = n66505 & n58125 ;
  assign n84087 = ~n58124 ;
  assign n58337 = x81 & n84087 ;
  assign n84088 = ~n58122 ;
  assign n58338 = n84088 & n58337 ;
  assign n58339 = n58126 | n58338 ;
  assign n84089 = ~n57713 ;
  assign n57715 = n57439 & n84089 ;
  assign n58127 = n57253 | n57439 ;
  assign n84090 = ~n58127 ;
  assign n58128 = n57435 & n84090 ;
  assign n58129 = n57715 | n58128 ;
  assign n58130 = n83972 & n58129 ;
  assign n58131 = n57244 & n83968 ;
  assign n58132 = n57818 & n58131 ;
  assign n58133 = n58130 | n58132 ;
  assign n58134 = n66379 & n58133 ;
  assign n84091 = ~n57430 ;
  assign n57434 = n84091 & n57433 ;
  assign n58135 = n57261 | n57433 ;
  assign n84092 = ~n58135 ;
  assign n58136 = n57709 & n84092 ;
  assign n58137 = n57434 | n58136 ;
  assign n58138 = n83972 & n58137 ;
  assign n58139 = n57252 & n83968 ;
  assign n58140 = n57818 & n58139 ;
  assign n58141 = n58138 | n58140 ;
  assign n58142 = n66299 & n58141 ;
  assign n84093 = ~n58140 ;
  assign n58327 = x79 & n84093 ;
  assign n84094 = ~n58138 ;
  assign n58328 = n84094 & n58327 ;
  assign n58329 = n58142 | n58328 ;
  assign n84095 = ~n57708 ;
  assign n57710 = n57428 & n84095 ;
  assign n58143 = n57269 | n57428 ;
  assign n84096 = ~n58143 ;
  assign n58144 = n57424 & n84096 ;
  assign n58145 = n57710 | n58144 ;
  assign n58146 = n83972 & n58145 ;
  assign n58147 = n57260 & n83968 ;
  assign n58148 = n57818 & n58147 ;
  assign n58149 = n58146 | n58148 ;
  assign n58150 = n66244 & n58149 ;
  assign n84097 = ~n57419 ;
  assign n57423 = n84097 & n57422 ;
  assign n58151 = n57277 | n57422 ;
  assign n84098 = ~n58151 ;
  assign n58152 = n57704 & n84098 ;
  assign n58153 = n57423 | n58152 ;
  assign n58154 = n83972 & n58153 ;
  assign n58155 = n57268 & n83968 ;
  assign n58156 = n57818 & n58155 ;
  assign n58157 = n58154 | n58156 ;
  assign n58158 = n66145 & n58157 ;
  assign n84099 = ~n58156 ;
  assign n58317 = x77 & n84099 ;
  assign n84100 = ~n58154 ;
  assign n58318 = n84100 & n58317 ;
  assign n58319 = n58158 | n58318 ;
  assign n84101 = ~n57703 ;
  assign n57705 = n57417 & n84101 ;
  assign n58159 = n57285 | n57417 ;
  assign n84102 = ~n58159 ;
  assign n58160 = n57413 & n84102 ;
  assign n58161 = n57705 | n58160 ;
  assign n58162 = n83972 & n58161 ;
  assign n58163 = n57276 & n83968 ;
  assign n58164 = n57818 & n58163 ;
  assign n58165 = n58162 | n58164 ;
  assign n58166 = n66081 & n58165 ;
  assign n84103 = ~n57408 ;
  assign n57412 = n84103 & n57411 ;
  assign n58167 = n57293 | n57411 ;
  assign n84104 = ~n58167 ;
  assign n58168 = n57699 & n84104 ;
  assign n58169 = n57412 | n58168 ;
  assign n58170 = n83972 & n58169 ;
  assign n58171 = n57284 & n83968 ;
  assign n58172 = n57818 & n58171 ;
  assign n58173 = n58170 | n58172 ;
  assign n58174 = n66043 & n58173 ;
  assign n84105 = ~n58172 ;
  assign n58307 = x75 & n84105 ;
  assign n84106 = ~n58170 ;
  assign n58308 = n84106 & n58307 ;
  assign n58309 = n58174 | n58308 ;
  assign n84107 = ~n57698 ;
  assign n57700 = n57406 & n84107 ;
  assign n58175 = n57301 | n57406 ;
  assign n84108 = ~n58175 ;
  assign n58176 = n57402 & n84108 ;
  assign n58177 = n57700 | n58176 ;
  assign n58178 = n83972 & n58177 ;
  assign n58179 = n57292 & n83968 ;
  assign n58180 = n57818 & n58179 ;
  assign n58181 = n58178 | n58180 ;
  assign n58182 = n65960 & n58181 ;
  assign n84109 = ~n57397 ;
  assign n57401 = n84109 & n57400 ;
  assign n58183 = n57309 | n57400 ;
  assign n84110 = ~n58183 ;
  assign n58184 = n57694 & n84110 ;
  assign n58185 = n57401 | n58184 ;
  assign n58186 = n83972 & n58185 ;
  assign n58187 = n57300 & n83968 ;
  assign n58188 = n57818 & n58187 ;
  assign n58189 = n58186 | n58188 ;
  assign n58190 = n65909 & n58189 ;
  assign n84111 = ~n58188 ;
  assign n58297 = x73 & n84111 ;
  assign n84112 = ~n58186 ;
  assign n58298 = n84112 & n58297 ;
  assign n58299 = n58190 | n58298 ;
  assign n84113 = ~n57693 ;
  assign n57695 = n57395 & n84113 ;
  assign n58191 = n57317 | n57395 ;
  assign n84114 = ~n58191 ;
  assign n58192 = n57391 & n84114 ;
  assign n58193 = n57695 | n58192 ;
  assign n58194 = n83972 & n58193 ;
  assign n58195 = n57308 & n83968 ;
  assign n58196 = n57818 & n58195 ;
  assign n58197 = n58194 | n58196 ;
  assign n58198 = n65877 & n58197 ;
  assign n84115 = ~n57386 ;
  assign n57390 = n84115 & n57389 ;
  assign n58199 = n57326 | n57389 ;
  assign n84116 = ~n58199 ;
  assign n58200 = n57690 & n84116 ;
  assign n58201 = n57390 | n58200 ;
  assign n58202 = n83972 & n58201 ;
  assign n58203 = n57316 & n83968 ;
  assign n58204 = n57818 & n58203 ;
  assign n58205 = n58202 | n58204 ;
  assign n58206 = n65820 & n58205 ;
  assign n84117 = ~n58204 ;
  assign n58287 = x71 & n84117 ;
  assign n84118 = ~n58202 ;
  assign n58288 = n84118 & n58287 ;
  assign n58289 = n58206 | n58288 ;
  assign n84119 = ~n57688 ;
  assign n57689 = n57384 & n84119 ;
  assign n58207 = n57335 | n57384 ;
  assign n84120 = ~n58207 ;
  assign n58208 = n57380 & n84120 ;
  assign n58209 = n57689 | n58208 ;
  assign n58210 = n83972 & n58209 ;
  assign n58211 = n57325 & n83968 ;
  assign n58212 = n57818 & n58211 ;
  assign n58213 = n58210 | n58212 ;
  assign n58214 = n65791 & n58213 ;
  assign n84121 = ~n57376 ;
  assign n57686 = n84121 & n57379 ;
  assign n58215 = n57374 | n57682 ;
  assign n58216 = n57343 | n57379 ;
  assign n84122 = ~n58216 ;
  assign n58217 = n58215 & n84122 ;
  assign n58218 = n57686 | n58217 ;
  assign n58219 = n83972 & n58218 ;
  assign n58220 = n57334 & n83968 ;
  assign n58221 = n57818 & n58220 ;
  assign n58222 = n58219 | n58221 ;
  assign n58223 = n65772 & n58222 ;
  assign n84123 = ~n58221 ;
  assign n58276 = x69 & n84123 ;
  assign n84124 = ~n58219 ;
  assign n58277 = n84124 & n58276 ;
  assign n58278 = n58223 | n58277 ;
  assign n84125 = ~n57682 ;
  assign n57684 = n57374 & n84125 ;
  assign n58224 = n57349 | n57374 ;
  assign n84126 = ~n58224 ;
  assign n58225 = n57681 & n84126 ;
  assign n58226 = n57684 | n58225 ;
  assign n58227 = n83972 & n58226 ;
  assign n58228 = n57342 & n83968 ;
  assign n58229 = n57818 & n58228 ;
  assign n58230 = n58227 | n58229 ;
  assign n58231 = n65746 & n58230 ;
  assign n84127 = ~n57367 ;
  assign n57680 = n84127 & n57679 ;
  assign n58232 = n57365 | n57679 ;
  assign n84128 = ~n58232 ;
  assign n58233 = n57366 & n84128 ;
  assign n58234 = n57680 | n58233 ;
  assign n58235 = n83972 & n58234 ;
  assign n58236 = n57348 & n83968 ;
  assign n58237 = n57818 & n58236 ;
  assign n58238 = n58235 | n58237 ;
  assign n58239 = n65721 & n58238 ;
  assign n84129 = ~n58237 ;
  assign n58266 = x67 & n84129 ;
  assign n84130 = ~n58235 ;
  assign n58267 = n84130 & n58266 ;
  assign n58268 = n58239 | n58267 ;
  assign n58240 = n25157 & n57363 ;
  assign n58241 = n83970 & n58240 ;
  assign n84131 = ~n58241 ;
  assign n58242 = n57366 & n84131 ;
  assign n58243 = n83972 & n58242 ;
  assign n58244 = n57360 & n83968 ;
  assign n58245 = n57818 & n58244 ;
  assign n58246 = n58243 | n58245 ;
  assign n58247 = n65686 & n58246 ;
  assign n57674 = n25157 & n83972 ;
  assign n58248 = n83968 & n57818 ;
  assign n84132 = ~n58248 ;
  assign n58249 = x64 & n84132 ;
  assign n84133 = ~n58249 ;
  assign n58250 = x8 & n84133 ;
  assign n58251 = n57674 | n58250 ;
  assign n58252 = x65 & n58251 ;
  assign n57673 = x64 & n83972 ;
  assign n84134 = ~n57673 ;
  assign n58253 = x8 & n84134 ;
  assign n58254 = n25157 & n84132 ;
  assign n58255 = x65 | n58254 ;
  assign n58256 = n58253 | n58255 ;
  assign n84135 = ~n58252 ;
  assign n58257 = n84135 & n58256 ;
  assign n58258 = n26052 | n58257 ;
  assign n58259 = n57674 | n58253 ;
  assign n58260 = n65670 & n58259 ;
  assign n84136 = ~n58260 ;
  assign n58261 = n58258 & n84136 ;
  assign n84137 = ~n58245 ;
  assign n58262 = x66 & n84137 ;
  assign n84138 = ~n58243 ;
  assign n58263 = n84138 & n58262 ;
  assign n58264 = n58247 | n58263 ;
  assign n58265 = n58261 | n58264 ;
  assign n84139 = ~n58247 ;
  assign n58269 = n84139 & n58265 ;
  assign n58270 = n58268 | n58269 ;
  assign n84140 = ~n58239 ;
  assign n58271 = n84140 & n58270 ;
  assign n84141 = ~n58229 ;
  assign n58272 = x68 & n84141 ;
  assign n84142 = ~n58227 ;
  assign n58273 = n84142 & n58272 ;
  assign n58274 = n58231 | n58273 ;
  assign n58275 = n58271 | n58274 ;
  assign n84143 = ~n58231 ;
  assign n58279 = n84143 & n58275 ;
  assign n58280 = n58278 | n58279 ;
  assign n84144 = ~n58223 ;
  assign n58281 = n84144 & n58280 ;
  assign n84145 = ~n58212 ;
  assign n58282 = x70 & n84145 ;
  assign n84146 = ~n58210 ;
  assign n58283 = n84146 & n58282 ;
  assign n58284 = n58214 | n58283 ;
  assign n58286 = n58281 | n58284 ;
  assign n84147 = ~n58214 ;
  assign n58290 = n84147 & n58286 ;
  assign n58291 = n58289 | n58290 ;
  assign n84148 = ~n58206 ;
  assign n58292 = n84148 & n58291 ;
  assign n84149 = ~n58196 ;
  assign n58293 = x72 & n84149 ;
  assign n84150 = ~n58194 ;
  assign n58294 = n84150 & n58293 ;
  assign n58295 = n58198 | n58294 ;
  assign n58296 = n58292 | n58295 ;
  assign n84151 = ~n58198 ;
  assign n58300 = n84151 & n58296 ;
  assign n58301 = n58299 | n58300 ;
  assign n84152 = ~n58190 ;
  assign n58302 = n84152 & n58301 ;
  assign n84153 = ~n58180 ;
  assign n58303 = x74 & n84153 ;
  assign n84154 = ~n58178 ;
  assign n58304 = n84154 & n58303 ;
  assign n58305 = n58182 | n58304 ;
  assign n58306 = n58302 | n58305 ;
  assign n84155 = ~n58182 ;
  assign n58310 = n84155 & n58306 ;
  assign n58311 = n58309 | n58310 ;
  assign n84156 = ~n58174 ;
  assign n58312 = n84156 & n58311 ;
  assign n84157 = ~n58164 ;
  assign n58313 = x76 & n84157 ;
  assign n84158 = ~n58162 ;
  assign n58314 = n84158 & n58313 ;
  assign n58315 = n58166 | n58314 ;
  assign n58316 = n58312 | n58315 ;
  assign n84159 = ~n58166 ;
  assign n58320 = n84159 & n58316 ;
  assign n58321 = n58319 | n58320 ;
  assign n84160 = ~n58158 ;
  assign n58322 = n84160 & n58321 ;
  assign n84161 = ~n58148 ;
  assign n58323 = x78 & n84161 ;
  assign n84162 = ~n58146 ;
  assign n58324 = n84162 & n58323 ;
  assign n58325 = n58150 | n58324 ;
  assign n58326 = n58322 | n58325 ;
  assign n84163 = ~n58150 ;
  assign n58330 = n84163 & n58326 ;
  assign n58331 = n58329 | n58330 ;
  assign n84164 = ~n58142 ;
  assign n58332 = n84164 & n58331 ;
  assign n84165 = ~n58132 ;
  assign n58333 = x80 & n84165 ;
  assign n84166 = ~n58130 ;
  assign n58334 = n84166 & n58333 ;
  assign n58335 = n58134 | n58334 ;
  assign n58336 = n58332 | n58335 ;
  assign n84167 = ~n58134 ;
  assign n58340 = n84167 & n58336 ;
  assign n58341 = n58339 | n58340 ;
  assign n84168 = ~n58126 ;
  assign n58342 = n84168 & n58341 ;
  assign n84169 = ~n58116 ;
  assign n58343 = x82 & n84169 ;
  assign n84170 = ~n58114 ;
  assign n58344 = n84170 & n58343 ;
  assign n58345 = n58118 | n58344 ;
  assign n58346 = n58342 | n58345 ;
  assign n84171 = ~n58118 ;
  assign n58350 = n84171 & n58346 ;
  assign n58351 = n58349 | n58350 ;
  assign n84172 = ~n58110 ;
  assign n58352 = n84172 & n58351 ;
  assign n84173 = ~n58100 ;
  assign n58353 = x84 & n84173 ;
  assign n84174 = ~n58098 ;
  assign n58354 = n84174 & n58353 ;
  assign n58355 = n58102 | n58354 ;
  assign n58356 = n58352 | n58355 ;
  assign n84175 = ~n58102 ;
  assign n58360 = n84175 & n58356 ;
  assign n58361 = n58359 | n58360 ;
  assign n84176 = ~n58094 ;
  assign n58362 = n84176 & n58361 ;
  assign n84177 = ~n58084 ;
  assign n58363 = x86 & n84177 ;
  assign n84178 = ~n58082 ;
  assign n58364 = n84178 & n58363 ;
  assign n58365 = n58086 | n58364 ;
  assign n58366 = n58362 | n58365 ;
  assign n84179 = ~n58086 ;
  assign n58370 = n84179 & n58366 ;
  assign n58371 = n58369 | n58370 ;
  assign n84180 = ~n58078 ;
  assign n58372 = n84180 & n58371 ;
  assign n84181 = ~n58068 ;
  assign n58373 = x88 & n84181 ;
  assign n84182 = ~n58066 ;
  assign n58374 = n84182 & n58373 ;
  assign n58375 = n58070 | n58374 ;
  assign n58376 = n58372 | n58375 ;
  assign n84183 = ~n58070 ;
  assign n58381 = n84183 & n58376 ;
  assign n58382 = n58379 | n58381 ;
  assign n84184 = ~n58062 ;
  assign n58383 = n84184 & n58382 ;
  assign n84185 = ~n58052 ;
  assign n58384 = x90 & n84185 ;
  assign n84186 = ~n58050 ;
  assign n58385 = n84186 & n58384 ;
  assign n58386 = n58054 | n58385 ;
  assign n58387 = n58383 | n58386 ;
  assign n84187 = ~n58054 ;
  assign n58391 = n84187 & n58387 ;
  assign n58392 = n58390 | n58391 ;
  assign n84188 = ~n58046 ;
  assign n58393 = n84188 & n58392 ;
  assign n84189 = ~n58036 ;
  assign n58394 = x92 & n84189 ;
  assign n84190 = ~n58034 ;
  assign n58395 = n84190 & n58394 ;
  assign n58396 = n58038 | n58395 ;
  assign n58397 = n58393 | n58396 ;
  assign n84191 = ~n58038 ;
  assign n58401 = n84191 & n58397 ;
  assign n58402 = n58400 | n58401 ;
  assign n84192 = ~n58030 ;
  assign n58403 = n84192 & n58402 ;
  assign n84193 = ~n58020 ;
  assign n58404 = x94 & n84193 ;
  assign n84194 = ~n58018 ;
  assign n58405 = n84194 & n58404 ;
  assign n58406 = n58022 | n58405 ;
  assign n58408 = n58403 | n58406 ;
  assign n84195 = ~n58022 ;
  assign n58412 = n84195 & n58408 ;
  assign n58413 = n58411 | n58412 ;
  assign n84196 = ~n58014 ;
  assign n58414 = n84196 & n58413 ;
  assign n84197 = ~n58004 ;
  assign n58415 = x96 & n84197 ;
  assign n84198 = ~n58002 ;
  assign n58416 = n84198 & n58415 ;
  assign n58417 = n58006 | n58416 ;
  assign n58418 = n58414 | n58417 ;
  assign n84199 = ~n58006 ;
  assign n58422 = n84199 & n58418 ;
  assign n58423 = n58421 | n58422 ;
  assign n84200 = ~n57998 ;
  assign n58424 = n84200 & n58423 ;
  assign n84201 = ~n57988 ;
  assign n58425 = x98 & n84201 ;
  assign n84202 = ~n57986 ;
  assign n58426 = n84202 & n58425 ;
  assign n58427 = n57990 | n58426 ;
  assign n58428 = n58424 | n58427 ;
  assign n84203 = ~n57990 ;
  assign n58433 = n84203 & n58428 ;
  assign n58434 = n58431 | n58433 ;
  assign n84204 = ~n57982 ;
  assign n58435 = n84204 & n58434 ;
  assign n84205 = ~n57972 ;
  assign n58436 = x100 & n84205 ;
  assign n84206 = ~n57970 ;
  assign n58437 = n84206 & n58436 ;
  assign n58438 = n57974 | n58437 ;
  assign n58439 = n58435 | n58438 ;
  assign n84207 = ~n57974 ;
  assign n58443 = n84207 & n58439 ;
  assign n58444 = n58442 | n58443 ;
  assign n84208 = ~n57966 ;
  assign n58445 = n84208 & n58444 ;
  assign n84209 = ~n57956 ;
  assign n58446 = x102 & n84209 ;
  assign n84210 = ~n57954 ;
  assign n58447 = n84210 & n58446 ;
  assign n58448 = n57958 | n58447 ;
  assign n58449 = n58445 | n58448 ;
  assign n84211 = ~n57958 ;
  assign n58453 = n84211 & n58449 ;
  assign n58454 = n58452 | n58453 ;
  assign n84212 = ~n57950 ;
  assign n58455 = n84212 & n58454 ;
  assign n84213 = ~n57940 ;
  assign n58456 = x104 & n84213 ;
  assign n84214 = ~n57938 ;
  assign n58457 = n84214 & n58456 ;
  assign n58458 = n57942 | n58457 ;
  assign n58459 = n58455 | n58458 ;
  assign n84215 = ~n57942 ;
  assign n58463 = n84215 & n58459 ;
  assign n58464 = n58462 | n58463 ;
  assign n84216 = ~n57934 ;
  assign n58465 = n84216 & n58464 ;
  assign n84217 = ~n57924 ;
  assign n58466 = x106 & n84217 ;
  assign n84218 = ~n57922 ;
  assign n58467 = n84218 & n58466 ;
  assign n58468 = n57926 | n58467 ;
  assign n58470 = n58465 | n58468 ;
  assign n84219 = ~n57926 ;
  assign n58474 = n84219 & n58470 ;
  assign n58475 = n58473 | n58474 ;
  assign n84220 = ~n57918 ;
  assign n58476 = n84220 & n58475 ;
  assign n84221 = ~n57908 ;
  assign n58477 = x108 & n84221 ;
  assign n84222 = ~n57906 ;
  assign n58478 = n84222 & n58477 ;
  assign n58479 = n57910 | n58478 ;
  assign n58480 = n58476 | n58479 ;
  assign n84223 = ~n57910 ;
  assign n58484 = n84223 & n58480 ;
  assign n58485 = n58483 | n58484 ;
  assign n84224 = ~n57902 ;
  assign n58486 = n84224 & n58485 ;
  assign n84225 = ~n57892 ;
  assign n58487 = x110 & n84225 ;
  assign n84226 = ~n57890 ;
  assign n58488 = n84226 & n58487 ;
  assign n58489 = n57894 | n58488 ;
  assign n58490 = n58486 | n58489 ;
  assign n84227 = ~n57894 ;
  assign n58494 = n84227 & n58490 ;
  assign n58495 = n58493 | n58494 ;
  assign n84228 = ~n57886 ;
  assign n58496 = n84228 & n58495 ;
  assign n84229 = ~n57876 ;
  assign n58497 = x112 & n84229 ;
  assign n84230 = ~n57874 ;
  assign n58498 = n84230 & n58497 ;
  assign n58499 = n57878 | n58498 ;
  assign n58500 = n58496 | n58499 ;
  assign n84231 = ~n57878 ;
  assign n58504 = n84231 & n58500 ;
  assign n58505 = n58503 | n58504 ;
  assign n84232 = ~n57870 ;
  assign n58506 = n84232 & n58505 ;
  assign n84233 = ~n57860 ;
  assign n58507 = x114 & n84233 ;
  assign n84234 = ~n57858 ;
  assign n58508 = n84234 & n58507 ;
  assign n58509 = n57862 | n58508 ;
  assign n58510 = n58506 | n58509 ;
  assign n84235 = ~n57862 ;
  assign n58514 = n84235 & n58510 ;
  assign n58515 = n58513 | n58514 ;
  assign n84236 = ~n57854 ;
  assign n58516 = n84236 & n58515 ;
  assign n84237 = ~n57844 ;
  assign n58517 = x116 & n84237 ;
  assign n84238 = ~n57842 ;
  assign n58518 = n84238 & n58517 ;
  assign n58519 = n57846 | n58518 ;
  assign n58520 = n58516 | n58519 ;
  assign n84239 = ~n57846 ;
  assign n58524 = n84239 & n58520 ;
  assign n58525 = n58523 | n58524 ;
  assign n84240 = ~n57838 ;
  assign n58526 = n84240 & n58525 ;
  assign n84241 = ~n57828 ;
  assign n58527 = x118 & n84241 ;
  assign n84242 = ~n57826 ;
  assign n58528 = n84242 & n58527 ;
  assign n58529 = n57830 | n58528 ;
  assign n58530 = n58526 | n58529 ;
  assign n84243 = ~n57830 ;
  assign n58534 = n84243 & n58530 ;
  assign n58535 = n58533 | n58534 ;
  assign n84244 = ~n57822 ;
  assign n58536 = n84244 & n58535 ;
  assign n58537 = n56933 | n57667 ;
  assign n58538 = n57663 | n58537 ;
  assign n84245 = ~n58538 ;
  assign n58539 = n57655 & n84245 ;
  assign n58540 = n57663 | n57667 ;
  assign n84246 = ~n57817 ;
  assign n58541 = n84246 & n58540 ;
  assign n58542 = n58539 | n58541 ;
  assign n58543 = n83972 & n58542 ;
  assign n58544 = n24576 & n56075 ;
  assign n58545 = n57818 & n58544 ;
  assign n58546 = n58543 | n58545 ;
  assign n58547 = n74021 & n58546 ;
  assign n84247 = ~n58545 ;
  assign n58548 = x120 & n84247 ;
  assign n84248 = ~n58543 ;
  assign n58549 = n84248 & n58548 ;
  assign n58550 = n278 | n58549 ;
  assign n58551 = n58547 | n58550 ;
  assign n58552 = n58536 | n58551 ;
  assign n58553 = n65681 & n58546 ;
  assign n84249 = ~n58553 ;
  assign n58554 = n58552 & n84249 ;
  assign n84250 = ~n58534 ;
  assign n58666 = n58533 & n84250 ;
  assign n58555 = x65 & n58259 ;
  assign n84251 = ~n58555 ;
  assign n58556 = n58256 & n84251 ;
  assign n58557 = n26052 | n58556 ;
  assign n58559 = n84136 & n58557 ;
  assign n58560 = n58264 | n58559 ;
  assign n58561 = n84139 & n58560 ;
  assign n58562 = n58268 | n58561 ;
  assign n58563 = n84140 & n58562 ;
  assign n58564 = n58274 | n58563 ;
  assign n58565 = n84143 & n58564 ;
  assign n58566 = n58278 | n58565 ;
  assign n58567 = n84144 & n58566 ;
  assign n58568 = n58284 | n58567 ;
  assign n58569 = n84147 & n58568 ;
  assign n58570 = n58289 | n58569 ;
  assign n58571 = n84148 & n58570 ;
  assign n58572 = n58295 | n58571 ;
  assign n58573 = n84151 & n58572 ;
  assign n58574 = n58299 | n58573 ;
  assign n58575 = n84152 & n58574 ;
  assign n58576 = n58305 | n58575 ;
  assign n58577 = n84155 & n58576 ;
  assign n58578 = n58309 | n58577 ;
  assign n58579 = n84156 & n58578 ;
  assign n58580 = n58315 | n58579 ;
  assign n58581 = n84159 & n58580 ;
  assign n58582 = n58319 | n58581 ;
  assign n58583 = n84160 & n58582 ;
  assign n58584 = n58325 | n58583 ;
  assign n58585 = n84163 & n58584 ;
  assign n58586 = n58329 | n58585 ;
  assign n58587 = n84164 & n58586 ;
  assign n58588 = n58335 | n58587 ;
  assign n58589 = n84167 & n58588 ;
  assign n58590 = n58339 | n58589 ;
  assign n58591 = n84168 & n58590 ;
  assign n58592 = n58345 | n58591 ;
  assign n58593 = n84171 & n58592 ;
  assign n58594 = n58349 | n58593 ;
  assign n58595 = n84172 & n58594 ;
  assign n58596 = n58355 | n58595 ;
  assign n58597 = n84175 & n58596 ;
  assign n58598 = n58359 | n58597 ;
  assign n58599 = n84176 & n58598 ;
  assign n58600 = n58365 | n58599 ;
  assign n58601 = n84179 & n58600 ;
  assign n58602 = n58369 | n58601 ;
  assign n58603 = n84180 & n58602 ;
  assign n58604 = n58375 | n58603 ;
  assign n58605 = n84183 & n58604 ;
  assign n58606 = n58379 | n58605 ;
  assign n58607 = n84184 & n58606 ;
  assign n58608 = n58386 | n58607 ;
  assign n58609 = n84187 & n58608 ;
  assign n58610 = n58390 | n58609 ;
  assign n58611 = n84188 & n58610 ;
  assign n58612 = n58396 | n58611 ;
  assign n58613 = n84191 & n58612 ;
  assign n58614 = n58400 | n58613 ;
  assign n58615 = n84192 & n58614 ;
  assign n58616 = n58406 | n58615 ;
  assign n58617 = n84195 & n58616 ;
  assign n58618 = n58411 | n58617 ;
  assign n58619 = n84196 & n58618 ;
  assign n58620 = n58417 | n58619 ;
  assign n58621 = n84199 & n58620 ;
  assign n58622 = n58421 | n58621 ;
  assign n58623 = n84200 & n58622 ;
  assign n58624 = n58427 | n58623 ;
  assign n58625 = n84203 & n58624 ;
  assign n58626 = n58431 | n58625 ;
  assign n58627 = n84204 & n58626 ;
  assign n58628 = n58438 | n58627 ;
  assign n58629 = n84207 & n58628 ;
  assign n58630 = n58442 | n58629 ;
  assign n58631 = n84208 & n58630 ;
  assign n58632 = n58448 | n58631 ;
  assign n58633 = n84211 & n58632 ;
  assign n58634 = n58452 | n58633 ;
  assign n58635 = n84212 & n58634 ;
  assign n58636 = n58458 | n58635 ;
  assign n58637 = n84215 & n58636 ;
  assign n58638 = n58462 | n58637 ;
  assign n58639 = n84216 & n58638 ;
  assign n58640 = n58468 | n58639 ;
  assign n58641 = n84219 & n58640 ;
  assign n58642 = n58473 | n58641 ;
  assign n58643 = n84220 & n58642 ;
  assign n58644 = n58479 | n58643 ;
  assign n58645 = n84223 & n58644 ;
  assign n58646 = n58483 | n58645 ;
  assign n58647 = n84224 & n58646 ;
  assign n58648 = n58489 | n58647 ;
  assign n58649 = n84227 & n58648 ;
  assign n58650 = n58493 | n58649 ;
  assign n58651 = n84228 & n58650 ;
  assign n58652 = n58499 | n58651 ;
  assign n58653 = n84231 & n58652 ;
  assign n58654 = n58503 | n58653 ;
  assign n58655 = n84232 & n58654 ;
  assign n58656 = n58509 | n58655 ;
  assign n58657 = n84235 & n58656 ;
  assign n58658 = n58513 | n58657 ;
  assign n58659 = n84236 & n58658 ;
  assign n58660 = n58519 | n58659 ;
  assign n58661 = n84239 & n58660 ;
  assign n58662 = n58523 | n58661 ;
  assign n58663 = n84240 & n58662 ;
  assign n58664 = n58529 | n58663 ;
  assign n58667 = n57830 | n58533 ;
  assign n84252 = ~n58667 ;
  assign n58668 = n58664 & n84252 ;
  assign n58669 = n58666 | n58668 ;
  assign n84253 = ~n58554 ;
  assign n58670 = n84253 & n58669 ;
  assign n58671 = n57821 & n84249 ;
  assign n58672 = n58552 & n58671 ;
  assign n58673 = n58670 | n58672 ;
  assign n58674 = n57822 | n58549 ;
  assign n58675 = n58547 | n58674 ;
  assign n84254 = ~n58675 ;
  assign n58676 = n58535 & n84254 ;
  assign n58665 = n84243 & n58664 ;
  assign n58677 = n58533 | n58665 ;
  assign n58678 = n84244 & n58677 ;
  assign n58679 = n58547 | n58549 ;
  assign n84255 = ~n58678 ;
  assign n58680 = n84255 & n58679 ;
  assign n58681 = n58676 | n58680 ;
  assign n58682 = n84253 & n58681 ;
  assign n58683 = n66655 & n58546 ;
  assign n58684 = n58552 & n58683 ;
  assign n58685 = n58682 | n58684 ;
  assign n58686 = n74029 & n58685 ;
  assign n58687 = n74021 & n58673 ;
  assign n84256 = ~n58663 ;
  assign n58688 = n58529 & n84256 ;
  assign n58689 = n57838 | n58529 ;
  assign n84257 = ~n58689 ;
  assign n58690 = n58525 & n84257 ;
  assign n58691 = n58688 | n58690 ;
  assign n58692 = n84253 & n58691 ;
  assign n58693 = n57829 & n84249 ;
  assign n58694 = n58552 & n58693 ;
  assign n58695 = n58692 | n58694 ;
  assign n58696 = n73617 & n58695 ;
  assign n84258 = ~n58524 ;
  assign n58697 = n58523 & n84258 ;
  assign n58698 = n57846 | n58523 ;
  assign n84259 = ~n58698 ;
  assign n58699 = n58660 & n84259 ;
  assign n58700 = n58697 | n58699 ;
  assign n58701 = n84253 & n58700 ;
  assign n58702 = n57837 & n84249 ;
  assign n58703 = n58552 & n58702 ;
  assign n58704 = n58701 | n58703 ;
  assign n58705 = n73188 & n58704 ;
  assign n84260 = ~n58659 ;
  assign n58707 = n58519 & n84260 ;
  assign n58708 = n57854 | n58519 ;
  assign n84261 = ~n58708 ;
  assign n58709 = n58515 & n84261 ;
  assign n58710 = n58707 | n58709 ;
  assign n58711 = n84253 & n58710 ;
  assign n58712 = n57845 & n84249 ;
  assign n58713 = n58552 & n58712 ;
  assign n58714 = n58711 | n58713 ;
  assign n58715 = n73177 & n58714 ;
  assign n84262 = ~n58514 ;
  assign n58716 = n58513 & n84262 ;
  assign n58717 = n57862 | n58513 ;
  assign n84263 = ~n58717 ;
  assign n58718 = n58656 & n84263 ;
  assign n58719 = n58716 | n58718 ;
  assign n58720 = n84253 & n58719 ;
  assign n58721 = n57853 & n84249 ;
  assign n58722 = n58552 & n58721 ;
  assign n58723 = n58720 | n58722 ;
  assign n58724 = n72752 & n58723 ;
  assign n84264 = ~n58655 ;
  assign n58725 = n58509 & n84264 ;
  assign n58726 = n57870 | n58509 ;
  assign n84265 = ~n58726 ;
  assign n58727 = n58505 & n84265 ;
  assign n58728 = n58725 | n58727 ;
  assign n58729 = n84253 & n58728 ;
  assign n58730 = n57861 & n84249 ;
  assign n58731 = n58552 & n58730 ;
  assign n58732 = n58729 | n58731 ;
  assign n58733 = n72393 & n58732 ;
  assign n84266 = ~n58504 ;
  assign n58734 = n58503 & n84266 ;
  assign n58735 = n57878 | n58503 ;
  assign n84267 = ~n58735 ;
  assign n58736 = n58652 & n84267 ;
  assign n58737 = n58734 | n58736 ;
  assign n58738 = n84253 & n58737 ;
  assign n58739 = n57869 & n84249 ;
  assign n58740 = n58552 & n58739 ;
  assign n58741 = n58738 | n58740 ;
  assign n58742 = n72385 & n58741 ;
  assign n84268 = ~n58651 ;
  assign n58743 = n58499 & n84268 ;
  assign n58744 = n57886 | n58499 ;
  assign n84269 = ~n58744 ;
  assign n58745 = n58495 & n84269 ;
  assign n58746 = n58743 | n58745 ;
  assign n58747 = n84253 & n58746 ;
  assign n58748 = n57877 & n84249 ;
  assign n58749 = n58552 & n58748 ;
  assign n58750 = n58747 | n58749 ;
  assign n58751 = n72025 & n58750 ;
  assign n84270 = ~n58494 ;
  assign n58752 = n58493 & n84270 ;
  assign n58753 = n57894 | n58493 ;
  assign n84271 = ~n58753 ;
  assign n58754 = n58648 & n84271 ;
  assign n58755 = n58752 | n58754 ;
  assign n58756 = n84253 & n58755 ;
  assign n58757 = n57885 & n84249 ;
  assign n58758 = n58552 & n58757 ;
  assign n58759 = n58756 | n58758 ;
  assign n58760 = n71645 & n58759 ;
  assign n84272 = ~n58647 ;
  assign n58761 = n58489 & n84272 ;
  assign n58762 = n57902 | n58489 ;
  assign n84273 = ~n58762 ;
  assign n58763 = n58485 & n84273 ;
  assign n58764 = n58761 | n58763 ;
  assign n58765 = n84253 & n58764 ;
  assign n58766 = n57893 & n84249 ;
  assign n58767 = n58552 & n58766 ;
  assign n58768 = n58765 | n58767 ;
  assign n58769 = n71633 & n58768 ;
  assign n84274 = ~n58484 ;
  assign n58770 = n58483 & n84274 ;
  assign n58771 = n57910 | n58483 ;
  assign n84275 = ~n58771 ;
  assign n58772 = n58644 & n84275 ;
  assign n58773 = n58770 | n58772 ;
  assign n58774 = n84253 & n58773 ;
  assign n58775 = n57901 & n84249 ;
  assign n58776 = n58552 & n58775 ;
  assign n58777 = n58774 | n58776 ;
  assign n58778 = n71253 & n58777 ;
  assign n84276 = ~n58643 ;
  assign n58779 = n58479 & n84276 ;
  assign n58780 = n57918 | n58479 ;
  assign n84277 = ~n58780 ;
  assign n58781 = n58475 & n84277 ;
  assign n58782 = n58779 | n58781 ;
  assign n58783 = n84253 & n58782 ;
  assign n58784 = n57909 & n84249 ;
  assign n58785 = n58552 & n58784 ;
  assign n58786 = n58783 | n58785 ;
  assign n58787 = n70935 & n58786 ;
  assign n84278 = ~n58474 ;
  assign n58788 = n58473 & n84278 ;
  assign n58789 = n57926 | n58473 ;
  assign n84279 = ~n58789 ;
  assign n58790 = n58640 & n84279 ;
  assign n58791 = n58788 | n58790 ;
  assign n58792 = n84253 & n58791 ;
  assign n58793 = n57917 & n84249 ;
  assign n58794 = n58552 & n58793 ;
  assign n58795 = n58792 | n58794 ;
  assign n58796 = n70927 & n58795 ;
  assign n84280 = ~n58639 ;
  assign n58797 = n58468 & n84280 ;
  assign n58469 = n57934 | n58468 ;
  assign n84281 = ~n58469 ;
  assign n58798 = n84281 & n58638 ;
  assign n58799 = n58797 | n58798 ;
  assign n58800 = n84253 & n58799 ;
  assign n58801 = n57925 & n84249 ;
  assign n58802 = n58552 & n58801 ;
  assign n58803 = n58800 | n58802 ;
  assign n58804 = n70609 & n58803 ;
  assign n84282 = ~n58463 ;
  assign n58805 = n58462 & n84282 ;
  assign n58806 = n57942 | n58462 ;
  assign n84283 = ~n58806 ;
  assign n58807 = n58636 & n84283 ;
  assign n58808 = n58805 | n58807 ;
  assign n58809 = n84253 & n58808 ;
  assign n58810 = n57933 & n84249 ;
  assign n58811 = n58552 & n58810 ;
  assign n58812 = n58809 | n58811 ;
  assign n58813 = n70276 & n58812 ;
  assign n84284 = ~n58635 ;
  assign n58814 = n58458 & n84284 ;
  assign n58815 = n57950 | n58458 ;
  assign n84285 = ~n58815 ;
  assign n58816 = n58454 & n84285 ;
  assign n58817 = n58814 | n58816 ;
  assign n58818 = n84253 & n58817 ;
  assign n58819 = n57941 & n84249 ;
  assign n58820 = n58552 & n58819 ;
  assign n58821 = n58818 | n58820 ;
  assign n58822 = n70176 & n58821 ;
  assign n84286 = ~n58453 ;
  assign n58823 = n58452 & n84286 ;
  assign n58824 = n57958 | n58452 ;
  assign n84287 = ~n58824 ;
  assign n58825 = n58632 & n84287 ;
  assign n58826 = n58823 | n58825 ;
  assign n58827 = n84253 & n58826 ;
  assign n58828 = n57949 & n84249 ;
  assign n58829 = n58552 & n58828 ;
  assign n58830 = n58827 | n58829 ;
  assign n58831 = n69857 & n58830 ;
  assign n84288 = ~n58631 ;
  assign n58832 = n58448 & n84288 ;
  assign n58833 = n57966 | n58448 ;
  assign n84289 = ~n58833 ;
  assign n58834 = n58444 & n84289 ;
  assign n58835 = n58832 | n58834 ;
  assign n58836 = n84253 & n58835 ;
  assign n58837 = n57957 & n84249 ;
  assign n58838 = n58552 & n58837 ;
  assign n58839 = n58836 | n58838 ;
  assign n58840 = n69656 & n58839 ;
  assign n84290 = ~n58443 ;
  assign n58841 = n58442 & n84290 ;
  assign n58842 = n57974 | n58442 ;
  assign n84291 = ~n58842 ;
  assign n58843 = n58628 & n84291 ;
  assign n58844 = n58841 | n58843 ;
  assign n58845 = n84253 & n58844 ;
  assign n58846 = n57965 & n84249 ;
  assign n58847 = n58552 & n58846 ;
  assign n58848 = n58845 | n58847 ;
  assign n58849 = n69528 & n58848 ;
  assign n84292 = ~n58627 ;
  assign n58850 = n58438 & n84292 ;
  assign n58851 = n57982 | n58438 ;
  assign n84293 = ~n58851 ;
  assign n58852 = n58434 & n84293 ;
  assign n58853 = n58850 | n58852 ;
  assign n58854 = n84253 & n58853 ;
  assign n58855 = n57973 & n84249 ;
  assign n58856 = n58552 & n58855 ;
  assign n58857 = n58854 | n58856 ;
  assign n58858 = n69261 & n58857 ;
  assign n84294 = ~n58433 ;
  assign n58859 = n58431 & n84294 ;
  assign n58432 = n57990 | n58431 ;
  assign n84295 = ~n58432 ;
  assign n58860 = n58428 & n84295 ;
  assign n58861 = n58859 | n58860 ;
  assign n58862 = n84253 & n58861 ;
  assign n58863 = n57981 & n84249 ;
  assign n58864 = n58552 & n58863 ;
  assign n58865 = n58862 | n58864 ;
  assign n58866 = n69075 & n58865 ;
  assign n84296 = ~n58623 ;
  assign n58867 = n58427 & n84296 ;
  assign n58868 = n57998 | n58427 ;
  assign n84297 = ~n58868 ;
  assign n58869 = n58423 & n84297 ;
  assign n58870 = n58867 | n58869 ;
  assign n58871 = n84253 & n58870 ;
  assign n58872 = n57989 & n84249 ;
  assign n58873 = n58552 & n58872 ;
  assign n58874 = n58871 | n58873 ;
  assign n58875 = n68993 & n58874 ;
  assign n84298 = ~n58422 ;
  assign n58876 = n58421 & n84298 ;
  assign n58877 = n58006 | n58421 ;
  assign n84299 = ~n58877 ;
  assign n58878 = n58620 & n84299 ;
  assign n58879 = n58876 | n58878 ;
  assign n58880 = n84253 & n58879 ;
  assign n58881 = n57997 & n84249 ;
  assign n58882 = n58552 & n58881 ;
  assign n58883 = n58880 | n58882 ;
  assign n58884 = n68716 & n58883 ;
  assign n84300 = ~n58619 ;
  assign n58885 = n58417 & n84300 ;
  assign n58886 = n58014 | n58417 ;
  assign n84301 = ~n58886 ;
  assign n58887 = n58413 & n84301 ;
  assign n58888 = n58885 | n58887 ;
  assign n58889 = n84253 & n58888 ;
  assign n58890 = n58005 & n84249 ;
  assign n58891 = n58552 & n58890 ;
  assign n58892 = n58889 | n58891 ;
  assign n58893 = n68545 & n58892 ;
  assign n84302 = ~n58412 ;
  assign n58894 = n58411 & n84302 ;
  assign n58895 = n58022 | n58411 ;
  assign n84303 = ~n58895 ;
  assign n58896 = n58616 & n84303 ;
  assign n58897 = n58894 | n58896 ;
  assign n58898 = n84253 & n58897 ;
  assign n58899 = n58013 & n84249 ;
  assign n58900 = n58552 & n58899 ;
  assign n58901 = n58898 | n58900 ;
  assign n58902 = n68438 & n58901 ;
  assign n84304 = ~n58615 ;
  assign n58903 = n58406 & n84304 ;
  assign n58407 = n58030 | n58406 ;
  assign n84305 = ~n58407 ;
  assign n58904 = n84305 & n58614 ;
  assign n58905 = n58903 | n58904 ;
  assign n58906 = n84253 & n58905 ;
  assign n58907 = n58021 & n84249 ;
  assign n58908 = n58552 & n58907 ;
  assign n58909 = n58906 | n58908 ;
  assign n58910 = n68214 & n58909 ;
  assign n84306 = ~n58401 ;
  assign n58911 = n58400 & n84306 ;
  assign n58912 = n58038 | n58400 ;
  assign n84307 = ~n58912 ;
  assign n58913 = n58612 & n84307 ;
  assign n58914 = n58911 | n58913 ;
  assign n58915 = n84253 & n58914 ;
  assign n58916 = n58029 & n84249 ;
  assign n58917 = n58552 & n58916 ;
  assign n58918 = n58915 | n58917 ;
  assign n58919 = n68058 & n58918 ;
  assign n84308 = ~n58611 ;
  assign n58920 = n58396 & n84308 ;
  assign n58921 = n58046 | n58396 ;
  assign n84309 = ~n58921 ;
  assign n58922 = n58392 & n84309 ;
  assign n58923 = n58920 | n58922 ;
  assign n58924 = n84253 & n58923 ;
  assign n58925 = n58037 & n84249 ;
  assign n58926 = n58552 & n58925 ;
  assign n58927 = n58924 | n58926 ;
  assign n58928 = n67986 & n58927 ;
  assign n84310 = ~n58391 ;
  assign n58929 = n58390 & n84310 ;
  assign n58930 = n58054 | n58390 ;
  assign n84311 = ~n58930 ;
  assign n58931 = n58608 & n84311 ;
  assign n58932 = n58929 | n58931 ;
  assign n58933 = n84253 & n58932 ;
  assign n58934 = n58045 & n84249 ;
  assign n58935 = n58552 & n58934 ;
  assign n58936 = n58933 | n58935 ;
  assign n58937 = n67763 & n58936 ;
  assign n84312 = ~n58607 ;
  assign n58938 = n58386 & n84312 ;
  assign n58939 = n58062 | n58386 ;
  assign n84313 = ~n58939 ;
  assign n58940 = n58382 & n84313 ;
  assign n58941 = n58938 | n58940 ;
  assign n58942 = n84253 & n58941 ;
  assign n58943 = n58053 & n84249 ;
  assign n58944 = n58552 & n58943 ;
  assign n58945 = n58942 | n58944 ;
  assign n58946 = n67622 & n58945 ;
  assign n84314 = ~n58381 ;
  assign n58947 = n58379 & n84314 ;
  assign n58380 = n58070 | n58379 ;
  assign n84315 = ~n58380 ;
  assign n58948 = n58376 & n84315 ;
  assign n58949 = n58947 | n58948 ;
  assign n58950 = n84253 & n58949 ;
  assign n58951 = n58061 & n84249 ;
  assign n58952 = n58552 & n58951 ;
  assign n58953 = n58950 | n58952 ;
  assign n58954 = n67531 & n58953 ;
  assign n84316 = ~n58603 ;
  assign n58955 = n58375 & n84316 ;
  assign n58956 = n58078 | n58375 ;
  assign n84317 = ~n58956 ;
  assign n58957 = n58371 & n84317 ;
  assign n58958 = n58955 | n58957 ;
  assign n58959 = n84253 & n58958 ;
  assign n58960 = n58069 & n84249 ;
  assign n58961 = n58552 & n58960 ;
  assign n58962 = n58959 | n58961 ;
  assign n58963 = n67348 & n58962 ;
  assign n84318 = ~n58370 ;
  assign n58964 = n58369 & n84318 ;
  assign n58965 = n58086 | n58369 ;
  assign n84319 = ~n58965 ;
  assign n58966 = n58600 & n84319 ;
  assign n58967 = n58964 | n58966 ;
  assign n58968 = n84253 & n58967 ;
  assign n58969 = n58077 & n84249 ;
  assign n58970 = n58552 & n58969 ;
  assign n58971 = n58968 | n58970 ;
  assign n58972 = n67222 & n58971 ;
  assign n84320 = ~n58599 ;
  assign n58973 = n58365 & n84320 ;
  assign n58974 = n58094 | n58365 ;
  assign n84321 = ~n58974 ;
  assign n58975 = n58361 & n84321 ;
  assign n58976 = n58973 | n58975 ;
  assign n58977 = n84253 & n58976 ;
  assign n58978 = n58085 & n84249 ;
  assign n58979 = n58552 & n58978 ;
  assign n58980 = n58977 | n58979 ;
  assign n58981 = n67164 & n58980 ;
  assign n84322 = ~n58360 ;
  assign n58982 = n58359 & n84322 ;
  assign n58983 = n58102 | n58359 ;
  assign n84323 = ~n58983 ;
  assign n58984 = n58596 & n84323 ;
  assign n58985 = n58982 | n58984 ;
  assign n58986 = n84253 & n58985 ;
  assign n58987 = n58093 & n84249 ;
  assign n58988 = n58552 & n58987 ;
  assign n58989 = n58986 | n58988 ;
  assign n58990 = n66979 & n58989 ;
  assign n84324 = ~n58595 ;
  assign n58991 = n58355 & n84324 ;
  assign n58992 = n58110 | n58355 ;
  assign n84325 = ~n58992 ;
  assign n58993 = n58351 & n84325 ;
  assign n58994 = n58991 | n58993 ;
  assign n58995 = n84253 & n58994 ;
  assign n58996 = n58101 & n84249 ;
  assign n58997 = n58552 & n58996 ;
  assign n58998 = n58995 | n58997 ;
  assign n58999 = n66868 & n58998 ;
  assign n84326 = ~n58350 ;
  assign n59000 = n58349 & n84326 ;
  assign n59001 = n58118 | n58349 ;
  assign n84327 = ~n59001 ;
  assign n59002 = n58592 & n84327 ;
  assign n59003 = n59000 | n59002 ;
  assign n59004 = n84253 & n59003 ;
  assign n59005 = n58109 & n84249 ;
  assign n59006 = n58552 & n59005 ;
  assign n59007 = n59004 | n59006 ;
  assign n59008 = n66797 & n59007 ;
  assign n84328 = ~n58591 ;
  assign n59009 = n58345 & n84328 ;
  assign n59010 = n58126 | n58345 ;
  assign n84329 = ~n59010 ;
  assign n59011 = n58341 & n84329 ;
  assign n59012 = n59009 | n59011 ;
  assign n59013 = n84253 & n59012 ;
  assign n59014 = n58117 & n84249 ;
  assign n59015 = n58552 & n59014 ;
  assign n59016 = n59013 | n59015 ;
  assign n59017 = n66654 & n59016 ;
  assign n84330 = ~n58340 ;
  assign n59018 = n58339 & n84330 ;
  assign n59019 = n58134 | n58339 ;
  assign n84331 = ~n59019 ;
  assign n59020 = n58588 & n84331 ;
  assign n59021 = n59018 | n59020 ;
  assign n59022 = n84253 & n59021 ;
  assign n59023 = n58125 & n84249 ;
  assign n59024 = n58552 & n59023 ;
  assign n59025 = n59022 | n59024 ;
  assign n59026 = n66560 & n59025 ;
  assign n84332 = ~n58587 ;
  assign n59027 = n58335 & n84332 ;
  assign n59028 = n58142 | n58335 ;
  assign n84333 = ~n59028 ;
  assign n59029 = n58331 & n84333 ;
  assign n59030 = n59027 | n59029 ;
  assign n59031 = n84253 & n59030 ;
  assign n59032 = n58133 & n84249 ;
  assign n59033 = n58552 & n59032 ;
  assign n59034 = n59031 | n59033 ;
  assign n59035 = n66505 & n59034 ;
  assign n84334 = ~n58330 ;
  assign n59036 = n58329 & n84334 ;
  assign n59037 = n58150 | n58329 ;
  assign n84335 = ~n59037 ;
  assign n59038 = n58584 & n84335 ;
  assign n59039 = n59036 | n59038 ;
  assign n59040 = n84253 & n59039 ;
  assign n59041 = n58141 & n84249 ;
  assign n59042 = n58552 & n59041 ;
  assign n59043 = n59040 | n59042 ;
  assign n59044 = n66379 & n59043 ;
  assign n84336 = ~n58583 ;
  assign n59045 = n58325 & n84336 ;
  assign n59046 = n58158 | n58325 ;
  assign n84337 = ~n59046 ;
  assign n59047 = n58321 & n84337 ;
  assign n59048 = n59045 | n59047 ;
  assign n59049 = n84253 & n59048 ;
  assign n59050 = n58149 & n84249 ;
  assign n59051 = n58552 & n59050 ;
  assign n59052 = n59049 | n59051 ;
  assign n59053 = n66299 & n59052 ;
  assign n84338 = ~n58320 ;
  assign n59054 = n58319 & n84338 ;
  assign n59055 = n58166 | n58319 ;
  assign n84339 = ~n59055 ;
  assign n59056 = n58580 & n84339 ;
  assign n59057 = n59054 | n59056 ;
  assign n59058 = n84253 & n59057 ;
  assign n59059 = n58157 & n84249 ;
  assign n59060 = n58552 & n59059 ;
  assign n59061 = n59058 | n59060 ;
  assign n59062 = n66244 & n59061 ;
  assign n84340 = ~n58579 ;
  assign n59063 = n58315 & n84340 ;
  assign n59064 = n58174 | n58315 ;
  assign n84341 = ~n59064 ;
  assign n59065 = n58311 & n84341 ;
  assign n59066 = n59063 | n59065 ;
  assign n59067 = n84253 & n59066 ;
  assign n59068 = n58165 & n84249 ;
  assign n59069 = n58552 & n59068 ;
  assign n59070 = n59067 | n59069 ;
  assign n59071 = n66145 & n59070 ;
  assign n84342 = ~n58310 ;
  assign n59072 = n58309 & n84342 ;
  assign n59073 = n58182 | n58309 ;
  assign n84343 = ~n59073 ;
  assign n59074 = n58576 & n84343 ;
  assign n59075 = n59072 | n59074 ;
  assign n59076 = n84253 & n59075 ;
  assign n59077 = n58173 & n84249 ;
  assign n59078 = n58552 & n59077 ;
  assign n59079 = n59076 | n59078 ;
  assign n59080 = n66081 & n59079 ;
  assign n84344 = ~n58575 ;
  assign n59081 = n58305 & n84344 ;
  assign n59082 = n58190 | n58305 ;
  assign n84345 = ~n59082 ;
  assign n59083 = n58301 & n84345 ;
  assign n59084 = n59081 | n59083 ;
  assign n59085 = n84253 & n59084 ;
  assign n59086 = n58181 & n84249 ;
  assign n59087 = n58552 & n59086 ;
  assign n59088 = n59085 | n59087 ;
  assign n59089 = n66043 & n59088 ;
  assign n84346 = ~n58300 ;
  assign n59090 = n58299 & n84346 ;
  assign n59091 = n58198 | n58299 ;
  assign n84347 = ~n59091 ;
  assign n59092 = n58572 & n84347 ;
  assign n59093 = n59090 | n59092 ;
  assign n59094 = n84253 & n59093 ;
  assign n59095 = n58189 & n84249 ;
  assign n59096 = n58552 & n59095 ;
  assign n59097 = n59094 | n59096 ;
  assign n59098 = n65960 & n59097 ;
  assign n84348 = ~n58571 ;
  assign n59099 = n58295 & n84348 ;
  assign n59100 = n58206 | n58295 ;
  assign n84349 = ~n59100 ;
  assign n59101 = n58291 & n84349 ;
  assign n59102 = n59099 | n59101 ;
  assign n59103 = n84253 & n59102 ;
  assign n59104 = n58197 & n84249 ;
  assign n59105 = n58552 & n59104 ;
  assign n59106 = n59103 | n59105 ;
  assign n59107 = n65909 & n59106 ;
  assign n84350 = ~n58290 ;
  assign n59108 = n58289 & n84350 ;
  assign n59109 = n58214 | n58289 ;
  assign n84351 = ~n59109 ;
  assign n59110 = n58568 & n84351 ;
  assign n59111 = n59108 | n59110 ;
  assign n59112 = n84253 & n59111 ;
  assign n59113 = n58205 & n84249 ;
  assign n59114 = n58552 & n59113 ;
  assign n59115 = n59112 | n59114 ;
  assign n59116 = n65877 & n59115 ;
  assign n84352 = ~n58567 ;
  assign n59117 = n58284 & n84352 ;
  assign n58285 = n58223 | n58284 ;
  assign n84353 = ~n58285 ;
  assign n59118 = n84353 & n58566 ;
  assign n59119 = n59117 | n59118 ;
  assign n59120 = n84253 & n59119 ;
  assign n59121 = n58213 & n84249 ;
  assign n59122 = n58552 & n59121 ;
  assign n59123 = n59120 | n59122 ;
  assign n59124 = n65820 & n59123 ;
  assign n84354 = ~n58279 ;
  assign n59125 = n58278 & n84354 ;
  assign n59126 = n58231 | n58278 ;
  assign n84355 = ~n59126 ;
  assign n59127 = n58564 & n84355 ;
  assign n59128 = n59125 | n59127 ;
  assign n59129 = n84253 & n59128 ;
  assign n59130 = n58222 & n84249 ;
  assign n59131 = n58552 & n59130 ;
  assign n59132 = n59129 | n59131 ;
  assign n59133 = n65791 & n59132 ;
  assign n84356 = ~n58563 ;
  assign n59134 = n58274 & n84356 ;
  assign n59135 = n58239 | n58274 ;
  assign n84357 = ~n59135 ;
  assign n59136 = n58270 & n84357 ;
  assign n59137 = n59134 | n59136 ;
  assign n59138 = n84253 & n59137 ;
  assign n59139 = n58230 & n84249 ;
  assign n59140 = n58552 & n59139 ;
  assign n59141 = n59138 | n59140 ;
  assign n59142 = n65772 & n59141 ;
  assign n84358 = ~n58269 ;
  assign n59144 = n58268 & n84358 ;
  assign n59143 = n58247 | n58268 ;
  assign n84359 = ~n59143 ;
  assign n59145 = n58265 & n84359 ;
  assign n59146 = n59144 | n59145 ;
  assign n59147 = n84253 & n59146 ;
  assign n59148 = n58238 & n84249 ;
  assign n59149 = n58552 & n59148 ;
  assign n59150 = n59147 | n59149 ;
  assign n59151 = n65746 & n59150 ;
  assign n84360 = ~n58559 ;
  assign n59152 = n58264 & n84360 ;
  assign n58558 = n58260 | n58264 ;
  assign n84361 = ~n58558 ;
  assign n59153 = n58557 & n84361 ;
  assign n59154 = n59152 | n59153 ;
  assign n59155 = n84253 & n59154 ;
  assign n59156 = n58246 & n84249 ;
  assign n59157 = n58552 & n59156 ;
  assign n59158 = n59155 | n59157 ;
  assign n59159 = n65721 & n59158 ;
  assign n59160 = n26052 & n58256 ;
  assign n59161 = n84251 & n59160 ;
  assign n84362 = ~n59161 ;
  assign n59162 = n58557 & n84362 ;
  assign n59163 = n84253 & n59162 ;
  assign n59164 = n58259 & n84249 ;
  assign n59165 = n58552 & n59164 ;
  assign n59166 = n59163 | n59165 ;
  assign n59167 = n65686 & n59166 ;
  assign n58706 = n26052 & n84253 ;
  assign n59172 = x64 & n84253 ;
  assign n84363 = ~n59172 ;
  assign n59173 = x7 & n84363 ;
  assign n59174 = n58706 | n59173 ;
  assign n59176 = x65 & n59174 ;
  assign n59168 = n58551 | n58678 ;
  assign n59169 = n84249 & n59168 ;
  assign n84364 = ~n59169 ;
  assign n59170 = x64 & n84364 ;
  assign n84365 = ~n59170 ;
  assign n59171 = x7 & n84365 ;
  assign n59175 = x65 | n58706 ;
  assign n59177 = n59171 | n59175 ;
  assign n84366 = ~n59176 ;
  assign n59178 = n84366 & n59177 ;
  assign n59179 = n26974 | n59178 ;
  assign n59180 = n65670 & n59174 ;
  assign n84367 = ~n59180 ;
  assign n59181 = n59179 & n84367 ;
  assign n84368 = ~n59165 ;
  assign n59182 = x66 & n84368 ;
  assign n84369 = ~n59163 ;
  assign n59183 = n84369 & n59182 ;
  assign n59184 = n59167 | n59183 ;
  assign n59185 = n59181 | n59184 ;
  assign n84370 = ~n59167 ;
  assign n59186 = n84370 & n59185 ;
  assign n84371 = ~n59157 ;
  assign n59187 = x67 & n84371 ;
  assign n84372 = ~n59155 ;
  assign n59188 = n84372 & n59187 ;
  assign n59189 = n59186 | n59188 ;
  assign n84373 = ~n59159 ;
  assign n59190 = n84373 & n59189 ;
  assign n84374 = ~n59149 ;
  assign n59191 = x68 & n84374 ;
  assign n84375 = ~n59147 ;
  assign n59192 = n84375 & n59191 ;
  assign n59193 = n59151 | n59192 ;
  assign n59194 = n59190 | n59193 ;
  assign n84376 = ~n59151 ;
  assign n59195 = n84376 & n59194 ;
  assign n84377 = ~n59140 ;
  assign n59196 = x69 & n84377 ;
  assign n84378 = ~n59138 ;
  assign n59197 = n84378 & n59196 ;
  assign n59198 = n59195 | n59197 ;
  assign n84379 = ~n59142 ;
  assign n59199 = n84379 & n59198 ;
  assign n84380 = ~n59131 ;
  assign n59200 = x70 & n84380 ;
  assign n84381 = ~n59129 ;
  assign n59201 = n84381 & n59200 ;
  assign n59202 = n59133 | n59201 ;
  assign n59203 = n59199 | n59202 ;
  assign n84382 = ~n59133 ;
  assign n59204 = n84382 & n59203 ;
  assign n84383 = ~n59122 ;
  assign n59205 = x71 & n84383 ;
  assign n84384 = ~n59120 ;
  assign n59206 = n84384 & n59205 ;
  assign n59207 = n59124 | n59206 ;
  assign n59209 = n59204 | n59207 ;
  assign n84385 = ~n59124 ;
  assign n59210 = n84385 & n59209 ;
  assign n84386 = ~n59114 ;
  assign n59211 = x72 & n84386 ;
  assign n84387 = ~n59112 ;
  assign n59212 = n84387 & n59211 ;
  assign n59213 = n59116 | n59212 ;
  assign n59214 = n59210 | n59213 ;
  assign n84388 = ~n59116 ;
  assign n59215 = n84388 & n59214 ;
  assign n84389 = ~n59105 ;
  assign n59216 = x73 & n84389 ;
  assign n84390 = ~n59103 ;
  assign n59217 = n84390 & n59216 ;
  assign n59218 = n59107 | n59217 ;
  assign n59220 = n59215 | n59218 ;
  assign n84391 = ~n59107 ;
  assign n59221 = n84391 & n59220 ;
  assign n84392 = ~n59096 ;
  assign n59222 = x74 & n84392 ;
  assign n84393 = ~n59094 ;
  assign n59223 = n84393 & n59222 ;
  assign n59224 = n59098 | n59223 ;
  assign n59225 = n59221 | n59224 ;
  assign n84394 = ~n59098 ;
  assign n59226 = n84394 & n59225 ;
  assign n84395 = ~n59087 ;
  assign n59227 = x75 & n84395 ;
  assign n84396 = ~n59085 ;
  assign n59228 = n84396 & n59227 ;
  assign n59229 = n59089 | n59228 ;
  assign n59231 = n59226 | n59229 ;
  assign n84397 = ~n59089 ;
  assign n59232 = n84397 & n59231 ;
  assign n84398 = ~n59078 ;
  assign n59233 = x76 & n84398 ;
  assign n84399 = ~n59076 ;
  assign n59234 = n84399 & n59233 ;
  assign n59235 = n59080 | n59234 ;
  assign n59236 = n59232 | n59235 ;
  assign n84400 = ~n59080 ;
  assign n59237 = n84400 & n59236 ;
  assign n84401 = ~n59069 ;
  assign n59238 = x77 & n84401 ;
  assign n84402 = ~n59067 ;
  assign n59239 = n84402 & n59238 ;
  assign n59240 = n59071 | n59239 ;
  assign n59242 = n59237 | n59240 ;
  assign n84403 = ~n59071 ;
  assign n59243 = n84403 & n59242 ;
  assign n84404 = ~n59060 ;
  assign n59244 = x78 & n84404 ;
  assign n84405 = ~n59058 ;
  assign n59245 = n84405 & n59244 ;
  assign n59246 = n59062 | n59245 ;
  assign n59247 = n59243 | n59246 ;
  assign n84406 = ~n59062 ;
  assign n59248 = n84406 & n59247 ;
  assign n84407 = ~n59051 ;
  assign n59249 = x79 & n84407 ;
  assign n84408 = ~n59049 ;
  assign n59250 = n84408 & n59249 ;
  assign n59251 = n59053 | n59250 ;
  assign n59253 = n59248 | n59251 ;
  assign n84409 = ~n59053 ;
  assign n59254 = n84409 & n59253 ;
  assign n84410 = ~n59042 ;
  assign n59255 = x80 & n84410 ;
  assign n84411 = ~n59040 ;
  assign n59256 = n84411 & n59255 ;
  assign n59257 = n59044 | n59256 ;
  assign n59258 = n59254 | n59257 ;
  assign n84412 = ~n59044 ;
  assign n59259 = n84412 & n59258 ;
  assign n84413 = ~n59033 ;
  assign n59260 = x81 & n84413 ;
  assign n84414 = ~n59031 ;
  assign n59261 = n84414 & n59260 ;
  assign n59262 = n59035 | n59261 ;
  assign n59264 = n59259 | n59262 ;
  assign n84415 = ~n59035 ;
  assign n59265 = n84415 & n59264 ;
  assign n84416 = ~n59024 ;
  assign n59266 = x82 & n84416 ;
  assign n84417 = ~n59022 ;
  assign n59267 = n84417 & n59266 ;
  assign n59268 = n59026 | n59267 ;
  assign n59269 = n59265 | n59268 ;
  assign n84418 = ~n59026 ;
  assign n59270 = n84418 & n59269 ;
  assign n84419 = ~n59015 ;
  assign n59271 = x83 & n84419 ;
  assign n84420 = ~n59013 ;
  assign n59272 = n84420 & n59271 ;
  assign n59273 = n59017 | n59272 ;
  assign n59275 = n59270 | n59273 ;
  assign n84421 = ~n59017 ;
  assign n59276 = n84421 & n59275 ;
  assign n84422 = ~n59006 ;
  assign n59277 = x84 & n84422 ;
  assign n84423 = ~n59004 ;
  assign n59278 = n84423 & n59277 ;
  assign n59279 = n59008 | n59278 ;
  assign n59280 = n59276 | n59279 ;
  assign n84424 = ~n59008 ;
  assign n59281 = n84424 & n59280 ;
  assign n84425 = ~n58997 ;
  assign n59282 = x85 & n84425 ;
  assign n84426 = ~n58995 ;
  assign n59283 = n84426 & n59282 ;
  assign n59284 = n58999 | n59283 ;
  assign n59286 = n59281 | n59284 ;
  assign n84427 = ~n58999 ;
  assign n59287 = n84427 & n59286 ;
  assign n84428 = ~n58988 ;
  assign n59288 = x86 & n84428 ;
  assign n84429 = ~n58986 ;
  assign n59289 = n84429 & n59288 ;
  assign n59290 = n58990 | n59289 ;
  assign n59291 = n59287 | n59290 ;
  assign n84430 = ~n58990 ;
  assign n59292 = n84430 & n59291 ;
  assign n84431 = ~n58979 ;
  assign n59293 = x87 & n84431 ;
  assign n84432 = ~n58977 ;
  assign n59294 = n84432 & n59293 ;
  assign n59295 = n58981 | n59294 ;
  assign n59297 = n59292 | n59295 ;
  assign n84433 = ~n58981 ;
  assign n59298 = n84433 & n59297 ;
  assign n84434 = ~n58970 ;
  assign n59299 = x88 & n84434 ;
  assign n84435 = ~n58968 ;
  assign n59300 = n84435 & n59299 ;
  assign n59301 = n58972 | n59300 ;
  assign n59302 = n59298 | n59301 ;
  assign n84436 = ~n58972 ;
  assign n59303 = n84436 & n59302 ;
  assign n84437 = ~n58961 ;
  assign n59304 = x89 & n84437 ;
  assign n84438 = ~n58959 ;
  assign n59305 = n84438 & n59304 ;
  assign n59306 = n58963 | n59305 ;
  assign n59308 = n59303 | n59306 ;
  assign n84439 = ~n58963 ;
  assign n59309 = n84439 & n59308 ;
  assign n84440 = ~n58952 ;
  assign n59310 = x90 & n84440 ;
  assign n84441 = ~n58950 ;
  assign n59311 = n84441 & n59310 ;
  assign n59312 = n58954 | n59311 ;
  assign n59313 = n59309 | n59312 ;
  assign n84442 = ~n58954 ;
  assign n59314 = n84442 & n59313 ;
  assign n84443 = ~n58944 ;
  assign n59315 = x91 & n84443 ;
  assign n84444 = ~n58942 ;
  assign n59316 = n84444 & n59315 ;
  assign n59317 = n58946 | n59316 ;
  assign n59319 = n59314 | n59317 ;
  assign n84445 = ~n58946 ;
  assign n59320 = n84445 & n59319 ;
  assign n84446 = ~n58935 ;
  assign n59321 = x92 & n84446 ;
  assign n84447 = ~n58933 ;
  assign n59322 = n84447 & n59321 ;
  assign n59323 = n58937 | n59322 ;
  assign n59324 = n59320 | n59323 ;
  assign n84448 = ~n58937 ;
  assign n59325 = n84448 & n59324 ;
  assign n84449 = ~n58926 ;
  assign n59326 = x93 & n84449 ;
  assign n84450 = ~n58924 ;
  assign n59327 = n84450 & n59326 ;
  assign n59328 = n58928 | n59327 ;
  assign n59330 = n59325 | n59328 ;
  assign n84451 = ~n58928 ;
  assign n59331 = n84451 & n59330 ;
  assign n84452 = ~n58917 ;
  assign n59332 = x94 & n84452 ;
  assign n84453 = ~n58915 ;
  assign n59333 = n84453 & n59332 ;
  assign n59334 = n58919 | n59333 ;
  assign n59335 = n59331 | n59334 ;
  assign n84454 = ~n58919 ;
  assign n59336 = n84454 & n59335 ;
  assign n84455 = ~n58908 ;
  assign n59337 = x95 & n84455 ;
  assign n84456 = ~n58906 ;
  assign n59338 = n84456 & n59337 ;
  assign n59339 = n58910 | n59338 ;
  assign n59341 = n59336 | n59339 ;
  assign n84457 = ~n58910 ;
  assign n59342 = n84457 & n59341 ;
  assign n84458 = ~n58900 ;
  assign n59343 = x96 & n84458 ;
  assign n84459 = ~n58898 ;
  assign n59344 = n84459 & n59343 ;
  assign n59345 = n58902 | n59344 ;
  assign n59346 = n59342 | n59345 ;
  assign n84460 = ~n58902 ;
  assign n59347 = n84460 & n59346 ;
  assign n84461 = ~n58891 ;
  assign n59348 = x97 & n84461 ;
  assign n84462 = ~n58889 ;
  assign n59349 = n84462 & n59348 ;
  assign n59350 = n58893 | n59349 ;
  assign n59352 = n59347 | n59350 ;
  assign n84463 = ~n58893 ;
  assign n59353 = n84463 & n59352 ;
  assign n84464 = ~n58882 ;
  assign n59354 = x98 & n84464 ;
  assign n84465 = ~n58880 ;
  assign n59355 = n84465 & n59354 ;
  assign n59356 = n58884 | n59355 ;
  assign n59357 = n59353 | n59356 ;
  assign n84466 = ~n58884 ;
  assign n59358 = n84466 & n59357 ;
  assign n84467 = ~n58873 ;
  assign n59359 = x99 & n84467 ;
  assign n84468 = ~n58871 ;
  assign n59360 = n84468 & n59359 ;
  assign n59361 = n58875 | n59360 ;
  assign n59363 = n59358 | n59361 ;
  assign n84469 = ~n58875 ;
  assign n59364 = n84469 & n59363 ;
  assign n84470 = ~n58864 ;
  assign n59365 = x100 & n84470 ;
  assign n84471 = ~n58862 ;
  assign n59366 = n84471 & n59365 ;
  assign n59367 = n58866 | n59366 ;
  assign n59368 = n59364 | n59367 ;
  assign n84472 = ~n58866 ;
  assign n59369 = n84472 & n59368 ;
  assign n84473 = ~n58856 ;
  assign n59370 = x101 & n84473 ;
  assign n84474 = ~n58854 ;
  assign n59371 = n84474 & n59370 ;
  assign n59372 = n58858 | n59371 ;
  assign n59374 = n59369 | n59372 ;
  assign n84475 = ~n58858 ;
  assign n59375 = n84475 & n59374 ;
  assign n84476 = ~n58847 ;
  assign n59376 = x102 & n84476 ;
  assign n84477 = ~n58845 ;
  assign n59377 = n84477 & n59376 ;
  assign n59378 = n58849 | n59377 ;
  assign n59379 = n59375 | n59378 ;
  assign n84478 = ~n58849 ;
  assign n59380 = n84478 & n59379 ;
  assign n84479 = ~n58838 ;
  assign n59381 = x103 & n84479 ;
  assign n84480 = ~n58836 ;
  assign n59382 = n84480 & n59381 ;
  assign n59383 = n58840 | n59382 ;
  assign n59385 = n59380 | n59383 ;
  assign n84481 = ~n58840 ;
  assign n59386 = n84481 & n59385 ;
  assign n84482 = ~n58829 ;
  assign n59387 = x104 & n84482 ;
  assign n84483 = ~n58827 ;
  assign n59388 = n84483 & n59387 ;
  assign n59389 = n58831 | n59388 ;
  assign n59390 = n59386 | n59389 ;
  assign n84484 = ~n58831 ;
  assign n59391 = n84484 & n59390 ;
  assign n84485 = ~n58820 ;
  assign n59392 = x105 & n84485 ;
  assign n84486 = ~n58818 ;
  assign n59393 = n84486 & n59392 ;
  assign n59394 = n58822 | n59393 ;
  assign n59396 = n59391 | n59394 ;
  assign n84487 = ~n58822 ;
  assign n59397 = n84487 & n59396 ;
  assign n84488 = ~n58811 ;
  assign n59398 = x106 & n84488 ;
  assign n84489 = ~n58809 ;
  assign n59399 = n84489 & n59398 ;
  assign n59400 = n58813 | n59399 ;
  assign n59401 = n59397 | n59400 ;
  assign n84490 = ~n58813 ;
  assign n59402 = n84490 & n59401 ;
  assign n84491 = ~n58802 ;
  assign n59403 = x107 & n84491 ;
  assign n84492 = ~n58800 ;
  assign n59404 = n84492 & n59403 ;
  assign n59405 = n58804 | n59404 ;
  assign n59407 = n59402 | n59405 ;
  assign n84493 = ~n58804 ;
  assign n59408 = n84493 & n59407 ;
  assign n84494 = ~n58794 ;
  assign n59409 = x108 & n84494 ;
  assign n84495 = ~n58792 ;
  assign n59410 = n84495 & n59409 ;
  assign n59411 = n58796 | n59410 ;
  assign n59412 = n59408 | n59411 ;
  assign n84496 = ~n58796 ;
  assign n59413 = n84496 & n59412 ;
  assign n84497 = ~n58785 ;
  assign n59414 = x109 & n84497 ;
  assign n84498 = ~n58783 ;
  assign n59415 = n84498 & n59414 ;
  assign n59416 = n58787 | n59415 ;
  assign n59418 = n59413 | n59416 ;
  assign n84499 = ~n58787 ;
  assign n59419 = n84499 & n59418 ;
  assign n84500 = ~n58776 ;
  assign n59420 = x110 & n84500 ;
  assign n84501 = ~n58774 ;
  assign n59421 = n84501 & n59420 ;
  assign n59422 = n58778 | n59421 ;
  assign n59423 = n59419 | n59422 ;
  assign n84502 = ~n58778 ;
  assign n59424 = n84502 & n59423 ;
  assign n84503 = ~n58767 ;
  assign n59425 = x111 & n84503 ;
  assign n84504 = ~n58765 ;
  assign n59426 = n84504 & n59425 ;
  assign n59427 = n58769 | n59426 ;
  assign n59429 = n59424 | n59427 ;
  assign n84505 = ~n58769 ;
  assign n59430 = n84505 & n59429 ;
  assign n84506 = ~n58758 ;
  assign n59431 = x112 & n84506 ;
  assign n84507 = ~n58756 ;
  assign n59432 = n84507 & n59431 ;
  assign n59433 = n58760 | n59432 ;
  assign n59434 = n59430 | n59433 ;
  assign n84508 = ~n58760 ;
  assign n59435 = n84508 & n59434 ;
  assign n84509 = ~n58749 ;
  assign n59436 = x113 & n84509 ;
  assign n84510 = ~n58747 ;
  assign n59437 = n84510 & n59436 ;
  assign n59438 = n58751 | n59437 ;
  assign n59440 = n59435 | n59438 ;
  assign n84511 = ~n58751 ;
  assign n59441 = n84511 & n59440 ;
  assign n84512 = ~n58740 ;
  assign n59442 = x114 & n84512 ;
  assign n84513 = ~n58738 ;
  assign n59443 = n84513 & n59442 ;
  assign n59444 = n58742 | n59443 ;
  assign n59445 = n59441 | n59444 ;
  assign n84514 = ~n58742 ;
  assign n59446 = n84514 & n59445 ;
  assign n84515 = ~n58731 ;
  assign n59447 = x115 & n84515 ;
  assign n84516 = ~n58729 ;
  assign n59448 = n84516 & n59447 ;
  assign n59449 = n58733 | n59448 ;
  assign n59451 = n59446 | n59449 ;
  assign n84517 = ~n58733 ;
  assign n59452 = n84517 & n59451 ;
  assign n84518 = ~n58722 ;
  assign n59453 = x116 & n84518 ;
  assign n84519 = ~n58720 ;
  assign n59454 = n84519 & n59453 ;
  assign n59455 = n58724 | n59454 ;
  assign n59456 = n59452 | n59455 ;
  assign n84520 = ~n58724 ;
  assign n59457 = n84520 & n59456 ;
  assign n84521 = ~n58713 ;
  assign n59458 = x117 & n84521 ;
  assign n84522 = ~n58711 ;
  assign n59459 = n84522 & n59458 ;
  assign n59460 = n58715 | n59459 ;
  assign n59462 = n59457 | n59460 ;
  assign n84523 = ~n58715 ;
  assign n59463 = n84523 & n59462 ;
  assign n84524 = ~n58703 ;
  assign n59464 = x118 & n84524 ;
  assign n84525 = ~n58701 ;
  assign n59465 = n84525 & n59464 ;
  assign n59466 = n58705 | n59465 ;
  assign n59467 = n59463 | n59466 ;
  assign n84526 = ~n58705 ;
  assign n59468 = n84526 & n59467 ;
  assign n84527 = ~n58694 ;
  assign n59469 = x119 & n84527 ;
  assign n84528 = ~n58692 ;
  assign n59470 = n84528 & n59469 ;
  assign n59471 = n58696 | n59470 ;
  assign n59473 = n59468 | n59471 ;
  assign n84529 = ~n58696 ;
  assign n59474 = n84529 & n59473 ;
  assign n84530 = ~n58672 ;
  assign n59475 = x120 & n84530 ;
  assign n84531 = ~n58670 ;
  assign n59476 = n84531 & n59475 ;
  assign n59477 = n58687 | n59476 ;
  assign n59478 = n59474 | n59477 ;
  assign n84532 = ~n58687 ;
  assign n59479 = n84532 & n59478 ;
  assign n84533 = ~n58684 ;
  assign n59480 = x121 & n84533 ;
  assign n84534 = ~n58682 ;
  assign n59481 = n84534 & n59480 ;
  assign n59482 = n58686 | n59481 ;
  assign n59484 = n59479 | n59482 ;
  assign n84535 = ~n58686 ;
  assign n59485 = n84535 & n59484 ;
  assign n59486 = n27311 | n59485 ;
  assign n59487 = n58673 & n59486 ;
  assign n59488 = n58706 | n59171 ;
  assign n59489 = x65 & n59488 ;
  assign n84536 = ~n59489 ;
  assign n59490 = n59177 & n84536 ;
  assign n59491 = n26974 | n59490 ;
  assign n59492 = n84367 & n59491 ;
  assign n59493 = n59184 | n59492 ;
  assign n59494 = n84370 & n59493 ;
  assign n59495 = n59159 | n59188 ;
  assign n59497 = n59494 | n59495 ;
  assign n59498 = n84373 & n59497 ;
  assign n59499 = n59192 | n59498 ;
  assign n59501 = n84376 & n59499 ;
  assign n59502 = n59142 | n59197 ;
  assign n59504 = n59501 | n59502 ;
  assign n59505 = n84379 & n59504 ;
  assign n59506 = n59201 | n59505 ;
  assign n59508 = n84382 & n59506 ;
  assign n59509 = n59207 | n59508 ;
  assign n59510 = n84385 & n59509 ;
  assign n59511 = n59213 | n59510 ;
  assign n59513 = n84388 & n59511 ;
  assign n59514 = n59218 | n59513 ;
  assign n59515 = n84391 & n59514 ;
  assign n59516 = n59224 | n59515 ;
  assign n59518 = n84394 & n59516 ;
  assign n59519 = n59229 | n59518 ;
  assign n59520 = n84397 & n59519 ;
  assign n59521 = n59235 | n59520 ;
  assign n59523 = n84400 & n59521 ;
  assign n59524 = n59240 | n59523 ;
  assign n59525 = n84403 & n59524 ;
  assign n59526 = n59246 | n59525 ;
  assign n59528 = n84406 & n59526 ;
  assign n59529 = n59251 | n59528 ;
  assign n59530 = n84409 & n59529 ;
  assign n59531 = n59257 | n59530 ;
  assign n59533 = n84412 & n59531 ;
  assign n59534 = n59262 | n59533 ;
  assign n59535 = n84415 & n59534 ;
  assign n59536 = n59268 | n59535 ;
  assign n59538 = n84418 & n59536 ;
  assign n59539 = n59273 | n59538 ;
  assign n59540 = n84421 & n59539 ;
  assign n59541 = n59279 | n59540 ;
  assign n59543 = n84424 & n59541 ;
  assign n59544 = n59284 | n59543 ;
  assign n59545 = n84427 & n59544 ;
  assign n59546 = n59290 | n59545 ;
  assign n59548 = n84430 & n59546 ;
  assign n59549 = n59295 | n59548 ;
  assign n59550 = n84433 & n59549 ;
  assign n59551 = n59301 | n59550 ;
  assign n59553 = n84436 & n59551 ;
  assign n59554 = n59306 | n59553 ;
  assign n59555 = n84439 & n59554 ;
  assign n59556 = n59312 | n59555 ;
  assign n59558 = n84442 & n59556 ;
  assign n59559 = n59317 | n59558 ;
  assign n59560 = n84445 & n59559 ;
  assign n59561 = n59323 | n59560 ;
  assign n59563 = n84448 & n59561 ;
  assign n59564 = n59328 | n59563 ;
  assign n59565 = n84451 & n59564 ;
  assign n59566 = n59334 | n59565 ;
  assign n59568 = n84454 & n59566 ;
  assign n59569 = n59339 | n59568 ;
  assign n59570 = n84457 & n59569 ;
  assign n59571 = n59345 | n59570 ;
  assign n59573 = n84460 & n59571 ;
  assign n59574 = n59350 | n59573 ;
  assign n59575 = n84463 & n59574 ;
  assign n59576 = n59356 | n59575 ;
  assign n59578 = n84466 & n59576 ;
  assign n59579 = n59361 | n59578 ;
  assign n59580 = n84469 & n59579 ;
  assign n59581 = n59367 | n59580 ;
  assign n59583 = n84472 & n59581 ;
  assign n59584 = n59372 | n59583 ;
  assign n59585 = n84475 & n59584 ;
  assign n59586 = n59378 | n59585 ;
  assign n59588 = n84478 & n59586 ;
  assign n59589 = n59383 | n59588 ;
  assign n59590 = n84481 & n59589 ;
  assign n59591 = n59389 | n59590 ;
  assign n59593 = n84484 & n59591 ;
  assign n59594 = n59394 | n59593 ;
  assign n59595 = n84487 & n59594 ;
  assign n59596 = n59400 | n59595 ;
  assign n59598 = n84490 & n59596 ;
  assign n59599 = n59405 | n59598 ;
  assign n59600 = n84493 & n59599 ;
  assign n59601 = n59411 | n59600 ;
  assign n59603 = n84496 & n59601 ;
  assign n59604 = n59416 | n59603 ;
  assign n59605 = n84499 & n59604 ;
  assign n59606 = n59422 | n59605 ;
  assign n59608 = n84502 & n59606 ;
  assign n59609 = n59427 | n59608 ;
  assign n59610 = n84505 & n59609 ;
  assign n59611 = n59433 | n59610 ;
  assign n59613 = n84508 & n59611 ;
  assign n59614 = n59438 | n59613 ;
  assign n59615 = n84511 & n59614 ;
  assign n59616 = n59444 | n59615 ;
  assign n59618 = n84514 & n59616 ;
  assign n59619 = n59449 | n59618 ;
  assign n59620 = n84517 & n59619 ;
  assign n59621 = n59455 | n59620 ;
  assign n59623 = n84520 & n59621 ;
  assign n59624 = n59460 | n59623 ;
  assign n59625 = n84523 & n59624 ;
  assign n59626 = n59466 | n59625 ;
  assign n59628 = n84526 & n59626 ;
  assign n59629 = n59471 | n59628 ;
  assign n59630 = n84529 & n59629 ;
  assign n84537 = ~n59630 ;
  assign n59631 = n59477 & n84537 ;
  assign n59633 = n58696 | n59477 ;
  assign n84538 = ~n59633 ;
  assign n59634 = n59473 & n84538 ;
  assign n59635 = n59631 | n59634 ;
  assign n59636 = n74318 & n59635 ;
  assign n84539 = ~n59485 ;
  assign n59637 = n84539 & n59636 ;
  assign n59638 = n59487 | n59637 ;
  assign n59639 = n74029 & n59638 ;
  assign n84540 = ~n59637 ;
  assign n60382 = x121 & n84540 ;
  assign n84541 = ~n59487 ;
  assign n60383 = n84541 & n60382 ;
  assign n60384 = n59639 | n60383 ;
  assign n59640 = n58695 & n59486 ;
  assign n84542 = ~n59468 ;
  assign n59472 = n84542 & n59471 ;
  assign n59641 = n58705 | n59471 ;
  assign n84543 = ~n59641 ;
  assign n59642 = n59626 & n84543 ;
  assign n59643 = n59472 | n59642 ;
  assign n59644 = n74318 & n59643 ;
  assign n59645 = n84539 & n59644 ;
  assign n59646 = n59640 | n59645 ;
  assign n59647 = n74021 & n59646 ;
  assign n59648 = n58704 & n59486 ;
  assign n84544 = ~n59625 ;
  assign n59627 = n59466 & n84544 ;
  assign n59649 = n58715 | n59466 ;
  assign n84545 = ~n59649 ;
  assign n59650 = n59462 & n84545 ;
  assign n59651 = n59627 | n59650 ;
  assign n59652 = n74318 & n59651 ;
  assign n59653 = n84539 & n59652 ;
  assign n59654 = n59648 | n59653 ;
  assign n59655 = n73617 & n59654 ;
  assign n84546 = ~n59653 ;
  assign n60372 = x119 & n84546 ;
  assign n84547 = ~n59648 ;
  assign n60373 = n84547 & n60372 ;
  assign n60374 = n59655 | n60373 ;
  assign n59656 = n58714 & n59486 ;
  assign n84548 = ~n59457 ;
  assign n59461 = n84548 & n59460 ;
  assign n59657 = n58724 | n59460 ;
  assign n84549 = ~n59657 ;
  assign n59658 = n59621 & n84549 ;
  assign n59659 = n59461 | n59658 ;
  assign n59660 = n74318 & n59659 ;
  assign n59661 = n84539 & n59660 ;
  assign n59662 = n59656 | n59661 ;
  assign n59663 = n73188 & n59662 ;
  assign n59664 = n58723 & n59486 ;
  assign n84550 = ~n59620 ;
  assign n59622 = n59455 & n84550 ;
  assign n59665 = n58733 | n59455 ;
  assign n84551 = ~n59665 ;
  assign n59666 = n59451 & n84551 ;
  assign n59667 = n59622 | n59666 ;
  assign n59668 = n74318 & n59667 ;
  assign n59669 = n84539 & n59668 ;
  assign n59670 = n59664 | n59669 ;
  assign n59671 = n73177 & n59670 ;
  assign n84552 = ~n59669 ;
  assign n60362 = x117 & n84552 ;
  assign n84553 = ~n59664 ;
  assign n60363 = n84553 & n60362 ;
  assign n60364 = n59671 | n60363 ;
  assign n59672 = n58732 & n59486 ;
  assign n84554 = ~n59446 ;
  assign n59450 = n84554 & n59449 ;
  assign n59673 = n58742 | n59449 ;
  assign n84555 = ~n59673 ;
  assign n59674 = n59616 & n84555 ;
  assign n59675 = n59450 | n59674 ;
  assign n59676 = n74318 & n59675 ;
  assign n59677 = n84539 & n59676 ;
  assign n59678 = n59672 | n59677 ;
  assign n59679 = n72752 & n59678 ;
  assign n59680 = n58741 & n59486 ;
  assign n84556 = ~n59615 ;
  assign n59617 = n59444 & n84556 ;
  assign n59681 = n58751 | n59444 ;
  assign n84557 = ~n59681 ;
  assign n59682 = n59440 & n84557 ;
  assign n59683 = n59617 | n59682 ;
  assign n59684 = n74318 & n59683 ;
  assign n59685 = n84539 & n59684 ;
  assign n59686 = n59680 | n59685 ;
  assign n59687 = n72393 & n59686 ;
  assign n84558 = ~n59685 ;
  assign n60351 = x115 & n84558 ;
  assign n84559 = ~n59680 ;
  assign n60352 = n84559 & n60351 ;
  assign n60353 = n59687 | n60352 ;
  assign n59688 = n58750 & n59486 ;
  assign n84560 = ~n59435 ;
  assign n59439 = n84560 & n59438 ;
  assign n59689 = n58760 | n59438 ;
  assign n84561 = ~n59689 ;
  assign n59690 = n59611 & n84561 ;
  assign n59691 = n59439 | n59690 ;
  assign n59692 = n74318 & n59691 ;
  assign n59693 = n84539 & n59692 ;
  assign n59694 = n59688 | n59693 ;
  assign n59695 = n72385 & n59694 ;
  assign n59696 = n58759 & n59486 ;
  assign n84562 = ~n59610 ;
  assign n59612 = n59433 & n84562 ;
  assign n59697 = n58769 | n59433 ;
  assign n84563 = ~n59697 ;
  assign n59698 = n59429 & n84563 ;
  assign n59699 = n59612 | n59698 ;
  assign n59700 = n74318 & n59699 ;
  assign n59701 = n84539 & n59700 ;
  assign n59702 = n59696 | n59701 ;
  assign n59703 = n72025 & n59702 ;
  assign n84564 = ~n59701 ;
  assign n60341 = x113 & n84564 ;
  assign n84565 = ~n59696 ;
  assign n60342 = n84565 & n60341 ;
  assign n60343 = n59703 | n60342 ;
  assign n59704 = n58768 & n59486 ;
  assign n84566 = ~n59424 ;
  assign n59428 = n84566 & n59427 ;
  assign n59705 = n58778 | n59427 ;
  assign n84567 = ~n59705 ;
  assign n59706 = n59606 & n84567 ;
  assign n59707 = n59428 | n59706 ;
  assign n59708 = n74318 & n59707 ;
  assign n59709 = n84539 & n59708 ;
  assign n59710 = n59704 | n59709 ;
  assign n59711 = n71645 & n59710 ;
  assign n59712 = n58777 & n59486 ;
  assign n84568 = ~n59605 ;
  assign n59607 = n59422 & n84568 ;
  assign n59713 = n58787 | n59422 ;
  assign n84569 = ~n59713 ;
  assign n59714 = n59418 & n84569 ;
  assign n59715 = n59607 | n59714 ;
  assign n59716 = n74318 & n59715 ;
  assign n59717 = n84539 & n59716 ;
  assign n59718 = n59712 | n59717 ;
  assign n59719 = n71633 & n59718 ;
  assign n84570 = ~n59717 ;
  assign n60331 = x111 & n84570 ;
  assign n84571 = ~n59712 ;
  assign n60332 = n84571 & n60331 ;
  assign n60333 = n59719 | n60332 ;
  assign n59720 = n58786 & n59486 ;
  assign n84572 = ~n59413 ;
  assign n59417 = n84572 & n59416 ;
  assign n59721 = n58796 | n59416 ;
  assign n84573 = ~n59721 ;
  assign n59722 = n59601 & n84573 ;
  assign n59723 = n59417 | n59722 ;
  assign n59724 = n74318 & n59723 ;
  assign n59725 = n84539 & n59724 ;
  assign n59726 = n59720 | n59725 ;
  assign n59727 = n71253 & n59726 ;
  assign n59728 = n58795 & n59486 ;
  assign n84574 = ~n59600 ;
  assign n59602 = n59411 & n84574 ;
  assign n59729 = n58804 | n59411 ;
  assign n84575 = ~n59729 ;
  assign n59730 = n59407 & n84575 ;
  assign n59731 = n59602 | n59730 ;
  assign n59732 = n74318 & n59731 ;
  assign n59733 = n84539 & n59732 ;
  assign n59734 = n59728 | n59733 ;
  assign n59735 = n70935 & n59734 ;
  assign n84576 = ~n59733 ;
  assign n60320 = x109 & n84576 ;
  assign n84577 = ~n59728 ;
  assign n60321 = n84577 & n60320 ;
  assign n60322 = n59735 | n60321 ;
  assign n59736 = n58803 & n59486 ;
  assign n84578 = ~n59402 ;
  assign n59406 = n84578 & n59405 ;
  assign n59737 = n58813 | n59405 ;
  assign n84579 = ~n59737 ;
  assign n59738 = n59596 & n84579 ;
  assign n59739 = n59406 | n59738 ;
  assign n59740 = n74318 & n59739 ;
  assign n59741 = n84539 & n59740 ;
  assign n59742 = n59736 | n59741 ;
  assign n59743 = n70927 & n59742 ;
  assign n59744 = n58812 & n59486 ;
  assign n84580 = ~n59595 ;
  assign n59597 = n59400 & n84580 ;
  assign n59745 = n58822 | n59400 ;
  assign n84581 = ~n59745 ;
  assign n59746 = n59396 & n84581 ;
  assign n59747 = n59597 | n59746 ;
  assign n59748 = n74318 & n59747 ;
  assign n59749 = n84539 & n59748 ;
  assign n59750 = n59744 | n59749 ;
  assign n59751 = n70609 & n59750 ;
  assign n84582 = ~n59749 ;
  assign n60310 = x107 & n84582 ;
  assign n84583 = ~n59744 ;
  assign n60311 = n84583 & n60310 ;
  assign n60312 = n59751 | n60311 ;
  assign n59752 = n58821 & n59486 ;
  assign n84584 = ~n59391 ;
  assign n59395 = n84584 & n59394 ;
  assign n59753 = n58831 | n59394 ;
  assign n84585 = ~n59753 ;
  assign n59754 = n59591 & n84585 ;
  assign n59755 = n59395 | n59754 ;
  assign n59756 = n74318 & n59755 ;
  assign n59757 = n84539 & n59756 ;
  assign n59758 = n59752 | n59757 ;
  assign n59759 = n70276 & n59758 ;
  assign n59760 = n58830 & n59486 ;
  assign n84586 = ~n59590 ;
  assign n59592 = n59389 & n84586 ;
  assign n59761 = n58840 | n59389 ;
  assign n84587 = ~n59761 ;
  assign n59762 = n59385 & n84587 ;
  assign n59763 = n59592 | n59762 ;
  assign n59764 = n74318 & n59763 ;
  assign n59765 = n84539 & n59764 ;
  assign n59766 = n59760 | n59765 ;
  assign n59767 = n70176 & n59766 ;
  assign n84588 = ~n59765 ;
  assign n60299 = x105 & n84588 ;
  assign n84589 = ~n59760 ;
  assign n60300 = n84589 & n60299 ;
  assign n60301 = n59767 | n60300 ;
  assign n59768 = n58839 & n59486 ;
  assign n84590 = ~n59380 ;
  assign n59384 = n84590 & n59383 ;
  assign n59769 = n58849 | n59383 ;
  assign n84591 = ~n59769 ;
  assign n59770 = n59586 & n84591 ;
  assign n59771 = n59384 | n59770 ;
  assign n59772 = n74318 & n59771 ;
  assign n59773 = n84539 & n59772 ;
  assign n59774 = n59768 | n59773 ;
  assign n59775 = n69857 & n59774 ;
  assign n59776 = n58848 & n59486 ;
  assign n84592 = ~n59585 ;
  assign n59587 = n59378 & n84592 ;
  assign n59777 = n58858 | n59378 ;
  assign n84593 = ~n59777 ;
  assign n59778 = n59374 & n84593 ;
  assign n59779 = n59587 | n59778 ;
  assign n59780 = n74318 & n59779 ;
  assign n59781 = n84539 & n59780 ;
  assign n59782 = n59776 | n59781 ;
  assign n59783 = n69656 & n59782 ;
  assign n84594 = ~n59781 ;
  assign n60289 = x103 & n84594 ;
  assign n84595 = ~n59776 ;
  assign n60290 = n84595 & n60289 ;
  assign n60291 = n59783 | n60290 ;
  assign n59784 = n58857 & n59486 ;
  assign n84596 = ~n59369 ;
  assign n59373 = n84596 & n59372 ;
  assign n59785 = n58866 | n59372 ;
  assign n84597 = ~n59785 ;
  assign n59786 = n59581 & n84597 ;
  assign n59787 = n59373 | n59786 ;
  assign n59788 = n74318 & n59787 ;
  assign n59789 = n84539 & n59788 ;
  assign n59790 = n59784 | n59789 ;
  assign n59791 = n69528 & n59790 ;
  assign n59792 = n58865 & n59486 ;
  assign n84598 = ~n59580 ;
  assign n59582 = n59367 & n84598 ;
  assign n59793 = n58875 | n59367 ;
  assign n84599 = ~n59793 ;
  assign n59794 = n59363 & n84599 ;
  assign n59795 = n59582 | n59794 ;
  assign n59796 = n74318 & n59795 ;
  assign n59797 = n84539 & n59796 ;
  assign n59798 = n59792 | n59797 ;
  assign n59799 = n69261 & n59798 ;
  assign n84600 = ~n59797 ;
  assign n60278 = x101 & n84600 ;
  assign n84601 = ~n59792 ;
  assign n60279 = n84601 & n60278 ;
  assign n60280 = n59799 | n60279 ;
  assign n59800 = n58874 & n59486 ;
  assign n84602 = ~n59358 ;
  assign n59362 = n84602 & n59361 ;
  assign n59801 = n58884 | n59361 ;
  assign n84603 = ~n59801 ;
  assign n59802 = n59576 & n84603 ;
  assign n59803 = n59362 | n59802 ;
  assign n59804 = n74318 & n59803 ;
  assign n59805 = n84539 & n59804 ;
  assign n59806 = n59800 | n59805 ;
  assign n59807 = n69075 & n59806 ;
  assign n59808 = n58883 & n59486 ;
  assign n84604 = ~n59575 ;
  assign n59577 = n59356 & n84604 ;
  assign n59809 = n58893 | n59356 ;
  assign n84605 = ~n59809 ;
  assign n59810 = n59352 & n84605 ;
  assign n59811 = n59577 | n59810 ;
  assign n59812 = n74318 & n59811 ;
  assign n59813 = n84539 & n59812 ;
  assign n59814 = n59808 | n59813 ;
  assign n59815 = n68993 & n59814 ;
  assign n84606 = ~n59813 ;
  assign n60268 = x99 & n84606 ;
  assign n84607 = ~n59808 ;
  assign n60269 = n84607 & n60268 ;
  assign n60270 = n59815 | n60269 ;
  assign n59816 = n58892 & n59486 ;
  assign n84608 = ~n59347 ;
  assign n59351 = n84608 & n59350 ;
  assign n59817 = n58902 | n59350 ;
  assign n84609 = ~n59817 ;
  assign n59818 = n59571 & n84609 ;
  assign n59819 = n59351 | n59818 ;
  assign n59820 = n74318 & n59819 ;
  assign n59821 = n84539 & n59820 ;
  assign n59822 = n59816 | n59821 ;
  assign n59823 = n68716 & n59822 ;
  assign n59824 = n58901 & n59486 ;
  assign n84610 = ~n59570 ;
  assign n59572 = n59345 & n84610 ;
  assign n59825 = n58910 | n59345 ;
  assign n84611 = ~n59825 ;
  assign n59826 = n59341 & n84611 ;
  assign n59827 = n59572 | n59826 ;
  assign n59828 = n74318 & n59827 ;
  assign n59829 = n84539 & n59828 ;
  assign n59830 = n59824 | n59829 ;
  assign n59831 = n68545 & n59830 ;
  assign n84612 = ~n59829 ;
  assign n60258 = x97 & n84612 ;
  assign n84613 = ~n59824 ;
  assign n60259 = n84613 & n60258 ;
  assign n60260 = n59831 | n60259 ;
  assign n59832 = n58909 & n59486 ;
  assign n84614 = ~n59336 ;
  assign n59340 = n84614 & n59339 ;
  assign n59833 = n58919 | n59339 ;
  assign n84615 = ~n59833 ;
  assign n59834 = n59566 & n84615 ;
  assign n59835 = n59340 | n59834 ;
  assign n59836 = n74318 & n59835 ;
  assign n59837 = n84539 & n59836 ;
  assign n59838 = n59832 | n59837 ;
  assign n59839 = n68438 & n59838 ;
  assign n59840 = n58918 & n59486 ;
  assign n84616 = ~n59565 ;
  assign n59567 = n59334 & n84616 ;
  assign n59841 = n58928 | n59334 ;
  assign n84617 = ~n59841 ;
  assign n59842 = n59330 & n84617 ;
  assign n59843 = n59567 | n59842 ;
  assign n59844 = n74318 & n59843 ;
  assign n59845 = n84539 & n59844 ;
  assign n59846 = n59840 | n59845 ;
  assign n59847 = n68214 & n59846 ;
  assign n84618 = ~n59845 ;
  assign n60248 = x95 & n84618 ;
  assign n84619 = ~n59840 ;
  assign n60249 = n84619 & n60248 ;
  assign n60250 = n59847 | n60249 ;
  assign n59848 = n58927 & n59486 ;
  assign n84620 = ~n59325 ;
  assign n59329 = n84620 & n59328 ;
  assign n59849 = n58937 | n59328 ;
  assign n84621 = ~n59849 ;
  assign n59850 = n59561 & n84621 ;
  assign n59851 = n59329 | n59850 ;
  assign n59852 = n74318 & n59851 ;
  assign n59853 = n84539 & n59852 ;
  assign n59854 = n59848 | n59853 ;
  assign n59855 = n68058 & n59854 ;
  assign n59856 = n58936 & n59486 ;
  assign n84622 = ~n59560 ;
  assign n59562 = n59323 & n84622 ;
  assign n59857 = n58946 | n59323 ;
  assign n84623 = ~n59857 ;
  assign n59858 = n59319 & n84623 ;
  assign n59859 = n59562 | n59858 ;
  assign n59860 = n74318 & n59859 ;
  assign n59861 = n84539 & n59860 ;
  assign n59862 = n59856 | n59861 ;
  assign n59863 = n67986 & n59862 ;
  assign n84624 = ~n59861 ;
  assign n60238 = x93 & n84624 ;
  assign n84625 = ~n59856 ;
  assign n60239 = n84625 & n60238 ;
  assign n60240 = n59863 | n60239 ;
  assign n59864 = n58945 & n59486 ;
  assign n84626 = ~n59314 ;
  assign n59318 = n84626 & n59317 ;
  assign n59865 = n58954 | n59317 ;
  assign n84627 = ~n59865 ;
  assign n59866 = n59556 & n84627 ;
  assign n59867 = n59318 | n59866 ;
  assign n59868 = n74318 & n59867 ;
  assign n59869 = n84539 & n59868 ;
  assign n59870 = n59864 | n59869 ;
  assign n59871 = n67763 & n59870 ;
  assign n59872 = n58953 & n59486 ;
  assign n84628 = ~n59555 ;
  assign n59557 = n59312 & n84628 ;
  assign n59873 = n58963 | n59312 ;
  assign n84629 = ~n59873 ;
  assign n59874 = n59308 & n84629 ;
  assign n59875 = n59557 | n59874 ;
  assign n59876 = n74318 & n59875 ;
  assign n59877 = n84539 & n59876 ;
  assign n59878 = n59872 | n59877 ;
  assign n59879 = n67622 & n59878 ;
  assign n84630 = ~n59877 ;
  assign n60228 = x91 & n84630 ;
  assign n84631 = ~n59872 ;
  assign n60229 = n84631 & n60228 ;
  assign n60230 = n59879 | n60229 ;
  assign n59880 = n58962 & n59486 ;
  assign n84632 = ~n59303 ;
  assign n59307 = n84632 & n59306 ;
  assign n59881 = n58972 | n59306 ;
  assign n84633 = ~n59881 ;
  assign n59882 = n59551 & n84633 ;
  assign n59883 = n59307 | n59882 ;
  assign n59884 = n74318 & n59883 ;
  assign n59885 = n84539 & n59884 ;
  assign n59886 = n59880 | n59885 ;
  assign n59887 = n67531 & n59886 ;
  assign n59888 = n58971 & n59486 ;
  assign n84634 = ~n59550 ;
  assign n59552 = n59301 & n84634 ;
  assign n59889 = n58981 | n59301 ;
  assign n84635 = ~n59889 ;
  assign n59890 = n59297 & n84635 ;
  assign n59891 = n59552 | n59890 ;
  assign n59892 = n74318 & n59891 ;
  assign n59893 = n84539 & n59892 ;
  assign n59894 = n59888 | n59893 ;
  assign n59895 = n67348 & n59894 ;
  assign n84636 = ~n59893 ;
  assign n60218 = x89 & n84636 ;
  assign n84637 = ~n59888 ;
  assign n60219 = n84637 & n60218 ;
  assign n60220 = n59895 | n60219 ;
  assign n59896 = n58980 & n59486 ;
  assign n84638 = ~n59292 ;
  assign n59296 = n84638 & n59295 ;
  assign n59897 = n58990 | n59295 ;
  assign n84639 = ~n59897 ;
  assign n59898 = n59546 & n84639 ;
  assign n59899 = n59296 | n59898 ;
  assign n59900 = n74318 & n59899 ;
  assign n59901 = n84539 & n59900 ;
  assign n59902 = n59896 | n59901 ;
  assign n59903 = n67222 & n59902 ;
  assign n59904 = n58989 & n59486 ;
  assign n84640 = ~n59545 ;
  assign n59547 = n59290 & n84640 ;
  assign n59905 = n58999 | n59290 ;
  assign n84641 = ~n59905 ;
  assign n59906 = n59286 & n84641 ;
  assign n59907 = n59547 | n59906 ;
  assign n59908 = n74318 & n59907 ;
  assign n59909 = n84539 & n59908 ;
  assign n59910 = n59904 | n59909 ;
  assign n59911 = n67164 & n59910 ;
  assign n84642 = ~n59909 ;
  assign n60208 = x87 & n84642 ;
  assign n84643 = ~n59904 ;
  assign n60209 = n84643 & n60208 ;
  assign n60210 = n59911 | n60209 ;
  assign n59912 = n58998 & n59486 ;
  assign n84644 = ~n59281 ;
  assign n59285 = n84644 & n59284 ;
  assign n59913 = n59008 | n59284 ;
  assign n84645 = ~n59913 ;
  assign n59914 = n59541 & n84645 ;
  assign n59915 = n59285 | n59914 ;
  assign n59916 = n74318 & n59915 ;
  assign n59917 = n84539 & n59916 ;
  assign n59918 = n59912 | n59917 ;
  assign n59919 = n66979 & n59918 ;
  assign n59920 = n59007 & n59486 ;
  assign n84646 = ~n59540 ;
  assign n59542 = n59279 & n84646 ;
  assign n59921 = n59017 | n59279 ;
  assign n84647 = ~n59921 ;
  assign n59922 = n59275 & n84647 ;
  assign n59923 = n59542 | n59922 ;
  assign n59924 = n74318 & n59923 ;
  assign n59925 = n84539 & n59924 ;
  assign n59926 = n59920 | n59925 ;
  assign n59927 = n66868 & n59926 ;
  assign n84648 = ~n59925 ;
  assign n60198 = x85 & n84648 ;
  assign n84649 = ~n59920 ;
  assign n60199 = n84649 & n60198 ;
  assign n60200 = n59927 | n60199 ;
  assign n59928 = n59016 & n59486 ;
  assign n84650 = ~n59270 ;
  assign n59274 = n84650 & n59273 ;
  assign n59929 = n59026 | n59273 ;
  assign n84651 = ~n59929 ;
  assign n59930 = n59536 & n84651 ;
  assign n59931 = n59274 | n59930 ;
  assign n59932 = n74318 & n59931 ;
  assign n59933 = n84539 & n59932 ;
  assign n59934 = n59928 | n59933 ;
  assign n59935 = n66797 & n59934 ;
  assign n59936 = n59025 & n59486 ;
  assign n84652 = ~n59535 ;
  assign n59537 = n59268 & n84652 ;
  assign n59937 = n59035 | n59268 ;
  assign n84653 = ~n59937 ;
  assign n59938 = n59264 & n84653 ;
  assign n59939 = n59537 | n59938 ;
  assign n59940 = n74318 & n59939 ;
  assign n59941 = n84539 & n59940 ;
  assign n59942 = n59936 | n59941 ;
  assign n59943 = n66654 & n59942 ;
  assign n84654 = ~n59941 ;
  assign n60188 = x83 & n84654 ;
  assign n84655 = ~n59936 ;
  assign n60189 = n84655 & n60188 ;
  assign n60190 = n59943 | n60189 ;
  assign n59944 = n59034 & n59486 ;
  assign n84656 = ~n59259 ;
  assign n59263 = n84656 & n59262 ;
  assign n59945 = n59044 | n59262 ;
  assign n84657 = ~n59945 ;
  assign n59946 = n59531 & n84657 ;
  assign n59947 = n59263 | n59946 ;
  assign n59948 = n74318 & n59947 ;
  assign n59949 = n84539 & n59948 ;
  assign n59950 = n59944 | n59949 ;
  assign n59951 = n66560 & n59950 ;
  assign n59952 = n59043 & n59486 ;
  assign n84658 = ~n59530 ;
  assign n59532 = n59257 & n84658 ;
  assign n59953 = n59053 | n59257 ;
  assign n84659 = ~n59953 ;
  assign n59954 = n59253 & n84659 ;
  assign n59955 = n59532 | n59954 ;
  assign n59956 = n74318 & n59955 ;
  assign n59957 = n84539 & n59956 ;
  assign n59958 = n59952 | n59957 ;
  assign n59959 = n66505 & n59958 ;
  assign n84660 = ~n59957 ;
  assign n60178 = x81 & n84660 ;
  assign n84661 = ~n59952 ;
  assign n60179 = n84661 & n60178 ;
  assign n60180 = n59959 | n60179 ;
  assign n59960 = n59052 & n59486 ;
  assign n84662 = ~n59248 ;
  assign n59252 = n84662 & n59251 ;
  assign n59961 = n59062 | n59251 ;
  assign n84663 = ~n59961 ;
  assign n59962 = n59526 & n84663 ;
  assign n59963 = n59252 | n59962 ;
  assign n59964 = n74318 & n59963 ;
  assign n59965 = n84539 & n59964 ;
  assign n59966 = n59960 | n59965 ;
  assign n59967 = n66379 & n59966 ;
  assign n59968 = n59061 & n59486 ;
  assign n84664 = ~n59525 ;
  assign n59527 = n59246 & n84664 ;
  assign n59969 = n59071 | n59246 ;
  assign n84665 = ~n59969 ;
  assign n59970 = n59242 & n84665 ;
  assign n59971 = n59527 | n59970 ;
  assign n59972 = n74318 & n59971 ;
  assign n59973 = n84539 & n59972 ;
  assign n59974 = n59968 | n59973 ;
  assign n59975 = n66299 & n59974 ;
  assign n84666 = ~n59973 ;
  assign n60168 = x79 & n84666 ;
  assign n84667 = ~n59968 ;
  assign n60169 = n84667 & n60168 ;
  assign n60170 = n59975 | n60169 ;
  assign n59976 = n59070 & n59486 ;
  assign n84668 = ~n59237 ;
  assign n59241 = n84668 & n59240 ;
  assign n59977 = n59080 | n59240 ;
  assign n84669 = ~n59977 ;
  assign n59978 = n59521 & n84669 ;
  assign n59979 = n59241 | n59978 ;
  assign n59980 = n74318 & n59979 ;
  assign n59981 = n84539 & n59980 ;
  assign n59982 = n59976 | n59981 ;
  assign n59983 = n66244 & n59982 ;
  assign n59984 = n59079 & n59486 ;
  assign n84670 = ~n59520 ;
  assign n59522 = n59235 & n84670 ;
  assign n59985 = n59089 | n59235 ;
  assign n84671 = ~n59985 ;
  assign n59986 = n59231 & n84671 ;
  assign n59987 = n59522 | n59986 ;
  assign n59988 = n74318 & n59987 ;
  assign n59989 = n84539 & n59988 ;
  assign n59990 = n59984 | n59989 ;
  assign n59991 = n66145 & n59990 ;
  assign n84672 = ~n59989 ;
  assign n60157 = x77 & n84672 ;
  assign n84673 = ~n59984 ;
  assign n60158 = n84673 & n60157 ;
  assign n60159 = n59991 | n60158 ;
  assign n59992 = n59088 & n59486 ;
  assign n84674 = ~n59226 ;
  assign n59230 = n84674 & n59229 ;
  assign n59993 = n59098 | n59229 ;
  assign n84675 = ~n59993 ;
  assign n59994 = n59516 & n84675 ;
  assign n59995 = n59230 | n59994 ;
  assign n59996 = n74318 & n59995 ;
  assign n59997 = n84539 & n59996 ;
  assign n59998 = n59992 | n59997 ;
  assign n59999 = n66081 & n59998 ;
  assign n60000 = n59097 & n59486 ;
  assign n84676 = ~n59515 ;
  assign n59517 = n59224 & n84676 ;
  assign n60001 = n59107 | n59224 ;
  assign n84677 = ~n60001 ;
  assign n60002 = n59220 & n84677 ;
  assign n60003 = n59517 | n60002 ;
  assign n60004 = n74318 & n60003 ;
  assign n60005 = n84539 & n60004 ;
  assign n60006 = n60000 | n60005 ;
  assign n60007 = n66043 & n60006 ;
  assign n84678 = ~n60005 ;
  assign n60146 = x75 & n84678 ;
  assign n84679 = ~n60000 ;
  assign n60147 = n84679 & n60146 ;
  assign n60148 = n60007 | n60147 ;
  assign n60008 = n59106 & n59486 ;
  assign n84680 = ~n59215 ;
  assign n59219 = n84680 & n59218 ;
  assign n60009 = n59116 | n59218 ;
  assign n84681 = ~n60009 ;
  assign n60010 = n59511 & n84681 ;
  assign n60011 = n59219 | n60010 ;
  assign n60012 = n74318 & n60011 ;
  assign n60013 = n84539 & n60012 ;
  assign n60014 = n60008 | n60013 ;
  assign n60015 = n65960 & n60014 ;
  assign n60016 = n59115 & n59486 ;
  assign n84682 = ~n59510 ;
  assign n59512 = n59213 & n84682 ;
  assign n60017 = n59124 | n59213 ;
  assign n84683 = ~n60017 ;
  assign n60018 = n59209 & n84683 ;
  assign n60019 = n59512 | n60018 ;
  assign n60020 = n74318 & n60019 ;
  assign n60021 = n84539 & n60020 ;
  assign n60022 = n60016 | n60021 ;
  assign n60023 = n65909 & n60022 ;
  assign n84684 = ~n60021 ;
  assign n60136 = x73 & n84684 ;
  assign n84685 = ~n60016 ;
  assign n60137 = n84685 & n60136 ;
  assign n60138 = n60023 | n60137 ;
  assign n60024 = n59123 & n59486 ;
  assign n84686 = ~n59204 ;
  assign n59208 = n84686 & n59207 ;
  assign n60025 = n59202 | n59505 ;
  assign n60026 = n59133 | n59207 ;
  assign n84687 = ~n60026 ;
  assign n60027 = n60025 & n84687 ;
  assign n60028 = n59208 | n60027 ;
  assign n60029 = n74318 & n60028 ;
  assign n60030 = n84539 & n60029 ;
  assign n60031 = n60024 | n60030 ;
  assign n60032 = n65877 & n60031 ;
  assign n60033 = n59132 & n59486 ;
  assign n84688 = ~n59505 ;
  assign n59507 = n59202 & n84688 ;
  assign n60034 = n59195 | n59502 ;
  assign n60035 = n59142 | n59202 ;
  assign n84689 = ~n60035 ;
  assign n60036 = n60034 & n84689 ;
  assign n60037 = n59507 | n60036 ;
  assign n60038 = n74318 & n60037 ;
  assign n60039 = n84539 & n60038 ;
  assign n60040 = n60033 | n60039 ;
  assign n60041 = n65820 & n60040 ;
  assign n84690 = ~n60039 ;
  assign n60126 = x71 & n84690 ;
  assign n84691 = ~n60033 ;
  assign n60127 = n84691 & n60126 ;
  assign n60128 = n60041 | n60127 ;
  assign n60042 = n59141 & n59486 ;
  assign n84692 = ~n59195 ;
  assign n59503 = n84692 & n59502 ;
  assign n60043 = n59193 | n59498 ;
  assign n60044 = n59151 | n59502 ;
  assign n84693 = ~n60044 ;
  assign n60045 = n60043 & n84693 ;
  assign n60046 = n59503 | n60045 ;
  assign n60047 = n74318 & n60046 ;
  assign n60048 = n84539 & n60047 ;
  assign n60049 = n60042 | n60048 ;
  assign n60050 = n65791 & n60049 ;
  assign n60051 = n59150 & n59486 ;
  assign n84694 = ~n59498 ;
  assign n59500 = n59193 & n84694 ;
  assign n60052 = n59186 | n59495 ;
  assign n60053 = n59159 | n59193 ;
  assign n84695 = ~n60053 ;
  assign n60054 = n60052 & n84695 ;
  assign n60055 = n59500 | n60054 ;
  assign n60056 = n74318 & n60055 ;
  assign n60057 = n84539 & n60056 ;
  assign n60058 = n60051 | n60057 ;
  assign n60059 = n65772 & n60058 ;
  assign n84696 = ~n60057 ;
  assign n60116 = x69 & n84696 ;
  assign n84697 = ~n60051 ;
  assign n60117 = n84697 & n60116 ;
  assign n60118 = n60059 | n60117 ;
  assign n60060 = n59158 & n59486 ;
  assign n84698 = ~n59186 ;
  assign n59496 = n84698 & n59495 ;
  assign n60061 = n59167 | n59495 ;
  assign n84699 = ~n60061 ;
  assign n60062 = n59185 & n84699 ;
  assign n60063 = n59496 | n60062 ;
  assign n60064 = n74318 & n60063 ;
  assign n60065 = n84539 & n60064 ;
  assign n60066 = n60060 | n60065 ;
  assign n60067 = n65746 & n60066 ;
  assign n60068 = n59166 & n59486 ;
  assign n60069 = n59180 | n59184 ;
  assign n84700 = ~n60069 ;
  assign n60070 = n59491 & n84700 ;
  assign n84701 = ~n59492 ;
  assign n60071 = n59184 & n84701 ;
  assign n60072 = n60070 | n60071 ;
  assign n60073 = n74318 & n60072 ;
  assign n60074 = n84539 & n60073 ;
  assign n60075 = n60068 | n60074 ;
  assign n60076 = n65721 & n60075 ;
  assign n84702 = ~n60074 ;
  assign n60106 = x67 & n84702 ;
  assign n84703 = ~n60068 ;
  assign n60107 = n84703 & n60106 ;
  assign n60108 = n60076 | n60107 ;
  assign n60077 = n59486 & n59488 ;
  assign n60078 = n26974 & n59177 ;
  assign n60079 = n84366 & n60078 ;
  assign n60080 = n27311 | n60079 ;
  assign n84704 = ~n60080 ;
  assign n60081 = n59491 & n84704 ;
  assign n60082 = n84539 & n60081 ;
  assign n60083 = n60077 | n60082 ;
  assign n60084 = n65686 & n60083 ;
  assign n60085 = n27880 & n84539 ;
  assign n84705 = ~n60085 ;
  assign n60086 = x6 & n84705 ;
  assign n60087 = n27890 & n84539 ;
  assign n60088 = n60086 | n60087 ;
  assign n60089 = x65 & n60088 ;
  assign n59632 = n59477 | n59630 ;
  assign n60090 = n84532 & n59632 ;
  assign n60091 = n59482 | n60090 ;
  assign n60092 = n84535 & n60091 ;
  assign n84706 = ~n60092 ;
  assign n60093 = n27880 & n84706 ;
  assign n84707 = ~n60093 ;
  assign n60094 = x6 & n84707 ;
  assign n60095 = x65 | n60087 ;
  assign n60096 = n60094 | n60095 ;
  assign n84708 = ~n60089 ;
  assign n60097 = n84708 & n60096 ;
  assign n60098 = n27897 | n60097 ;
  assign n60099 = n60087 | n60094 ;
  assign n60100 = n65670 & n60099 ;
  assign n84709 = ~n60100 ;
  assign n60101 = n60098 & n84709 ;
  assign n84710 = ~n60082 ;
  assign n60102 = x66 & n84710 ;
  assign n84711 = ~n60077 ;
  assign n60103 = n84711 & n60102 ;
  assign n60104 = n60084 | n60103 ;
  assign n60105 = n60101 | n60104 ;
  assign n84712 = ~n60084 ;
  assign n60109 = n84712 & n60105 ;
  assign n60110 = n60108 | n60109 ;
  assign n84713 = ~n60076 ;
  assign n60111 = n84713 & n60110 ;
  assign n84714 = ~n60065 ;
  assign n60112 = x68 & n84714 ;
  assign n84715 = ~n60060 ;
  assign n60113 = n84715 & n60112 ;
  assign n60114 = n60067 | n60113 ;
  assign n60115 = n60111 | n60114 ;
  assign n84716 = ~n60067 ;
  assign n60119 = n84716 & n60115 ;
  assign n60120 = n60118 | n60119 ;
  assign n84717 = ~n60059 ;
  assign n60121 = n84717 & n60120 ;
  assign n84718 = ~n60048 ;
  assign n60122 = x70 & n84718 ;
  assign n84719 = ~n60042 ;
  assign n60123 = n84719 & n60122 ;
  assign n60124 = n60050 | n60123 ;
  assign n60125 = n60121 | n60124 ;
  assign n84720 = ~n60050 ;
  assign n60129 = n84720 & n60125 ;
  assign n60130 = n60128 | n60129 ;
  assign n84721 = ~n60041 ;
  assign n60131 = n84721 & n60130 ;
  assign n84722 = ~n60030 ;
  assign n60132 = x72 & n84722 ;
  assign n84723 = ~n60024 ;
  assign n60133 = n84723 & n60132 ;
  assign n60134 = n60032 | n60133 ;
  assign n60135 = n60131 | n60134 ;
  assign n84724 = ~n60032 ;
  assign n60139 = n84724 & n60135 ;
  assign n60140 = n60138 | n60139 ;
  assign n84725 = ~n60023 ;
  assign n60141 = n84725 & n60140 ;
  assign n84726 = ~n60013 ;
  assign n60142 = x74 & n84726 ;
  assign n84727 = ~n60008 ;
  assign n60143 = n84727 & n60142 ;
  assign n60144 = n60015 | n60143 ;
  assign n60145 = n60141 | n60144 ;
  assign n84728 = ~n60015 ;
  assign n60150 = n84728 & n60145 ;
  assign n60151 = n60148 | n60150 ;
  assign n84729 = ~n60007 ;
  assign n60152 = n84729 & n60151 ;
  assign n84730 = ~n59997 ;
  assign n60153 = x76 & n84730 ;
  assign n84731 = ~n59992 ;
  assign n60154 = n84731 & n60153 ;
  assign n60155 = n59999 | n60154 ;
  assign n60156 = n60152 | n60155 ;
  assign n84732 = ~n59999 ;
  assign n60161 = n84732 & n60156 ;
  assign n60162 = n60159 | n60161 ;
  assign n84733 = ~n59991 ;
  assign n60163 = n84733 & n60162 ;
  assign n84734 = ~n59981 ;
  assign n60164 = x78 & n84734 ;
  assign n84735 = ~n59976 ;
  assign n60165 = n84735 & n60164 ;
  assign n60166 = n59983 | n60165 ;
  assign n60167 = n60163 | n60166 ;
  assign n84736 = ~n59983 ;
  assign n60171 = n84736 & n60167 ;
  assign n60172 = n60170 | n60171 ;
  assign n84737 = ~n59975 ;
  assign n60173 = n84737 & n60172 ;
  assign n84738 = ~n59965 ;
  assign n60174 = x80 & n84738 ;
  assign n84739 = ~n59960 ;
  assign n60175 = n84739 & n60174 ;
  assign n60176 = n59967 | n60175 ;
  assign n60177 = n60173 | n60176 ;
  assign n84740 = ~n59967 ;
  assign n60181 = n84740 & n60177 ;
  assign n60182 = n60180 | n60181 ;
  assign n84741 = ~n59959 ;
  assign n60183 = n84741 & n60182 ;
  assign n84742 = ~n59949 ;
  assign n60184 = x82 & n84742 ;
  assign n84743 = ~n59944 ;
  assign n60185 = n84743 & n60184 ;
  assign n60186 = n59951 | n60185 ;
  assign n60187 = n60183 | n60186 ;
  assign n84744 = ~n59951 ;
  assign n60191 = n84744 & n60187 ;
  assign n60192 = n60190 | n60191 ;
  assign n84745 = ~n59943 ;
  assign n60193 = n84745 & n60192 ;
  assign n84746 = ~n59933 ;
  assign n60194 = x84 & n84746 ;
  assign n84747 = ~n59928 ;
  assign n60195 = n84747 & n60194 ;
  assign n60196 = n59935 | n60195 ;
  assign n60197 = n60193 | n60196 ;
  assign n84748 = ~n59935 ;
  assign n60201 = n84748 & n60197 ;
  assign n60202 = n60200 | n60201 ;
  assign n84749 = ~n59927 ;
  assign n60203 = n84749 & n60202 ;
  assign n84750 = ~n59917 ;
  assign n60204 = x86 & n84750 ;
  assign n84751 = ~n59912 ;
  assign n60205 = n84751 & n60204 ;
  assign n60206 = n59919 | n60205 ;
  assign n60207 = n60203 | n60206 ;
  assign n84752 = ~n59919 ;
  assign n60211 = n84752 & n60207 ;
  assign n60212 = n60210 | n60211 ;
  assign n84753 = ~n59911 ;
  assign n60213 = n84753 & n60212 ;
  assign n84754 = ~n59901 ;
  assign n60214 = x88 & n84754 ;
  assign n84755 = ~n59896 ;
  assign n60215 = n84755 & n60214 ;
  assign n60216 = n59903 | n60215 ;
  assign n60217 = n60213 | n60216 ;
  assign n84756 = ~n59903 ;
  assign n60221 = n84756 & n60217 ;
  assign n60222 = n60220 | n60221 ;
  assign n84757 = ~n59895 ;
  assign n60223 = n84757 & n60222 ;
  assign n84758 = ~n59885 ;
  assign n60224 = x90 & n84758 ;
  assign n84759 = ~n59880 ;
  assign n60225 = n84759 & n60224 ;
  assign n60226 = n59887 | n60225 ;
  assign n60227 = n60223 | n60226 ;
  assign n84760 = ~n59887 ;
  assign n60231 = n84760 & n60227 ;
  assign n60232 = n60230 | n60231 ;
  assign n84761 = ~n59879 ;
  assign n60233 = n84761 & n60232 ;
  assign n84762 = ~n59869 ;
  assign n60234 = x92 & n84762 ;
  assign n84763 = ~n59864 ;
  assign n60235 = n84763 & n60234 ;
  assign n60236 = n59871 | n60235 ;
  assign n60237 = n60233 | n60236 ;
  assign n84764 = ~n59871 ;
  assign n60241 = n84764 & n60237 ;
  assign n60242 = n60240 | n60241 ;
  assign n84765 = ~n59863 ;
  assign n60243 = n84765 & n60242 ;
  assign n84766 = ~n59853 ;
  assign n60244 = x94 & n84766 ;
  assign n84767 = ~n59848 ;
  assign n60245 = n84767 & n60244 ;
  assign n60246 = n59855 | n60245 ;
  assign n60247 = n60243 | n60246 ;
  assign n84768 = ~n59855 ;
  assign n60251 = n84768 & n60247 ;
  assign n60252 = n60250 | n60251 ;
  assign n84769 = ~n59847 ;
  assign n60253 = n84769 & n60252 ;
  assign n84770 = ~n59837 ;
  assign n60254 = x96 & n84770 ;
  assign n84771 = ~n59832 ;
  assign n60255 = n84771 & n60254 ;
  assign n60256 = n59839 | n60255 ;
  assign n60257 = n60253 | n60256 ;
  assign n84772 = ~n59839 ;
  assign n60261 = n84772 & n60257 ;
  assign n60262 = n60260 | n60261 ;
  assign n84773 = ~n59831 ;
  assign n60263 = n84773 & n60262 ;
  assign n84774 = ~n59821 ;
  assign n60264 = x98 & n84774 ;
  assign n84775 = ~n59816 ;
  assign n60265 = n84775 & n60264 ;
  assign n60266 = n59823 | n60265 ;
  assign n60267 = n60263 | n60266 ;
  assign n84776 = ~n59823 ;
  assign n60271 = n84776 & n60267 ;
  assign n60272 = n60270 | n60271 ;
  assign n84777 = ~n59815 ;
  assign n60273 = n84777 & n60272 ;
  assign n84778 = ~n59805 ;
  assign n60274 = x100 & n84778 ;
  assign n84779 = ~n59800 ;
  assign n60275 = n84779 & n60274 ;
  assign n60276 = n59807 | n60275 ;
  assign n60277 = n60273 | n60276 ;
  assign n84780 = ~n59807 ;
  assign n60281 = n84780 & n60277 ;
  assign n60282 = n60280 | n60281 ;
  assign n84781 = ~n59799 ;
  assign n60283 = n84781 & n60282 ;
  assign n84782 = ~n59789 ;
  assign n60284 = x102 & n84782 ;
  assign n84783 = ~n59784 ;
  assign n60285 = n84783 & n60284 ;
  assign n60286 = n59791 | n60285 ;
  assign n60288 = n60283 | n60286 ;
  assign n84784 = ~n59791 ;
  assign n60292 = n84784 & n60288 ;
  assign n60293 = n60291 | n60292 ;
  assign n84785 = ~n59783 ;
  assign n60294 = n84785 & n60293 ;
  assign n84786 = ~n59773 ;
  assign n60295 = x104 & n84786 ;
  assign n84787 = ~n59768 ;
  assign n60296 = n84787 & n60295 ;
  assign n60297 = n59775 | n60296 ;
  assign n60298 = n60294 | n60297 ;
  assign n84788 = ~n59775 ;
  assign n60303 = n84788 & n60298 ;
  assign n60304 = n60301 | n60303 ;
  assign n84789 = ~n59767 ;
  assign n60305 = n84789 & n60304 ;
  assign n84790 = ~n59757 ;
  assign n60306 = x106 & n84790 ;
  assign n84791 = ~n59752 ;
  assign n60307 = n84791 & n60306 ;
  assign n60308 = n59759 | n60307 ;
  assign n60309 = n60305 | n60308 ;
  assign n84792 = ~n59759 ;
  assign n60313 = n84792 & n60309 ;
  assign n60314 = n60312 | n60313 ;
  assign n84793 = ~n59751 ;
  assign n60315 = n84793 & n60314 ;
  assign n84794 = ~n59741 ;
  assign n60316 = x108 & n84794 ;
  assign n84795 = ~n59736 ;
  assign n60317 = n84795 & n60316 ;
  assign n60318 = n59743 | n60317 ;
  assign n60319 = n60315 | n60318 ;
  assign n84796 = ~n59743 ;
  assign n60323 = n84796 & n60319 ;
  assign n60324 = n60322 | n60323 ;
  assign n84797 = ~n59735 ;
  assign n60325 = n84797 & n60324 ;
  assign n84798 = ~n59725 ;
  assign n60326 = x110 & n84798 ;
  assign n84799 = ~n59720 ;
  assign n60327 = n84799 & n60326 ;
  assign n60328 = n59727 | n60327 ;
  assign n60330 = n60325 | n60328 ;
  assign n84800 = ~n59727 ;
  assign n60334 = n84800 & n60330 ;
  assign n60335 = n60333 | n60334 ;
  assign n84801 = ~n59719 ;
  assign n60336 = n84801 & n60335 ;
  assign n84802 = ~n59709 ;
  assign n60337 = x112 & n84802 ;
  assign n84803 = ~n59704 ;
  assign n60338 = n84803 & n60337 ;
  assign n60339 = n59711 | n60338 ;
  assign n60340 = n60336 | n60339 ;
  assign n84804 = ~n59711 ;
  assign n60344 = n84804 & n60340 ;
  assign n60345 = n60343 | n60344 ;
  assign n84805 = ~n59703 ;
  assign n60346 = n84805 & n60345 ;
  assign n84806 = ~n59693 ;
  assign n60347 = x114 & n84806 ;
  assign n84807 = ~n59688 ;
  assign n60348 = n84807 & n60347 ;
  assign n60349 = n59695 | n60348 ;
  assign n60350 = n60346 | n60349 ;
  assign n84808 = ~n59695 ;
  assign n60355 = n84808 & n60350 ;
  assign n60356 = n60353 | n60355 ;
  assign n84809 = ~n59687 ;
  assign n60357 = n84809 & n60356 ;
  assign n84810 = ~n59677 ;
  assign n60358 = x116 & n84810 ;
  assign n84811 = ~n59672 ;
  assign n60359 = n84811 & n60358 ;
  assign n60360 = n59679 | n60359 ;
  assign n60361 = n60357 | n60360 ;
  assign n84812 = ~n59679 ;
  assign n60365 = n84812 & n60361 ;
  assign n60366 = n60364 | n60365 ;
  assign n84813 = ~n59671 ;
  assign n60367 = n84813 & n60366 ;
  assign n84814 = ~n59661 ;
  assign n60368 = x118 & n84814 ;
  assign n84815 = ~n59656 ;
  assign n60369 = n84815 & n60368 ;
  assign n60370 = n59663 | n60369 ;
  assign n60371 = n60367 | n60370 ;
  assign n84816 = ~n59663 ;
  assign n60375 = n84816 & n60371 ;
  assign n60376 = n60374 | n60375 ;
  assign n84817 = ~n59655 ;
  assign n60377 = n84817 & n60376 ;
  assign n84818 = ~n59645 ;
  assign n60378 = x120 & n84818 ;
  assign n84819 = ~n59640 ;
  assign n60379 = n84819 & n60378 ;
  assign n60380 = n59647 | n60379 ;
  assign n60381 = n60377 | n60380 ;
  assign n84820 = ~n59647 ;
  assign n60386 = n84820 & n60381 ;
  assign n60387 = n60384 | n60386 ;
  assign n84821 = ~n59639 ;
  assign n60388 = n84821 & n60387 ;
  assign n84822 = ~n59479 ;
  assign n59483 = n84822 & n59482 ;
  assign n60389 = n58687 | n59482 ;
  assign n84823 = ~n60389 ;
  assign n60390 = n59632 & n84823 ;
  assign n60391 = n59483 | n60390 ;
  assign n60392 = n59486 | n60391 ;
  assign n84824 = ~n58685 ;
  assign n60393 = n84824 & n59486 ;
  assign n84825 = ~n60393 ;
  assign n60394 = n60392 & n84825 ;
  assign n60395 = n74431 & n60394 ;
  assign n84826 = ~n59486 ;
  assign n60396 = n84826 & n60391 ;
  assign n60397 = n58685 & n59486 ;
  assign n84827 = ~n60397 ;
  assign n60398 = x122 & n84827 ;
  assign n84828 = ~n60396 ;
  assign n60399 = n84828 & n60398 ;
  assign n60400 = n28217 | n60399 ;
  assign n60401 = n60395 | n60400 ;
  assign n60402 = n60388 | n60401 ;
  assign n60403 = n74318 & n60394 ;
  assign n84829 = ~n60403 ;
  assign n60404 = n60402 & n84829 ;
  assign n61354 = n59639 | n60399 ;
  assign n61355 = n60395 | n61354 ;
  assign n84830 = ~n61355 ;
  assign n61356 = n60387 & n84830 ;
  assign n60414 = x65 & n60099 ;
  assign n84831 = ~n60414 ;
  assign n60415 = n60096 & n84831 ;
  assign n60416 = n27897 | n60415 ;
  assign n60417 = n84709 & n60416 ;
  assign n60418 = n60104 | n60417 ;
  assign n60419 = n84712 & n60418 ;
  assign n60420 = n60108 | n60419 ;
  assign n60421 = n84713 & n60420 ;
  assign n60422 = n60114 | n60421 ;
  assign n60423 = n84716 & n60422 ;
  assign n60424 = n60118 | n60423 ;
  assign n60425 = n84717 & n60424 ;
  assign n60426 = n60124 | n60425 ;
  assign n60427 = n84720 & n60426 ;
  assign n60428 = n60128 | n60427 ;
  assign n60429 = n84721 & n60428 ;
  assign n60430 = n60134 | n60429 ;
  assign n60431 = n84724 & n60430 ;
  assign n60432 = n60138 | n60431 ;
  assign n60433 = n84725 & n60432 ;
  assign n60434 = n60144 | n60433 ;
  assign n60435 = n84728 & n60434 ;
  assign n60436 = n60148 | n60435 ;
  assign n60437 = n84729 & n60436 ;
  assign n60438 = n60155 | n60437 ;
  assign n60439 = n84732 & n60438 ;
  assign n60440 = n60159 | n60439 ;
  assign n60441 = n84733 & n60440 ;
  assign n60442 = n60166 | n60441 ;
  assign n60443 = n84736 & n60442 ;
  assign n60444 = n60170 | n60443 ;
  assign n60445 = n84737 & n60444 ;
  assign n60446 = n60176 | n60445 ;
  assign n60447 = n84740 & n60446 ;
  assign n60448 = n60180 | n60447 ;
  assign n60449 = n84741 & n60448 ;
  assign n60450 = n60186 | n60449 ;
  assign n60451 = n84744 & n60450 ;
  assign n60452 = n60190 | n60451 ;
  assign n60453 = n84745 & n60452 ;
  assign n60454 = n60196 | n60453 ;
  assign n60455 = n84748 & n60454 ;
  assign n60456 = n60200 | n60455 ;
  assign n60457 = n84749 & n60456 ;
  assign n60458 = n60206 | n60457 ;
  assign n60459 = n84752 & n60458 ;
  assign n60460 = n60210 | n60459 ;
  assign n60461 = n84753 & n60460 ;
  assign n60462 = n60216 | n60461 ;
  assign n60463 = n84756 & n60462 ;
  assign n60464 = n60220 | n60463 ;
  assign n60465 = n84757 & n60464 ;
  assign n60466 = n60226 | n60465 ;
  assign n60467 = n84760 & n60466 ;
  assign n60468 = n60230 | n60467 ;
  assign n60469 = n84761 & n60468 ;
  assign n60470 = n60236 | n60469 ;
  assign n60471 = n84764 & n60470 ;
  assign n60472 = n60240 | n60471 ;
  assign n60473 = n84765 & n60472 ;
  assign n60474 = n60246 | n60473 ;
  assign n60475 = n84768 & n60474 ;
  assign n60476 = n60250 | n60475 ;
  assign n60477 = n84769 & n60476 ;
  assign n60478 = n60256 | n60477 ;
  assign n60479 = n84772 & n60478 ;
  assign n60480 = n60260 | n60479 ;
  assign n60481 = n84773 & n60480 ;
  assign n60482 = n60266 | n60481 ;
  assign n60483 = n84776 & n60482 ;
  assign n60484 = n60270 | n60483 ;
  assign n60485 = n84777 & n60484 ;
  assign n60486 = n60276 | n60485 ;
  assign n60487 = n84780 & n60486 ;
  assign n60488 = n60280 | n60487 ;
  assign n60489 = n84781 & n60488 ;
  assign n60490 = n60286 | n60489 ;
  assign n60491 = n84784 & n60490 ;
  assign n60492 = n60291 | n60491 ;
  assign n60493 = n84785 & n60492 ;
  assign n60494 = n60297 | n60493 ;
  assign n60495 = n84788 & n60494 ;
  assign n60496 = n60301 | n60495 ;
  assign n60497 = n84789 & n60496 ;
  assign n60498 = n60308 | n60497 ;
  assign n60499 = n84792 & n60498 ;
  assign n60500 = n60312 | n60499 ;
  assign n60501 = n84793 & n60500 ;
  assign n60502 = n60318 | n60501 ;
  assign n60503 = n84796 & n60502 ;
  assign n60504 = n60322 | n60503 ;
  assign n60505 = n84797 & n60504 ;
  assign n60506 = n60328 | n60505 ;
  assign n60507 = n84800 & n60506 ;
  assign n60508 = n60333 | n60507 ;
  assign n60509 = n84801 & n60508 ;
  assign n60510 = n60339 | n60509 ;
  assign n60511 = n84804 & n60510 ;
  assign n60512 = n60343 | n60511 ;
  assign n60513 = n84805 & n60512 ;
  assign n60514 = n60349 | n60513 ;
  assign n60515 = n84808 & n60514 ;
  assign n60516 = n60353 | n60515 ;
  assign n60517 = n84809 & n60516 ;
  assign n60518 = n60360 | n60517 ;
  assign n60519 = n84812 & n60518 ;
  assign n60520 = n60364 | n60519 ;
  assign n60521 = n84813 & n60520 ;
  assign n60522 = n60370 | n60521 ;
  assign n60523 = n84816 & n60522 ;
  assign n60524 = n60374 | n60523 ;
  assign n60525 = n84817 & n60524 ;
  assign n61026 = n60380 | n60525 ;
  assign n61027 = n84820 & n61026 ;
  assign n61028 = n60384 | n61027 ;
  assign n61029 = n84821 & n61028 ;
  assign n61357 = n60395 | n60399 ;
  assign n84832 = ~n61029 ;
  assign n61358 = n84832 & n61357 ;
  assign n61359 = n61356 | n61358 ;
  assign n84833 = ~n60404 ;
  assign n61360 = n84833 & n61359 ;
  assign n61361 = n27311 & n58685 ;
  assign n61362 = n60402 & n61361 ;
  assign n61363 = n61360 | n61362 ;
  assign n61369 = n74908 & n61363 ;
  assign n84834 = ~n60386 ;
  assign n60406 = n60384 & n84834 ;
  assign n60385 = n59647 | n60384 ;
  assign n84835 = ~n60385 ;
  assign n60407 = n60381 & n84835 ;
  assign n60408 = n60406 | n60407 ;
  assign n60409 = n84833 & n60408 ;
  assign n60410 = n59638 & n84829 ;
  assign n60411 = n60402 & n60410 ;
  assign n60412 = n60409 | n60411 ;
  assign n60413 = n74431 & n60412 ;
  assign n84836 = ~n60525 ;
  assign n60526 = n60380 & n84836 ;
  assign n60527 = n59655 | n60380 ;
  assign n84837 = ~n60527 ;
  assign n60528 = n60376 & n84837 ;
  assign n60529 = n60526 | n60528 ;
  assign n60530 = n84833 & n60529 ;
  assign n60531 = n59646 & n84829 ;
  assign n60532 = n60402 & n60531 ;
  assign n60533 = n60530 | n60532 ;
  assign n60534 = n74029 & n60533 ;
  assign n84838 = ~n60375 ;
  assign n60535 = n60374 & n84838 ;
  assign n60536 = n59663 | n60374 ;
  assign n84839 = ~n60536 ;
  assign n60537 = n60522 & n84839 ;
  assign n60538 = n60535 | n60537 ;
  assign n60539 = n84833 & n60538 ;
  assign n60540 = n59654 & n84829 ;
  assign n60541 = n60402 & n60540 ;
  assign n60542 = n60539 | n60541 ;
  assign n60543 = n74021 & n60542 ;
  assign n84840 = ~n60521 ;
  assign n60544 = n60370 & n84840 ;
  assign n60545 = n59671 | n60370 ;
  assign n84841 = ~n60545 ;
  assign n60546 = n60366 & n84841 ;
  assign n60547 = n60544 | n60546 ;
  assign n60548 = n84833 & n60547 ;
  assign n60549 = n59662 & n84829 ;
  assign n60550 = n60402 & n60549 ;
  assign n60551 = n60548 | n60550 ;
  assign n60552 = n73617 & n60551 ;
  assign n84842 = ~n60365 ;
  assign n60553 = n60364 & n84842 ;
  assign n60554 = n59679 | n60364 ;
  assign n84843 = ~n60554 ;
  assign n60555 = n60518 & n84843 ;
  assign n60556 = n60553 | n60555 ;
  assign n60557 = n84833 & n60556 ;
  assign n60558 = n59670 & n84829 ;
  assign n60559 = n60402 & n60558 ;
  assign n60560 = n60557 | n60559 ;
  assign n60561 = n73188 & n60560 ;
  assign n84844 = ~n60517 ;
  assign n60562 = n60360 & n84844 ;
  assign n60563 = n59687 | n60360 ;
  assign n84845 = ~n60563 ;
  assign n60564 = n60356 & n84845 ;
  assign n60565 = n60562 | n60564 ;
  assign n60566 = n84833 & n60565 ;
  assign n60567 = n59678 & n84829 ;
  assign n60568 = n60402 & n60567 ;
  assign n60569 = n60566 | n60568 ;
  assign n60570 = n73177 & n60569 ;
  assign n84846 = ~n60355 ;
  assign n60571 = n60353 & n84846 ;
  assign n60354 = n59695 | n60353 ;
  assign n84847 = ~n60354 ;
  assign n60572 = n60350 & n84847 ;
  assign n60573 = n60571 | n60572 ;
  assign n60574 = n84833 & n60573 ;
  assign n60575 = n59686 & n84829 ;
  assign n60576 = n60402 & n60575 ;
  assign n60577 = n60574 | n60576 ;
  assign n60578 = n72752 & n60577 ;
  assign n84848 = ~n60513 ;
  assign n60579 = n60349 & n84848 ;
  assign n60580 = n59703 | n60349 ;
  assign n84849 = ~n60580 ;
  assign n60581 = n60345 & n84849 ;
  assign n60582 = n60579 | n60581 ;
  assign n60583 = n84833 & n60582 ;
  assign n60584 = n59694 & n84829 ;
  assign n60585 = n60402 & n60584 ;
  assign n60586 = n60583 | n60585 ;
  assign n60587 = n72393 & n60586 ;
  assign n84850 = ~n60344 ;
  assign n60588 = n60343 & n84850 ;
  assign n60589 = n59711 | n60343 ;
  assign n84851 = ~n60589 ;
  assign n60590 = n60510 & n84851 ;
  assign n60591 = n60588 | n60590 ;
  assign n60592 = n84833 & n60591 ;
  assign n60593 = n59702 & n84829 ;
  assign n60594 = n60402 & n60593 ;
  assign n60595 = n60592 | n60594 ;
  assign n60596 = n72385 & n60595 ;
  assign n84852 = ~n60509 ;
  assign n60597 = n60339 & n84852 ;
  assign n60598 = n59719 | n60339 ;
  assign n84853 = ~n60598 ;
  assign n60599 = n60335 & n84853 ;
  assign n60600 = n60597 | n60599 ;
  assign n60601 = n84833 & n60600 ;
  assign n60602 = n59710 & n84829 ;
  assign n60603 = n60402 & n60602 ;
  assign n60604 = n60601 | n60603 ;
  assign n60605 = n72025 & n60604 ;
  assign n84854 = ~n60334 ;
  assign n60606 = n60333 & n84854 ;
  assign n60607 = n59727 | n60333 ;
  assign n84855 = ~n60607 ;
  assign n60608 = n60506 & n84855 ;
  assign n60609 = n60606 | n60608 ;
  assign n60610 = n84833 & n60609 ;
  assign n60611 = n59718 & n84829 ;
  assign n60612 = n60402 & n60611 ;
  assign n60613 = n60610 | n60612 ;
  assign n60614 = n71645 & n60613 ;
  assign n84856 = ~n60505 ;
  assign n60615 = n60328 & n84856 ;
  assign n60329 = n59735 | n60328 ;
  assign n84857 = ~n60329 ;
  assign n60616 = n84857 & n60504 ;
  assign n60617 = n60615 | n60616 ;
  assign n60618 = n84833 & n60617 ;
  assign n60619 = n59726 & n84829 ;
  assign n60620 = n60402 & n60619 ;
  assign n60621 = n60618 | n60620 ;
  assign n60622 = n71633 & n60621 ;
  assign n84858 = ~n60323 ;
  assign n60623 = n60322 & n84858 ;
  assign n60624 = n59743 | n60322 ;
  assign n84859 = ~n60624 ;
  assign n60625 = n60502 & n84859 ;
  assign n60626 = n60623 | n60625 ;
  assign n60627 = n84833 & n60626 ;
  assign n60628 = n59734 & n84829 ;
  assign n60629 = n60402 & n60628 ;
  assign n60630 = n60627 | n60629 ;
  assign n60631 = n71253 & n60630 ;
  assign n84860 = ~n60501 ;
  assign n60632 = n60318 & n84860 ;
  assign n60633 = n59751 | n60318 ;
  assign n84861 = ~n60633 ;
  assign n60634 = n60314 & n84861 ;
  assign n60635 = n60632 | n60634 ;
  assign n60636 = n84833 & n60635 ;
  assign n60637 = n59742 & n84829 ;
  assign n60638 = n60402 & n60637 ;
  assign n60639 = n60636 | n60638 ;
  assign n60640 = n70935 & n60639 ;
  assign n84862 = ~n60313 ;
  assign n60641 = n60312 & n84862 ;
  assign n60642 = n59759 | n60312 ;
  assign n84863 = ~n60642 ;
  assign n60643 = n60498 & n84863 ;
  assign n60644 = n60641 | n60643 ;
  assign n60645 = n84833 & n60644 ;
  assign n60646 = n59750 & n84829 ;
  assign n60647 = n60402 & n60646 ;
  assign n60648 = n60645 | n60647 ;
  assign n60649 = n70927 & n60648 ;
  assign n84864 = ~n60497 ;
  assign n60650 = n60308 & n84864 ;
  assign n60651 = n59767 | n60308 ;
  assign n84865 = ~n60651 ;
  assign n60652 = n60304 & n84865 ;
  assign n60653 = n60650 | n60652 ;
  assign n60654 = n84833 & n60653 ;
  assign n60655 = n59758 & n84829 ;
  assign n60656 = n60402 & n60655 ;
  assign n60657 = n60654 | n60656 ;
  assign n60658 = n70609 & n60657 ;
  assign n84866 = ~n60303 ;
  assign n60659 = n60301 & n84866 ;
  assign n60302 = n59775 | n60301 ;
  assign n84867 = ~n60302 ;
  assign n60660 = n60298 & n84867 ;
  assign n60661 = n60659 | n60660 ;
  assign n60662 = n84833 & n60661 ;
  assign n60663 = n59766 & n84829 ;
  assign n60664 = n60402 & n60663 ;
  assign n60665 = n60662 | n60664 ;
  assign n60666 = n70276 & n60665 ;
  assign n84868 = ~n60493 ;
  assign n60667 = n60297 & n84868 ;
  assign n60668 = n59783 | n60297 ;
  assign n84869 = ~n60668 ;
  assign n60669 = n60293 & n84869 ;
  assign n60670 = n60667 | n60669 ;
  assign n60671 = n84833 & n60670 ;
  assign n60672 = n59774 & n84829 ;
  assign n60673 = n60402 & n60672 ;
  assign n60674 = n60671 | n60673 ;
  assign n60675 = n70176 & n60674 ;
  assign n84870 = ~n60292 ;
  assign n60676 = n60291 & n84870 ;
  assign n60677 = n59791 | n60291 ;
  assign n84871 = ~n60677 ;
  assign n60678 = n60490 & n84871 ;
  assign n60679 = n60676 | n60678 ;
  assign n60680 = n84833 & n60679 ;
  assign n60681 = n59782 & n84829 ;
  assign n60682 = n60402 & n60681 ;
  assign n60683 = n60680 | n60682 ;
  assign n60684 = n69857 & n60683 ;
  assign n84872 = ~n60489 ;
  assign n60685 = n60286 & n84872 ;
  assign n60287 = n59799 | n60286 ;
  assign n84873 = ~n60287 ;
  assign n60686 = n84873 & n60488 ;
  assign n60687 = n60685 | n60686 ;
  assign n60688 = n84833 & n60687 ;
  assign n60689 = n59790 & n84829 ;
  assign n60690 = n60402 & n60689 ;
  assign n60691 = n60688 | n60690 ;
  assign n60692 = n69656 & n60691 ;
  assign n84874 = ~n60281 ;
  assign n60693 = n60280 & n84874 ;
  assign n60694 = n59807 | n60280 ;
  assign n84875 = ~n60694 ;
  assign n60695 = n60486 & n84875 ;
  assign n60696 = n60693 | n60695 ;
  assign n60697 = n84833 & n60696 ;
  assign n60698 = n59798 & n84829 ;
  assign n60699 = n60402 & n60698 ;
  assign n60700 = n60697 | n60699 ;
  assign n60701 = n69528 & n60700 ;
  assign n84876 = ~n60485 ;
  assign n60702 = n60276 & n84876 ;
  assign n60703 = n59815 | n60276 ;
  assign n84877 = ~n60703 ;
  assign n60704 = n60272 & n84877 ;
  assign n60705 = n60702 | n60704 ;
  assign n60706 = n84833 & n60705 ;
  assign n60707 = n59806 & n84829 ;
  assign n60708 = n60402 & n60707 ;
  assign n60709 = n60706 | n60708 ;
  assign n60710 = n69261 & n60709 ;
  assign n84878 = ~n60271 ;
  assign n60711 = n60270 & n84878 ;
  assign n60712 = n59823 | n60270 ;
  assign n84879 = ~n60712 ;
  assign n60713 = n60482 & n84879 ;
  assign n60714 = n60711 | n60713 ;
  assign n60715 = n84833 & n60714 ;
  assign n60716 = n59814 & n84829 ;
  assign n60717 = n60402 & n60716 ;
  assign n60718 = n60715 | n60717 ;
  assign n60719 = n69075 & n60718 ;
  assign n84880 = ~n60481 ;
  assign n60720 = n60266 & n84880 ;
  assign n60721 = n59831 | n60266 ;
  assign n84881 = ~n60721 ;
  assign n60722 = n60262 & n84881 ;
  assign n60723 = n60720 | n60722 ;
  assign n60724 = n84833 & n60723 ;
  assign n60725 = n59822 & n84829 ;
  assign n60726 = n60402 & n60725 ;
  assign n60727 = n60724 | n60726 ;
  assign n60728 = n68993 & n60727 ;
  assign n84882 = ~n60261 ;
  assign n60729 = n60260 & n84882 ;
  assign n60730 = n59839 | n60260 ;
  assign n84883 = ~n60730 ;
  assign n60731 = n60478 & n84883 ;
  assign n60732 = n60729 | n60731 ;
  assign n60733 = n84833 & n60732 ;
  assign n60734 = n59830 & n84829 ;
  assign n60735 = n60402 & n60734 ;
  assign n60736 = n60733 | n60735 ;
  assign n60737 = n68716 & n60736 ;
  assign n84884 = ~n60477 ;
  assign n60738 = n60256 & n84884 ;
  assign n60739 = n59847 | n60256 ;
  assign n84885 = ~n60739 ;
  assign n60740 = n60252 & n84885 ;
  assign n60741 = n60738 | n60740 ;
  assign n60742 = n84833 & n60741 ;
  assign n60743 = n59838 & n84829 ;
  assign n60744 = n60402 & n60743 ;
  assign n60745 = n60742 | n60744 ;
  assign n60746 = n68545 & n60745 ;
  assign n84886 = ~n60251 ;
  assign n60747 = n60250 & n84886 ;
  assign n60748 = n59855 | n60250 ;
  assign n84887 = ~n60748 ;
  assign n60749 = n60474 & n84887 ;
  assign n60750 = n60747 | n60749 ;
  assign n60751 = n84833 & n60750 ;
  assign n60752 = n59846 & n84829 ;
  assign n60753 = n60402 & n60752 ;
  assign n60754 = n60751 | n60753 ;
  assign n60755 = n68438 & n60754 ;
  assign n84888 = ~n60473 ;
  assign n60756 = n60246 & n84888 ;
  assign n60757 = n59863 | n60246 ;
  assign n84889 = ~n60757 ;
  assign n60758 = n60242 & n84889 ;
  assign n60759 = n60756 | n60758 ;
  assign n60760 = n84833 & n60759 ;
  assign n60761 = n59854 & n84829 ;
  assign n60762 = n60402 & n60761 ;
  assign n60763 = n60760 | n60762 ;
  assign n60764 = n68214 & n60763 ;
  assign n84890 = ~n60241 ;
  assign n60765 = n60240 & n84890 ;
  assign n60766 = n59871 | n60240 ;
  assign n84891 = ~n60766 ;
  assign n60767 = n60470 & n84891 ;
  assign n60768 = n60765 | n60767 ;
  assign n60769 = n84833 & n60768 ;
  assign n60770 = n59862 & n84829 ;
  assign n60771 = n60402 & n60770 ;
  assign n60772 = n60769 | n60771 ;
  assign n60773 = n68058 & n60772 ;
  assign n84892 = ~n60469 ;
  assign n60774 = n60236 & n84892 ;
  assign n60775 = n59879 | n60236 ;
  assign n84893 = ~n60775 ;
  assign n60776 = n60232 & n84893 ;
  assign n60777 = n60774 | n60776 ;
  assign n60778 = n84833 & n60777 ;
  assign n60779 = n59870 & n84829 ;
  assign n60780 = n60402 & n60779 ;
  assign n60781 = n60778 | n60780 ;
  assign n60782 = n67986 & n60781 ;
  assign n84894 = ~n60231 ;
  assign n60783 = n60230 & n84894 ;
  assign n60784 = n59887 | n60230 ;
  assign n84895 = ~n60784 ;
  assign n60785 = n60466 & n84895 ;
  assign n60786 = n60783 | n60785 ;
  assign n60787 = n84833 & n60786 ;
  assign n60788 = n59878 & n84829 ;
  assign n60789 = n60402 & n60788 ;
  assign n60790 = n60787 | n60789 ;
  assign n60791 = n67763 & n60790 ;
  assign n84896 = ~n60465 ;
  assign n60792 = n60226 & n84896 ;
  assign n60793 = n59895 | n60226 ;
  assign n84897 = ~n60793 ;
  assign n60794 = n60222 & n84897 ;
  assign n60795 = n60792 | n60794 ;
  assign n60796 = n84833 & n60795 ;
  assign n60797 = n59886 & n84829 ;
  assign n60798 = n60402 & n60797 ;
  assign n60799 = n60796 | n60798 ;
  assign n60800 = n67622 & n60799 ;
  assign n84898 = ~n60221 ;
  assign n60801 = n60220 & n84898 ;
  assign n60802 = n59903 | n60220 ;
  assign n84899 = ~n60802 ;
  assign n60803 = n60462 & n84899 ;
  assign n60804 = n60801 | n60803 ;
  assign n60805 = n84833 & n60804 ;
  assign n60806 = n59894 & n84829 ;
  assign n60807 = n60402 & n60806 ;
  assign n60808 = n60805 | n60807 ;
  assign n60809 = n67531 & n60808 ;
  assign n84900 = ~n60461 ;
  assign n60810 = n60216 & n84900 ;
  assign n60811 = n59911 | n60216 ;
  assign n84901 = ~n60811 ;
  assign n60812 = n60212 & n84901 ;
  assign n60813 = n60810 | n60812 ;
  assign n60814 = n84833 & n60813 ;
  assign n60815 = n59902 & n84829 ;
  assign n60816 = n60402 & n60815 ;
  assign n60817 = n60814 | n60816 ;
  assign n60818 = n67348 & n60817 ;
  assign n84902 = ~n60211 ;
  assign n60819 = n60210 & n84902 ;
  assign n60820 = n59919 | n60210 ;
  assign n84903 = ~n60820 ;
  assign n60821 = n60458 & n84903 ;
  assign n60822 = n60819 | n60821 ;
  assign n60823 = n84833 & n60822 ;
  assign n60824 = n59910 & n84829 ;
  assign n60825 = n60402 & n60824 ;
  assign n60826 = n60823 | n60825 ;
  assign n60827 = n67222 & n60826 ;
  assign n84904 = ~n60457 ;
  assign n60828 = n60206 & n84904 ;
  assign n60829 = n59927 | n60206 ;
  assign n84905 = ~n60829 ;
  assign n60830 = n60202 & n84905 ;
  assign n60831 = n60828 | n60830 ;
  assign n60832 = n84833 & n60831 ;
  assign n60833 = n59918 & n84829 ;
  assign n60834 = n60402 & n60833 ;
  assign n60835 = n60832 | n60834 ;
  assign n60836 = n67164 & n60835 ;
  assign n84906 = ~n60201 ;
  assign n60837 = n60200 & n84906 ;
  assign n60838 = n59935 | n60200 ;
  assign n84907 = ~n60838 ;
  assign n60839 = n60454 & n84907 ;
  assign n60840 = n60837 | n60839 ;
  assign n60841 = n84833 & n60840 ;
  assign n60842 = n59926 & n84829 ;
  assign n60843 = n60402 & n60842 ;
  assign n60844 = n60841 | n60843 ;
  assign n60845 = n66979 & n60844 ;
  assign n84908 = ~n60453 ;
  assign n60846 = n60196 & n84908 ;
  assign n60847 = n59943 | n60196 ;
  assign n84909 = ~n60847 ;
  assign n60848 = n60192 & n84909 ;
  assign n60849 = n60846 | n60848 ;
  assign n60850 = n84833 & n60849 ;
  assign n60851 = n59934 & n84829 ;
  assign n60852 = n60402 & n60851 ;
  assign n60853 = n60850 | n60852 ;
  assign n60854 = n66868 & n60853 ;
  assign n84910 = ~n60191 ;
  assign n60855 = n60190 & n84910 ;
  assign n60856 = n59951 | n60190 ;
  assign n84911 = ~n60856 ;
  assign n60857 = n60450 & n84911 ;
  assign n60858 = n60855 | n60857 ;
  assign n60859 = n84833 & n60858 ;
  assign n60860 = n59942 & n84829 ;
  assign n60861 = n60402 & n60860 ;
  assign n60862 = n60859 | n60861 ;
  assign n60863 = n66797 & n60862 ;
  assign n84912 = ~n60449 ;
  assign n60864 = n60186 & n84912 ;
  assign n60865 = n59959 | n60186 ;
  assign n84913 = ~n60865 ;
  assign n60866 = n60182 & n84913 ;
  assign n60867 = n60864 | n60866 ;
  assign n60868 = n84833 & n60867 ;
  assign n60869 = n59950 & n84829 ;
  assign n60870 = n60402 & n60869 ;
  assign n60871 = n60868 | n60870 ;
  assign n60872 = n66654 & n60871 ;
  assign n84914 = ~n60181 ;
  assign n60873 = n60180 & n84914 ;
  assign n60874 = n59967 | n60180 ;
  assign n84915 = ~n60874 ;
  assign n60875 = n60446 & n84915 ;
  assign n60876 = n60873 | n60875 ;
  assign n60877 = n84833 & n60876 ;
  assign n60878 = n59958 & n84829 ;
  assign n60879 = n60402 & n60878 ;
  assign n60880 = n60877 | n60879 ;
  assign n60881 = n66560 & n60880 ;
  assign n84916 = ~n60445 ;
  assign n60882 = n60176 & n84916 ;
  assign n60883 = n59975 | n60176 ;
  assign n84917 = ~n60883 ;
  assign n60884 = n60172 & n84917 ;
  assign n60885 = n60882 | n60884 ;
  assign n60886 = n84833 & n60885 ;
  assign n60887 = n59966 & n84829 ;
  assign n60888 = n60402 & n60887 ;
  assign n60889 = n60886 | n60888 ;
  assign n60890 = n66505 & n60889 ;
  assign n84918 = ~n60171 ;
  assign n60891 = n60170 & n84918 ;
  assign n60892 = n59983 | n60170 ;
  assign n84919 = ~n60892 ;
  assign n60893 = n60442 & n84919 ;
  assign n60894 = n60891 | n60893 ;
  assign n60895 = n84833 & n60894 ;
  assign n60896 = n59974 & n84829 ;
  assign n60897 = n60402 & n60896 ;
  assign n60898 = n60895 | n60897 ;
  assign n60899 = n66379 & n60898 ;
  assign n84920 = ~n60441 ;
  assign n60900 = n60166 & n84920 ;
  assign n60901 = n59991 | n60166 ;
  assign n84921 = ~n60901 ;
  assign n60902 = n60162 & n84921 ;
  assign n60903 = n60900 | n60902 ;
  assign n60904 = n84833 & n60903 ;
  assign n60905 = n59982 & n84829 ;
  assign n60906 = n60402 & n60905 ;
  assign n60907 = n60904 | n60906 ;
  assign n60908 = n66299 & n60907 ;
  assign n84922 = ~n60161 ;
  assign n60909 = n60159 & n84922 ;
  assign n60160 = n59999 | n60159 ;
  assign n84923 = ~n60160 ;
  assign n60910 = n60156 & n84923 ;
  assign n60911 = n60909 | n60910 ;
  assign n60912 = n84833 & n60911 ;
  assign n60913 = n59990 & n84829 ;
  assign n60914 = n60402 & n60913 ;
  assign n60915 = n60912 | n60914 ;
  assign n60916 = n66244 & n60915 ;
  assign n84924 = ~n60437 ;
  assign n60917 = n60155 & n84924 ;
  assign n60918 = n60007 | n60155 ;
  assign n84925 = ~n60918 ;
  assign n60919 = n60151 & n84925 ;
  assign n60920 = n60917 | n60919 ;
  assign n60921 = n84833 & n60920 ;
  assign n60922 = n59998 & n84829 ;
  assign n60923 = n60402 & n60922 ;
  assign n60924 = n60921 | n60923 ;
  assign n60925 = n66145 & n60924 ;
  assign n84926 = ~n60150 ;
  assign n60926 = n60148 & n84926 ;
  assign n60149 = n60015 | n60148 ;
  assign n84927 = ~n60149 ;
  assign n60927 = n60145 & n84927 ;
  assign n60928 = n60926 | n60927 ;
  assign n60929 = n84833 & n60928 ;
  assign n60930 = n60006 & n84829 ;
  assign n60931 = n60402 & n60930 ;
  assign n60932 = n60929 | n60931 ;
  assign n60933 = n66081 & n60932 ;
  assign n84928 = ~n60433 ;
  assign n60934 = n60144 & n84928 ;
  assign n60935 = n60023 | n60144 ;
  assign n84929 = ~n60935 ;
  assign n60936 = n60140 & n84929 ;
  assign n60937 = n60934 | n60936 ;
  assign n60938 = n84833 & n60937 ;
  assign n60939 = n60014 & n84829 ;
  assign n60940 = n60402 & n60939 ;
  assign n60941 = n60938 | n60940 ;
  assign n60942 = n66043 & n60941 ;
  assign n84930 = ~n60139 ;
  assign n60943 = n60138 & n84930 ;
  assign n60944 = n60032 | n60138 ;
  assign n84931 = ~n60944 ;
  assign n60945 = n60430 & n84931 ;
  assign n60946 = n60943 | n60945 ;
  assign n60947 = n84833 & n60946 ;
  assign n60948 = n60022 & n84829 ;
  assign n60949 = n60402 & n60948 ;
  assign n60950 = n60947 | n60949 ;
  assign n60951 = n65960 & n60950 ;
  assign n84932 = ~n60429 ;
  assign n60952 = n60134 & n84932 ;
  assign n60953 = n60041 | n60134 ;
  assign n84933 = ~n60953 ;
  assign n60954 = n60130 & n84933 ;
  assign n60955 = n60952 | n60954 ;
  assign n60956 = n84833 & n60955 ;
  assign n60957 = n60031 & n84829 ;
  assign n60958 = n60402 & n60957 ;
  assign n60959 = n60956 | n60958 ;
  assign n60960 = n65909 & n60959 ;
  assign n84934 = ~n60129 ;
  assign n60961 = n60128 & n84934 ;
  assign n60962 = n60050 | n60128 ;
  assign n84935 = ~n60962 ;
  assign n60963 = n60426 & n84935 ;
  assign n60964 = n60961 | n60963 ;
  assign n60965 = n84833 & n60964 ;
  assign n60966 = n60040 & n84829 ;
  assign n60967 = n60402 & n60966 ;
  assign n60968 = n60965 | n60967 ;
  assign n60969 = n65877 & n60968 ;
  assign n84936 = ~n60425 ;
  assign n60970 = n60124 & n84936 ;
  assign n60971 = n60059 | n60124 ;
  assign n84937 = ~n60971 ;
  assign n60972 = n60120 & n84937 ;
  assign n60973 = n60970 | n60972 ;
  assign n60974 = n84833 & n60973 ;
  assign n60975 = n60049 & n84829 ;
  assign n60976 = n60402 & n60975 ;
  assign n60977 = n60974 | n60976 ;
  assign n60978 = n65820 & n60977 ;
  assign n84938 = ~n60119 ;
  assign n60979 = n60118 & n84938 ;
  assign n60980 = n60067 | n60118 ;
  assign n84939 = ~n60980 ;
  assign n60981 = n60422 & n84939 ;
  assign n60982 = n60979 | n60981 ;
  assign n60983 = n84833 & n60982 ;
  assign n60984 = n60058 & n84829 ;
  assign n60985 = n60402 & n60984 ;
  assign n60986 = n60983 | n60985 ;
  assign n60987 = n65791 & n60986 ;
  assign n84940 = ~n60421 ;
  assign n60989 = n60114 & n84940 ;
  assign n60988 = n60076 | n60114 ;
  assign n84941 = ~n60988 ;
  assign n60990 = n60420 & n84941 ;
  assign n60991 = n60989 | n60990 ;
  assign n60992 = n84833 & n60991 ;
  assign n60993 = n60066 & n84829 ;
  assign n60994 = n60402 & n60993 ;
  assign n60995 = n60992 | n60994 ;
  assign n60996 = n65772 & n60995 ;
  assign n84942 = ~n60109 ;
  assign n60998 = n60108 & n84942 ;
  assign n60997 = n60084 | n60108 ;
  assign n84943 = ~n60997 ;
  assign n60999 = n60105 & n84943 ;
  assign n61000 = n60998 | n60999 ;
  assign n61001 = n84833 & n61000 ;
  assign n61002 = n60075 & n84829 ;
  assign n61003 = n60402 & n61002 ;
  assign n61004 = n61001 | n61003 ;
  assign n61005 = n65746 & n61004 ;
  assign n84944 = ~n60417 ;
  assign n61007 = n60104 & n84944 ;
  assign n61006 = n60100 | n60104 ;
  assign n84945 = ~n61006 ;
  assign n61008 = n60416 & n84945 ;
  assign n61009 = n61007 | n61008 ;
  assign n61010 = n84833 & n61009 ;
  assign n61011 = n60083 & n84829 ;
  assign n61012 = n60402 & n61011 ;
  assign n61013 = n61010 | n61012 ;
  assign n61014 = n65721 & n61013 ;
  assign n61015 = n27897 & n60096 ;
  assign n61016 = n84831 & n61015 ;
  assign n84946 = ~n61016 ;
  assign n61017 = n60416 & n84946 ;
  assign n61018 = n84833 & n61017 ;
  assign n61019 = n60099 & n84829 ;
  assign n61020 = n60402 & n61019 ;
  assign n61021 = n61018 | n61020 ;
  assign n61022 = n65686 & n61021 ;
  assign n60405 = n27897 & n84833 ;
  assign n61023 = x64 & n84833 ;
  assign n84947 = ~n61023 ;
  assign n61024 = x5 & n84947 ;
  assign n61025 = n60405 | n61024 ;
  assign n61039 = n65670 & n61025 ;
  assign n61030 = n60401 | n61029 ;
  assign n61031 = n84829 & n61030 ;
  assign n84948 = ~n61031 ;
  assign n61032 = x64 & n84948 ;
  assign n84949 = ~n61032 ;
  assign n61033 = x5 & n84949 ;
  assign n61034 = n60405 | n61033 ;
  assign n61035 = x65 & n61034 ;
  assign n61036 = x65 | n60405 ;
  assign n61037 = n61033 | n61036 ;
  assign n84950 = ~n61035 ;
  assign n61038 = n84950 & n61037 ;
  assign n61040 = n28839 | n61038 ;
  assign n84951 = ~n61039 ;
  assign n61041 = n84951 & n61040 ;
  assign n84952 = ~n61020 ;
  assign n61042 = x66 & n84952 ;
  assign n84953 = ~n61018 ;
  assign n61043 = n84953 & n61042 ;
  assign n61044 = n61022 | n61043 ;
  assign n61045 = n61041 | n61044 ;
  assign n84954 = ~n61022 ;
  assign n61046 = n84954 & n61045 ;
  assign n84955 = ~n61012 ;
  assign n61047 = x67 & n84955 ;
  assign n84956 = ~n61010 ;
  assign n61048 = n84956 & n61047 ;
  assign n61049 = n61014 | n61048 ;
  assign n61050 = n61046 | n61049 ;
  assign n84957 = ~n61014 ;
  assign n61051 = n84957 & n61050 ;
  assign n84958 = ~n61003 ;
  assign n61052 = x68 & n84958 ;
  assign n84959 = ~n61001 ;
  assign n61053 = n84959 & n61052 ;
  assign n61054 = n61005 | n61053 ;
  assign n61055 = n61051 | n61054 ;
  assign n84960 = ~n61005 ;
  assign n61056 = n84960 & n61055 ;
  assign n84961 = ~n60994 ;
  assign n61057 = x69 & n84961 ;
  assign n84962 = ~n60992 ;
  assign n61058 = n84962 & n61057 ;
  assign n61059 = n60996 | n61058 ;
  assign n61060 = n61056 | n61059 ;
  assign n84963 = ~n60996 ;
  assign n61061 = n84963 & n61060 ;
  assign n84964 = ~n60985 ;
  assign n61062 = x70 & n84964 ;
  assign n84965 = ~n60983 ;
  assign n61063 = n84965 & n61062 ;
  assign n61064 = n60987 | n61063 ;
  assign n61066 = n61061 | n61064 ;
  assign n84966 = ~n60987 ;
  assign n61067 = n84966 & n61066 ;
  assign n84967 = ~n60976 ;
  assign n61068 = x71 & n84967 ;
  assign n84968 = ~n60974 ;
  assign n61069 = n84968 & n61068 ;
  assign n61070 = n60978 | n61069 ;
  assign n61071 = n61067 | n61070 ;
  assign n84969 = ~n60978 ;
  assign n61072 = n84969 & n61071 ;
  assign n84970 = ~n60967 ;
  assign n61073 = x72 & n84970 ;
  assign n84971 = ~n60965 ;
  assign n61074 = n84971 & n61073 ;
  assign n61075 = n60969 | n61074 ;
  assign n61077 = n61072 | n61075 ;
  assign n84972 = ~n60969 ;
  assign n61078 = n84972 & n61077 ;
  assign n84973 = ~n60958 ;
  assign n61079 = x73 & n84973 ;
  assign n84974 = ~n60956 ;
  assign n61080 = n84974 & n61079 ;
  assign n61081 = n60960 | n61080 ;
  assign n61082 = n61078 | n61081 ;
  assign n84975 = ~n60960 ;
  assign n61083 = n84975 & n61082 ;
  assign n84976 = ~n60949 ;
  assign n61084 = x74 & n84976 ;
  assign n84977 = ~n60947 ;
  assign n61085 = n84977 & n61084 ;
  assign n61086 = n60951 | n61085 ;
  assign n61088 = n61083 | n61086 ;
  assign n84978 = ~n60951 ;
  assign n61089 = n84978 & n61088 ;
  assign n84979 = ~n60940 ;
  assign n61090 = x75 & n84979 ;
  assign n84980 = ~n60938 ;
  assign n61091 = n84980 & n61090 ;
  assign n61092 = n60942 | n61091 ;
  assign n61093 = n61089 | n61092 ;
  assign n84981 = ~n60942 ;
  assign n61094 = n84981 & n61093 ;
  assign n84982 = ~n60931 ;
  assign n61095 = x76 & n84982 ;
  assign n84983 = ~n60929 ;
  assign n61096 = n84983 & n61095 ;
  assign n61097 = n60933 | n61096 ;
  assign n61099 = n61094 | n61097 ;
  assign n84984 = ~n60933 ;
  assign n61100 = n84984 & n61099 ;
  assign n84985 = ~n60923 ;
  assign n61101 = x77 & n84985 ;
  assign n84986 = ~n60921 ;
  assign n61102 = n84986 & n61101 ;
  assign n61103 = n60925 | n61102 ;
  assign n61104 = n61100 | n61103 ;
  assign n84987 = ~n60925 ;
  assign n61105 = n84987 & n61104 ;
  assign n84988 = ~n60914 ;
  assign n61106 = x78 & n84988 ;
  assign n84989 = ~n60912 ;
  assign n61107 = n84989 & n61106 ;
  assign n61108 = n60916 | n61107 ;
  assign n61110 = n61105 | n61108 ;
  assign n84990 = ~n60916 ;
  assign n61111 = n84990 & n61110 ;
  assign n84991 = ~n60906 ;
  assign n61112 = x79 & n84991 ;
  assign n84992 = ~n60904 ;
  assign n61113 = n84992 & n61112 ;
  assign n61114 = n60908 | n61113 ;
  assign n61115 = n61111 | n61114 ;
  assign n84993 = ~n60908 ;
  assign n61116 = n84993 & n61115 ;
  assign n84994 = ~n60897 ;
  assign n61117 = x80 & n84994 ;
  assign n84995 = ~n60895 ;
  assign n61118 = n84995 & n61117 ;
  assign n61119 = n60899 | n61118 ;
  assign n61121 = n61116 | n61119 ;
  assign n84996 = ~n60899 ;
  assign n61122 = n84996 & n61121 ;
  assign n84997 = ~n60888 ;
  assign n61123 = x81 & n84997 ;
  assign n84998 = ~n60886 ;
  assign n61124 = n84998 & n61123 ;
  assign n61125 = n60890 | n61124 ;
  assign n61126 = n61122 | n61125 ;
  assign n84999 = ~n60890 ;
  assign n61127 = n84999 & n61126 ;
  assign n85000 = ~n60879 ;
  assign n61128 = x82 & n85000 ;
  assign n85001 = ~n60877 ;
  assign n61129 = n85001 & n61128 ;
  assign n61130 = n60881 | n61129 ;
  assign n61132 = n61127 | n61130 ;
  assign n85002 = ~n60881 ;
  assign n61133 = n85002 & n61132 ;
  assign n85003 = ~n60870 ;
  assign n61134 = x83 & n85003 ;
  assign n85004 = ~n60868 ;
  assign n61135 = n85004 & n61134 ;
  assign n61136 = n60872 | n61135 ;
  assign n61137 = n61133 | n61136 ;
  assign n85005 = ~n60872 ;
  assign n61138 = n85005 & n61137 ;
  assign n85006 = ~n60861 ;
  assign n61139 = x84 & n85006 ;
  assign n85007 = ~n60859 ;
  assign n61140 = n85007 & n61139 ;
  assign n61141 = n60863 | n61140 ;
  assign n61143 = n61138 | n61141 ;
  assign n85008 = ~n60863 ;
  assign n61144 = n85008 & n61143 ;
  assign n85009 = ~n60852 ;
  assign n61145 = x85 & n85009 ;
  assign n85010 = ~n60850 ;
  assign n61146 = n85010 & n61145 ;
  assign n61147 = n60854 | n61146 ;
  assign n61148 = n61144 | n61147 ;
  assign n85011 = ~n60854 ;
  assign n61149 = n85011 & n61148 ;
  assign n85012 = ~n60843 ;
  assign n61150 = x86 & n85012 ;
  assign n85013 = ~n60841 ;
  assign n61151 = n85013 & n61150 ;
  assign n61152 = n60845 | n61151 ;
  assign n61154 = n61149 | n61152 ;
  assign n85014 = ~n60845 ;
  assign n61155 = n85014 & n61154 ;
  assign n85015 = ~n60834 ;
  assign n61156 = x87 & n85015 ;
  assign n85016 = ~n60832 ;
  assign n61157 = n85016 & n61156 ;
  assign n61158 = n60836 | n61157 ;
  assign n61159 = n61155 | n61158 ;
  assign n85017 = ~n60836 ;
  assign n61160 = n85017 & n61159 ;
  assign n85018 = ~n60825 ;
  assign n61161 = x88 & n85018 ;
  assign n85019 = ~n60823 ;
  assign n61162 = n85019 & n61161 ;
  assign n61163 = n60827 | n61162 ;
  assign n61165 = n61160 | n61163 ;
  assign n85020 = ~n60827 ;
  assign n61166 = n85020 & n61165 ;
  assign n85021 = ~n60816 ;
  assign n61167 = x89 & n85021 ;
  assign n85022 = ~n60814 ;
  assign n61168 = n85022 & n61167 ;
  assign n61169 = n60818 | n61168 ;
  assign n61170 = n61166 | n61169 ;
  assign n85023 = ~n60818 ;
  assign n61171 = n85023 & n61170 ;
  assign n85024 = ~n60807 ;
  assign n61172 = x90 & n85024 ;
  assign n85025 = ~n60805 ;
  assign n61173 = n85025 & n61172 ;
  assign n61174 = n60809 | n61173 ;
  assign n61176 = n61171 | n61174 ;
  assign n85026 = ~n60809 ;
  assign n61177 = n85026 & n61176 ;
  assign n85027 = ~n60798 ;
  assign n61178 = x91 & n85027 ;
  assign n85028 = ~n60796 ;
  assign n61179 = n85028 & n61178 ;
  assign n61180 = n60800 | n61179 ;
  assign n61181 = n61177 | n61180 ;
  assign n85029 = ~n60800 ;
  assign n61182 = n85029 & n61181 ;
  assign n85030 = ~n60789 ;
  assign n61183 = x92 & n85030 ;
  assign n85031 = ~n60787 ;
  assign n61184 = n85031 & n61183 ;
  assign n61185 = n60791 | n61184 ;
  assign n61187 = n61182 | n61185 ;
  assign n85032 = ~n60791 ;
  assign n61188 = n85032 & n61187 ;
  assign n85033 = ~n60780 ;
  assign n61189 = x93 & n85033 ;
  assign n85034 = ~n60778 ;
  assign n61190 = n85034 & n61189 ;
  assign n61191 = n60782 | n61190 ;
  assign n61192 = n61188 | n61191 ;
  assign n85035 = ~n60782 ;
  assign n61193 = n85035 & n61192 ;
  assign n85036 = ~n60771 ;
  assign n61194 = x94 & n85036 ;
  assign n85037 = ~n60769 ;
  assign n61195 = n85037 & n61194 ;
  assign n61196 = n60773 | n61195 ;
  assign n61198 = n61193 | n61196 ;
  assign n85038 = ~n60773 ;
  assign n61199 = n85038 & n61198 ;
  assign n85039 = ~n60762 ;
  assign n61200 = x95 & n85039 ;
  assign n85040 = ~n60760 ;
  assign n61201 = n85040 & n61200 ;
  assign n61202 = n60764 | n61201 ;
  assign n61203 = n61199 | n61202 ;
  assign n85041 = ~n60764 ;
  assign n61204 = n85041 & n61203 ;
  assign n85042 = ~n60753 ;
  assign n61205 = x96 & n85042 ;
  assign n85043 = ~n60751 ;
  assign n61206 = n85043 & n61205 ;
  assign n61207 = n60755 | n61206 ;
  assign n61209 = n61204 | n61207 ;
  assign n85044 = ~n60755 ;
  assign n61210 = n85044 & n61209 ;
  assign n85045 = ~n60744 ;
  assign n61211 = x97 & n85045 ;
  assign n85046 = ~n60742 ;
  assign n61212 = n85046 & n61211 ;
  assign n61213 = n60746 | n61212 ;
  assign n61214 = n61210 | n61213 ;
  assign n85047 = ~n60746 ;
  assign n61215 = n85047 & n61214 ;
  assign n85048 = ~n60735 ;
  assign n61216 = x98 & n85048 ;
  assign n85049 = ~n60733 ;
  assign n61217 = n85049 & n61216 ;
  assign n61218 = n60737 | n61217 ;
  assign n61220 = n61215 | n61218 ;
  assign n85050 = ~n60737 ;
  assign n61221 = n85050 & n61220 ;
  assign n85051 = ~n60726 ;
  assign n61222 = x99 & n85051 ;
  assign n85052 = ~n60724 ;
  assign n61223 = n85052 & n61222 ;
  assign n61224 = n60728 | n61223 ;
  assign n61225 = n61221 | n61224 ;
  assign n85053 = ~n60728 ;
  assign n61226 = n85053 & n61225 ;
  assign n85054 = ~n60717 ;
  assign n61227 = x100 & n85054 ;
  assign n85055 = ~n60715 ;
  assign n61228 = n85055 & n61227 ;
  assign n61229 = n60719 | n61228 ;
  assign n61231 = n61226 | n61229 ;
  assign n85056 = ~n60719 ;
  assign n61232 = n85056 & n61231 ;
  assign n85057 = ~n60708 ;
  assign n61233 = x101 & n85057 ;
  assign n85058 = ~n60706 ;
  assign n61234 = n85058 & n61233 ;
  assign n61235 = n60710 | n61234 ;
  assign n61236 = n61232 | n61235 ;
  assign n85059 = ~n60710 ;
  assign n61237 = n85059 & n61236 ;
  assign n85060 = ~n60699 ;
  assign n61238 = x102 & n85060 ;
  assign n85061 = ~n60697 ;
  assign n61239 = n85061 & n61238 ;
  assign n61240 = n60701 | n61239 ;
  assign n61242 = n61237 | n61240 ;
  assign n85062 = ~n60701 ;
  assign n61243 = n85062 & n61242 ;
  assign n85063 = ~n60690 ;
  assign n61244 = x103 & n85063 ;
  assign n85064 = ~n60688 ;
  assign n61245 = n85064 & n61244 ;
  assign n61246 = n60692 | n61245 ;
  assign n61247 = n61243 | n61246 ;
  assign n85065 = ~n60692 ;
  assign n61248 = n85065 & n61247 ;
  assign n85066 = ~n60682 ;
  assign n61249 = x104 & n85066 ;
  assign n85067 = ~n60680 ;
  assign n61250 = n85067 & n61249 ;
  assign n61251 = n60684 | n61250 ;
  assign n61253 = n61248 | n61251 ;
  assign n85068 = ~n60684 ;
  assign n61254 = n85068 & n61253 ;
  assign n85069 = ~n60673 ;
  assign n61255 = x105 & n85069 ;
  assign n85070 = ~n60671 ;
  assign n61256 = n85070 & n61255 ;
  assign n61257 = n60675 | n61256 ;
  assign n61258 = n61254 | n61257 ;
  assign n85071 = ~n60675 ;
  assign n61259 = n85071 & n61258 ;
  assign n85072 = ~n60664 ;
  assign n61260 = x106 & n85072 ;
  assign n85073 = ~n60662 ;
  assign n61261 = n85073 & n61260 ;
  assign n61262 = n60666 | n61261 ;
  assign n61264 = n61259 | n61262 ;
  assign n85074 = ~n60666 ;
  assign n61265 = n85074 & n61264 ;
  assign n85075 = ~n60656 ;
  assign n61266 = x107 & n85075 ;
  assign n85076 = ~n60654 ;
  assign n61267 = n85076 & n61266 ;
  assign n61268 = n60658 | n61267 ;
  assign n61269 = n61265 | n61268 ;
  assign n85077 = ~n60658 ;
  assign n61270 = n85077 & n61269 ;
  assign n85078 = ~n60647 ;
  assign n61271 = x108 & n85078 ;
  assign n85079 = ~n60645 ;
  assign n61272 = n85079 & n61271 ;
  assign n61273 = n60649 | n61272 ;
  assign n61275 = n61270 | n61273 ;
  assign n85080 = ~n60649 ;
  assign n61276 = n85080 & n61275 ;
  assign n85081 = ~n60638 ;
  assign n61277 = x109 & n85081 ;
  assign n85082 = ~n60636 ;
  assign n61278 = n85082 & n61277 ;
  assign n61279 = n60640 | n61278 ;
  assign n61280 = n61276 | n61279 ;
  assign n85083 = ~n60640 ;
  assign n61281 = n85083 & n61280 ;
  assign n85084 = ~n60629 ;
  assign n61282 = x110 & n85084 ;
  assign n85085 = ~n60627 ;
  assign n61283 = n85085 & n61282 ;
  assign n61284 = n60631 | n61283 ;
  assign n61286 = n61281 | n61284 ;
  assign n85086 = ~n60631 ;
  assign n61287 = n85086 & n61286 ;
  assign n85087 = ~n60620 ;
  assign n61288 = x111 & n85087 ;
  assign n85088 = ~n60618 ;
  assign n61289 = n85088 & n61288 ;
  assign n61290 = n60622 | n61289 ;
  assign n61291 = n61287 | n61290 ;
  assign n85089 = ~n60622 ;
  assign n61292 = n85089 & n61291 ;
  assign n85090 = ~n60612 ;
  assign n61293 = x112 & n85090 ;
  assign n85091 = ~n60610 ;
  assign n61294 = n85091 & n61293 ;
  assign n61295 = n60614 | n61294 ;
  assign n61297 = n61292 | n61295 ;
  assign n85092 = ~n60614 ;
  assign n61298 = n85092 & n61297 ;
  assign n85093 = ~n60603 ;
  assign n61299 = x113 & n85093 ;
  assign n85094 = ~n60601 ;
  assign n61300 = n85094 & n61299 ;
  assign n61301 = n60605 | n61300 ;
  assign n61302 = n61298 | n61301 ;
  assign n85095 = ~n60605 ;
  assign n61303 = n85095 & n61302 ;
  assign n85096 = ~n60594 ;
  assign n61304 = x114 & n85096 ;
  assign n85097 = ~n60592 ;
  assign n61305 = n85097 & n61304 ;
  assign n61306 = n60596 | n61305 ;
  assign n61308 = n61303 | n61306 ;
  assign n85098 = ~n60596 ;
  assign n61309 = n85098 & n61308 ;
  assign n85099 = ~n60585 ;
  assign n61310 = x115 & n85099 ;
  assign n85100 = ~n60583 ;
  assign n61311 = n85100 & n61310 ;
  assign n61312 = n60587 | n61311 ;
  assign n61313 = n61309 | n61312 ;
  assign n85101 = ~n60587 ;
  assign n61314 = n85101 & n61313 ;
  assign n85102 = ~n60576 ;
  assign n61315 = x116 & n85102 ;
  assign n85103 = ~n60574 ;
  assign n61316 = n85103 & n61315 ;
  assign n61317 = n60578 | n61316 ;
  assign n61319 = n61314 | n61317 ;
  assign n85104 = ~n60578 ;
  assign n61320 = n85104 & n61319 ;
  assign n85105 = ~n60568 ;
  assign n61321 = x117 & n85105 ;
  assign n85106 = ~n60566 ;
  assign n61322 = n85106 & n61321 ;
  assign n61323 = n60570 | n61322 ;
  assign n61324 = n61320 | n61323 ;
  assign n85107 = ~n60570 ;
  assign n61325 = n85107 & n61324 ;
  assign n85108 = ~n60559 ;
  assign n61326 = x118 & n85108 ;
  assign n85109 = ~n60557 ;
  assign n61327 = n85109 & n61326 ;
  assign n61328 = n60561 | n61327 ;
  assign n61330 = n61325 | n61328 ;
  assign n85110 = ~n60561 ;
  assign n61331 = n85110 & n61330 ;
  assign n85111 = ~n60550 ;
  assign n61332 = x119 & n85111 ;
  assign n85112 = ~n60548 ;
  assign n61333 = n85112 & n61332 ;
  assign n61334 = n60552 | n61333 ;
  assign n61335 = n61331 | n61334 ;
  assign n85113 = ~n60552 ;
  assign n61336 = n85113 & n61335 ;
  assign n85114 = ~n60541 ;
  assign n61337 = x120 & n85114 ;
  assign n85115 = ~n60539 ;
  assign n61338 = n85115 & n61337 ;
  assign n61339 = n60543 | n61338 ;
  assign n61341 = n61336 | n61339 ;
  assign n85116 = ~n60543 ;
  assign n61342 = n85116 & n61341 ;
  assign n85117 = ~n60532 ;
  assign n61343 = x121 & n85117 ;
  assign n85118 = ~n60530 ;
  assign n61344 = n85118 & n61343 ;
  assign n61345 = n60534 | n61344 ;
  assign n61346 = n61342 | n61345 ;
  assign n85119 = ~n60534 ;
  assign n61347 = n85119 & n61346 ;
  assign n85120 = ~n60411 ;
  assign n61348 = x122 & n85120 ;
  assign n85121 = ~n60409 ;
  assign n61349 = n85121 & n61348 ;
  assign n61350 = n60413 | n61349 ;
  assign n61352 = n61347 | n61350 ;
  assign n85122 = ~n60413 ;
  assign n61353 = n85122 & n61352 ;
  assign n61364 = n74905 & n61363 ;
  assign n85123 = ~n61362 ;
  assign n61365 = x123 & n85123 ;
  assign n85124 = ~n61360 ;
  assign n61366 = n85124 & n61365 ;
  assign n61367 = n65369 | n61366 ;
  assign n61368 = n61364 | n61367 ;
  assign n61370 = n61353 | n61368 ;
  assign n85125 = ~n61369 ;
  assign n61371 = n85125 & n61370 ;
  assign n85126 = ~n61347 ;
  assign n61351 = n85126 & n61350 ;
  assign n61374 = x65 & n61025 ;
  assign n85127 = ~n61374 ;
  assign n61375 = n61037 & n85127 ;
  assign n61376 = n28839 | n61375 ;
  assign n61377 = n84951 & n61376 ;
  assign n61378 = n61044 | n61377 ;
  assign n61379 = n84954 & n61378 ;
  assign n61381 = n61049 | n61379 ;
  assign n61382 = n84957 & n61381 ;
  assign n61384 = n61054 | n61382 ;
  assign n61385 = n84960 & n61384 ;
  assign n61386 = n61059 | n61385 ;
  assign n61388 = n84963 & n61386 ;
  assign n61389 = n61064 | n61388 ;
  assign n61390 = n84966 & n61389 ;
  assign n61391 = n61070 | n61390 ;
  assign n61393 = n84969 & n61391 ;
  assign n61394 = n61075 | n61393 ;
  assign n61395 = n84972 & n61394 ;
  assign n61396 = n61081 | n61395 ;
  assign n61398 = n84975 & n61396 ;
  assign n61399 = n61086 | n61398 ;
  assign n61400 = n84978 & n61399 ;
  assign n61401 = n61092 | n61400 ;
  assign n61403 = n84981 & n61401 ;
  assign n61404 = n61097 | n61403 ;
  assign n61405 = n84984 & n61404 ;
  assign n61406 = n61103 | n61405 ;
  assign n61408 = n84987 & n61406 ;
  assign n61409 = n61108 | n61408 ;
  assign n61410 = n84990 & n61409 ;
  assign n61411 = n61114 | n61410 ;
  assign n61413 = n84993 & n61411 ;
  assign n61414 = n61119 | n61413 ;
  assign n61415 = n84996 & n61414 ;
  assign n61416 = n61125 | n61415 ;
  assign n61418 = n84999 & n61416 ;
  assign n61419 = n61130 | n61418 ;
  assign n61420 = n85002 & n61419 ;
  assign n61421 = n61136 | n61420 ;
  assign n61423 = n85005 & n61421 ;
  assign n61424 = n61141 | n61423 ;
  assign n61425 = n85008 & n61424 ;
  assign n61426 = n61147 | n61425 ;
  assign n61428 = n85011 & n61426 ;
  assign n61429 = n61152 | n61428 ;
  assign n61430 = n85014 & n61429 ;
  assign n61431 = n61158 | n61430 ;
  assign n61433 = n85017 & n61431 ;
  assign n61434 = n61163 | n61433 ;
  assign n61435 = n85020 & n61434 ;
  assign n61436 = n61169 | n61435 ;
  assign n61438 = n85023 & n61436 ;
  assign n61439 = n61174 | n61438 ;
  assign n61440 = n85026 & n61439 ;
  assign n61441 = n61180 | n61440 ;
  assign n61443 = n85029 & n61441 ;
  assign n61444 = n61185 | n61443 ;
  assign n61445 = n85032 & n61444 ;
  assign n61446 = n61191 | n61445 ;
  assign n61448 = n85035 & n61446 ;
  assign n61449 = n61196 | n61448 ;
  assign n61450 = n85038 & n61449 ;
  assign n61451 = n61202 | n61450 ;
  assign n61453 = n85041 & n61451 ;
  assign n61454 = n61207 | n61453 ;
  assign n61455 = n85044 & n61454 ;
  assign n61456 = n61213 | n61455 ;
  assign n61458 = n85047 & n61456 ;
  assign n61459 = n61218 | n61458 ;
  assign n61460 = n85050 & n61459 ;
  assign n61461 = n61224 | n61460 ;
  assign n61463 = n85053 & n61461 ;
  assign n61464 = n61229 | n61463 ;
  assign n61465 = n85056 & n61464 ;
  assign n61466 = n61235 | n61465 ;
  assign n61468 = n85059 & n61466 ;
  assign n61469 = n61240 | n61468 ;
  assign n61470 = n85062 & n61469 ;
  assign n61471 = n61246 | n61470 ;
  assign n61473 = n85065 & n61471 ;
  assign n61474 = n61251 | n61473 ;
  assign n61475 = n85068 & n61474 ;
  assign n61476 = n61257 | n61475 ;
  assign n61478 = n85071 & n61476 ;
  assign n61479 = n61262 | n61478 ;
  assign n61480 = n85074 & n61479 ;
  assign n61481 = n61268 | n61480 ;
  assign n61483 = n85077 & n61481 ;
  assign n61484 = n61273 | n61483 ;
  assign n61485 = n85080 & n61484 ;
  assign n61486 = n61279 | n61485 ;
  assign n61488 = n85083 & n61486 ;
  assign n61489 = n61284 | n61488 ;
  assign n61490 = n85086 & n61489 ;
  assign n61491 = n61290 | n61490 ;
  assign n61493 = n85089 & n61491 ;
  assign n61494 = n61295 | n61493 ;
  assign n61495 = n85092 & n61494 ;
  assign n61496 = n61301 | n61495 ;
  assign n61498 = n85095 & n61496 ;
  assign n61499 = n61306 | n61498 ;
  assign n61500 = n85098 & n61499 ;
  assign n61501 = n61312 | n61500 ;
  assign n61503 = n85101 & n61501 ;
  assign n61504 = n61317 | n61503 ;
  assign n61505 = n85104 & n61504 ;
  assign n61506 = n61323 | n61505 ;
  assign n61508 = n85107 & n61506 ;
  assign n61509 = n61328 | n61508 ;
  assign n61510 = n85110 & n61509 ;
  assign n61511 = n61334 | n61510 ;
  assign n61513 = n85113 & n61511 ;
  assign n61514 = n61339 | n61513 ;
  assign n61515 = n85116 & n61514 ;
  assign n61516 = n61345 | n61515 ;
  assign n61518 = n60534 | n61350 ;
  assign n85128 = ~n61518 ;
  assign n61519 = n61516 & n85128 ;
  assign n61520 = n61351 | n61519 ;
  assign n85129 = ~n61371 ;
  assign n61521 = n85129 & n61520 ;
  assign n61522 = n85119 & n61516 ;
  assign n61523 = n61350 | n61522 ;
  assign n61524 = n85122 & n61523 ;
  assign n61525 = n61368 | n61524 ;
  assign n61526 = n60412 & n85125 ;
  assign n61527 = n61525 & n61526 ;
  assign n61528 = n61521 | n61527 ;
  assign n61529 = n74905 & n61528 ;
  assign n85130 = ~n61527 ;
  assign n62290 = x123 & n85130 ;
  assign n85131 = ~n61521 ;
  assign n62291 = n85131 & n62290 ;
  assign n62292 = n61529 | n62291 ;
  assign n85132 = ~n61515 ;
  assign n61517 = n61345 & n85132 ;
  assign n61530 = n60543 | n61345 ;
  assign n85133 = ~n61530 ;
  assign n61531 = n61341 & n85133 ;
  assign n61532 = n61517 | n61531 ;
  assign n61533 = n85129 & n61532 ;
  assign n61534 = n60533 & n85125 ;
  assign n61535 = n61525 & n61534 ;
  assign n61536 = n61533 | n61535 ;
  assign n61537 = n74431 & n61536 ;
  assign n85134 = ~n61336 ;
  assign n61340 = n85134 & n61339 ;
  assign n61538 = n60552 | n61339 ;
  assign n85135 = ~n61538 ;
  assign n61539 = n61511 & n85135 ;
  assign n61540 = n61340 | n61539 ;
  assign n61541 = n85129 & n61540 ;
  assign n61542 = n60542 & n85125 ;
  assign n61543 = n61525 & n61542 ;
  assign n61544 = n61541 | n61543 ;
  assign n61545 = n74029 & n61544 ;
  assign n85136 = ~n61543 ;
  assign n62279 = x121 & n85136 ;
  assign n85137 = ~n61541 ;
  assign n62280 = n85137 & n62279 ;
  assign n62281 = n61545 | n62280 ;
  assign n85138 = ~n61510 ;
  assign n61512 = n61334 & n85138 ;
  assign n61546 = n60561 | n61334 ;
  assign n85139 = ~n61546 ;
  assign n61547 = n61330 & n85139 ;
  assign n61548 = n61512 | n61547 ;
  assign n61549 = n85129 & n61548 ;
  assign n61550 = n60551 & n85125 ;
  assign n61551 = n61525 & n61550 ;
  assign n61552 = n61549 | n61551 ;
  assign n61553 = n74021 & n61552 ;
  assign n85140 = ~n61325 ;
  assign n61329 = n85140 & n61328 ;
  assign n61554 = n60570 | n61328 ;
  assign n85141 = ~n61554 ;
  assign n61555 = n61506 & n85141 ;
  assign n61556 = n61329 | n61555 ;
  assign n61557 = n85129 & n61556 ;
  assign n61558 = n60560 & n85125 ;
  assign n61559 = n61525 & n61558 ;
  assign n61560 = n61557 | n61559 ;
  assign n61561 = n73617 & n61560 ;
  assign n85142 = ~n61559 ;
  assign n62268 = x119 & n85142 ;
  assign n85143 = ~n61557 ;
  assign n62269 = n85143 & n62268 ;
  assign n62270 = n61561 | n62269 ;
  assign n85144 = ~n61505 ;
  assign n61507 = n61323 & n85144 ;
  assign n61562 = n60578 | n61323 ;
  assign n85145 = ~n61562 ;
  assign n61563 = n61319 & n85145 ;
  assign n61564 = n61507 | n61563 ;
  assign n61565 = n85129 & n61564 ;
  assign n61566 = n60569 & n85125 ;
  assign n61567 = n61525 & n61566 ;
  assign n61568 = n61565 | n61567 ;
  assign n61569 = n73188 & n61568 ;
  assign n85146 = ~n61314 ;
  assign n61318 = n85146 & n61317 ;
  assign n61570 = n60587 | n61317 ;
  assign n85147 = ~n61570 ;
  assign n61571 = n61501 & n85147 ;
  assign n61572 = n61318 | n61571 ;
  assign n61573 = n85129 & n61572 ;
  assign n61574 = n60577 & n85125 ;
  assign n61575 = n61525 & n61574 ;
  assign n61576 = n61573 | n61575 ;
  assign n61577 = n73177 & n61576 ;
  assign n85148 = ~n61575 ;
  assign n62258 = x117 & n85148 ;
  assign n85149 = ~n61573 ;
  assign n62259 = n85149 & n62258 ;
  assign n62260 = n61577 | n62259 ;
  assign n85150 = ~n61500 ;
  assign n61502 = n61312 & n85150 ;
  assign n61578 = n60596 | n61312 ;
  assign n85151 = ~n61578 ;
  assign n61579 = n61308 & n85151 ;
  assign n61580 = n61502 | n61579 ;
  assign n61581 = n85129 & n61580 ;
  assign n61582 = n60586 & n85125 ;
  assign n61583 = n61525 & n61582 ;
  assign n61584 = n61581 | n61583 ;
  assign n61585 = n72752 & n61584 ;
  assign n85152 = ~n61303 ;
  assign n61307 = n85152 & n61306 ;
  assign n61586 = n60605 | n61306 ;
  assign n85153 = ~n61586 ;
  assign n61587 = n61496 & n85153 ;
  assign n61588 = n61307 | n61587 ;
  assign n61589 = n85129 & n61588 ;
  assign n61590 = n60595 & n85125 ;
  assign n61591 = n61525 & n61590 ;
  assign n61592 = n61589 | n61591 ;
  assign n61593 = n72393 & n61592 ;
  assign n85154 = ~n61591 ;
  assign n62248 = x115 & n85154 ;
  assign n85155 = ~n61589 ;
  assign n62249 = n85155 & n62248 ;
  assign n62250 = n61593 | n62249 ;
  assign n85156 = ~n61495 ;
  assign n61497 = n61301 & n85156 ;
  assign n61594 = n60614 | n61301 ;
  assign n85157 = ~n61594 ;
  assign n61595 = n61297 & n85157 ;
  assign n61596 = n61497 | n61595 ;
  assign n61597 = n85129 & n61596 ;
  assign n61598 = n60604 & n85125 ;
  assign n61599 = n61525 & n61598 ;
  assign n61600 = n61597 | n61599 ;
  assign n61601 = n72385 & n61600 ;
  assign n85158 = ~n61292 ;
  assign n61296 = n85158 & n61295 ;
  assign n61602 = n60622 | n61295 ;
  assign n85159 = ~n61602 ;
  assign n61603 = n61491 & n85159 ;
  assign n61604 = n61296 | n61603 ;
  assign n61605 = n85129 & n61604 ;
  assign n61606 = n60613 & n85125 ;
  assign n61607 = n61525 & n61606 ;
  assign n61608 = n61605 | n61607 ;
  assign n61609 = n72025 & n61608 ;
  assign n85160 = ~n61607 ;
  assign n62238 = x113 & n85160 ;
  assign n85161 = ~n61605 ;
  assign n62239 = n85161 & n62238 ;
  assign n62240 = n61609 | n62239 ;
  assign n85162 = ~n61490 ;
  assign n61492 = n61290 & n85162 ;
  assign n61610 = n60631 | n61290 ;
  assign n85163 = ~n61610 ;
  assign n61611 = n61286 & n85163 ;
  assign n61612 = n61492 | n61611 ;
  assign n61613 = n85129 & n61612 ;
  assign n61614 = n60621 & n85125 ;
  assign n61615 = n61525 & n61614 ;
  assign n61616 = n61613 | n61615 ;
  assign n61617 = n71645 & n61616 ;
  assign n85164 = ~n61281 ;
  assign n61285 = n85164 & n61284 ;
  assign n61618 = n60640 | n61284 ;
  assign n85165 = ~n61618 ;
  assign n61619 = n61486 & n85165 ;
  assign n61620 = n61285 | n61619 ;
  assign n61621 = n85129 & n61620 ;
  assign n61622 = n60630 & n85125 ;
  assign n61623 = n61525 & n61622 ;
  assign n61624 = n61621 | n61623 ;
  assign n61625 = n71633 & n61624 ;
  assign n85166 = ~n61623 ;
  assign n62228 = x111 & n85166 ;
  assign n85167 = ~n61621 ;
  assign n62229 = n85167 & n62228 ;
  assign n62230 = n61625 | n62229 ;
  assign n85168 = ~n61485 ;
  assign n61487 = n61279 & n85168 ;
  assign n61626 = n60649 | n61279 ;
  assign n85169 = ~n61626 ;
  assign n61627 = n61275 & n85169 ;
  assign n61628 = n61487 | n61627 ;
  assign n61629 = n85129 & n61628 ;
  assign n61630 = n60639 & n85125 ;
  assign n61631 = n61525 & n61630 ;
  assign n61632 = n61629 | n61631 ;
  assign n61633 = n71253 & n61632 ;
  assign n85170 = ~n61270 ;
  assign n61274 = n85170 & n61273 ;
  assign n61634 = n60658 | n61273 ;
  assign n85171 = ~n61634 ;
  assign n61635 = n61481 & n85171 ;
  assign n61636 = n61274 | n61635 ;
  assign n61637 = n85129 & n61636 ;
  assign n61638 = n60648 & n85125 ;
  assign n61639 = n61525 & n61638 ;
  assign n61640 = n61637 | n61639 ;
  assign n61641 = n70935 & n61640 ;
  assign n85172 = ~n61639 ;
  assign n62218 = x109 & n85172 ;
  assign n85173 = ~n61637 ;
  assign n62219 = n85173 & n62218 ;
  assign n62220 = n61641 | n62219 ;
  assign n85174 = ~n61480 ;
  assign n61482 = n61268 & n85174 ;
  assign n61642 = n60666 | n61268 ;
  assign n85175 = ~n61642 ;
  assign n61643 = n61264 & n85175 ;
  assign n61644 = n61482 | n61643 ;
  assign n61645 = n85129 & n61644 ;
  assign n61646 = n60657 & n85125 ;
  assign n61647 = n61525 & n61646 ;
  assign n61648 = n61645 | n61647 ;
  assign n61649 = n70927 & n61648 ;
  assign n85176 = ~n61259 ;
  assign n61263 = n85176 & n61262 ;
  assign n61650 = n60675 | n61262 ;
  assign n85177 = ~n61650 ;
  assign n61651 = n61476 & n85177 ;
  assign n61652 = n61263 | n61651 ;
  assign n61653 = n85129 & n61652 ;
  assign n61654 = n60665 & n85125 ;
  assign n61655 = n61525 & n61654 ;
  assign n61656 = n61653 | n61655 ;
  assign n61657 = n70609 & n61656 ;
  assign n85178 = ~n61655 ;
  assign n62207 = x107 & n85178 ;
  assign n85179 = ~n61653 ;
  assign n62208 = n85179 & n62207 ;
  assign n62209 = n61657 | n62208 ;
  assign n85180 = ~n61475 ;
  assign n61477 = n61257 & n85180 ;
  assign n61658 = n60684 | n61257 ;
  assign n85181 = ~n61658 ;
  assign n61659 = n61253 & n85181 ;
  assign n61660 = n61477 | n61659 ;
  assign n61661 = n85129 & n61660 ;
  assign n61662 = n60674 & n85125 ;
  assign n61663 = n61525 & n61662 ;
  assign n61664 = n61661 | n61663 ;
  assign n61665 = n70276 & n61664 ;
  assign n85182 = ~n61248 ;
  assign n61252 = n85182 & n61251 ;
  assign n61666 = n60692 | n61251 ;
  assign n85183 = ~n61666 ;
  assign n61667 = n61471 & n85183 ;
  assign n61668 = n61252 | n61667 ;
  assign n61669 = n85129 & n61668 ;
  assign n61670 = n60683 & n85125 ;
  assign n61671 = n61525 & n61670 ;
  assign n61672 = n61669 | n61671 ;
  assign n61673 = n70176 & n61672 ;
  assign n85184 = ~n61671 ;
  assign n62197 = x105 & n85184 ;
  assign n85185 = ~n61669 ;
  assign n62198 = n85185 & n62197 ;
  assign n62199 = n61673 | n62198 ;
  assign n85186 = ~n61470 ;
  assign n61472 = n61246 & n85186 ;
  assign n61674 = n60701 | n61246 ;
  assign n85187 = ~n61674 ;
  assign n61675 = n61242 & n85187 ;
  assign n61676 = n61472 | n61675 ;
  assign n61677 = n85129 & n61676 ;
  assign n61678 = n60691 & n85125 ;
  assign n61679 = n61525 & n61678 ;
  assign n61680 = n61677 | n61679 ;
  assign n61681 = n69857 & n61680 ;
  assign n85188 = ~n61237 ;
  assign n61241 = n85188 & n61240 ;
  assign n61682 = n60710 | n61240 ;
  assign n85189 = ~n61682 ;
  assign n61683 = n61466 & n85189 ;
  assign n61684 = n61241 | n61683 ;
  assign n61685 = n85129 & n61684 ;
  assign n61686 = n60700 & n85125 ;
  assign n61687 = n61525 & n61686 ;
  assign n61688 = n61685 | n61687 ;
  assign n61689 = n69656 & n61688 ;
  assign n85190 = ~n61687 ;
  assign n62187 = x103 & n85190 ;
  assign n85191 = ~n61685 ;
  assign n62188 = n85191 & n62187 ;
  assign n62189 = n61689 | n62188 ;
  assign n85192 = ~n61465 ;
  assign n61467 = n61235 & n85192 ;
  assign n61690 = n60719 | n61235 ;
  assign n85193 = ~n61690 ;
  assign n61691 = n61231 & n85193 ;
  assign n61692 = n61467 | n61691 ;
  assign n61693 = n85129 & n61692 ;
  assign n61694 = n60709 & n85125 ;
  assign n61695 = n61525 & n61694 ;
  assign n61696 = n61693 | n61695 ;
  assign n61697 = n69528 & n61696 ;
  assign n85194 = ~n61226 ;
  assign n61230 = n85194 & n61229 ;
  assign n61698 = n60728 | n61229 ;
  assign n85195 = ~n61698 ;
  assign n61699 = n61461 & n85195 ;
  assign n61700 = n61230 | n61699 ;
  assign n61701 = n85129 & n61700 ;
  assign n61702 = n60718 & n85125 ;
  assign n61703 = n61525 & n61702 ;
  assign n61704 = n61701 | n61703 ;
  assign n61705 = n69261 & n61704 ;
  assign n85196 = ~n61703 ;
  assign n62177 = x101 & n85196 ;
  assign n85197 = ~n61701 ;
  assign n62178 = n85197 & n62177 ;
  assign n62179 = n61705 | n62178 ;
  assign n85198 = ~n61460 ;
  assign n61462 = n61224 & n85198 ;
  assign n61706 = n60737 | n61224 ;
  assign n85199 = ~n61706 ;
  assign n61707 = n61220 & n85199 ;
  assign n61708 = n61462 | n61707 ;
  assign n61709 = n85129 & n61708 ;
  assign n61710 = n60727 & n85125 ;
  assign n61711 = n61525 & n61710 ;
  assign n61712 = n61709 | n61711 ;
  assign n61713 = n69075 & n61712 ;
  assign n85200 = ~n61215 ;
  assign n61219 = n85200 & n61218 ;
  assign n61714 = n60746 | n61218 ;
  assign n85201 = ~n61714 ;
  assign n61715 = n61456 & n85201 ;
  assign n61716 = n61219 | n61715 ;
  assign n61717 = n85129 & n61716 ;
  assign n61718 = n60736 & n85125 ;
  assign n61719 = n61525 & n61718 ;
  assign n61720 = n61717 | n61719 ;
  assign n61721 = n68993 & n61720 ;
  assign n85202 = ~n61719 ;
  assign n62167 = x99 & n85202 ;
  assign n85203 = ~n61717 ;
  assign n62168 = n85203 & n62167 ;
  assign n62169 = n61721 | n62168 ;
  assign n85204 = ~n61455 ;
  assign n61457 = n61213 & n85204 ;
  assign n61722 = n60755 | n61213 ;
  assign n85205 = ~n61722 ;
  assign n61723 = n61209 & n85205 ;
  assign n61724 = n61457 | n61723 ;
  assign n61725 = n85129 & n61724 ;
  assign n61726 = n60745 & n85125 ;
  assign n61727 = n61525 & n61726 ;
  assign n61728 = n61725 | n61727 ;
  assign n61729 = n68716 & n61728 ;
  assign n85206 = ~n61204 ;
  assign n61208 = n85206 & n61207 ;
  assign n61730 = n60764 | n61207 ;
  assign n85207 = ~n61730 ;
  assign n61731 = n61451 & n85207 ;
  assign n61732 = n61208 | n61731 ;
  assign n61733 = n85129 & n61732 ;
  assign n61734 = n60754 & n85125 ;
  assign n61735 = n61525 & n61734 ;
  assign n61736 = n61733 | n61735 ;
  assign n61737 = n68545 & n61736 ;
  assign n85208 = ~n61735 ;
  assign n62157 = x97 & n85208 ;
  assign n85209 = ~n61733 ;
  assign n62158 = n85209 & n62157 ;
  assign n62159 = n61737 | n62158 ;
  assign n85210 = ~n61450 ;
  assign n61452 = n61202 & n85210 ;
  assign n61738 = n60773 | n61202 ;
  assign n85211 = ~n61738 ;
  assign n61739 = n61198 & n85211 ;
  assign n61740 = n61452 | n61739 ;
  assign n61741 = n85129 & n61740 ;
  assign n61742 = n60763 & n85125 ;
  assign n61743 = n61525 & n61742 ;
  assign n61744 = n61741 | n61743 ;
  assign n61745 = n68438 & n61744 ;
  assign n85212 = ~n61193 ;
  assign n61197 = n85212 & n61196 ;
  assign n61746 = n60782 | n61196 ;
  assign n85213 = ~n61746 ;
  assign n61747 = n61446 & n85213 ;
  assign n61748 = n61197 | n61747 ;
  assign n61749 = n85129 & n61748 ;
  assign n61750 = n60772 & n85125 ;
  assign n61751 = n61525 & n61750 ;
  assign n61752 = n61749 | n61751 ;
  assign n61753 = n68214 & n61752 ;
  assign n85214 = ~n61751 ;
  assign n62147 = x95 & n85214 ;
  assign n85215 = ~n61749 ;
  assign n62148 = n85215 & n62147 ;
  assign n62149 = n61753 | n62148 ;
  assign n85216 = ~n61445 ;
  assign n61447 = n61191 & n85216 ;
  assign n61754 = n60791 | n61191 ;
  assign n85217 = ~n61754 ;
  assign n61755 = n61187 & n85217 ;
  assign n61756 = n61447 | n61755 ;
  assign n61757 = n85129 & n61756 ;
  assign n61758 = n60781 & n85125 ;
  assign n61759 = n61525 & n61758 ;
  assign n61760 = n61757 | n61759 ;
  assign n61761 = n68058 & n61760 ;
  assign n85218 = ~n61182 ;
  assign n61186 = n85218 & n61185 ;
  assign n61762 = n60800 | n61185 ;
  assign n85219 = ~n61762 ;
  assign n61763 = n61441 & n85219 ;
  assign n61764 = n61186 | n61763 ;
  assign n61765 = n85129 & n61764 ;
  assign n61766 = n60790 & n85125 ;
  assign n61767 = n61525 & n61766 ;
  assign n61768 = n61765 | n61767 ;
  assign n61769 = n67986 & n61768 ;
  assign n85220 = ~n61767 ;
  assign n62137 = x93 & n85220 ;
  assign n85221 = ~n61765 ;
  assign n62138 = n85221 & n62137 ;
  assign n62139 = n61769 | n62138 ;
  assign n85222 = ~n61440 ;
  assign n61442 = n61180 & n85222 ;
  assign n61770 = n60809 | n61180 ;
  assign n85223 = ~n61770 ;
  assign n61771 = n61176 & n85223 ;
  assign n61772 = n61442 | n61771 ;
  assign n61773 = n85129 & n61772 ;
  assign n61774 = n60799 & n85125 ;
  assign n61775 = n61525 & n61774 ;
  assign n61776 = n61773 | n61775 ;
  assign n61777 = n67763 & n61776 ;
  assign n85224 = ~n61171 ;
  assign n61175 = n85224 & n61174 ;
  assign n61778 = n60818 | n61174 ;
  assign n85225 = ~n61778 ;
  assign n61779 = n61436 & n85225 ;
  assign n61780 = n61175 | n61779 ;
  assign n61781 = n85129 & n61780 ;
  assign n61782 = n60808 & n85125 ;
  assign n61783 = n61525 & n61782 ;
  assign n61784 = n61781 | n61783 ;
  assign n61785 = n67622 & n61784 ;
  assign n85226 = ~n61783 ;
  assign n62126 = x91 & n85226 ;
  assign n85227 = ~n61781 ;
  assign n62127 = n85227 & n62126 ;
  assign n62128 = n61785 | n62127 ;
  assign n85228 = ~n61435 ;
  assign n61437 = n61169 & n85228 ;
  assign n61786 = n60827 | n61169 ;
  assign n85229 = ~n61786 ;
  assign n61787 = n61165 & n85229 ;
  assign n61788 = n61437 | n61787 ;
  assign n61789 = n85129 & n61788 ;
  assign n61790 = n60817 & n85125 ;
  assign n61791 = n61525 & n61790 ;
  assign n61792 = n61789 | n61791 ;
  assign n61793 = n67531 & n61792 ;
  assign n85230 = ~n61160 ;
  assign n61164 = n85230 & n61163 ;
  assign n61794 = n60836 | n61163 ;
  assign n85231 = ~n61794 ;
  assign n61795 = n61431 & n85231 ;
  assign n61796 = n61164 | n61795 ;
  assign n61797 = n85129 & n61796 ;
  assign n61798 = n60826 & n85125 ;
  assign n61799 = n61525 & n61798 ;
  assign n61800 = n61797 | n61799 ;
  assign n61801 = n67348 & n61800 ;
  assign n85232 = ~n61799 ;
  assign n62116 = x89 & n85232 ;
  assign n85233 = ~n61797 ;
  assign n62117 = n85233 & n62116 ;
  assign n62118 = n61801 | n62117 ;
  assign n85234 = ~n61430 ;
  assign n61432 = n61158 & n85234 ;
  assign n61802 = n60845 | n61158 ;
  assign n85235 = ~n61802 ;
  assign n61803 = n61154 & n85235 ;
  assign n61804 = n61432 | n61803 ;
  assign n61805 = n85129 & n61804 ;
  assign n61806 = n60835 & n85125 ;
  assign n61807 = n61525 & n61806 ;
  assign n61808 = n61805 | n61807 ;
  assign n61809 = n67222 & n61808 ;
  assign n85236 = ~n61149 ;
  assign n61153 = n85236 & n61152 ;
  assign n61810 = n60854 | n61152 ;
  assign n85237 = ~n61810 ;
  assign n61811 = n61426 & n85237 ;
  assign n61812 = n61153 | n61811 ;
  assign n61813 = n85129 & n61812 ;
  assign n61814 = n60844 & n85125 ;
  assign n61815 = n61525 & n61814 ;
  assign n61816 = n61813 | n61815 ;
  assign n61817 = n67164 & n61816 ;
  assign n85238 = ~n61815 ;
  assign n62106 = x87 & n85238 ;
  assign n85239 = ~n61813 ;
  assign n62107 = n85239 & n62106 ;
  assign n62108 = n61817 | n62107 ;
  assign n85240 = ~n61425 ;
  assign n61427 = n61147 & n85240 ;
  assign n61818 = n60863 | n61147 ;
  assign n85241 = ~n61818 ;
  assign n61819 = n61143 & n85241 ;
  assign n61820 = n61427 | n61819 ;
  assign n61821 = n85129 & n61820 ;
  assign n61822 = n60853 & n85125 ;
  assign n61823 = n61525 & n61822 ;
  assign n61824 = n61821 | n61823 ;
  assign n61825 = n66979 & n61824 ;
  assign n85242 = ~n61138 ;
  assign n61142 = n85242 & n61141 ;
  assign n61826 = n60872 | n61141 ;
  assign n85243 = ~n61826 ;
  assign n61827 = n61421 & n85243 ;
  assign n61828 = n61142 | n61827 ;
  assign n61829 = n85129 & n61828 ;
  assign n61830 = n60862 & n85125 ;
  assign n61831 = n61525 & n61830 ;
  assign n61832 = n61829 | n61831 ;
  assign n61833 = n66868 & n61832 ;
  assign n85244 = ~n61831 ;
  assign n62096 = x85 & n85244 ;
  assign n85245 = ~n61829 ;
  assign n62097 = n85245 & n62096 ;
  assign n62098 = n61833 | n62097 ;
  assign n85246 = ~n61420 ;
  assign n61422 = n61136 & n85246 ;
  assign n61834 = n60881 | n61136 ;
  assign n85247 = ~n61834 ;
  assign n61835 = n61132 & n85247 ;
  assign n61836 = n61422 | n61835 ;
  assign n61837 = n85129 & n61836 ;
  assign n61838 = n60871 & n85125 ;
  assign n61839 = n61525 & n61838 ;
  assign n61840 = n61837 | n61839 ;
  assign n61841 = n66797 & n61840 ;
  assign n85248 = ~n61127 ;
  assign n61131 = n85248 & n61130 ;
  assign n61842 = n60890 | n61130 ;
  assign n85249 = ~n61842 ;
  assign n61843 = n61416 & n85249 ;
  assign n61844 = n61131 | n61843 ;
  assign n61845 = n85129 & n61844 ;
  assign n61846 = n60880 & n85125 ;
  assign n61847 = n61525 & n61846 ;
  assign n61848 = n61845 | n61847 ;
  assign n61849 = n66654 & n61848 ;
  assign n85250 = ~n61847 ;
  assign n62086 = x83 & n85250 ;
  assign n85251 = ~n61845 ;
  assign n62087 = n85251 & n62086 ;
  assign n62088 = n61849 | n62087 ;
  assign n85252 = ~n61415 ;
  assign n61417 = n61125 & n85252 ;
  assign n61850 = n60899 | n61125 ;
  assign n85253 = ~n61850 ;
  assign n61851 = n61121 & n85253 ;
  assign n61852 = n61417 | n61851 ;
  assign n61853 = n85129 & n61852 ;
  assign n61854 = n60889 & n85125 ;
  assign n61855 = n61525 & n61854 ;
  assign n61856 = n61853 | n61855 ;
  assign n61857 = n66560 & n61856 ;
  assign n85254 = ~n61116 ;
  assign n61120 = n85254 & n61119 ;
  assign n61858 = n60908 | n61119 ;
  assign n85255 = ~n61858 ;
  assign n61859 = n61411 & n85255 ;
  assign n61860 = n61120 | n61859 ;
  assign n61861 = n85129 & n61860 ;
  assign n61862 = n60898 & n85125 ;
  assign n61863 = n61525 & n61862 ;
  assign n61864 = n61861 | n61863 ;
  assign n61865 = n66505 & n61864 ;
  assign n85256 = ~n61863 ;
  assign n62076 = x81 & n85256 ;
  assign n85257 = ~n61861 ;
  assign n62077 = n85257 & n62076 ;
  assign n62078 = n61865 | n62077 ;
  assign n85258 = ~n61410 ;
  assign n61412 = n61114 & n85258 ;
  assign n61866 = n60916 | n61114 ;
  assign n85259 = ~n61866 ;
  assign n61867 = n61110 & n85259 ;
  assign n61868 = n61412 | n61867 ;
  assign n61869 = n85129 & n61868 ;
  assign n61870 = n60907 & n85125 ;
  assign n61871 = n61525 & n61870 ;
  assign n61872 = n61869 | n61871 ;
  assign n61873 = n66379 & n61872 ;
  assign n85260 = ~n61105 ;
  assign n61109 = n85260 & n61108 ;
  assign n61874 = n60925 | n61108 ;
  assign n85261 = ~n61874 ;
  assign n61875 = n61406 & n85261 ;
  assign n61876 = n61109 | n61875 ;
  assign n61877 = n85129 & n61876 ;
  assign n61878 = n60915 & n85125 ;
  assign n61879 = n61525 & n61878 ;
  assign n61880 = n61877 | n61879 ;
  assign n61881 = n66299 & n61880 ;
  assign n85262 = ~n61879 ;
  assign n62066 = x79 & n85262 ;
  assign n85263 = ~n61877 ;
  assign n62067 = n85263 & n62066 ;
  assign n62068 = n61881 | n62067 ;
  assign n85264 = ~n61405 ;
  assign n61407 = n61103 & n85264 ;
  assign n61882 = n60933 | n61103 ;
  assign n85265 = ~n61882 ;
  assign n61883 = n61099 & n85265 ;
  assign n61884 = n61407 | n61883 ;
  assign n61885 = n85129 & n61884 ;
  assign n61886 = n60924 & n85125 ;
  assign n61887 = n61525 & n61886 ;
  assign n61888 = n61885 | n61887 ;
  assign n61889 = n66244 & n61888 ;
  assign n85266 = ~n61094 ;
  assign n61098 = n85266 & n61097 ;
  assign n61890 = n60942 | n61097 ;
  assign n85267 = ~n61890 ;
  assign n61891 = n61401 & n85267 ;
  assign n61892 = n61098 | n61891 ;
  assign n61893 = n85129 & n61892 ;
  assign n61894 = n60932 & n85125 ;
  assign n61895 = n61525 & n61894 ;
  assign n61896 = n61893 | n61895 ;
  assign n61897 = n66145 & n61896 ;
  assign n85268 = ~n61895 ;
  assign n62056 = x77 & n85268 ;
  assign n85269 = ~n61893 ;
  assign n62057 = n85269 & n62056 ;
  assign n62058 = n61897 | n62057 ;
  assign n85270 = ~n61400 ;
  assign n61402 = n61092 & n85270 ;
  assign n61898 = n60951 | n61092 ;
  assign n85271 = ~n61898 ;
  assign n61899 = n61088 & n85271 ;
  assign n61900 = n61402 | n61899 ;
  assign n61901 = n85129 & n61900 ;
  assign n61902 = n60941 & n85125 ;
  assign n61903 = n61525 & n61902 ;
  assign n61904 = n61901 | n61903 ;
  assign n61905 = n66081 & n61904 ;
  assign n85272 = ~n61083 ;
  assign n61087 = n85272 & n61086 ;
  assign n61906 = n60960 | n61086 ;
  assign n85273 = ~n61906 ;
  assign n61907 = n61396 & n85273 ;
  assign n61908 = n61087 | n61907 ;
  assign n61909 = n85129 & n61908 ;
  assign n61910 = n60950 & n85125 ;
  assign n61911 = n61525 & n61910 ;
  assign n61912 = n61909 | n61911 ;
  assign n61913 = n66043 & n61912 ;
  assign n85274 = ~n61911 ;
  assign n62045 = x75 & n85274 ;
  assign n85275 = ~n61909 ;
  assign n62046 = n85275 & n62045 ;
  assign n62047 = n61913 | n62046 ;
  assign n85276 = ~n61395 ;
  assign n61397 = n61081 & n85276 ;
  assign n61914 = n60969 | n61081 ;
  assign n85277 = ~n61914 ;
  assign n61915 = n61077 & n85277 ;
  assign n61916 = n61397 | n61915 ;
  assign n61917 = n85129 & n61916 ;
  assign n61918 = n60959 & n85125 ;
  assign n61919 = n61525 & n61918 ;
  assign n61920 = n61917 | n61919 ;
  assign n61921 = n65960 & n61920 ;
  assign n85278 = ~n61072 ;
  assign n61076 = n85278 & n61075 ;
  assign n61922 = n60978 | n61075 ;
  assign n85279 = ~n61922 ;
  assign n61923 = n61391 & n85279 ;
  assign n61924 = n61076 | n61923 ;
  assign n61925 = n85129 & n61924 ;
  assign n61926 = n60968 & n85125 ;
  assign n61927 = n61525 & n61926 ;
  assign n61928 = n61925 | n61927 ;
  assign n61929 = n65909 & n61928 ;
  assign n85280 = ~n61927 ;
  assign n62035 = x73 & n85280 ;
  assign n85281 = ~n61925 ;
  assign n62036 = n85281 & n62035 ;
  assign n62037 = n61929 | n62036 ;
  assign n85282 = ~n61390 ;
  assign n61392 = n61070 & n85282 ;
  assign n61930 = n60987 | n61070 ;
  assign n85283 = ~n61930 ;
  assign n61931 = n61066 & n85283 ;
  assign n61932 = n61392 | n61931 ;
  assign n61933 = n85129 & n61932 ;
  assign n61934 = n60977 & n85125 ;
  assign n61935 = n61525 & n61934 ;
  assign n61936 = n61933 | n61935 ;
  assign n61937 = n65877 & n61936 ;
  assign n85284 = ~n61061 ;
  assign n61065 = n85284 & n61064 ;
  assign n61938 = n60996 | n61064 ;
  assign n85285 = ~n61938 ;
  assign n61939 = n61386 & n85285 ;
  assign n61940 = n61065 | n61939 ;
  assign n61941 = n85129 & n61940 ;
  assign n61942 = n60986 & n85125 ;
  assign n61943 = n61525 & n61942 ;
  assign n61944 = n61941 | n61943 ;
  assign n61945 = n65820 & n61944 ;
  assign n85286 = ~n61943 ;
  assign n62025 = x71 & n85286 ;
  assign n85287 = ~n61941 ;
  assign n62026 = n85287 & n62025 ;
  assign n62027 = n61945 | n62026 ;
  assign n85288 = ~n61385 ;
  assign n61387 = n61059 & n85288 ;
  assign n61946 = n61005 | n61059 ;
  assign n85289 = ~n61946 ;
  assign n61947 = n61055 & n85289 ;
  assign n61948 = n61387 | n61947 ;
  assign n61949 = n85129 & n61948 ;
  assign n61950 = n60995 & n85125 ;
  assign n61951 = n61525 & n61950 ;
  assign n61952 = n61949 | n61951 ;
  assign n61953 = n65791 & n61952 ;
  assign n85290 = ~n61051 ;
  assign n61383 = n85290 & n61054 ;
  assign n61954 = n61014 | n61054 ;
  assign n85291 = ~n61954 ;
  assign n61955 = n61381 & n85291 ;
  assign n61956 = n61383 | n61955 ;
  assign n61957 = n85129 & n61956 ;
  assign n61958 = n61004 & n85125 ;
  assign n61959 = n61525 & n61958 ;
  assign n61960 = n61957 | n61959 ;
  assign n61961 = n65772 & n61960 ;
  assign n85292 = ~n61959 ;
  assign n62015 = x69 & n85292 ;
  assign n85293 = ~n61957 ;
  assign n62016 = n85293 & n62015 ;
  assign n62017 = n61961 | n62016 ;
  assign n85294 = ~n61379 ;
  assign n61380 = n61049 & n85294 ;
  assign n61962 = n61022 | n61049 ;
  assign n85295 = ~n61962 ;
  assign n61963 = n61378 & n85295 ;
  assign n61964 = n61380 | n61963 ;
  assign n61965 = n85129 & n61964 ;
  assign n61966 = n61013 & n85125 ;
  assign n61967 = n61525 & n61966 ;
  assign n61968 = n61965 | n61967 ;
  assign n61969 = n65746 & n61968 ;
  assign n85296 = ~n61377 ;
  assign n61971 = n61044 & n85296 ;
  assign n61970 = n61039 | n61044 ;
  assign n85297 = ~n61970 ;
  assign n61972 = n61040 & n85297 ;
  assign n61973 = n61971 | n61972 ;
  assign n61974 = n85129 & n61973 ;
  assign n61975 = n61021 & n85125 ;
  assign n61976 = n61525 & n61975 ;
  assign n61977 = n61974 | n61976 ;
  assign n61978 = n65721 & n61977 ;
  assign n85298 = ~n61976 ;
  assign n62005 = x67 & n85298 ;
  assign n85299 = ~n61974 ;
  assign n62006 = n85299 & n62005 ;
  assign n62007 = n61978 | n62006 ;
  assign n61979 = n28839 & n61037 ;
  assign n61980 = n85127 & n61979 ;
  assign n85300 = ~n61980 ;
  assign n61981 = n61040 & n85300 ;
  assign n61982 = n85129 & n61981 ;
  assign n61983 = n61025 & n85125 ;
  assign n61984 = n61525 & n61983 ;
  assign n61985 = n61982 | n61984 ;
  assign n61986 = n65686 & n61985 ;
  assign n61372 = n28839 & n85129 ;
  assign n61987 = n85125 & n61525 ;
  assign n85301 = ~n61987 ;
  assign n61988 = x64 & n85301 ;
  assign n85302 = ~n61988 ;
  assign n61989 = x4 & n85302 ;
  assign n61990 = n61372 | n61989 ;
  assign n61991 = x65 & n61990 ;
  assign n61373 = x64 & n85129 ;
  assign n85303 = ~n61373 ;
  assign n61992 = x4 & n85303 ;
  assign n61993 = n28839 & n85301 ;
  assign n61994 = x65 | n61993 ;
  assign n61995 = n61992 | n61994 ;
  assign n85304 = ~n61991 ;
  assign n61996 = n85304 & n61995 ;
  assign n61997 = n29800 | n61996 ;
  assign n61998 = n61372 | n61992 ;
  assign n61999 = n65670 & n61998 ;
  assign n85305 = ~n61999 ;
  assign n62000 = n61997 & n85305 ;
  assign n85306 = ~n61984 ;
  assign n62001 = x66 & n85306 ;
  assign n85307 = ~n61982 ;
  assign n62002 = n85307 & n62001 ;
  assign n62003 = n61986 | n62002 ;
  assign n62004 = n62000 | n62003 ;
  assign n85308 = ~n61986 ;
  assign n62008 = n85308 & n62004 ;
  assign n62009 = n62007 | n62008 ;
  assign n85309 = ~n61978 ;
  assign n62010 = n85309 & n62009 ;
  assign n85310 = ~n61967 ;
  assign n62011 = x68 & n85310 ;
  assign n85311 = ~n61965 ;
  assign n62012 = n85311 & n62011 ;
  assign n62013 = n61969 | n62012 ;
  assign n62014 = n62010 | n62013 ;
  assign n85312 = ~n61969 ;
  assign n62018 = n85312 & n62014 ;
  assign n62019 = n62017 | n62018 ;
  assign n85313 = ~n61961 ;
  assign n62020 = n85313 & n62019 ;
  assign n85314 = ~n61951 ;
  assign n62021 = x70 & n85314 ;
  assign n85315 = ~n61949 ;
  assign n62022 = n85315 & n62021 ;
  assign n62023 = n61953 | n62022 ;
  assign n62024 = n62020 | n62023 ;
  assign n85316 = ~n61953 ;
  assign n62028 = n85316 & n62024 ;
  assign n62029 = n62027 | n62028 ;
  assign n85317 = ~n61945 ;
  assign n62030 = n85317 & n62029 ;
  assign n85318 = ~n61935 ;
  assign n62031 = x72 & n85318 ;
  assign n85319 = ~n61933 ;
  assign n62032 = n85319 & n62031 ;
  assign n62033 = n61937 | n62032 ;
  assign n62034 = n62030 | n62033 ;
  assign n85320 = ~n61937 ;
  assign n62038 = n85320 & n62034 ;
  assign n62039 = n62037 | n62038 ;
  assign n85321 = ~n61929 ;
  assign n62040 = n85321 & n62039 ;
  assign n85322 = ~n61919 ;
  assign n62041 = x74 & n85322 ;
  assign n85323 = ~n61917 ;
  assign n62042 = n85323 & n62041 ;
  assign n62043 = n61921 | n62042 ;
  assign n62044 = n62040 | n62043 ;
  assign n85324 = ~n61921 ;
  assign n62048 = n85324 & n62044 ;
  assign n62049 = n62047 | n62048 ;
  assign n85325 = ~n61913 ;
  assign n62050 = n85325 & n62049 ;
  assign n85326 = ~n61903 ;
  assign n62051 = x76 & n85326 ;
  assign n85327 = ~n61901 ;
  assign n62052 = n85327 & n62051 ;
  assign n62053 = n61905 | n62052 ;
  assign n62055 = n62050 | n62053 ;
  assign n85328 = ~n61905 ;
  assign n62059 = n85328 & n62055 ;
  assign n62060 = n62058 | n62059 ;
  assign n85329 = ~n61897 ;
  assign n62061 = n85329 & n62060 ;
  assign n85330 = ~n61887 ;
  assign n62062 = x78 & n85330 ;
  assign n85331 = ~n61885 ;
  assign n62063 = n85331 & n62062 ;
  assign n62064 = n61889 | n62063 ;
  assign n62065 = n62061 | n62064 ;
  assign n85332 = ~n61889 ;
  assign n62069 = n85332 & n62065 ;
  assign n62070 = n62068 | n62069 ;
  assign n85333 = ~n61881 ;
  assign n62071 = n85333 & n62070 ;
  assign n85334 = ~n61871 ;
  assign n62072 = x80 & n85334 ;
  assign n85335 = ~n61869 ;
  assign n62073 = n85335 & n62072 ;
  assign n62074 = n61873 | n62073 ;
  assign n62075 = n62071 | n62074 ;
  assign n85336 = ~n61873 ;
  assign n62079 = n85336 & n62075 ;
  assign n62080 = n62078 | n62079 ;
  assign n85337 = ~n61865 ;
  assign n62081 = n85337 & n62080 ;
  assign n85338 = ~n61855 ;
  assign n62082 = x82 & n85338 ;
  assign n85339 = ~n61853 ;
  assign n62083 = n85339 & n62082 ;
  assign n62084 = n61857 | n62083 ;
  assign n62085 = n62081 | n62084 ;
  assign n85340 = ~n61857 ;
  assign n62089 = n85340 & n62085 ;
  assign n62090 = n62088 | n62089 ;
  assign n85341 = ~n61849 ;
  assign n62091 = n85341 & n62090 ;
  assign n85342 = ~n61839 ;
  assign n62092 = x84 & n85342 ;
  assign n85343 = ~n61837 ;
  assign n62093 = n85343 & n62092 ;
  assign n62094 = n61841 | n62093 ;
  assign n62095 = n62091 | n62094 ;
  assign n85344 = ~n61841 ;
  assign n62099 = n85344 & n62095 ;
  assign n62100 = n62098 | n62099 ;
  assign n85345 = ~n61833 ;
  assign n62101 = n85345 & n62100 ;
  assign n85346 = ~n61823 ;
  assign n62102 = x86 & n85346 ;
  assign n85347 = ~n61821 ;
  assign n62103 = n85347 & n62102 ;
  assign n62104 = n61825 | n62103 ;
  assign n62105 = n62101 | n62104 ;
  assign n85348 = ~n61825 ;
  assign n62109 = n85348 & n62105 ;
  assign n62110 = n62108 | n62109 ;
  assign n85349 = ~n61817 ;
  assign n62111 = n85349 & n62110 ;
  assign n85350 = ~n61807 ;
  assign n62112 = x88 & n85350 ;
  assign n85351 = ~n61805 ;
  assign n62113 = n85351 & n62112 ;
  assign n62114 = n61809 | n62113 ;
  assign n62115 = n62111 | n62114 ;
  assign n85352 = ~n61809 ;
  assign n62119 = n85352 & n62115 ;
  assign n62120 = n62118 | n62119 ;
  assign n85353 = ~n61801 ;
  assign n62121 = n85353 & n62120 ;
  assign n85354 = ~n61791 ;
  assign n62122 = x90 & n85354 ;
  assign n85355 = ~n61789 ;
  assign n62123 = n85355 & n62122 ;
  assign n62124 = n61793 | n62123 ;
  assign n62125 = n62121 | n62124 ;
  assign n85356 = ~n61793 ;
  assign n62130 = n85356 & n62125 ;
  assign n62131 = n62128 | n62130 ;
  assign n85357 = ~n61785 ;
  assign n62132 = n85357 & n62131 ;
  assign n85358 = ~n61775 ;
  assign n62133 = x92 & n85358 ;
  assign n85359 = ~n61773 ;
  assign n62134 = n85359 & n62133 ;
  assign n62135 = n61777 | n62134 ;
  assign n62136 = n62132 | n62135 ;
  assign n85360 = ~n61777 ;
  assign n62140 = n85360 & n62136 ;
  assign n62141 = n62139 | n62140 ;
  assign n85361 = ~n61769 ;
  assign n62142 = n85361 & n62141 ;
  assign n85362 = ~n61759 ;
  assign n62143 = x94 & n85362 ;
  assign n85363 = ~n61757 ;
  assign n62144 = n85363 & n62143 ;
  assign n62145 = n61761 | n62144 ;
  assign n62146 = n62142 | n62145 ;
  assign n85364 = ~n61761 ;
  assign n62150 = n85364 & n62146 ;
  assign n62151 = n62149 | n62150 ;
  assign n85365 = ~n61753 ;
  assign n62152 = n85365 & n62151 ;
  assign n85366 = ~n61743 ;
  assign n62153 = x96 & n85366 ;
  assign n85367 = ~n61741 ;
  assign n62154 = n85367 & n62153 ;
  assign n62155 = n61745 | n62154 ;
  assign n62156 = n62152 | n62155 ;
  assign n85368 = ~n61745 ;
  assign n62160 = n85368 & n62156 ;
  assign n62161 = n62159 | n62160 ;
  assign n85369 = ~n61737 ;
  assign n62162 = n85369 & n62161 ;
  assign n85370 = ~n61727 ;
  assign n62163 = x98 & n85370 ;
  assign n85371 = ~n61725 ;
  assign n62164 = n85371 & n62163 ;
  assign n62165 = n61729 | n62164 ;
  assign n62166 = n62162 | n62165 ;
  assign n85372 = ~n61729 ;
  assign n62170 = n85372 & n62166 ;
  assign n62171 = n62169 | n62170 ;
  assign n85373 = ~n61721 ;
  assign n62172 = n85373 & n62171 ;
  assign n85374 = ~n61711 ;
  assign n62173 = x100 & n85374 ;
  assign n85375 = ~n61709 ;
  assign n62174 = n85375 & n62173 ;
  assign n62175 = n61713 | n62174 ;
  assign n62176 = n62172 | n62175 ;
  assign n85376 = ~n61713 ;
  assign n62180 = n85376 & n62176 ;
  assign n62181 = n62179 | n62180 ;
  assign n85377 = ~n61705 ;
  assign n62182 = n85377 & n62181 ;
  assign n85378 = ~n61695 ;
  assign n62183 = x102 & n85378 ;
  assign n85379 = ~n61693 ;
  assign n62184 = n85379 & n62183 ;
  assign n62185 = n61697 | n62184 ;
  assign n62186 = n62182 | n62185 ;
  assign n85380 = ~n61697 ;
  assign n62190 = n85380 & n62186 ;
  assign n62191 = n62189 | n62190 ;
  assign n85381 = ~n61689 ;
  assign n62192 = n85381 & n62191 ;
  assign n85382 = ~n61679 ;
  assign n62193 = x104 & n85382 ;
  assign n85383 = ~n61677 ;
  assign n62194 = n85383 & n62193 ;
  assign n62195 = n61681 | n62194 ;
  assign n62196 = n62192 | n62195 ;
  assign n85384 = ~n61681 ;
  assign n62200 = n85384 & n62196 ;
  assign n62201 = n62199 | n62200 ;
  assign n85385 = ~n61673 ;
  assign n62202 = n85385 & n62201 ;
  assign n85386 = ~n61663 ;
  assign n62203 = x106 & n85386 ;
  assign n85387 = ~n61661 ;
  assign n62204 = n85387 & n62203 ;
  assign n62205 = n61665 | n62204 ;
  assign n62206 = n62202 | n62205 ;
  assign n85388 = ~n61665 ;
  assign n62211 = n85388 & n62206 ;
  assign n62212 = n62209 | n62211 ;
  assign n85389 = ~n61657 ;
  assign n62213 = n85389 & n62212 ;
  assign n85390 = ~n61647 ;
  assign n62214 = x108 & n85390 ;
  assign n85391 = ~n61645 ;
  assign n62215 = n85391 & n62214 ;
  assign n62216 = n61649 | n62215 ;
  assign n62217 = n62213 | n62216 ;
  assign n85392 = ~n61649 ;
  assign n62221 = n85392 & n62217 ;
  assign n62222 = n62220 | n62221 ;
  assign n85393 = ~n61641 ;
  assign n62223 = n85393 & n62222 ;
  assign n85394 = ~n61631 ;
  assign n62224 = x110 & n85394 ;
  assign n85395 = ~n61629 ;
  assign n62225 = n85395 & n62224 ;
  assign n62226 = n61633 | n62225 ;
  assign n62227 = n62223 | n62226 ;
  assign n85396 = ~n61633 ;
  assign n62231 = n85396 & n62227 ;
  assign n62232 = n62230 | n62231 ;
  assign n85397 = ~n61625 ;
  assign n62233 = n85397 & n62232 ;
  assign n85398 = ~n61615 ;
  assign n62234 = x112 & n85398 ;
  assign n85399 = ~n61613 ;
  assign n62235 = n85399 & n62234 ;
  assign n62236 = n61617 | n62235 ;
  assign n62237 = n62233 | n62236 ;
  assign n85400 = ~n61617 ;
  assign n62241 = n85400 & n62237 ;
  assign n62242 = n62240 | n62241 ;
  assign n85401 = ~n61609 ;
  assign n62243 = n85401 & n62242 ;
  assign n85402 = ~n61599 ;
  assign n62244 = x114 & n85402 ;
  assign n85403 = ~n61597 ;
  assign n62245 = n85403 & n62244 ;
  assign n62246 = n61601 | n62245 ;
  assign n62247 = n62243 | n62246 ;
  assign n85404 = ~n61601 ;
  assign n62251 = n85404 & n62247 ;
  assign n62252 = n62250 | n62251 ;
  assign n85405 = ~n61593 ;
  assign n62253 = n85405 & n62252 ;
  assign n85406 = ~n61583 ;
  assign n62254 = x116 & n85406 ;
  assign n85407 = ~n61581 ;
  assign n62255 = n85407 & n62254 ;
  assign n62256 = n61585 | n62255 ;
  assign n62257 = n62253 | n62256 ;
  assign n85408 = ~n61585 ;
  assign n62261 = n85408 & n62257 ;
  assign n62262 = n62260 | n62261 ;
  assign n85409 = ~n61577 ;
  assign n62263 = n85409 & n62262 ;
  assign n85410 = ~n61567 ;
  assign n62264 = x118 & n85410 ;
  assign n85411 = ~n61565 ;
  assign n62265 = n85411 & n62264 ;
  assign n62266 = n61569 | n62265 ;
  assign n62267 = n62263 | n62266 ;
  assign n85412 = ~n61569 ;
  assign n62272 = n85412 & n62267 ;
  assign n62273 = n62270 | n62272 ;
  assign n85413 = ~n61561 ;
  assign n62274 = n85413 & n62273 ;
  assign n85414 = ~n61551 ;
  assign n62275 = x120 & n85414 ;
  assign n85415 = ~n61549 ;
  assign n62276 = n85415 & n62275 ;
  assign n62277 = n61553 | n62276 ;
  assign n62278 = n62274 | n62277 ;
  assign n85416 = ~n61553 ;
  assign n62283 = n85416 & n62278 ;
  assign n62284 = n62281 | n62283 ;
  assign n85417 = ~n61545 ;
  assign n62285 = n85417 & n62284 ;
  assign n85418 = ~n61535 ;
  assign n62286 = x122 & n85418 ;
  assign n85419 = ~n61533 ;
  assign n62287 = n85419 & n62286 ;
  assign n62288 = n61537 | n62287 ;
  assign n62289 = n62285 | n62288 ;
  assign n85420 = ~n61537 ;
  assign n62293 = n85420 & n62289 ;
  assign n62294 = n62292 | n62293 ;
  assign n85421 = ~n61529 ;
  assign n62295 = n85421 & n62294 ;
  assign n62296 = n60413 | n61366 ;
  assign n62297 = n61364 | n62296 ;
  assign n85422 = ~n62297 ;
  assign n62298 = n61352 & n85422 ;
  assign n62299 = n61364 | n61366 ;
  assign n85423 = ~n61524 ;
  assign n62300 = n85423 & n62299 ;
  assign n62301 = n62298 | n62300 ;
  assign n62302 = n85129 & n62301 ;
  assign n62303 = n28217 & n61363 ;
  assign n62304 = n61525 & n62303 ;
  assign n62305 = n62302 | n62304 ;
  assign n62306 = n75210 & n62305 ;
  assign n85424 = ~n62304 ;
  assign n62307 = x124 & n85424 ;
  assign n85425 = ~n62302 ;
  assign n62308 = n85425 & n62307 ;
  assign n62309 = n274 | n62308 ;
  assign n62310 = n62306 | n62309 ;
  assign n62311 = n62295 | n62310 ;
  assign n62312 = n73619 & n62305 ;
  assign n85426 = ~n62312 ;
  assign n62313 = n62311 & n85426 ;
  assign n63298 = n61529 | n62308 ;
  assign n63299 = n62306 | n63298 ;
  assign n85427 = ~n63299 ;
  assign n63300 = n62294 & n85427 ;
  assign n62314 = x65 & n61998 ;
  assign n85428 = ~n62314 ;
  assign n62315 = n61995 & n85428 ;
  assign n62316 = n29800 | n62315 ;
  assign n62318 = n85305 & n62316 ;
  assign n62319 = n62003 | n62318 ;
  assign n62320 = n85308 & n62319 ;
  assign n62321 = n62007 | n62320 ;
  assign n62322 = n85309 & n62321 ;
  assign n62323 = n62013 | n62322 ;
  assign n62324 = n85312 & n62323 ;
  assign n62325 = n62017 | n62324 ;
  assign n62326 = n85313 & n62325 ;
  assign n62327 = n62023 | n62326 ;
  assign n62328 = n85316 & n62327 ;
  assign n62329 = n62027 | n62328 ;
  assign n62330 = n85317 & n62329 ;
  assign n62331 = n62033 | n62330 ;
  assign n62332 = n85320 & n62331 ;
  assign n62333 = n62037 | n62332 ;
  assign n62334 = n85321 & n62333 ;
  assign n62335 = n62043 | n62334 ;
  assign n62336 = n85324 & n62335 ;
  assign n62337 = n62047 | n62336 ;
  assign n62338 = n85325 & n62337 ;
  assign n62339 = n62053 | n62338 ;
  assign n62340 = n85328 & n62339 ;
  assign n62341 = n62058 | n62340 ;
  assign n62342 = n85329 & n62341 ;
  assign n62343 = n62064 | n62342 ;
  assign n62344 = n85332 & n62343 ;
  assign n62345 = n62068 | n62344 ;
  assign n62346 = n85333 & n62345 ;
  assign n62347 = n62074 | n62346 ;
  assign n62348 = n85336 & n62347 ;
  assign n62349 = n62078 | n62348 ;
  assign n62350 = n85337 & n62349 ;
  assign n62351 = n62084 | n62350 ;
  assign n62352 = n85340 & n62351 ;
  assign n62353 = n62088 | n62352 ;
  assign n62354 = n85341 & n62353 ;
  assign n62355 = n62094 | n62354 ;
  assign n62356 = n85344 & n62355 ;
  assign n62357 = n62098 | n62356 ;
  assign n62358 = n85345 & n62357 ;
  assign n62359 = n62104 | n62358 ;
  assign n62360 = n85348 & n62359 ;
  assign n62361 = n62108 | n62360 ;
  assign n62362 = n85349 & n62361 ;
  assign n62363 = n62114 | n62362 ;
  assign n62364 = n85352 & n62363 ;
  assign n62365 = n62118 | n62364 ;
  assign n62366 = n85353 & n62365 ;
  assign n62367 = n62124 | n62366 ;
  assign n62368 = n85356 & n62367 ;
  assign n62369 = n62128 | n62368 ;
  assign n62370 = n85357 & n62369 ;
  assign n62371 = n62135 | n62370 ;
  assign n62372 = n85360 & n62371 ;
  assign n62373 = n62139 | n62372 ;
  assign n62374 = n85361 & n62373 ;
  assign n62375 = n62145 | n62374 ;
  assign n62376 = n85364 & n62375 ;
  assign n62377 = n62149 | n62376 ;
  assign n62378 = n85365 & n62377 ;
  assign n62379 = n62155 | n62378 ;
  assign n62380 = n85368 & n62379 ;
  assign n62381 = n62159 | n62380 ;
  assign n62382 = n85369 & n62381 ;
  assign n62383 = n62165 | n62382 ;
  assign n62384 = n85372 & n62383 ;
  assign n62385 = n62169 | n62384 ;
  assign n62386 = n85373 & n62385 ;
  assign n62387 = n62175 | n62386 ;
  assign n62388 = n85376 & n62387 ;
  assign n62389 = n62179 | n62388 ;
  assign n62390 = n85377 & n62389 ;
  assign n62391 = n62185 | n62390 ;
  assign n62392 = n85380 & n62391 ;
  assign n62393 = n62189 | n62392 ;
  assign n62394 = n85381 & n62393 ;
  assign n62395 = n62195 | n62394 ;
  assign n62396 = n85384 & n62395 ;
  assign n62397 = n62199 | n62396 ;
  assign n62398 = n85385 & n62397 ;
  assign n62399 = n62205 | n62398 ;
  assign n62400 = n85388 & n62399 ;
  assign n62401 = n62209 | n62400 ;
  assign n62402 = n85389 & n62401 ;
  assign n62403 = n62216 | n62402 ;
  assign n62404 = n85392 & n62403 ;
  assign n62405 = n62220 | n62404 ;
  assign n62406 = n85393 & n62405 ;
  assign n62407 = n62226 | n62406 ;
  assign n62408 = n85396 & n62407 ;
  assign n62409 = n62230 | n62408 ;
  assign n62410 = n85397 & n62409 ;
  assign n62411 = n62236 | n62410 ;
  assign n62412 = n85400 & n62411 ;
  assign n62413 = n62240 | n62412 ;
  assign n62414 = n85401 & n62413 ;
  assign n62415 = n62246 | n62414 ;
  assign n62416 = n85404 & n62415 ;
  assign n62417 = n62250 | n62416 ;
  assign n62418 = n85405 & n62417 ;
  assign n62419 = n62256 | n62418 ;
  assign n62420 = n85408 & n62419 ;
  assign n62421 = n62260 | n62420 ;
  assign n62422 = n85409 & n62421 ;
  assign n62423 = n62266 | n62422 ;
  assign n62424 = n85412 & n62423 ;
  assign n62425 = n62270 | n62424 ;
  assign n62426 = n85413 & n62425 ;
  assign n62427 = n62277 | n62426 ;
  assign n62428 = n85416 & n62427 ;
  assign n62429 = n62281 | n62428 ;
  assign n62430 = n85417 & n62429 ;
  assign n62431 = n62288 | n62430 ;
  assign n62432 = n85420 & n62431 ;
  assign n62961 = n62292 | n62432 ;
  assign n62962 = n85421 & n62961 ;
  assign n63301 = n62306 | n62308 ;
  assign n85429 = ~n62962 ;
  assign n63302 = n85429 & n63301 ;
  assign n63303 = n63300 | n63302 ;
  assign n85430 = ~n62313 ;
  assign n63304 = n85430 & n63303 ;
  assign n63305 = n65369 & n62305 ;
  assign n63306 = n62311 & n63305 ;
  assign n63307 = n63304 | n63306 ;
  assign n63313 = n73624 & n63307 ;
  assign n85431 = ~n62293 ;
  assign n62433 = n62292 & n85431 ;
  assign n62434 = n61537 | n62292 ;
  assign n85432 = ~n62434 ;
  assign n62435 = n62431 & n85432 ;
  assign n62436 = n62433 | n62435 ;
  assign n62437 = n85430 & n62436 ;
  assign n62438 = n61528 & n85426 ;
  assign n62439 = n62311 & n62438 ;
  assign n62440 = n62437 | n62439 ;
  assign n62441 = n75210 & n62440 ;
  assign n85433 = ~n62430 ;
  assign n62442 = n62288 & n85433 ;
  assign n62443 = n61545 | n62288 ;
  assign n85434 = ~n62443 ;
  assign n62444 = n62284 & n85434 ;
  assign n62445 = n62442 | n62444 ;
  assign n62446 = n85430 & n62445 ;
  assign n62447 = n61536 & n85426 ;
  assign n62448 = n62311 & n62447 ;
  assign n62449 = n62446 | n62448 ;
  assign n62450 = n74905 & n62449 ;
  assign n85435 = ~n62283 ;
  assign n62452 = n62281 & n85435 ;
  assign n62282 = n61553 | n62281 ;
  assign n85436 = ~n62282 ;
  assign n62453 = n62278 & n85436 ;
  assign n62454 = n62452 | n62453 ;
  assign n62455 = n85430 & n62454 ;
  assign n62456 = n61544 & n85426 ;
  assign n62457 = n62311 & n62456 ;
  assign n62458 = n62455 | n62457 ;
  assign n62459 = n74431 & n62458 ;
  assign n85437 = ~n62426 ;
  assign n62460 = n62277 & n85437 ;
  assign n62461 = n61561 | n62277 ;
  assign n85438 = ~n62461 ;
  assign n62462 = n62273 & n85438 ;
  assign n62463 = n62460 | n62462 ;
  assign n62464 = n85430 & n62463 ;
  assign n62465 = n61552 & n85426 ;
  assign n62466 = n62311 & n62465 ;
  assign n62467 = n62464 | n62466 ;
  assign n62468 = n74029 & n62467 ;
  assign n85439 = ~n62272 ;
  assign n62469 = n62270 & n85439 ;
  assign n62271 = n61569 | n62270 ;
  assign n85440 = ~n62271 ;
  assign n62470 = n62267 & n85440 ;
  assign n62471 = n62469 | n62470 ;
  assign n62472 = n85430 & n62471 ;
  assign n62473 = n61560 & n85426 ;
  assign n62474 = n62311 & n62473 ;
  assign n62475 = n62472 | n62474 ;
  assign n62476 = n74021 & n62475 ;
  assign n85441 = ~n62422 ;
  assign n62477 = n62266 & n85441 ;
  assign n62478 = n61577 | n62266 ;
  assign n85442 = ~n62478 ;
  assign n62479 = n62262 & n85442 ;
  assign n62480 = n62477 | n62479 ;
  assign n62481 = n85430 & n62480 ;
  assign n62482 = n61568 & n85426 ;
  assign n62483 = n62311 & n62482 ;
  assign n62484 = n62481 | n62483 ;
  assign n62485 = n73617 & n62484 ;
  assign n85443 = ~n62261 ;
  assign n62486 = n62260 & n85443 ;
  assign n62487 = n61585 | n62260 ;
  assign n85444 = ~n62487 ;
  assign n62488 = n62419 & n85444 ;
  assign n62489 = n62486 | n62488 ;
  assign n62490 = n85430 & n62489 ;
  assign n62491 = n61576 & n85426 ;
  assign n62492 = n62311 & n62491 ;
  assign n62493 = n62490 | n62492 ;
  assign n62494 = n73188 & n62493 ;
  assign n85445 = ~n62418 ;
  assign n62495 = n62256 & n85445 ;
  assign n62496 = n61593 | n62256 ;
  assign n85446 = ~n62496 ;
  assign n62497 = n62252 & n85446 ;
  assign n62498 = n62495 | n62497 ;
  assign n62499 = n85430 & n62498 ;
  assign n62500 = n61584 & n85426 ;
  assign n62501 = n62311 & n62500 ;
  assign n62502 = n62499 | n62501 ;
  assign n62503 = n73177 & n62502 ;
  assign n85447 = ~n62251 ;
  assign n62504 = n62250 & n85447 ;
  assign n62505 = n61601 | n62250 ;
  assign n85448 = ~n62505 ;
  assign n62506 = n62415 & n85448 ;
  assign n62507 = n62504 | n62506 ;
  assign n62508 = n85430 & n62507 ;
  assign n62509 = n61592 & n85426 ;
  assign n62510 = n62311 & n62509 ;
  assign n62511 = n62508 | n62510 ;
  assign n62512 = n72752 & n62511 ;
  assign n85449 = ~n62414 ;
  assign n62513 = n62246 & n85449 ;
  assign n62514 = n61609 | n62246 ;
  assign n85450 = ~n62514 ;
  assign n62515 = n62242 & n85450 ;
  assign n62516 = n62513 | n62515 ;
  assign n62517 = n85430 & n62516 ;
  assign n62518 = n61600 & n85426 ;
  assign n62519 = n62311 & n62518 ;
  assign n62520 = n62517 | n62519 ;
  assign n62521 = n72393 & n62520 ;
  assign n85451 = ~n62241 ;
  assign n62522 = n62240 & n85451 ;
  assign n62523 = n61617 | n62240 ;
  assign n85452 = ~n62523 ;
  assign n62524 = n62411 & n85452 ;
  assign n62525 = n62522 | n62524 ;
  assign n62526 = n85430 & n62525 ;
  assign n62527 = n61608 & n85426 ;
  assign n62528 = n62311 & n62527 ;
  assign n62529 = n62526 | n62528 ;
  assign n62530 = n72385 & n62529 ;
  assign n85453 = ~n62410 ;
  assign n62531 = n62236 & n85453 ;
  assign n62532 = n61625 | n62236 ;
  assign n85454 = ~n62532 ;
  assign n62533 = n62232 & n85454 ;
  assign n62534 = n62531 | n62533 ;
  assign n62535 = n85430 & n62534 ;
  assign n62536 = n61616 & n85426 ;
  assign n62537 = n62311 & n62536 ;
  assign n62538 = n62535 | n62537 ;
  assign n62539 = n72025 & n62538 ;
  assign n85455 = ~n62231 ;
  assign n62540 = n62230 & n85455 ;
  assign n62541 = n61633 | n62230 ;
  assign n85456 = ~n62541 ;
  assign n62542 = n62407 & n85456 ;
  assign n62543 = n62540 | n62542 ;
  assign n62544 = n85430 & n62543 ;
  assign n62545 = n61624 & n85426 ;
  assign n62546 = n62311 & n62545 ;
  assign n62547 = n62544 | n62546 ;
  assign n62548 = n71645 & n62547 ;
  assign n85457 = ~n62406 ;
  assign n62549 = n62226 & n85457 ;
  assign n62550 = n61641 | n62226 ;
  assign n85458 = ~n62550 ;
  assign n62551 = n62222 & n85458 ;
  assign n62552 = n62549 | n62551 ;
  assign n62553 = n85430 & n62552 ;
  assign n62554 = n61632 & n85426 ;
  assign n62555 = n62311 & n62554 ;
  assign n62556 = n62553 | n62555 ;
  assign n62557 = n71633 & n62556 ;
  assign n85459 = ~n62221 ;
  assign n62558 = n62220 & n85459 ;
  assign n62559 = n61649 | n62220 ;
  assign n85460 = ~n62559 ;
  assign n62560 = n62403 & n85460 ;
  assign n62561 = n62558 | n62560 ;
  assign n62562 = n85430 & n62561 ;
  assign n62563 = n61640 & n85426 ;
  assign n62564 = n62311 & n62563 ;
  assign n62565 = n62562 | n62564 ;
  assign n62566 = n71253 & n62565 ;
  assign n85461 = ~n62402 ;
  assign n62567 = n62216 & n85461 ;
  assign n62568 = n61657 | n62216 ;
  assign n85462 = ~n62568 ;
  assign n62569 = n62212 & n85462 ;
  assign n62570 = n62567 | n62569 ;
  assign n62571 = n85430 & n62570 ;
  assign n62572 = n61648 & n85426 ;
  assign n62573 = n62311 & n62572 ;
  assign n62574 = n62571 | n62573 ;
  assign n62575 = n70935 & n62574 ;
  assign n85463 = ~n62211 ;
  assign n62576 = n62209 & n85463 ;
  assign n62210 = n61665 | n62209 ;
  assign n85464 = ~n62210 ;
  assign n62577 = n62206 & n85464 ;
  assign n62578 = n62576 | n62577 ;
  assign n62579 = n85430 & n62578 ;
  assign n62580 = n61656 & n85426 ;
  assign n62581 = n62311 & n62580 ;
  assign n62582 = n62579 | n62581 ;
  assign n62583 = n70927 & n62582 ;
  assign n85465 = ~n62398 ;
  assign n62584 = n62205 & n85465 ;
  assign n62585 = n61673 | n62205 ;
  assign n85466 = ~n62585 ;
  assign n62586 = n62201 & n85466 ;
  assign n62587 = n62584 | n62586 ;
  assign n62588 = n85430 & n62587 ;
  assign n62589 = n61664 & n85426 ;
  assign n62590 = n62311 & n62589 ;
  assign n62591 = n62588 | n62590 ;
  assign n62592 = n70609 & n62591 ;
  assign n85467 = ~n62200 ;
  assign n62593 = n62199 & n85467 ;
  assign n62594 = n61681 | n62199 ;
  assign n85468 = ~n62594 ;
  assign n62595 = n62395 & n85468 ;
  assign n62596 = n62593 | n62595 ;
  assign n62597 = n85430 & n62596 ;
  assign n62598 = n61672 & n85426 ;
  assign n62599 = n62311 & n62598 ;
  assign n62600 = n62597 | n62599 ;
  assign n62601 = n70276 & n62600 ;
  assign n85469 = ~n62394 ;
  assign n62602 = n62195 & n85469 ;
  assign n62603 = n61689 | n62195 ;
  assign n85470 = ~n62603 ;
  assign n62604 = n62191 & n85470 ;
  assign n62605 = n62602 | n62604 ;
  assign n62606 = n85430 & n62605 ;
  assign n62607 = n61680 & n85426 ;
  assign n62608 = n62311 & n62607 ;
  assign n62609 = n62606 | n62608 ;
  assign n62610 = n70176 & n62609 ;
  assign n85471 = ~n62190 ;
  assign n62611 = n62189 & n85471 ;
  assign n62612 = n61697 | n62189 ;
  assign n85472 = ~n62612 ;
  assign n62613 = n62391 & n85472 ;
  assign n62614 = n62611 | n62613 ;
  assign n62615 = n85430 & n62614 ;
  assign n62616 = n61688 & n85426 ;
  assign n62617 = n62311 & n62616 ;
  assign n62618 = n62615 | n62617 ;
  assign n62619 = n69857 & n62618 ;
  assign n85473 = ~n62390 ;
  assign n62620 = n62185 & n85473 ;
  assign n62621 = n61705 | n62185 ;
  assign n85474 = ~n62621 ;
  assign n62622 = n62181 & n85474 ;
  assign n62623 = n62620 | n62622 ;
  assign n62624 = n85430 & n62623 ;
  assign n62625 = n61696 & n85426 ;
  assign n62626 = n62311 & n62625 ;
  assign n62627 = n62624 | n62626 ;
  assign n62628 = n69656 & n62627 ;
  assign n85475 = ~n62180 ;
  assign n62629 = n62179 & n85475 ;
  assign n62630 = n61713 | n62179 ;
  assign n85476 = ~n62630 ;
  assign n62631 = n62387 & n85476 ;
  assign n62632 = n62629 | n62631 ;
  assign n62633 = n85430 & n62632 ;
  assign n62634 = n61704 & n85426 ;
  assign n62635 = n62311 & n62634 ;
  assign n62636 = n62633 | n62635 ;
  assign n62637 = n69528 & n62636 ;
  assign n85477 = ~n62386 ;
  assign n62638 = n62175 & n85477 ;
  assign n62639 = n61721 | n62175 ;
  assign n85478 = ~n62639 ;
  assign n62640 = n62171 & n85478 ;
  assign n62641 = n62638 | n62640 ;
  assign n62642 = n85430 & n62641 ;
  assign n62643 = n61712 & n85426 ;
  assign n62644 = n62311 & n62643 ;
  assign n62645 = n62642 | n62644 ;
  assign n62646 = n69261 & n62645 ;
  assign n85479 = ~n62170 ;
  assign n62647 = n62169 & n85479 ;
  assign n62648 = n61729 | n62169 ;
  assign n85480 = ~n62648 ;
  assign n62649 = n62383 & n85480 ;
  assign n62650 = n62647 | n62649 ;
  assign n62651 = n85430 & n62650 ;
  assign n62652 = n61720 & n85426 ;
  assign n62653 = n62311 & n62652 ;
  assign n62654 = n62651 | n62653 ;
  assign n62655 = n69075 & n62654 ;
  assign n85481 = ~n62382 ;
  assign n62656 = n62165 & n85481 ;
  assign n62657 = n61737 | n62165 ;
  assign n85482 = ~n62657 ;
  assign n62658 = n62161 & n85482 ;
  assign n62659 = n62656 | n62658 ;
  assign n62660 = n85430 & n62659 ;
  assign n62661 = n61728 & n85426 ;
  assign n62662 = n62311 & n62661 ;
  assign n62663 = n62660 | n62662 ;
  assign n62664 = n68993 & n62663 ;
  assign n85483 = ~n62160 ;
  assign n62665 = n62159 & n85483 ;
  assign n62666 = n61745 | n62159 ;
  assign n85484 = ~n62666 ;
  assign n62667 = n62379 & n85484 ;
  assign n62668 = n62665 | n62667 ;
  assign n62669 = n85430 & n62668 ;
  assign n62670 = n61736 & n85426 ;
  assign n62671 = n62311 & n62670 ;
  assign n62672 = n62669 | n62671 ;
  assign n62673 = n68716 & n62672 ;
  assign n85485 = ~n62378 ;
  assign n62674 = n62155 & n85485 ;
  assign n62675 = n61753 | n62155 ;
  assign n85486 = ~n62675 ;
  assign n62676 = n62151 & n85486 ;
  assign n62677 = n62674 | n62676 ;
  assign n62678 = n85430 & n62677 ;
  assign n62679 = n61744 & n85426 ;
  assign n62680 = n62311 & n62679 ;
  assign n62681 = n62678 | n62680 ;
  assign n62682 = n68545 & n62681 ;
  assign n85487 = ~n62150 ;
  assign n62683 = n62149 & n85487 ;
  assign n62684 = n61761 | n62149 ;
  assign n85488 = ~n62684 ;
  assign n62685 = n62375 & n85488 ;
  assign n62686 = n62683 | n62685 ;
  assign n62687 = n85430 & n62686 ;
  assign n62688 = n61752 & n85426 ;
  assign n62689 = n62311 & n62688 ;
  assign n62690 = n62687 | n62689 ;
  assign n62691 = n68438 & n62690 ;
  assign n85489 = ~n62374 ;
  assign n62692 = n62145 & n85489 ;
  assign n62693 = n61769 | n62145 ;
  assign n85490 = ~n62693 ;
  assign n62694 = n62141 & n85490 ;
  assign n62695 = n62692 | n62694 ;
  assign n62696 = n85430 & n62695 ;
  assign n62697 = n61760 & n85426 ;
  assign n62698 = n62311 & n62697 ;
  assign n62699 = n62696 | n62698 ;
  assign n62700 = n68214 & n62699 ;
  assign n85491 = ~n62140 ;
  assign n62701 = n62139 & n85491 ;
  assign n62702 = n61777 | n62139 ;
  assign n85492 = ~n62702 ;
  assign n62703 = n62371 & n85492 ;
  assign n62704 = n62701 | n62703 ;
  assign n62705 = n85430 & n62704 ;
  assign n62706 = n61768 & n85426 ;
  assign n62707 = n62311 & n62706 ;
  assign n62708 = n62705 | n62707 ;
  assign n62709 = n68058 & n62708 ;
  assign n85493 = ~n62370 ;
  assign n62710 = n62135 & n85493 ;
  assign n62711 = n61785 | n62135 ;
  assign n85494 = ~n62711 ;
  assign n62712 = n62131 & n85494 ;
  assign n62713 = n62710 | n62712 ;
  assign n62714 = n85430 & n62713 ;
  assign n62715 = n61776 & n85426 ;
  assign n62716 = n62311 & n62715 ;
  assign n62717 = n62714 | n62716 ;
  assign n62718 = n67986 & n62717 ;
  assign n85495 = ~n62130 ;
  assign n62719 = n62128 & n85495 ;
  assign n62129 = n61793 | n62128 ;
  assign n85496 = ~n62129 ;
  assign n62720 = n62125 & n85496 ;
  assign n62721 = n62719 | n62720 ;
  assign n62722 = n85430 & n62721 ;
  assign n62723 = n61784 & n85426 ;
  assign n62724 = n62311 & n62723 ;
  assign n62725 = n62722 | n62724 ;
  assign n62726 = n67763 & n62725 ;
  assign n85497 = ~n62366 ;
  assign n62727 = n62124 & n85497 ;
  assign n62728 = n61801 | n62124 ;
  assign n85498 = ~n62728 ;
  assign n62729 = n62120 & n85498 ;
  assign n62730 = n62727 | n62729 ;
  assign n62731 = n85430 & n62730 ;
  assign n62732 = n61792 & n85426 ;
  assign n62733 = n62311 & n62732 ;
  assign n62734 = n62731 | n62733 ;
  assign n62735 = n67622 & n62734 ;
  assign n85499 = ~n62119 ;
  assign n62736 = n62118 & n85499 ;
  assign n62737 = n61809 | n62118 ;
  assign n85500 = ~n62737 ;
  assign n62738 = n62363 & n85500 ;
  assign n62739 = n62736 | n62738 ;
  assign n62740 = n85430 & n62739 ;
  assign n62741 = n61800 & n85426 ;
  assign n62742 = n62311 & n62741 ;
  assign n62743 = n62740 | n62742 ;
  assign n62744 = n67531 & n62743 ;
  assign n85501 = ~n62362 ;
  assign n62745 = n62114 & n85501 ;
  assign n62746 = n61817 | n62114 ;
  assign n85502 = ~n62746 ;
  assign n62747 = n62110 & n85502 ;
  assign n62748 = n62745 | n62747 ;
  assign n62749 = n85430 & n62748 ;
  assign n62750 = n61808 & n85426 ;
  assign n62751 = n62311 & n62750 ;
  assign n62752 = n62749 | n62751 ;
  assign n62753 = n67348 & n62752 ;
  assign n85503 = ~n62109 ;
  assign n62754 = n62108 & n85503 ;
  assign n62755 = n61825 | n62108 ;
  assign n85504 = ~n62755 ;
  assign n62756 = n62359 & n85504 ;
  assign n62757 = n62754 | n62756 ;
  assign n62758 = n85430 & n62757 ;
  assign n62759 = n61816 & n85426 ;
  assign n62760 = n62311 & n62759 ;
  assign n62761 = n62758 | n62760 ;
  assign n62762 = n67222 & n62761 ;
  assign n85505 = ~n62358 ;
  assign n62763 = n62104 & n85505 ;
  assign n62764 = n61833 | n62104 ;
  assign n85506 = ~n62764 ;
  assign n62765 = n62100 & n85506 ;
  assign n62766 = n62763 | n62765 ;
  assign n62767 = n85430 & n62766 ;
  assign n62768 = n61824 & n85426 ;
  assign n62769 = n62311 & n62768 ;
  assign n62770 = n62767 | n62769 ;
  assign n62771 = n67164 & n62770 ;
  assign n85507 = ~n62099 ;
  assign n62772 = n62098 & n85507 ;
  assign n62773 = n61841 | n62098 ;
  assign n85508 = ~n62773 ;
  assign n62774 = n62355 & n85508 ;
  assign n62775 = n62772 | n62774 ;
  assign n62776 = n85430 & n62775 ;
  assign n62777 = n61832 & n85426 ;
  assign n62778 = n62311 & n62777 ;
  assign n62779 = n62776 | n62778 ;
  assign n62780 = n66979 & n62779 ;
  assign n85509 = ~n62354 ;
  assign n62781 = n62094 & n85509 ;
  assign n62782 = n61849 | n62094 ;
  assign n85510 = ~n62782 ;
  assign n62783 = n62090 & n85510 ;
  assign n62784 = n62781 | n62783 ;
  assign n62785 = n85430 & n62784 ;
  assign n62786 = n61840 & n85426 ;
  assign n62787 = n62311 & n62786 ;
  assign n62788 = n62785 | n62787 ;
  assign n62789 = n66868 & n62788 ;
  assign n85511 = ~n62089 ;
  assign n62790 = n62088 & n85511 ;
  assign n62791 = n61857 | n62088 ;
  assign n85512 = ~n62791 ;
  assign n62792 = n62351 & n85512 ;
  assign n62793 = n62790 | n62792 ;
  assign n62794 = n85430 & n62793 ;
  assign n62795 = n61848 & n85426 ;
  assign n62796 = n62311 & n62795 ;
  assign n62797 = n62794 | n62796 ;
  assign n62798 = n66797 & n62797 ;
  assign n85513 = ~n62350 ;
  assign n62799 = n62084 & n85513 ;
  assign n62800 = n61865 | n62084 ;
  assign n85514 = ~n62800 ;
  assign n62801 = n62080 & n85514 ;
  assign n62802 = n62799 | n62801 ;
  assign n62803 = n85430 & n62802 ;
  assign n62804 = n61856 & n85426 ;
  assign n62805 = n62311 & n62804 ;
  assign n62806 = n62803 | n62805 ;
  assign n62807 = n66654 & n62806 ;
  assign n85515 = ~n62079 ;
  assign n62808 = n62078 & n85515 ;
  assign n62809 = n61873 | n62078 ;
  assign n85516 = ~n62809 ;
  assign n62810 = n62347 & n85516 ;
  assign n62811 = n62808 | n62810 ;
  assign n62812 = n85430 & n62811 ;
  assign n62813 = n61864 & n85426 ;
  assign n62814 = n62311 & n62813 ;
  assign n62815 = n62812 | n62814 ;
  assign n62816 = n66560 & n62815 ;
  assign n85517 = ~n62346 ;
  assign n62817 = n62074 & n85517 ;
  assign n62818 = n61881 | n62074 ;
  assign n85518 = ~n62818 ;
  assign n62819 = n62070 & n85518 ;
  assign n62820 = n62817 | n62819 ;
  assign n62821 = n85430 & n62820 ;
  assign n62822 = n61872 & n85426 ;
  assign n62823 = n62311 & n62822 ;
  assign n62824 = n62821 | n62823 ;
  assign n62825 = n66505 & n62824 ;
  assign n85519 = ~n62069 ;
  assign n62826 = n62068 & n85519 ;
  assign n62827 = n61889 | n62068 ;
  assign n85520 = ~n62827 ;
  assign n62828 = n62343 & n85520 ;
  assign n62829 = n62826 | n62828 ;
  assign n62830 = n85430 & n62829 ;
  assign n62831 = n61880 & n85426 ;
  assign n62832 = n62311 & n62831 ;
  assign n62833 = n62830 | n62832 ;
  assign n62834 = n66379 & n62833 ;
  assign n85521 = ~n62342 ;
  assign n62835 = n62064 & n85521 ;
  assign n62836 = n61897 | n62064 ;
  assign n85522 = ~n62836 ;
  assign n62837 = n62060 & n85522 ;
  assign n62838 = n62835 | n62837 ;
  assign n62839 = n85430 & n62838 ;
  assign n62840 = n61888 & n85426 ;
  assign n62841 = n62311 & n62840 ;
  assign n62842 = n62839 | n62841 ;
  assign n62843 = n66299 & n62842 ;
  assign n85523 = ~n62059 ;
  assign n62844 = n62058 & n85523 ;
  assign n62845 = n61905 | n62058 ;
  assign n85524 = ~n62845 ;
  assign n62846 = n62339 & n85524 ;
  assign n62847 = n62844 | n62846 ;
  assign n62848 = n85430 & n62847 ;
  assign n62849 = n61896 & n85426 ;
  assign n62850 = n62311 & n62849 ;
  assign n62851 = n62848 | n62850 ;
  assign n62852 = n66244 & n62851 ;
  assign n85525 = ~n62338 ;
  assign n62853 = n62053 & n85525 ;
  assign n62054 = n61913 | n62053 ;
  assign n85526 = ~n62054 ;
  assign n62854 = n85526 & n62337 ;
  assign n62855 = n62853 | n62854 ;
  assign n62856 = n85430 & n62855 ;
  assign n62857 = n61904 & n85426 ;
  assign n62858 = n62311 & n62857 ;
  assign n62859 = n62856 | n62858 ;
  assign n62860 = n66145 & n62859 ;
  assign n85527 = ~n62048 ;
  assign n62861 = n62047 & n85527 ;
  assign n62862 = n61921 | n62047 ;
  assign n85528 = ~n62862 ;
  assign n62863 = n62335 & n85528 ;
  assign n62864 = n62861 | n62863 ;
  assign n62865 = n85430 & n62864 ;
  assign n62866 = n61912 & n85426 ;
  assign n62867 = n62311 & n62866 ;
  assign n62868 = n62865 | n62867 ;
  assign n62869 = n66081 & n62868 ;
  assign n85529 = ~n62334 ;
  assign n62870 = n62043 & n85529 ;
  assign n62871 = n61929 | n62043 ;
  assign n85530 = ~n62871 ;
  assign n62872 = n62039 & n85530 ;
  assign n62873 = n62870 | n62872 ;
  assign n62874 = n85430 & n62873 ;
  assign n62875 = n61920 & n85426 ;
  assign n62876 = n62311 & n62875 ;
  assign n62877 = n62874 | n62876 ;
  assign n62878 = n66043 & n62877 ;
  assign n85531 = ~n62038 ;
  assign n62879 = n62037 & n85531 ;
  assign n62880 = n61937 | n62037 ;
  assign n85532 = ~n62880 ;
  assign n62881 = n62331 & n85532 ;
  assign n62882 = n62879 | n62881 ;
  assign n62883 = n85430 & n62882 ;
  assign n62884 = n61928 & n85426 ;
  assign n62885 = n62311 & n62884 ;
  assign n62886 = n62883 | n62885 ;
  assign n62887 = n65960 & n62886 ;
  assign n85533 = ~n62330 ;
  assign n62888 = n62033 & n85533 ;
  assign n62889 = n61945 | n62033 ;
  assign n85534 = ~n62889 ;
  assign n62890 = n62029 & n85534 ;
  assign n62891 = n62888 | n62890 ;
  assign n62892 = n85430 & n62891 ;
  assign n62893 = n61936 & n85426 ;
  assign n62894 = n62311 & n62893 ;
  assign n62895 = n62892 | n62894 ;
  assign n62896 = n65909 & n62895 ;
  assign n85535 = ~n62028 ;
  assign n62897 = n62027 & n85535 ;
  assign n62898 = n61953 | n62027 ;
  assign n85536 = ~n62898 ;
  assign n62899 = n62327 & n85536 ;
  assign n62900 = n62897 | n62899 ;
  assign n62901 = n85430 & n62900 ;
  assign n62902 = n61944 & n85426 ;
  assign n62903 = n62311 & n62902 ;
  assign n62904 = n62901 | n62903 ;
  assign n62905 = n65877 & n62904 ;
  assign n85537 = ~n62326 ;
  assign n62906 = n62023 & n85537 ;
  assign n62907 = n61961 | n62023 ;
  assign n85538 = ~n62907 ;
  assign n62908 = n62019 & n85538 ;
  assign n62909 = n62906 | n62908 ;
  assign n62910 = n85430 & n62909 ;
  assign n62911 = n61952 & n85426 ;
  assign n62912 = n62311 & n62911 ;
  assign n62913 = n62910 | n62912 ;
  assign n62914 = n65820 & n62913 ;
  assign n85539 = ~n62018 ;
  assign n62915 = n62017 & n85539 ;
  assign n62916 = n61969 | n62017 ;
  assign n85540 = ~n62916 ;
  assign n62917 = n62323 & n85540 ;
  assign n62918 = n62915 | n62917 ;
  assign n62919 = n85430 & n62918 ;
  assign n62920 = n61960 & n85426 ;
  assign n62921 = n62311 & n62920 ;
  assign n62922 = n62919 | n62921 ;
  assign n62923 = n65791 & n62922 ;
  assign n85541 = ~n62322 ;
  assign n62925 = n62013 & n85541 ;
  assign n62924 = n61978 | n62013 ;
  assign n85542 = ~n62924 ;
  assign n62926 = n62321 & n85542 ;
  assign n62927 = n62925 | n62926 ;
  assign n62928 = n85430 & n62927 ;
  assign n62929 = n61968 & n85426 ;
  assign n62930 = n62311 & n62929 ;
  assign n62931 = n62928 | n62930 ;
  assign n62932 = n65772 & n62931 ;
  assign n85543 = ~n62008 ;
  assign n62934 = n62007 & n85543 ;
  assign n62933 = n61986 | n62007 ;
  assign n85544 = ~n62933 ;
  assign n62935 = n62004 & n85544 ;
  assign n62936 = n62934 | n62935 ;
  assign n62937 = n85430 & n62936 ;
  assign n62938 = n61977 & n85426 ;
  assign n62939 = n62311 & n62938 ;
  assign n62940 = n62937 | n62939 ;
  assign n62941 = n65746 & n62940 ;
  assign n85545 = ~n62318 ;
  assign n62942 = n62003 & n85545 ;
  assign n62317 = n61999 | n62003 ;
  assign n85546 = ~n62317 ;
  assign n62943 = n62316 & n85546 ;
  assign n62944 = n62942 | n62943 ;
  assign n62945 = n85430 & n62944 ;
  assign n62946 = n61985 & n85426 ;
  assign n62947 = n62311 & n62946 ;
  assign n62948 = n62945 | n62947 ;
  assign n62949 = n65721 & n62948 ;
  assign n62950 = n29800 & n61995 ;
  assign n62951 = n85428 & n62950 ;
  assign n85547 = ~n62951 ;
  assign n62952 = n62316 & n85547 ;
  assign n62953 = n85430 & n62952 ;
  assign n62954 = n61998 & n85426 ;
  assign n62955 = n62311 & n62954 ;
  assign n62956 = n62953 | n62955 ;
  assign n62957 = n65686 & n62956 ;
  assign n62451 = n29800 & n85430 ;
  assign n62958 = x64 & n85430 ;
  assign n85548 = ~n62958 ;
  assign n62959 = x3 & n85548 ;
  assign n62960 = n62451 | n62959 ;
  assign n62972 = n65670 & n62960 ;
  assign n62963 = n62310 | n62962 ;
  assign n62964 = n85426 & n62963 ;
  assign n85549 = ~n62964 ;
  assign n62965 = x64 & n85549 ;
  assign n85550 = ~n62965 ;
  assign n62966 = x3 & n85550 ;
  assign n62967 = n62451 | n62966 ;
  assign n62968 = x65 & n62967 ;
  assign n62969 = x65 | n62451 ;
  assign n62970 = n62966 | n62969 ;
  assign n85551 = ~n62968 ;
  assign n62971 = n85551 & n62970 ;
  assign n62973 = n30774 | n62971 ;
  assign n85552 = ~n62972 ;
  assign n62974 = n85552 & n62973 ;
  assign n85553 = ~n62955 ;
  assign n62975 = x66 & n85553 ;
  assign n85554 = ~n62953 ;
  assign n62976 = n85554 & n62975 ;
  assign n62977 = n62957 | n62976 ;
  assign n62978 = n62974 | n62977 ;
  assign n85555 = ~n62957 ;
  assign n62979 = n85555 & n62978 ;
  assign n85556 = ~n62947 ;
  assign n62980 = x67 & n85556 ;
  assign n85557 = ~n62945 ;
  assign n62981 = n85557 & n62980 ;
  assign n62982 = n62949 | n62981 ;
  assign n62983 = n62979 | n62982 ;
  assign n85558 = ~n62949 ;
  assign n62984 = n85558 & n62983 ;
  assign n85559 = ~n62939 ;
  assign n62985 = x68 & n85559 ;
  assign n85560 = ~n62937 ;
  assign n62986 = n85560 & n62985 ;
  assign n62987 = n62941 | n62986 ;
  assign n62988 = n62984 | n62987 ;
  assign n85561 = ~n62941 ;
  assign n62989 = n85561 & n62988 ;
  assign n85562 = ~n62930 ;
  assign n62990 = x69 & n85562 ;
  assign n85563 = ~n62928 ;
  assign n62991 = n85563 & n62990 ;
  assign n62992 = n62932 | n62991 ;
  assign n62993 = n62989 | n62992 ;
  assign n85564 = ~n62932 ;
  assign n62994 = n85564 & n62993 ;
  assign n85565 = ~n62921 ;
  assign n62995 = x70 & n85565 ;
  assign n85566 = ~n62919 ;
  assign n62996 = n85566 & n62995 ;
  assign n62997 = n62923 | n62996 ;
  assign n62999 = n62994 | n62997 ;
  assign n85567 = ~n62923 ;
  assign n63000 = n85567 & n62999 ;
  assign n85568 = ~n62912 ;
  assign n63001 = x71 & n85568 ;
  assign n85569 = ~n62910 ;
  assign n63002 = n85569 & n63001 ;
  assign n63003 = n62914 | n63002 ;
  assign n63004 = n63000 | n63003 ;
  assign n85570 = ~n62914 ;
  assign n63005 = n85570 & n63004 ;
  assign n85571 = ~n62903 ;
  assign n63006 = x72 & n85571 ;
  assign n85572 = ~n62901 ;
  assign n63007 = n85572 & n63006 ;
  assign n63008 = n62905 | n63007 ;
  assign n63010 = n63005 | n63008 ;
  assign n85573 = ~n62905 ;
  assign n63011 = n85573 & n63010 ;
  assign n85574 = ~n62894 ;
  assign n63012 = x73 & n85574 ;
  assign n85575 = ~n62892 ;
  assign n63013 = n85575 & n63012 ;
  assign n63014 = n62896 | n63013 ;
  assign n63015 = n63011 | n63014 ;
  assign n85576 = ~n62896 ;
  assign n63016 = n85576 & n63015 ;
  assign n85577 = ~n62885 ;
  assign n63017 = x74 & n85577 ;
  assign n85578 = ~n62883 ;
  assign n63018 = n85578 & n63017 ;
  assign n63019 = n62887 | n63018 ;
  assign n63021 = n63016 | n63019 ;
  assign n85579 = ~n62887 ;
  assign n63022 = n85579 & n63021 ;
  assign n85580 = ~n62876 ;
  assign n63023 = x75 & n85580 ;
  assign n85581 = ~n62874 ;
  assign n63024 = n85581 & n63023 ;
  assign n63025 = n62878 | n63024 ;
  assign n63026 = n63022 | n63025 ;
  assign n85582 = ~n62878 ;
  assign n63027 = n85582 & n63026 ;
  assign n85583 = ~n62867 ;
  assign n63028 = x76 & n85583 ;
  assign n85584 = ~n62865 ;
  assign n63029 = n85584 & n63028 ;
  assign n63030 = n62869 | n63029 ;
  assign n63032 = n63027 | n63030 ;
  assign n85585 = ~n62869 ;
  assign n63033 = n85585 & n63032 ;
  assign n85586 = ~n62858 ;
  assign n63034 = x77 & n85586 ;
  assign n85587 = ~n62856 ;
  assign n63035 = n85587 & n63034 ;
  assign n63036 = n62860 | n63035 ;
  assign n63037 = n63033 | n63036 ;
  assign n85588 = ~n62860 ;
  assign n63038 = n85588 & n63037 ;
  assign n85589 = ~n62850 ;
  assign n63039 = x78 & n85589 ;
  assign n85590 = ~n62848 ;
  assign n63040 = n85590 & n63039 ;
  assign n63041 = n62852 | n63040 ;
  assign n63043 = n63038 | n63041 ;
  assign n85591 = ~n62852 ;
  assign n63044 = n85591 & n63043 ;
  assign n85592 = ~n62841 ;
  assign n63045 = x79 & n85592 ;
  assign n85593 = ~n62839 ;
  assign n63046 = n85593 & n63045 ;
  assign n63047 = n62843 | n63046 ;
  assign n63048 = n63044 | n63047 ;
  assign n85594 = ~n62843 ;
  assign n63049 = n85594 & n63048 ;
  assign n85595 = ~n62832 ;
  assign n63050 = x80 & n85595 ;
  assign n85596 = ~n62830 ;
  assign n63051 = n85596 & n63050 ;
  assign n63052 = n62834 | n63051 ;
  assign n63054 = n63049 | n63052 ;
  assign n85597 = ~n62834 ;
  assign n63055 = n85597 & n63054 ;
  assign n85598 = ~n62823 ;
  assign n63056 = x81 & n85598 ;
  assign n85599 = ~n62821 ;
  assign n63057 = n85599 & n63056 ;
  assign n63058 = n62825 | n63057 ;
  assign n63059 = n63055 | n63058 ;
  assign n85600 = ~n62825 ;
  assign n63060 = n85600 & n63059 ;
  assign n85601 = ~n62814 ;
  assign n63061 = x82 & n85601 ;
  assign n85602 = ~n62812 ;
  assign n63062 = n85602 & n63061 ;
  assign n63063 = n62816 | n63062 ;
  assign n63065 = n63060 | n63063 ;
  assign n85603 = ~n62816 ;
  assign n63066 = n85603 & n63065 ;
  assign n85604 = ~n62805 ;
  assign n63067 = x83 & n85604 ;
  assign n85605 = ~n62803 ;
  assign n63068 = n85605 & n63067 ;
  assign n63069 = n62807 | n63068 ;
  assign n63070 = n63066 | n63069 ;
  assign n85606 = ~n62807 ;
  assign n63071 = n85606 & n63070 ;
  assign n85607 = ~n62796 ;
  assign n63072 = x84 & n85607 ;
  assign n85608 = ~n62794 ;
  assign n63073 = n85608 & n63072 ;
  assign n63074 = n62798 | n63073 ;
  assign n63076 = n63071 | n63074 ;
  assign n85609 = ~n62798 ;
  assign n63077 = n85609 & n63076 ;
  assign n85610 = ~n62787 ;
  assign n63078 = x85 & n85610 ;
  assign n85611 = ~n62785 ;
  assign n63079 = n85611 & n63078 ;
  assign n63080 = n62789 | n63079 ;
  assign n63081 = n63077 | n63080 ;
  assign n85612 = ~n62789 ;
  assign n63082 = n85612 & n63081 ;
  assign n85613 = ~n62778 ;
  assign n63083 = x86 & n85613 ;
  assign n85614 = ~n62776 ;
  assign n63084 = n85614 & n63083 ;
  assign n63085 = n62780 | n63084 ;
  assign n63087 = n63082 | n63085 ;
  assign n85615 = ~n62780 ;
  assign n63088 = n85615 & n63087 ;
  assign n85616 = ~n62769 ;
  assign n63089 = x87 & n85616 ;
  assign n85617 = ~n62767 ;
  assign n63090 = n85617 & n63089 ;
  assign n63091 = n62771 | n63090 ;
  assign n63092 = n63088 | n63091 ;
  assign n85618 = ~n62771 ;
  assign n63093 = n85618 & n63092 ;
  assign n85619 = ~n62760 ;
  assign n63094 = x88 & n85619 ;
  assign n85620 = ~n62758 ;
  assign n63095 = n85620 & n63094 ;
  assign n63096 = n62762 | n63095 ;
  assign n63098 = n63093 | n63096 ;
  assign n85621 = ~n62762 ;
  assign n63099 = n85621 & n63098 ;
  assign n85622 = ~n62751 ;
  assign n63100 = x89 & n85622 ;
  assign n85623 = ~n62749 ;
  assign n63101 = n85623 & n63100 ;
  assign n63102 = n62753 | n63101 ;
  assign n63103 = n63099 | n63102 ;
  assign n85624 = ~n62753 ;
  assign n63104 = n85624 & n63103 ;
  assign n85625 = ~n62742 ;
  assign n63105 = x90 & n85625 ;
  assign n85626 = ~n62740 ;
  assign n63106 = n85626 & n63105 ;
  assign n63107 = n62744 | n63106 ;
  assign n63109 = n63104 | n63107 ;
  assign n85627 = ~n62744 ;
  assign n63110 = n85627 & n63109 ;
  assign n85628 = ~n62733 ;
  assign n63111 = x91 & n85628 ;
  assign n85629 = ~n62731 ;
  assign n63112 = n85629 & n63111 ;
  assign n63113 = n62735 | n63112 ;
  assign n63114 = n63110 | n63113 ;
  assign n85630 = ~n62735 ;
  assign n63115 = n85630 & n63114 ;
  assign n85631 = ~n62724 ;
  assign n63116 = x92 & n85631 ;
  assign n85632 = ~n62722 ;
  assign n63117 = n85632 & n63116 ;
  assign n63118 = n62726 | n63117 ;
  assign n63120 = n63115 | n63118 ;
  assign n85633 = ~n62726 ;
  assign n63121 = n85633 & n63120 ;
  assign n85634 = ~n62716 ;
  assign n63122 = x93 & n85634 ;
  assign n85635 = ~n62714 ;
  assign n63123 = n85635 & n63122 ;
  assign n63124 = n62718 | n63123 ;
  assign n63125 = n63121 | n63124 ;
  assign n85636 = ~n62718 ;
  assign n63126 = n85636 & n63125 ;
  assign n85637 = ~n62707 ;
  assign n63127 = x94 & n85637 ;
  assign n85638 = ~n62705 ;
  assign n63128 = n85638 & n63127 ;
  assign n63129 = n62709 | n63128 ;
  assign n63131 = n63126 | n63129 ;
  assign n85639 = ~n62709 ;
  assign n63132 = n85639 & n63131 ;
  assign n85640 = ~n62698 ;
  assign n63133 = x95 & n85640 ;
  assign n85641 = ~n62696 ;
  assign n63134 = n85641 & n63133 ;
  assign n63135 = n62700 | n63134 ;
  assign n63136 = n63132 | n63135 ;
  assign n85642 = ~n62700 ;
  assign n63137 = n85642 & n63136 ;
  assign n85643 = ~n62689 ;
  assign n63138 = x96 & n85643 ;
  assign n85644 = ~n62687 ;
  assign n63139 = n85644 & n63138 ;
  assign n63140 = n62691 | n63139 ;
  assign n63142 = n63137 | n63140 ;
  assign n85645 = ~n62691 ;
  assign n63143 = n85645 & n63142 ;
  assign n85646 = ~n62680 ;
  assign n63144 = x97 & n85646 ;
  assign n85647 = ~n62678 ;
  assign n63145 = n85647 & n63144 ;
  assign n63146 = n62682 | n63145 ;
  assign n63147 = n63143 | n63146 ;
  assign n85648 = ~n62682 ;
  assign n63148 = n85648 & n63147 ;
  assign n85649 = ~n62671 ;
  assign n63149 = x98 & n85649 ;
  assign n85650 = ~n62669 ;
  assign n63150 = n85650 & n63149 ;
  assign n63151 = n62673 | n63150 ;
  assign n63153 = n63148 | n63151 ;
  assign n85651 = ~n62673 ;
  assign n63154 = n85651 & n63153 ;
  assign n85652 = ~n62662 ;
  assign n63155 = x99 & n85652 ;
  assign n85653 = ~n62660 ;
  assign n63156 = n85653 & n63155 ;
  assign n63157 = n62664 | n63156 ;
  assign n63158 = n63154 | n63157 ;
  assign n85654 = ~n62664 ;
  assign n63159 = n85654 & n63158 ;
  assign n85655 = ~n62653 ;
  assign n63160 = x100 & n85655 ;
  assign n85656 = ~n62651 ;
  assign n63161 = n85656 & n63160 ;
  assign n63162 = n62655 | n63161 ;
  assign n63164 = n63159 | n63162 ;
  assign n85657 = ~n62655 ;
  assign n63165 = n85657 & n63164 ;
  assign n85658 = ~n62644 ;
  assign n63166 = x101 & n85658 ;
  assign n85659 = ~n62642 ;
  assign n63167 = n85659 & n63166 ;
  assign n63168 = n62646 | n63167 ;
  assign n63169 = n63165 | n63168 ;
  assign n85660 = ~n62646 ;
  assign n63170 = n85660 & n63169 ;
  assign n85661 = ~n62635 ;
  assign n63171 = x102 & n85661 ;
  assign n85662 = ~n62633 ;
  assign n63172 = n85662 & n63171 ;
  assign n63173 = n62637 | n63172 ;
  assign n63175 = n63170 | n63173 ;
  assign n85663 = ~n62637 ;
  assign n63176 = n85663 & n63175 ;
  assign n85664 = ~n62626 ;
  assign n63177 = x103 & n85664 ;
  assign n85665 = ~n62624 ;
  assign n63178 = n85665 & n63177 ;
  assign n63179 = n62628 | n63178 ;
  assign n63180 = n63176 | n63179 ;
  assign n85666 = ~n62628 ;
  assign n63181 = n85666 & n63180 ;
  assign n85667 = ~n62617 ;
  assign n63182 = x104 & n85667 ;
  assign n85668 = ~n62615 ;
  assign n63183 = n85668 & n63182 ;
  assign n63184 = n62619 | n63183 ;
  assign n63186 = n63181 | n63184 ;
  assign n85669 = ~n62619 ;
  assign n63187 = n85669 & n63186 ;
  assign n85670 = ~n62608 ;
  assign n63188 = x105 & n85670 ;
  assign n85671 = ~n62606 ;
  assign n63189 = n85671 & n63188 ;
  assign n63190 = n62610 | n63189 ;
  assign n63191 = n63187 | n63190 ;
  assign n85672 = ~n62610 ;
  assign n63192 = n85672 & n63191 ;
  assign n85673 = ~n62599 ;
  assign n63193 = x106 & n85673 ;
  assign n85674 = ~n62597 ;
  assign n63194 = n85674 & n63193 ;
  assign n63195 = n62601 | n63194 ;
  assign n63197 = n63192 | n63195 ;
  assign n85675 = ~n62601 ;
  assign n63198 = n85675 & n63197 ;
  assign n85676 = ~n62590 ;
  assign n63199 = x107 & n85676 ;
  assign n85677 = ~n62588 ;
  assign n63200 = n85677 & n63199 ;
  assign n63201 = n62592 | n63200 ;
  assign n63202 = n63198 | n63201 ;
  assign n85678 = ~n62592 ;
  assign n63203 = n85678 & n63202 ;
  assign n85679 = ~n62581 ;
  assign n63204 = x108 & n85679 ;
  assign n85680 = ~n62579 ;
  assign n63205 = n85680 & n63204 ;
  assign n63206 = n62583 | n63205 ;
  assign n63208 = n63203 | n63206 ;
  assign n85681 = ~n62583 ;
  assign n63209 = n85681 & n63208 ;
  assign n85682 = ~n62573 ;
  assign n63210 = x109 & n85682 ;
  assign n85683 = ~n62571 ;
  assign n63211 = n85683 & n63210 ;
  assign n63212 = n62575 | n63211 ;
  assign n63213 = n63209 | n63212 ;
  assign n85684 = ~n62575 ;
  assign n63214 = n85684 & n63213 ;
  assign n85685 = ~n62564 ;
  assign n63215 = x110 & n85685 ;
  assign n85686 = ~n62562 ;
  assign n63216 = n85686 & n63215 ;
  assign n63217 = n62566 | n63216 ;
  assign n63219 = n63214 | n63217 ;
  assign n85687 = ~n62566 ;
  assign n63220 = n85687 & n63219 ;
  assign n85688 = ~n62555 ;
  assign n63221 = x111 & n85688 ;
  assign n85689 = ~n62553 ;
  assign n63222 = n85689 & n63221 ;
  assign n63223 = n62557 | n63222 ;
  assign n63224 = n63220 | n63223 ;
  assign n85690 = ~n62557 ;
  assign n63225 = n85690 & n63224 ;
  assign n85691 = ~n62546 ;
  assign n63226 = x112 & n85691 ;
  assign n85692 = ~n62544 ;
  assign n63227 = n85692 & n63226 ;
  assign n63228 = n62548 | n63227 ;
  assign n63230 = n63225 | n63228 ;
  assign n85693 = ~n62548 ;
  assign n63231 = n85693 & n63230 ;
  assign n85694 = ~n62537 ;
  assign n63232 = x113 & n85694 ;
  assign n85695 = ~n62535 ;
  assign n63233 = n85695 & n63232 ;
  assign n63234 = n62539 | n63233 ;
  assign n63235 = n63231 | n63234 ;
  assign n85696 = ~n62539 ;
  assign n63236 = n85696 & n63235 ;
  assign n85697 = ~n62528 ;
  assign n63237 = x114 & n85697 ;
  assign n85698 = ~n62526 ;
  assign n63238 = n85698 & n63237 ;
  assign n63239 = n62530 | n63238 ;
  assign n63241 = n63236 | n63239 ;
  assign n85699 = ~n62530 ;
  assign n63242 = n85699 & n63241 ;
  assign n85700 = ~n62519 ;
  assign n63243 = x115 & n85700 ;
  assign n85701 = ~n62517 ;
  assign n63244 = n85701 & n63243 ;
  assign n63245 = n62521 | n63244 ;
  assign n63246 = n63242 | n63245 ;
  assign n85702 = ~n62521 ;
  assign n63247 = n85702 & n63246 ;
  assign n85703 = ~n62510 ;
  assign n63248 = x116 & n85703 ;
  assign n85704 = ~n62508 ;
  assign n63249 = n85704 & n63248 ;
  assign n63250 = n62512 | n63249 ;
  assign n63252 = n63247 | n63250 ;
  assign n85705 = ~n62512 ;
  assign n63253 = n85705 & n63252 ;
  assign n85706 = ~n62501 ;
  assign n63254 = x117 & n85706 ;
  assign n85707 = ~n62499 ;
  assign n63255 = n85707 & n63254 ;
  assign n63256 = n62503 | n63255 ;
  assign n63257 = n63253 | n63256 ;
  assign n85708 = ~n62503 ;
  assign n63258 = n85708 & n63257 ;
  assign n85709 = ~n62492 ;
  assign n63259 = x118 & n85709 ;
  assign n85710 = ~n62490 ;
  assign n63260 = n85710 & n63259 ;
  assign n63261 = n62494 | n63260 ;
  assign n63263 = n63258 | n63261 ;
  assign n85711 = ~n62494 ;
  assign n63264 = n85711 & n63263 ;
  assign n85712 = ~n62483 ;
  assign n63265 = x119 & n85712 ;
  assign n85713 = ~n62481 ;
  assign n63266 = n85713 & n63265 ;
  assign n63267 = n62485 | n63266 ;
  assign n63268 = n63264 | n63267 ;
  assign n85714 = ~n62485 ;
  assign n63269 = n85714 & n63268 ;
  assign n85715 = ~n62474 ;
  assign n63270 = x120 & n85715 ;
  assign n85716 = ~n62472 ;
  assign n63271 = n85716 & n63270 ;
  assign n63272 = n62476 | n63271 ;
  assign n63274 = n63269 | n63272 ;
  assign n85717 = ~n62476 ;
  assign n63275 = n85717 & n63274 ;
  assign n85718 = ~n62466 ;
  assign n63276 = x121 & n85718 ;
  assign n85719 = ~n62464 ;
  assign n63277 = n85719 & n63276 ;
  assign n63278 = n62468 | n63277 ;
  assign n63279 = n63275 | n63278 ;
  assign n85720 = ~n62468 ;
  assign n63280 = n85720 & n63279 ;
  assign n85721 = ~n62457 ;
  assign n63281 = x122 & n85721 ;
  assign n85722 = ~n62455 ;
  assign n63282 = n85722 & n63281 ;
  assign n63283 = n62459 | n63282 ;
  assign n63285 = n63280 | n63283 ;
  assign n85723 = ~n62459 ;
  assign n63286 = n85723 & n63285 ;
  assign n85724 = ~n62448 ;
  assign n63287 = x123 & n85724 ;
  assign n85725 = ~n62446 ;
  assign n63288 = n85725 & n63287 ;
  assign n63289 = n62450 | n63288 ;
  assign n63290 = n63286 | n63289 ;
  assign n85726 = ~n62450 ;
  assign n63291 = n85726 & n63290 ;
  assign n85727 = ~n62439 ;
  assign n63292 = x124 & n85727 ;
  assign n85728 = ~n62437 ;
  assign n63293 = n85728 & n63292 ;
  assign n63294 = n62441 | n63293 ;
  assign n63296 = n63291 | n63294 ;
  assign n85729 = ~n62441 ;
  assign n63297 = n85729 & n63296 ;
  assign n63308 = n75517 & n63307 ;
  assign n85730 = ~n63306 ;
  assign n63309 = x125 & n85730 ;
  assign n85731 = ~n63304 ;
  assign n63310 = n85731 & n63309 ;
  assign n63311 = n65362 | n63310 ;
  assign n63312 = n63308 | n63311 ;
  assign n63314 = n63297 | n63312 ;
  assign n85732 = ~n63313 ;
  assign n63315 = n85732 & n63314 ;
  assign n85733 = ~n63291 ;
  assign n63295 = n85733 & n63294 ;
  assign n63318 = x65 & n62960 ;
  assign n85734 = ~n63318 ;
  assign n63319 = n62970 & n85734 ;
  assign n63320 = n30774 | n63319 ;
  assign n63321 = n85552 & n63320 ;
  assign n63322 = n62977 | n63321 ;
  assign n63323 = n85555 & n63322 ;
  assign n63325 = n62982 | n63323 ;
  assign n63326 = n85558 & n63325 ;
  assign n63328 = n62987 | n63326 ;
  assign n63329 = n85561 & n63328 ;
  assign n63330 = n62992 | n63329 ;
  assign n63332 = n85564 & n63330 ;
  assign n63333 = n62997 | n63332 ;
  assign n63334 = n85567 & n63333 ;
  assign n63335 = n63003 | n63334 ;
  assign n63337 = n85570 & n63335 ;
  assign n63338 = n63008 | n63337 ;
  assign n63339 = n85573 & n63338 ;
  assign n63340 = n63014 | n63339 ;
  assign n63342 = n85576 & n63340 ;
  assign n63343 = n63019 | n63342 ;
  assign n63344 = n85579 & n63343 ;
  assign n63345 = n63025 | n63344 ;
  assign n63347 = n85582 & n63345 ;
  assign n63348 = n63030 | n63347 ;
  assign n63349 = n85585 & n63348 ;
  assign n63350 = n63036 | n63349 ;
  assign n63352 = n85588 & n63350 ;
  assign n63353 = n63041 | n63352 ;
  assign n63354 = n85591 & n63353 ;
  assign n63355 = n63047 | n63354 ;
  assign n63357 = n85594 & n63355 ;
  assign n63358 = n63052 | n63357 ;
  assign n63359 = n85597 & n63358 ;
  assign n63360 = n63058 | n63359 ;
  assign n63362 = n85600 & n63360 ;
  assign n63363 = n63063 | n63362 ;
  assign n63364 = n85603 & n63363 ;
  assign n63365 = n63069 | n63364 ;
  assign n63367 = n85606 & n63365 ;
  assign n63368 = n63074 | n63367 ;
  assign n63369 = n85609 & n63368 ;
  assign n63370 = n63080 | n63369 ;
  assign n63372 = n85612 & n63370 ;
  assign n63373 = n63085 | n63372 ;
  assign n63374 = n85615 & n63373 ;
  assign n63375 = n63091 | n63374 ;
  assign n63377 = n85618 & n63375 ;
  assign n63378 = n63096 | n63377 ;
  assign n63379 = n85621 & n63378 ;
  assign n63380 = n63102 | n63379 ;
  assign n63382 = n85624 & n63380 ;
  assign n63383 = n63107 | n63382 ;
  assign n63384 = n85627 & n63383 ;
  assign n63385 = n63113 | n63384 ;
  assign n63387 = n85630 & n63385 ;
  assign n63388 = n63118 | n63387 ;
  assign n63389 = n85633 & n63388 ;
  assign n63390 = n63124 | n63389 ;
  assign n63392 = n85636 & n63390 ;
  assign n63393 = n63129 | n63392 ;
  assign n63394 = n85639 & n63393 ;
  assign n63395 = n63135 | n63394 ;
  assign n63397 = n85642 & n63395 ;
  assign n63398 = n63140 | n63397 ;
  assign n63399 = n85645 & n63398 ;
  assign n63400 = n63146 | n63399 ;
  assign n63402 = n85648 & n63400 ;
  assign n63403 = n63151 | n63402 ;
  assign n63404 = n85651 & n63403 ;
  assign n63405 = n63157 | n63404 ;
  assign n63407 = n85654 & n63405 ;
  assign n63408 = n63162 | n63407 ;
  assign n63409 = n85657 & n63408 ;
  assign n63410 = n63168 | n63409 ;
  assign n63412 = n85660 & n63410 ;
  assign n63413 = n63173 | n63412 ;
  assign n63414 = n85663 & n63413 ;
  assign n63415 = n63179 | n63414 ;
  assign n63417 = n85666 & n63415 ;
  assign n63418 = n63184 | n63417 ;
  assign n63419 = n85669 & n63418 ;
  assign n63420 = n63190 | n63419 ;
  assign n63422 = n85672 & n63420 ;
  assign n63423 = n63195 | n63422 ;
  assign n63424 = n85675 & n63423 ;
  assign n63425 = n63201 | n63424 ;
  assign n63427 = n85678 & n63425 ;
  assign n63428 = n63206 | n63427 ;
  assign n63429 = n85681 & n63428 ;
  assign n63430 = n63212 | n63429 ;
  assign n63432 = n85684 & n63430 ;
  assign n63433 = n63217 | n63432 ;
  assign n63434 = n85687 & n63433 ;
  assign n63435 = n63223 | n63434 ;
  assign n63437 = n85690 & n63435 ;
  assign n63438 = n63228 | n63437 ;
  assign n63439 = n85693 & n63438 ;
  assign n63440 = n63234 | n63439 ;
  assign n63442 = n85696 & n63440 ;
  assign n63443 = n63239 | n63442 ;
  assign n63444 = n85699 & n63443 ;
  assign n63445 = n63245 | n63444 ;
  assign n63447 = n85702 & n63445 ;
  assign n63448 = n63250 | n63447 ;
  assign n63449 = n85705 & n63448 ;
  assign n63450 = n63256 | n63449 ;
  assign n63452 = n85708 & n63450 ;
  assign n63453 = n63261 | n63452 ;
  assign n63454 = n85711 & n63453 ;
  assign n63455 = n63267 | n63454 ;
  assign n63457 = n85714 & n63455 ;
  assign n63458 = n63272 | n63457 ;
  assign n63459 = n85717 & n63458 ;
  assign n63460 = n63278 | n63459 ;
  assign n63462 = n85720 & n63460 ;
  assign n63463 = n63283 | n63462 ;
  assign n63464 = n85723 & n63463 ;
  assign n63465 = n63289 | n63464 ;
  assign n63467 = n62450 | n63294 ;
  assign n85735 = ~n63467 ;
  assign n63468 = n63465 & n85735 ;
  assign n63469 = n63295 | n63468 ;
  assign n85736 = ~n63315 ;
  assign n63470 = n85736 & n63469 ;
  assign n63471 = n85726 & n63465 ;
  assign n63472 = n63294 | n63471 ;
  assign n63473 = n85729 & n63472 ;
  assign n63474 = n63312 | n63473 ;
  assign n63475 = n62440 & n85732 ;
  assign n63476 = n63474 & n63475 ;
  assign n63477 = n63470 | n63476 ;
  assign n63478 = n75517 & n63477 ;
  assign n85737 = ~n63476 ;
  assign n64271 = x125 & n85737 ;
  assign n85738 = ~n63470 ;
  assign n64272 = n85738 & n64271 ;
  assign n64273 = n63478 | n64272 ;
  assign n85739 = ~n63464 ;
  assign n63466 = n63289 & n85739 ;
  assign n63479 = n62459 | n63289 ;
  assign n85740 = ~n63479 ;
  assign n63480 = n63285 & n85740 ;
  assign n63481 = n63466 | n63480 ;
  assign n63482 = n85736 & n63481 ;
  assign n63483 = n62449 & n85732 ;
  assign n63484 = n63474 & n63483 ;
  assign n63485 = n63482 | n63484 ;
  assign n63486 = n75210 & n63485 ;
  assign n85741 = ~n63280 ;
  assign n63284 = n85741 & n63283 ;
  assign n63487 = n62468 | n63283 ;
  assign n85742 = ~n63487 ;
  assign n63488 = n63460 & n85742 ;
  assign n63489 = n63284 | n63488 ;
  assign n63490 = n85736 & n63489 ;
  assign n63491 = n62458 & n85732 ;
  assign n63492 = n63474 & n63491 ;
  assign n63493 = n63490 | n63492 ;
  assign n63494 = n74905 & n63493 ;
  assign n85743 = ~n63492 ;
  assign n64260 = x123 & n85743 ;
  assign n85744 = ~n63490 ;
  assign n64261 = n85744 & n64260 ;
  assign n64262 = n63494 | n64261 ;
  assign n85745 = ~n63459 ;
  assign n63461 = n63278 & n85745 ;
  assign n63495 = n62476 | n63278 ;
  assign n85746 = ~n63495 ;
  assign n63496 = n63274 & n85746 ;
  assign n63497 = n63461 | n63496 ;
  assign n63498 = n85736 & n63497 ;
  assign n63499 = n62467 & n85732 ;
  assign n63500 = n63474 & n63499 ;
  assign n63501 = n63498 | n63500 ;
  assign n63502 = n74431 & n63501 ;
  assign n85747 = ~n63269 ;
  assign n63273 = n85747 & n63272 ;
  assign n63503 = n62485 | n63272 ;
  assign n85748 = ~n63503 ;
  assign n63504 = n63455 & n85748 ;
  assign n63505 = n63273 | n63504 ;
  assign n63506 = n85736 & n63505 ;
  assign n63507 = n62475 & n85732 ;
  assign n63508 = n63474 & n63507 ;
  assign n63509 = n63506 | n63508 ;
  assign n63510 = n74029 & n63509 ;
  assign n85749 = ~n63508 ;
  assign n64250 = x121 & n85749 ;
  assign n85750 = ~n63506 ;
  assign n64251 = n85750 & n64250 ;
  assign n64252 = n63510 | n64251 ;
  assign n85751 = ~n63454 ;
  assign n63456 = n63267 & n85751 ;
  assign n63511 = n62494 | n63267 ;
  assign n85752 = ~n63511 ;
  assign n63512 = n63263 & n85752 ;
  assign n63513 = n63456 | n63512 ;
  assign n63514 = n85736 & n63513 ;
  assign n63515 = n62484 & n85732 ;
  assign n63516 = n63474 & n63515 ;
  assign n63517 = n63514 | n63516 ;
  assign n63518 = n74021 & n63517 ;
  assign n85753 = ~n63258 ;
  assign n63262 = n85753 & n63261 ;
  assign n63519 = n62503 | n63261 ;
  assign n85754 = ~n63519 ;
  assign n63520 = n63450 & n85754 ;
  assign n63521 = n63262 | n63520 ;
  assign n63522 = n85736 & n63521 ;
  assign n63523 = n62493 & n85732 ;
  assign n63524 = n63474 & n63523 ;
  assign n63525 = n63522 | n63524 ;
  assign n63526 = n73617 & n63525 ;
  assign n85755 = ~n63524 ;
  assign n64239 = x119 & n85755 ;
  assign n85756 = ~n63522 ;
  assign n64240 = n85756 & n64239 ;
  assign n64241 = n63526 | n64240 ;
  assign n85757 = ~n63449 ;
  assign n63451 = n63256 & n85757 ;
  assign n63527 = n62512 | n63256 ;
  assign n85758 = ~n63527 ;
  assign n63528 = n63252 & n85758 ;
  assign n63529 = n63451 | n63528 ;
  assign n63530 = n85736 & n63529 ;
  assign n63531 = n62502 & n85732 ;
  assign n63532 = n63474 & n63531 ;
  assign n63533 = n63530 | n63532 ;
  assign n63534 = n73188 & n63533 ;
  assign n85759 = ~n63247 ;
  assign n63251 = n85759 & n63250 ;
  assign n63535 = n62521 | n63250 ;
  assign n85760 = ~n63535 ;
  assign n63536 = n63445 & n85760 ;
  assign n63537 = n63251 | n63536 ;
  assign n63538 = n85736 & n63537 ;
  assign n63539 = n62511 & n85732 ;
  assign n63540 = n63474 & n63539 ;
  assign n63541 = n63538 | n63540 ;
  assign n63542 = n73177 & n63541 ;
  assign n85761 = ~n63540 ;
  assign n64229 = x117 & n85761 ;
  assign n85762 = ~n63538 ;
  assign n64230 = n85762 & n64229 ;
  assign n64231 = n63542 | n64230 ;
  assign n85763 = ~n63444 ;
  assign n63446 = n63245 & n85763 ;
  assign n63543 = n62530 | n63245 ;
  assign n85764 = ~n63543 ;
  assign n63544 = n63241 & n85764 ;
  assign n63545 = n63446 | n63544 ;
  assign n63546 = n85736 & n63545 ;
  assign n63547 = n62520 & n85732 ;
  assign n63548 = n63474 & n63547 ;
  assign n63549 = n63546 | n63548 ;
  assign n63550 = n72752 & n63549 ;
  assign n85765 = ~n63236 ;
  assign n63240 = n85765 & n63239 ;
  assign n63551 = n62539 | n63239 ;
  assign n85766 = ~n63551 ;
  assign n63552 = n63440 & n85766 ;
  assign n63553 = n63240 | n63552 ;
  assign n63554 = n85736 & n63553 ;
  assign n63555 = n62529 & n85732 ;
  assign n63556 = n63474 & n63555 ;
  assign n63557 = n63554 | n63556 ;
  assign n63558 = n72393 & n63557 ;
  assign n85767 = ~n63556 ;
  assign n64218 = x115 & n85767 ;
  assign n85768 = ~n63554 ;
  assign n64219 = n85768 & n64218 ;
  assign n64220 = n63558 | n64219 ;
  assign n85769 = ~n63439 ;
  assign n63441 = n63234 & n85769 ;
  assign n63559 = n62548 | n63234 ;
  assign n85770 = ~n63559 ;
  assign n63560 = n63230 & n85770 ;
  assign n63561 = n63441 | n63560 ;
  assign n63562 = n85736 & n63561 ;
  assign n63563 = n62538 & n85732 ;
  assign n63564 = n63474 & n63563 ;
  assign n63565 = n63562 | n63564 ;
  assign n63566 = n72385 & n63565 ;
  assign n85771 = ~n63225 ;
  assign n63229 = n85771 & n63228 ;
  assign n63567 = n62557 | n63228 ;
  assign n85772 = ~n63567 ;
  assign n63568 = n63435 & n85772 ;
  assign n63569 = n63229 | n63568 ;
  assign n63570 = n85736 & n63569 ;
  assign n63571 = n62547 & n85732 ;
  assign n63572 = n63474 & n63571 ;
  assign n63573 = n63570 | n63572 ;
  assign n63574 = n72025 & n63573 ;
  assign n85773 = ~n63572 ;
  assign n64207 = x113 & n85773 ;
  assign n85774 = ~n63570 ;
  assign n64208 = n85774 & n64207 ;
  assign n64209 = n63574 | n64208 ;
  assign n85775 = ~n63434 ;
  assign n63436 = n63223 & n85775 ;
  assign n63575 = n62566 | n63223 ;
  assign n85776 = ~n63575 ;
  assign n63576 = n63219 & n85776 ;
  assign n63577 = n63436 | n63576 ;
  assign n63578 = n85736 & n63577 ;
  assign n63579 = n62556 & n85732 ;
  assign n63580 = n63474 & n63579 ;
  assign n63581 = n63578 | n63580 ;
  assign n63582 = n71645 & n63581 ;
  assign n85777 = ~n63214 ;
  assign n63218 = n85777 & n63217 ;
  assign n63583 = n62575 | n63217 ;
  assign n85778 = ~n63583 ;
  assign n63584 = n63430 & n85778 ;
  assign n63585 = n63218 | n63584 ;
  assign n63586 = n85736 & n63585 ;
  assign n63587 = n62565 & n85732 ;
  assign n63588 = n63474 & n63587 ;
  assign n63589 = n63586 | n63588 ;
  assign n63590 = n71633 & n63589 ;
  assign n85779 = ~n63588 ;
  assign n64197 = x111 & n85779 ;
  assign n85780 = ~n63586 ;
  assign n64198 = n85780 & n64197 ;
  assign n64199 = n63590 | n64198 ;
  assign n85781 = ~n63429 ;
  assign n63431 = n63212 & n85781 ;
  assign n63591 = n62583 | n63212 ;
  assign n85782 = ~n63591 ;
  assign n63592 = n63208 & n85782 ;
  assign n63593 = n63431 | n63592 ;
  assign n63594 = n85736 & n63593 ;
  assign n63595 = n62574 & n85732 ;
  assign n63596 = n63474 & n63595 ;
  assign n63597 = n63594 | n63596 ;
  assign n63598 = n71253 & n63597 ;
  assign n85783 = ~n63203 ;
  assign n63207 = n85783 & n63206 ;
  assign n63599 = n62592 | n63206 ;
  assign n85784 = ~n63599 ;
  assign n63600 = n63425 & n85784 ;
  assign n63601 = n63207 | n63600 ;
  assign n63602 = n85736 & n63601 ;
  assign n63603 = n62582 & n85732 ;
  assign n63604 = n63474 & n63603 ;
  assign n63605 = n63602 | n63604 ;
  assign n63606 = n70935 & n63605 ;
  assign n85785 = ~n63604 ;
  assign n64185 = x109 & n85785 ;
  assign n85786 = ~n63602 ;
  assign n64186 = n85786 & n64185 ;
  assign n64187 = n63606 | n64186 ;
  assign n85787 = ~n63424 ;
  assign n63426 = n63201 & n85787 ;
  assign n63607 = n62601 | n63201 ;
  assign n85788 = ~n63607 ;
  assign n63608 = n63197 & n85788 ;
  assign n63609 = n63426 | n63608 ;
  assign n63610 = n85736 & n63609 ;
  assign n63611 = n62591 & n85732 ;
  assign n63612 = n63474 & n63611 ;
  assign n63613 = n63610 | n63612 ;
  assign n63614 = n70927 & n63613 ;
  assign n85789 = ~n63192 ;
  assign n63196 = n85789 & n63195 ;
  assign n63615 = n62610 | n63195 ;
  assign n85790 = ~n63615 ;
  assign n63616 = n63420 & n85790 ;
  assign n63617 = n63196 | n63616 ;
  assign n63618 = n85736 & n63617 ;
  assign n63619 = n62600 & n85732 ;
  assign n63620 = n63474 & n63619 ;
  assign n63621 = n63618 | n63620 ;
  assign n63622 = n70609 & n63621 ;
  assign n85791 = ~n63620 ;
  assign n64175 = x107 & n85791 ;
  assign n85792 = ~n63618 ;
  assign n64176 = n85792 & n64175 ;
  assign n64177 = n63622 | n64176 ;
  assign n85793 = ~n63419 ;
  assign n63421 = n63190 & n85793 ;
  assign n63623 = n62619 | n63190 ;
  assign n85794 = ~n63623 ;
  assign n63624 = n63186 & n85794 ;
  assign n63625 = n63421 | n63624 ;
  assign n63626 = n85736 & n63625 ;
  assign n63627 = n62609 & n85732 ;
  assign n63628 = n63474 & n63627 ;
  assign n63629 = n63626 | n63628 ;
  assign n63630 = n70276 & n63629 ;
  assign n85795 = ~n63181 ;
  assign n63185 = n85795 & n63184 ;
  assign n63631 = n62628 | n63184 ;
  assign n85796 = ~n63631 ;
  assign n63632 = n63415 & n85796 ;
  assign n63633 = n63185 | n63632 ;
  assign n63634 = n85736 & n63633 ;
  assign n63635 = n62618 & n85732 ;
  assign n63636 = n63474 & n63635 ;
  assign n63637 = n63634 | n63636 ;
  assign n63638 = n70176 & n63637 ;
  assign n85797 = ~n63636 ;
  assign n64164 = x105 & n85797 ;
  assign n85798 = ~n63634 ;
  assign n64165 = n85798 & n64164 ;
  assign n64166 = n63638 | n64165 ;
  assign n85799 = ~n63414 ;
  assign n63416 = n63179 & n85799 ;
  assign n63639 = n62637 | n63179 ;
  assign n85800 = ~n63639 ;
  assign n63640 = n63175 & n85800 ;
  assign n63641 = n63416 | n63640 ;
  assign n63642 = n85736 & n63641 ;
  assign n63643 = n62627 & n85732 ;
  assign n63644 = n63474 & n63643 ;
  assign n63645 = n63642 | n63644 ;
  assign n63646 = n69857 & n63645 ;
  assign n85801 = ~n63170 ;
  assign n63174 = n85801 & n63173 ;
  assign n63647 = n62646 | n63173 ;
  assign n85802 = ~n63647 ;
  assign n63648 = n63410 & n85802 ;
  assign n63649 = n63174 | n63648 ;
  assign n63650 = n85736 & n63649 ;
  assign n63651 = n62636 & n85732 ;
  assign n63652 = n63474 & n63651 ;
  assign n63653 = n63650 | n63652 ;
  assign n63654 = n69656 & n63653 ;
  assign n85803 = ~n63652 ;
  assign n64154 = x103 & n85803 ;
  assign n85804 = ~n63650 ;
  assign n64155 = n85804 & n64154 ;
  assign n64156 = n63654 | n64155 ;
  assign n85805 = ~n63409 ;
  assign n63411 = n63168 & n85805 ;
  assign n63655 = n62655 | n63168 ;
  assign n85806 = ~n63655 ;
  assign n63656 = n63164 & n85806 ;
  assign n63657 = n63411 | n63656 ;
  assign n63658 = n85736 & n63657 ;
  assign n63659 = n62645 & n85732 ;
  assign n63660 = n63474 & n63659 ;
  assign n63661 = n63658 | n63660 ;
  assign n63662 = n69528 & n63661 ;
  assign n85807 = ~n63159 ;
  assign n63163 = n85807 & n63162 ;
  assign n63663 = n62664 | n63162 ;
  assign n85808 = ~n63663 ;
  assign n63664 = n63405 & n85808 ;
  assign n63665 = n63163 | n63664 ;
  assign n63666 = n85736 & n63665 ;
  assign n63667 = n62654 & n85732 ;
  assign n63668 = n63474 & n63667 ;
  assign n63669 = n63666 | n63668 ;
  assign n63670 = n69261 & n63669 ;
  assign n85809 = ~n63668 ;
  assign n64144 = x101 & n85809 ;
  assign n85810 = ~n63666 ;
  assign n64145 = n85810 & n64144 ;
  assign n64146 = n63670 | n64145 ;
  assign n85811 = ~n63404 ;
  assign n63406 = n63157 & n85811 ;
  assign n63671 = n62673 | n63157 ;
  assign n85812 = ~n63671 ;
  assign n63672 = n63153 & n85812 ;
  assign n63673 = n63406 | n63672 ;
  assign n63674 = n85736 & n63673 ;
  assign n63675 = n62663 & n85732 ;
  assign n63676 = n63474 & n63675 ;
  assign n63677 = n63674 | n63676 ;
  assign n63678 = n69075 & n63677 ;
  assign n85813 = ~n63148 ;
  assign n63152 = n85813 & n63151 ;
  assign n63679 = n62682 | n63151 ;
  assign n85814 = ~n63679 ;
  assign n63680 = n63400 & n85814 ;
  assign n63681 = n63152 | n63680 ;
  assign n63682 = n85736 & n63681 ;
  assign n63683 = n62672 & n85732 ;
  assign n63684 = n63474 & n63683 ;
  assign n63685 = n63682 | n63684 ;
  assign n63686 = n68993 & n63685 ;
  assign n85815 = ~n63684 ;
  assign n64134 = x99 & n85815 ;
  assign n85816 = ~n63682 ;
  assign n64135 = n85816 & n64134 ;
  assign n64136 = n63686 | n64135 ;
  assign n85817 = ~n63399 ;
  assign n63401 = n63146 & n85817 ;
  assign n63687 = n62691 | n63146 ;
  assign n85818 = ~n63687 ;
  assign n63688 = n63142 & n85818 ;
  assign n63689 = n63401 | n63688 ;
  assign n63690 = n85736 & n63689 ;
  assign n63691 = n62681 & n85732 ;
  assign n63692 = n63474 & n63691 ;
  assign n63693 = n63690 | n63692 ;
  assign n63694 = n68716 & n63693 ;
  assign n85819 = ~n63137 ;
  assign n63141 = n85819 & n63140 ;
  assign n63695 = n62700 | n63140 ;
  assign n85820 = ~n63695 ;
  assign n63696 = n63395 & n85820 ;
  assign n63697 = n63141 | n63696 ;
  assign n63698 = n85736 & n63697 ;
  assign n63699 = n62690 & n85732 ;
  assign n63700 = n63474 & n63699 ;
  assign n63701 = n63698 | n63700 ;
  assign n63702 = n68545 & n63701 ;
  assign n85821 = ~n63700 ;
  assign n64124 = x97 & n85821 ;
  assign n85822 = ~n63698 ;
  assign n64125 = n85822 & n64124 ;
  assign n64126 = n63702 | n64125 ;
  assign n85823 = ~n63394 ;
  assign n63396 = n63135 & n85823 ;
  assign n63703 = n62709 | n63135 ;
  assign n85824 = ~n63703 ;
  assign n63704 = n63131 & n85824 ;
  assign n63705 = n63396 | n63704 ;
  assign n63706 = n85736 & n63705 ;
  assign n63707 = n62699 & n85732 ;
  assign n63708 = n63474 & n63707 ;
  assign n63709 = n63706 | n63708 ;
  assign n63710 = n68438 & n63709 ;
  assign n85825 = ~n63126 ;
  assign n63130 = n85825 & n63129 ;
  assign n63711 = n62718 | n63129 ;
  assign n85826 = ~n63711 ;
  assign n63712 = n63390 & n85826 ;
  assign n63713 = n63130 | n63712 ;
  assign n63714 = n85736 & n63713 ;
  assign n63715 = n62708 & n85732 ;
  assign n63716 = n63474 & n63715 ;
  assign n63717 = n63714 | n63716 ;
  assign n63718 = n68214 & n63717 ;
  assign n85827 = ~n63716 ;
  assign n64114 = x95 & n85827 ;
  assign n85828 = ~n63714 ;
  assign n64115 = n85828 & n64114 ;
  assign n64116 = n63718 | n64115 ;
  assign n85829 = ~n63389 ;
  assign n63391 = n63124 & n85829 ;
  assign n63719 = n62726 | n63124 ;
  assign n85830 = ~n63719 ;
  assign n63720 = n63120 & n85830 ;
  assign n63721 = n63391 | n63720 ;
  assign n63722 = n85736 & n63721 ;
  assign n63723 = n62717 & n85732 ;
  assign n63724 = n63474 & n63723 ;
  assign n63725 = n63722 | n63724 ;
  assign n63726 = n68058 & n63725 ;
  assign n85831 = ~n63115 ;
  assign n63119 = n85831 & n63118 ;
  assign n63727 = n62735 | n63118 ;
  assign n85832 = ~n63727 ;
  assign n63728 = n63385 & n85832 ;
  assign n63729 = n63119 | n63728 ;
  assign n63730 = n85736 & n63729 ;
  assign n63731 = n62725 & n85732 ;
  assign n63732 = n63474 & n63731 ;
  assign n63733 = n63730 | n63732 ;
  assign n63734 = n67986 & n63733 ;
  assign n85833 = ~n63732 ;
  assign n64104 = x93 & n85833 ;
  assign n85834 = ~n63730 ;
  assign n64105 = n85834 & n64104 ;
  assign n64106 = n63734 | n64105 ;
  assign n85835 = ~n63384 ;
  assign n63386 = n63113 & n85835 ;
  assign n63735 = n62744 | n63113 ;
  assign n85836 = ~n63735 ;
  assign n63736 = n63109 & n85836 ;
  assign n63737 = n63386 | n63736 ;
  assign n63738 = n85736 & n63737 ;
  assign n63739 = n62734 & n85732 ;
  assign n63740 = n63474 & n63739 ;
  assign n63741 = n63738 | n63740 ;
  assign n63742 = n67763 & n63741 ;
  assign n85837 = ~n63104 ;
  assign n63108 = n85837 & n63107 ;
  assign n63743 = n62753 | n63107 ;
  assign n85838 = ~n63743 ;
  assign n63744 = n63380 & n85838 ;
  assign n63745 = n63108 | n63744 ;
  assign n63746 = n85736 & n63745 ;
  assign n63747 = n62743 & n85732 ;
  assign n63748 = n63474 & n63747 ;
  assign n63749 = n63746 | n63748 ;
  assign n63750 = n67622 & n63749 ;
  assign n85839 = ~n63748 ;
  assign n64094 = x91 & n85839 ;
  assign n85840 = ~n63746 ;
  assign n64095 = n85840 & n64094 ;
  assign n64096 = n63750 | n64095 ;
  assign n85841 = ~n63379 ;
  assign n63381 = n63102 & n85841 ;
  assign n63751 = n62762 | n63102 ;
  assign n85842 = ~n63751 ;
  assign n63752 = n63098 & n85842 ;
  assign n63753 = n63381 | n63752 ;
  assign n63754 = n85736 & n63753 ;
  assign n63755 = n62752 & n85732 ;
  assign n63756 = n63474 & n63755 ;
  assign n63757 = n63754 | n63756 ;
  assign n63758 = n67531 & n63757 ;
  assign n85843 = ~n63093 ;
  assign n63097 = n85843 & n63096 ;
  assign n63759 = n62771 | n63096 ;
  assign n85844 = ~n63759 ;
  assign n63760 = n63375 & n85844 ;
  assign n63761 = n63097 | n63760 ;
  assign n63762 = n85736 & n63761 ;
  assign n63763 = n62761 & n85732 ;
  assign n63764 = n63474 & n63763 ;
  assign n63765 = n63762 | n63764 ;
  assign n63766 = n67348 & n63765 ;
  assign n85845 = ~n63764 ;
  assign n64083 = x89 & n85845 ;
  assign n85846 = ~n63762 ;
  assign n64084 = n85846 & n64083 ;
  assign n64085 = n63766 | n64084 ;
  assign n85847 = ~n63374 ;
  assign n63376 = n63091 & n85847 ;
  assign n63767 = n62780 | n63091 ;
  assign n85848 = ~n63767 ;
  assign n63768 = n63087 & n85848 ;
  assign n63769 = n63376 | n63768 ;
  assign n63770 = n85736 & n63769 ;
  assign n63771 = n62770 & n85732 ;
  assign n63772 = n63474 & n63771 ;
  assign n63773 = n63770 | n63772 ;
  assign n63774 = n67222 & n63773 ;
  assign n85849 = ~n63082 ;
  assign n63086 = n85849 & n63085 ;
  assign n63775 = n62789 | n63085 ;
  assign n85850 = ~n63775 ;
  assign n63776 = n63370 & n85850 ;
  assign n63777 = n63086 | n63776 ;
  assign n63778 = n85736 & n63777 ;
  assign n63779 = n62779 & n85732 ;
  assign n63780 = n63474 & n63779 ;
  assign n63781 = n63778 | n63780 ;
  assign n63782 = n67164 & n63781 ;
  assign n85851 = ~n63780 ;
  assign n64073 = x87 & n85851 ;
  assign n85852 = ~n63778 ;
  assign n64074 = n85852 & n64073 ;
  assign n64075 = n63782 | n64074 ;
  assign n85853 = ~n63369 ;
  assign n63371 = n63080 & n85853 ;
  assign n63783 = n62798 | n63080 ;
  assign n85854 = ~n63783 ;
  assign n63784 = n63076 & n85854 ;
  assign n63785 = n63371 | n63784 ;
  assign n63786 = n85736 & n63785 ;
  assign n63787 = n62788 & n85732 ;
  assign n63788 = n63474 & n63787 ;
  assign n63789 = n63786 | n63788 ;
  assign n63790 = n66979 & n63789 ;
  assign n85855 = ~n63071 ;
  assign n63075 = n85855 & n63074 ;
  assign n63791 = n62807 | n63074 ;
  assign n85856 = ~n63791 ;
  assign n63792 = n63365 & n85856 ;
  assign n63793 = n63075 | n63792 ;
  assign n63794 = n85736 & n63793 ;
  assign n63795 = n62797 & n85732 ;
  assign n63796 = n63474 & n63795 ;
  assign n63797 = n63794 | n63796 ;
  assign n63798 = n66868 & n63797 ;
  assign n85857 = ~n63796 ;
  assign n64063 = x85 & n85857 ;
  assign n85858 = ~n63794 ;
  assign n64064 = n85858 & n64063 ;
  assign n64065 = n63798 | n64064 ;
  assign n85859 = ~n63364 ;
  assign n63366 = n63069 & n85859 ;
  assign n63799 = n62816 | n63069 ;
  assign n85860 = ~n63799 ;
  assign n63800 = n63065 & n85860 ;
  assign n63801 = n63366 | n63800 ;
  assign n63802 = n85736 & n63801 ;
  assign n63803 = n62806 & n85732 ;
  assign n63804 = n63474 & n63803 ;
  assign n63805 = n63802 | n63804 ;
  assign n63806 = n66797 & n63805 ;
  assign n85861 = ~n63060 ;
  assign n63064 = n85861 & n63063 ;
  assign n63807 = n62825 | n63063 ;
  assign n85862 = ~n63807 ;
  assign n63808 = n63360 & n85862 ;
  assign n63809 = n63064 | n63808 ;
  assign n63810 = n85736 & n63809 ;
  assign n63811 = n62815 & n85732 ;
  assign n63812 = n63474 & n63811 ;
  assign n63813 = n63810 | n63812 ;
  assign n63814 = n66654 & n63813 ;
  assign n85863 = ~n63812 ;
  assign n64053 = x83 & n85863 ;
  assign n85864 = ~n63810 ;
  assign n64054 = n85864 & n64053 ;
  assign n64055 = n63814 | n64054 ;
  assign n85865 = ~n63359 ;
  assign n63361 = n63058 & n85865 ;
  assign n63815 = n62834 | n63058 ;
  assign n85866 = ~n63815 ;
  assign n63816 = n63054 & n85866 ;
  assign n63817 = n63361 | n63816 ;
  assign n63818 = n85736 & n63817 ;
  assign n63819 = n62824 & n85732 ;
  assign n63820 = n63474 & n63819 ;
  assign n63821 = n63818 | n63820 ;
  assign n63822 = n66560 & n63821 ;
  assign n85867 = ~n63049 ;
  assign n63053 = n85867 & n63052 ;
  assign n63823 = n62843 | n63052 ;
  assign n85868 = ~n63823 ;
  assign n63824 = n63355 & n85868 ;
  assign n63825 = n63053 | n63824 ;
  assign n63826 = n85736 & n63825 ;
  assign n63827 = n62833 & n85732 ;
  assign n63828 = n63474 & n63827 ;
  assign n63829 = n63826 | n63828 ;
  assign n63830 = n66505 & n63829 ;
  assign n85869 = ~n63828 ;
  assign n64043 = x81 & n85869 ;
  assign n85870 = ~n63826 ;
  assign n64044 = n85870 & n64043 ;
  assign n64045 = n63830 | n64044 ;
  assign n85871 = ~n63354 ;
  assign n63356 = n63047 & n85871 ;
  assign n63831 = n62852 | n63047 ;
  assign n85872 = ~n63831 ;
  assign n63832 = n63043 & n85872 ;
  assign n63833 = n63356 | n63832 ;
  assign n63834 = n85736 & n63833 ;
  assign n63835 = n62842 & n85732 ;
  assign n63836 = n63474 & n63835 ;
  assign n63837 = n63834 | n63836 ;
  assign n63838 = n66379 & n63837 ;
  assign n85873 = ~n63038 ;
  assign n63042 = n85873 & n63041 ;
  assign n63839 = n62860 | n63041 ;
  assign n85874 = ~n63839 ;
  assign n63840 = n63350 & n85874 ;
  assign n63841 = n63042 | n63840 ;
  assign n63842 = n85736 & n63841 ;
  assign n63843 = n62851 & n85732 ;
  assign n63844 = n63474 & n63843 ;
  assign n63845 = n63842 | n63844 ;
  assign n63846 = n66299 & n63845 ;
  assign n85875 = ~n63844 ;
  assign n64032 = x79 & n85875 ;
  assign n85876 = ~n63842 ;
  assign n64033 = n85876 & n64032 ;
  assign n64034 = n63846 | n64033 ;
  assign n85877 = ~n63349 ;
  assign n63351 = n63036 & n85877 ;
  assign n63847 = n62869 | n63036 ;
  assign n85878 = ~n63847 ;
  assign n63848 = n63032 & n85878 ;
  assign n63849 = n63351 | n63848 ;
  assign n63850 = n85736 & n63849 ;
  assign n63851 = n62859 & n85732 ;
  assign n63852 = n63474 & n63851 ;
  assign n63853 = n63850 | n63852 ;
  assign n63854 = n66244 & n63853 ;
  assign n85879 = ~n63027 ;
  assign n63031 = n85879 & n63030 ;
  assign n63855 = n62878 | n63030 ;
  assign n85880 = ~n63855 ;
  assign n63856 = n63345 & n85880 ;
  assign n63857 = n63031 | n63856 ;
  assign n63858 = n85736 & n63857 ;
  assign n63859 = n62868 & n85732 ;
  assign n63860 = n63474 & n63859 ;
  assign n63861 = n63858 | n63860 ;
  assign n63862 = n66145 & n63861 ;
  assign n85881 = ~n63860 ;
  assign n64022 = x77 & n85881 ;
  assign n85882 = ~n63858 ;
  assign n64023 = n85882 & n64022 ;
  assign n64024 = n63862 | n64023 ;
  assign n85883 = ~n63344 ;
  assign n63346 = n63025 & n85883 ;
  assign n63863 = n62887 | n63025 ;
  assign n85884 = ~n63863 ;
  assign n63864 = n63021 & n85884 ;
  assign n63865 = n63346 | n63864 ;
  assign n63866 = n85736 & n63865 ;
  assign n63867 = n62877 & n85732 ;
  assign n63868 = n63474 & n63867 ;
  assign n63869 = n63866 | n63868 ;
  assign n63870 = n66081 & n63869 ;
  assign n85885 = ~n63016 ;
  assign n63020 = n85885 & n63019 ;
  assign n63871 = n62896 | n63019 ;
  assign n85886 = ~n63871 ;
  assign n63872 = n63340 & n85886 ;
  assign n63873 = n63020 | n63872 ;
  assign n63874 = n85736 & n63873 ;
  assign n63875 = n62886 & n85732 ;
  assign n63876 = n63474 & n63875 ;
  assign n63877 = n63874 | n63876 ;
  assign n63878 = n66043 & n63877 ;
  assign n85887 = ~n63876 ;
  assign n64011 = x75 & n85887 ;
  assign n85888 = ~n63874 ;
  assign n64012 = n85888 & n64011 ;
  assign n64013 = n63878 | n64012 ;
  assign n85889 = ~n63339 ;
  assign n63341 = n63014 & n85889 ;
  assign n63879 = n62905 | n63014 ;
  assign n85890 = ~n63879 ;
  assign n63880 = n63010 & n85890 ;
  assign n63881 = n63341 | n63880 ;
  assign n63882 = n85736 & n63881 ;
  assign n63883 = n62895 & n85732 ;
  assign n63884 = n63474 & n63883 ;
  assign n63885 = n63882 | n63884 ;
  assign n63886 = n65960 & n63885 ;
  assign n85891 = ~n63005 ;
  assign n63009 = n85891 & n63008 ;
  assign n63887 = n62914 | n63008 ;
  assign n85892 = ~n63887 ;
  assign n63888 = n63335 & n85892 ;
  assign n63889 = n63009 | n63888 ;
  assign n63890 = n85736 & n63889 ;
  assign n63891 = n62904 & n85732 ;
  assign n63892 = n63474 & n63891 ;
  assign n63893 = n63890 | n63892 ;
  assign n63894 = n65909 & n63893 ;
  assign n85893 = ~n63892 ;
  assign n64001 = x73 & n85893 ;
  assign n85894 = ~n63890 ;
  assign n64002 = n85894 & n64001 ;
  assign n64003 = n63894 | n64002 ;
  assign n85895 = ~n63334 ;
  assign n63336 = n63003 & n85895 ;
  assign n63895 = n62923 | n63003 ;
  assign n85896 = ~n63895 ;
  assign n63896 = n62999 & n85896 ;
  assign n63897 = n63336 | n63896 ;
  assign n63898 = n85736 & n63897 ;
  assign n63899 = n62913 & n85732 ;
  assign n63900 = n63474 & n63899 ;
  assign n63901 = n63898 | n63900 ;
  assign n63902 = n65877 & n63901 ;
  assign n85897 = ~n62994 ;
  assign n62998 = n85897 & n62997 ;
  assign n63903 = n62932 | n62997 ;
  assign n85898 = ~n63903 ;
  assign n63904 = n63330 & n85898 ;
  assign n63905 = n62998 | n63904 ;
  assign n63906 = n85736 & n63905 ;
  assign n63907 = n62922 & n85732 ;
  assign n63908 = n63474 & n63907 ;
  assign n63909 = n63906 | n63908 ;
  assign n63910 = n65820 & n63909 ;
  assign n85899 = ~n63908 ;
  assign n63991 = x71 & n85899 ;
  assign n85900 = ~n63906 ;
  assign n63992 = n85900 & n63991 ;
  assign n63993 = n63910 | n63992 ;
  assign n85901 = ~n63329 ;
  assign n63331 = n62992 & n85901 ;
  assign n63911 = n62941 | n62992 ;
  assign n85902 = ~n63911 ;
  assign n63912 = n62988 & n85902 ;
  assign n63913 = n63331 | n63912 ;
  assign n63914 = n85736 & n63913 ;
  assign n63915 = n62931 & n85732 ;
  assign n63916 = n63474 & n63915 ;
  assign n63917 = n63914 | n63916 ;
  assign n63918 = n65791 & n63917 ;
  assign n85903 = ~n62984 ;
  assign n63327 = n85903 & n62987 ;
  assign n63919 = n62949 | n62987 ;
  assign n85904 = ~n63919 ;
  assign n63920 = n63325 & n85904 ;
  assign n63921 = n63327 | n63920 ;
  assign n63922 = n85736 & n63921 ;
  assign n63923 = n62940 & n85732 ;
  assign n63924 = n63474 & n63923 ;
  assign n63925 = n63922 | n63924 ;
  assign n63926 = n65772 & n63925 ;
  assign n85905 = ~n63924 ;
  assign n63980 = x69 & n85905 ;
  assign n85906 = ~n63922 ;
  assign n63981 = n85906 & n63980 ;
  assign n63982 = n63926 | n63981 ;
  assign n85907 = ~n63323 ;
  assign n63324 = n62982 & n85907 ;
  assign n63927 = n62957 | n62982 ;
  assign n85908 = ~n63927 ;
  assign n63928 = n63322 & n85908 ;
  assign n63929 = n63324 | n63928 ;
  assign n63930 = n85736 & n63929 ;
  assign n63931 = n62948 & n85732 ;
  assign n63932 = n63474 & n63931 ;
  assign n63933 = n63930 | n63932 ;
  assign n63934 = n65746 & n63933 ;
  assign n85909 = ~n63321 ;
  assign n63936 = n62977 & n85909 ;
  assign n63935 = n62972 | n62977 ;
  assign n85910 = ~n63935 ;
  assign n63937 = n62973 & n85910 ;
  assign n63938 = n63936 | n63937 ;
  assign n63939 = n85736 & n63938 ;
  assign n63940 = n62956 & n85732 ;
  assign n63941 = n63474 & n63940 ;
  assign n63942 = n63939 | n63941 ;
  assign n63943 = n65721 & n63942 ;
  assign n85911 = ~n63941 ;
  assign n63970 = x67 & n85911 ;
  assign n85912 = ~n63939 ;
  assign n63971 = n85912 & n63970 ;
  assign n63972 = n63943 | n63971 ;
  assign n63944 = n30774 & n62970 ;
  assign n63945 = n85734 & n63944 ;
  assign n85913 = ~n63945 ;
  assign n63946 = n62973 & n85913 ;
  assign n63947 = n85736 & n63946 ;
  assign n63948 = n62960 & n85732 ;
  assign n63949 = n63474 & n63948 ;
  assign n63950 = n63947 | n63949 ;
  assign n63951 = n65686 & n63950 ;
  assign n63316 = n30774 & n85736 ;
  assign n63952 = n85732 & n63474 ;
  assign n85914 = ~n63952 ;
  assign n63953 = x64 & n85914 ;
  assign n85915 = ~n63953 ;
  assign n63954 = x2 & n85915 ;
  assign n63955 = n63316 | n63954 ;
  assign n63956 = x65 & n63955 ;
  assign n63317 = x64 & n85736 ;
  assign n85916 = ~n63317 ;
  assign n63957 = x2 & n85916 ;
  assign n63958 = n30774 & n85914 ;
  assign n63959 = x65 | n63958 ;
  assign n63960 = n63957 | n63959 ;
  assign n85917 = ~n63956 ;
  assign n63961 = n85917 & n63960 ;
  assign n63962 = n31770 | n63961 ;
  assign n63963 = n63316 | n63957 ;
  assign n63964 = n65670 & n63963 ;
  assign n85918 = ~n63964 ;
  assign n63965 = n63962 & n85918 ;
  assign n85919 = ~n63949 ;
  assign n63966 = x66 & n85919 ;
  assign n85920 = ~n63947 ;
  assign n63967 = n85920 & n63966 ;
  assign n63968 = n63951 | n63967 ;
  assign n63969 = n63965 | n63968 ;
  assign n85921 = ~n63951 ;
  assign n63973 = n85921 & n63969 ;
  assign n63974 = n63972 | n63973 ;
  assign n85922 = ~n63943 ;
  assign n63975 = n85922 & n63974 ;
  assign n85923 = ~n63932 ;
  assign n63976 = x68 & n85923 ;
  assign n85924 = ~n63930 ;
  assign n63977 = n85924 & n63976 ;
  assign n63978 = n63934 | n63977 ;
  assign n63979 = n63975 | n63978 ;
  assign n85925 = ~n63934 ;
  assign n63984 = n85925 & n63979 ;
  assign n63985 = n63982 | n63984 ;
  assign n85926 = ~n63926 ;
  assign n63986 = n85926 & n63985 ;
  assign n85927 = ~n63916 ;
  assign n63987 = x70 & n85927 ;
  assign n85928 = ~n63914 ;
  assign n63988 = n85928 & n63987 ;
  assign n63989 = n63918 | n63988 ;
  assign n63990 = n63986 | n63989 ;
  assign n85929 = ~n63918 ;
  assign n63994 = n85929 & n63990 ;
  assign n63995 = n63993 | n63994 ;
  assign n85930 = ~n63910 ;
  assign n63996 = n85930 & n63995 ;
  assign n85931 = ~n63900 ;
  assign n63997 = x72 & n85931 ;
  assign n85932 = ~n63898 ;
  assign n63998 = n85932 & n63997 ;
  assign n63999 = n63902 | n63998 ;
  assign n64000 = n63996 | n63999 ;
  assign n85933 = ~n63902 ;
  assign n64004 = n85933 & n64000 ;
  assign n64005 = n64003 | n64004 ;
  assign n85934 = ~n63894 ;
  assign n64006 = n85934 & n64005 ;
  assign n85935 = ~n63884 ;
  assign n64007 = x74 & n85935 ;
  assign n85936 = ~n63882 ;
  assign n64008 = n85936 & n64007 ;
  assign n64009 = n63886 | n64008 ;
  assign n64010 = n64006 | n64009 ;
  assign n85937 = ~n63886 ;
  assign n64014 = n85937 & n64010 ;
  assign n64015 = n64013 | n64014 ;
  assign n85938 = ~n63878 ;
  assign n64016 = n85938 & n64015 ;
  assign n85939 = ~n63868 ;
  assign n64017 = x76 & n85939 ;
  assign n85940 = ~n63866 ;
  assign n64018 = n85940 & n64017 ;
  assign n64019 = n63870 | n64018 ;
  assign n64021 = n64016 | n64019 ;
  assign n85941 = ~n63870 ;
  assign n64025 = n85941 & n64021 ;
  assign n64026 = n64024 | n64025 ;
  assign n85942 = ~n63862 ;
  assign n64027 = n85942 & n64026 ;
  assign n85943 = ~n63852 ;
  assign n64028 = x78 & n85943 ;
  assign n85944 = ~n63850 ;
  assign n64029 = n85944 & n64028 ;
  assign n64030 = n63854 | n64029 ;
  assign n64031 = n64027 | n64030 ;
  assign n85945 = ~n63854 ;
  assign n64035 = n85945 & n64031 ;
  assign n64036 = n64034 | n64035 ;
  assign n85946 = ~n63846 ;
  assign n64037 = n85946 & n64036 ;
  assign n85947 = ~n63836 ;
  assign n64038 = x80 & n85947 ;
  assign n85948 = ~n63834 ;
  assign n64039 = n85948 & n64038 ;
  assign n64040 = n63838 | n64039 ;
  assign n64042 = n64037 | n64040 ;
  assign n85949 = ~n63838 ;
  assign n64046 = n85949 & n64042 ;
  assign n64047 = n64045 | n64046 ;
  assign n85950 = ~n63830 ;
  assign n64048 = n85950 & n64047 ;
  assign n85951 = ~n63820 ;
  assign n64049 = x82 & n85951 ;
  assign n85952 = ~n63818 ;
  assign n64050 = n85952 & n64049 ;
  assign n64051 = n63822 | n64050 ;
  assign n64052 = n64048 | n64051 ;
  assign n85953 = ~n63822 ;
  assign n64056 = n85953 & n64052 ;
  assign n64057 = n64055 | n64056 ;
  assign n85954 = ~n63814 ;
  assign n64058 = n85954 & n64057 ;
  assign n85955 = ~n63804 ;
  assign n64059 = x84 & n85955 ;
  assign n85956 = ~n63802 ;
  assign n64060 = n85956 & n64059 ;
  assign n64061 = n63806 | n64060 ;
  assign n64062 = n64058 | n64061 ;
  assign n85957 = ~n63806 ;
  assign n64066 = n85957 & n64062 ;
  assign n64067 = n64065 | n64066 ;
  assign n85958 = ~n63798 ;
  assign n64068 = n85958 & n64067 ;
  assign n85959 = ~n63788 ;
  assign n64069 = x86 & n85959 ;
  assign n85960 = ~n63786 ;
  assign n64070 = n85960 & n64069 ;
  assign n64071 = n63790 | n64070 ;
  assign n64072 = n64068 | n64071 ;
  assign n85961 = ~n63790 ;
  assign n64076 = n85961 & n64072 ;
  assign n64077 = n64075 | n64076 ;
  assign n85962 = ~n63782 ;
  assign n64078 = n85962 & n64077 ;
  assign n85963 = ~n63772 ;
  assign n64079 = x88 & n85963 ;
  assign n85964 = ~n63770 ;
  assign n64080 = n85964 & n64079 ;
  assign n64081 = n63774 | n64080 ;
  assign n64082 = n64078 | n64081 ;
  assign n85965 = ~n63774 ;
  assign n64087 = n85965 & n64082 ;
  assign n64088 = n64085 | n64087 ;
  assign n85966 = ~n63766 ;
  assign n64089 = n85966 & n64088 ;
  assign n85967 = ~n63756 ;
  assign n64090 = x90 & n85967 ;
  assign n85968 = ~n63754 ;
  assign n64091 = n85968 & n64090 ;
  assign n64092 = n63758 | n64091 ;
  assign n64093 = n64089 | n64092 ;
  assign n85969 = ~n63758 ;
  assign n64097 = n85969 & n64093 ;
  assign n64098 = n64096 | n64097 ;
  assign n85970 = ~n63750 ;
  assign n64099 = n85970 & n64098 ;
  assign n85971 = ~n63740 ;
  assign n64100 = x92 & n85971 ;
  assign n85972 = ~n63738 ;
  assign n64101 = n85972 & n64100 ;
  assign n64102 = n63742 | n64101 ;
  assign n64103 = n64099 | n64102 ;
  assign n85973 = ~n63742 ;
  assign n64107 = n85973 & n64103 ;
  assign n64108 = n64106 | n64107 ;
  assign n85974 = ~n63734 ;
  assign n64109 = n85974 & n64108 ;
  assign n85975 = ~n63724 ;
  assign n64110 = x94 & n85975 ;
  assign n85976 = ~n63722 ;
  assign n64111 = n85976 & n64110 ;
  assign n64112 = n63726 | n64111 ;
  assign n64113 = n64109 | n64112 ;
  assign n85977 = ~n63726 ;
  assign n64117 = n85977 & n64113 ;
  assign n64118 = n64116 | n64117 ;
  assign n85978 = ~n63718 ;
  assign n64119 = n85978 & n64118 ;
  assign n85979 = ~n63708 ;
  assign n64120 = x96 & n85979 ;
  assign n85980 = ~n63706 ;
  assign n64121 = n85980 & n64120 ;
  assign n64122 = n63710 | n64121 ;
  assign n64123 = n64119 | n64122 ;
  assign n85981 = ~n63710 ;
  assign n64127 = n85981 & n64123 ;
  assign n64128 = n64126 | n64127 ;
  assign n85982 = ~n63702 ;
  assign n64129 = n85982 & n64128 ;
  assign n85983 = ~n63692 ;
  assign n64130 = x98 & n85983 ;
  assign n85984 = ~n63690 ;
  assign n64131 = n85984 & n64130 ;
  assign n64132 = n63694 | n64131 ;
  assign n64133 = n64129 | n64132 ;
  assign n85985 = ~n63694 ;
  assign n64137 = n85985 & n64133 ;
  assign n64138 = n64136 | n64137 ;
  assign n85986 = ~n63686 ;
  assign n64139 = n85986 & n64138 ;
  assign n85987 = ~n63676 ;
  assign n64140 = x100 & n85987 ;
  assign n85988 = ~n63674 ;
  assign n64141 = n85988 & n64140 ;
  assign n64142 = n63678 | n64141 ;
  assign n64143 = n64139 | n64142 ;
  assign n85989 = ~n63678 ;
  assign n64147 = n85989 & n64143 ;
  assign n64148 = n64146 | n64147 ;
  assign n85990 = ~n63670 ;
  assign n64149 = n85990 & n64148 ;
  assign n85991 = ~n63660 ;
  assign n64150 = x102 & n85991 ;
  assign n85992 = ~n63658 ;
  assign n64151 = n85992 & n64150 ;
  assign n64152 = n63662 | n64151 ;
  assign n64153 = n64149 | n64152 ;
  assign n85993 = ~n63662 ;
  assign n64157 = n85993 & n64153 ;
  assign n64158 = n64156 | n64157 ;
  assign n85994 = ~n63654 ;
  assign n64159 = n85994 & n64158 ;
  assign n85995 = ~n63644 ;
  assign n64160 = x104 & n85995 ;
  assign n85996 = ~n63642 ;
  assign n64161 = n85996 & n64160 ;
  assign n64162 = n63646 | n64161 ;
  assign n64163 = n64159 | n64162 ;
  assign n85997 = ~n63646 ;
  assign n64167 = n85997 & n64163 ;
  assign n64168 = n64166 | n64167 ;
  assign n85998 = ~n63638 ;
  assign n64169 = n85998 & n64168 ;
  assign n85999 = ~n63628 ;
  assign n64170 = x106 & n85999 ;
  assign n86000 = ~n63626 ;
  assign n64171 = n86000 & n64170 ;
  assign n64172 = n63630 | n64171 ;
  assign n64174 = n64169 | n64172 ;
  assign n86001 = ~n63630 ;
  assign n64178 = n86001 & n64174 ;
  assign n64179 = n64177 | n64178 ;
  assign n86002 = ~n63622 ;
  assign n64180 = n86002 & n64179 ;
  assign n86003 = ~n63612 ;
  assign n64181 = x108 & n86003 ;
  assign n86004 = ~n63610 ;
  assign n64182 = n86004 & n64181 ;
  assign n64183 = n63614 | n64182 ;
  assign n64184 = n64180 | n64183 ;
  assign n86005 = ~n63614 ;
  assign n64189 = n86005 & n64184 ;
  assign n64190 = n64187 | n64189 ;
  assign n86006 = ~n63606 ;
  assign n64191 = n86006 & n64190 ;
  assign n86007 = ~n63596 ;
  assign n64192 = x110 & n86007 ;
  assign n86008 = ~n63594 ;
  assign n64193 = n86008 & n64192 ;
  assign n64194 = n63598 | n64193 ;
  assign n64196 = n64191 | n64194 ;
  assign n86009 = ~n63598 ;
  assign n64200 = n86009 & n64196 ;
  assign n64201 = n64199 | n64200 ;
  assign n86010 = ~n63590 ;
  assign n64202 = n86010 & n64201 ;
  assign n86011 = ~n63580 ;
  assign n64203 = x112 & n86011 ;
  assign n86012 = ~n63578 ;
  assign n64204 = n86012 & n64203 ;
  assign n64205 = n63582 | n64204 ;
  assign n64206 = n64202 | n64205 ;
  assign n86013 = ~n63582 ;
  assign n64210 = n86013 & n64206 ;
  assign n64211 = n64209 | n64210 ;
  assign n86014 = ~n63574 ;
  assign n64212 = n86014 & n64211 ;
  assign n86015 = ~n63564 ;
  assign n64213 = x114 & n86015 ;
  assign n86016 = ~n63562 ;
  assign n64214 = n86016 & n64213 ;
  assign n64215 = n63566 | n64214 ;
  assign n64217 = n64212 | n64215 ;
  assign n86017 = ~n63566 ;
  assign n64222 = n86017 & n64217 ;
  assign n64223 = n64220 | n64222 ;
  assign n86018 = ~n63558 ;
  assign n64224 = n86018 & n64223 ;
  assign n86019 = ~n63548 ;
  assign n64225 = x116 & n86019 ;
  assign n86020 = ~n63546 ;
  assign n64226 = n86020 & n64225 ;
  assign n64227 = n63550 | n64226 ;
  assign n64228 = n64224 | n64227 ;
  assign n86021 = ~n63550 ;
  assign n64232 = n86021 & n64228 ;
  assign n64233 = n64231 | n64232 ;
  assign n86022 = ~n63542 ;
  assign n64234 = n86022 & n64233 ;
  assign n86023 = ~n63532 ;
  assign n64235 = x118 & n86023 ;
  assign n86024 = ~n63530 ;
  assign n64236 = n86024 & n64235 ;
  assign n64237 = n63534 | n64236 ;
  assign n64238 = n64234 | n64237 ;
  assign n86025 = ~n63534 ;
  assign n64243 = n86025 & n64238 ;
  assign n64244 = n64241 | n64243 ;
  assign n86026 = ~n63526 ;
  assign n64245 = n86026 & n64244 ;
  assign n86027 = ~n63516 ;
  assign n64246 = x120 & n86027 ;
  assign n86028 = ~n63514 ;
  assign n64247 = n86028 & n64246 ;
  assign n64248 = n63518 | n64247 ;
  assign n64249 = n64245 | n64248 ;
  assign n86029 = ~n63518 ;
  assign n64253 = n86029 & n64249 ;
  assign n64254 = n64252 | n64253 ;
  assign n86030 = ~n63510 ;
  assign n64255 = n86030 & n64254 ;
  assign n86031 = ~n63500 ;
  assign n64256 = x122 & n86031 ;
  assign n86032 = ~n63498 ;
  assign n64257 = n86032 & n64256 ;
  assign n64258 = n63502 | n64257 ;
  assign n64259 = n64255 | n64258 ;
  assign n86033 = ~n63502 ;
  assign n64263 = n86033 & n64259 ;
  assign n64264 = n64262 | n64263 ;
  assign n86034 = ~n63494 ;
  assign n64265 = n86034 & n64264 ;
  assign n86035 = ~n63484 ;
  assign n64266 = x124 & n86035 ;
  assign n86036 = ~n63482 ;
  assign n64267 = n86036 & n64266 ;
  assign n64268 = n63486 | n64267 ;
  assign n64270 = n64265 | n64268 ;
  assign n86037 = ~n63486 ;
  assign n64274 = n86037 & n64270 ;
  assign n64275 = n64273 | n64274 ;
  assign n86038 = ~n63478 ;
  assign n64276 = n86038 & n64275 ;
  assign n64277 = n62441 | n63310 ;
  assign n64278 = n63308 | n64277 ;
  assign n86039 = ~n64278 ;
  assign n64279 = n63296 & n86039 ;
  assign n64280 = n63308 | n63310 ;
  assign n86040 = ~n63473 ;
  assign n64281 = n86040 & n64280 ;
  assign n64282 = n64279 | n64281 ;
  assign n64283 = n85736 & n64282 ;
  assign n64284 = n274 & n63307 ;
  assign n64285 = n63474 & n64284 ;
  assign n64286 = n64283 | n64285 ;
  assign n64287 = n75832 & n64286 ;
  assign n86041 = ~n64285 ;
  assign n64288 = x126 & n86041 ;
  assign n86042 = ~n64283 ;
  assign n64289 = n86042 & n64288 ;
  assign n64290 = x127 | n64289 ;
  assign n64291 = n64287 | n64290 ;
  assign n64292 = n64276 | n64291 ;
  assign n64293 = n75526 & n64286 ;
  assign n86043 = ~n64293 ;
  assign n64294 = n64292 & n86043 ;
  assign n64295 = n63478 | n64289 ;
  assign n64296 = n64287 | n64295 ;
  assign n86044 = ~n64296 ;
  assign n64297 = n64275 & n86044 ;
  assign n64298 = n64287 | n64289 ;
  assign n86045 = ~n64276 ;
  assign n64299 = n86045 & n64298 ;
  assign n64300 = n64297 | n64299 ;
  assign n86046 = ~n64294 ;
  assign n64301 = n86046 & n64300 ;
  assign n64302 = n65362 & n64286 ;
  assign n64303 = n64292 & n64302 ;
  assign n64304 = n64301 | n64303 ;
  assign n86047 = ~x127 ;
  assign n64305 = n86047 & n64304 ;
  assign n64307 = n63486 | n64273 ;
  assign n86048 = ~n64307 ;
  assign n64308 = n64270 & n86048 ;
  assign n86049 = ~n64274 ;
  assign n64309 = n64273 & n86049 ;
  assign n64310 = n64308 | n64309 ;
  assign n64311 = n86046 & n64310 ;
  assign n64312 = n63477 & n86043 ;
  assign n64313 = n64292 & n64312 ;
  assign n64314 = n64311 | n64313 ;
  assign n64315 = n75832 & n64314 ;
  assign n64269 = n63494 | n64268 ;
  assign n86050 = ~n64269 ;
  assign n64316 = n64264 & n86050 ;
  assign n86051 = ~n64265 ;
  assign n64317 = n86051 & n64268 ;
  assign n64318 = n64316 | n64317 ;
  assign n64319 = n86046 & n64318 ;
  assign n64320 = n63485 & n86043 ;
  assign n64321 = n64292 & n64320 ;
  assign n64322 = n64319 | n64321 ;
  assign n64323 = n75517 & n64322 ;
  assign n64324 = n63502 | n64262 ;
  assign n86052 = ~n64324 ;
  assign n64325 = n64259 & n86052 ;
  assign n86053 = ~n64263 ;
  assign n64326 = n64262 & n86053 ;
  assign n64327 = n64325 | n64326 ;
  assign n64328 = n86046 & n64327 ;
  assign n64329 = n63493 & n86043 ;
  assign n64330 = n64292 & n64329 ;
  assign n64331 = n64328 | n64330 ;
  assign n64332 = n75210 & n64331 ;
  assign n86054 = ~n64255 ;
  assign n64333 = n86054 & n64258 ;
  assign n64334 = n63510 | n64258 ;
  assign n86055 = ~n64334 ;
  assign n64335 = n64254 & n86055 ;
  assign n64336 = n64333 | n64335 ;
  assign n64337 = n86046 & n64336 ;
  assign n64338 = n63501 & n86043 ;
  assign n64339 = n64292 & n64338 ;
  assign n64340 = n64337 | n64339 ;
  assign n64341 = n74905 & n64340 ;
  assign n64342 = n63518 | n64252 ;
  assign n86056 = ~n64342 ;
  assign n64343 = n64249 & n86056 ;
  assign n86057 = ~n64253 ;
  assign n64344 = n64252 & n86057 ;
  assign n64345 = n64343 | n64344 ;
  assign n64346 = n86046 & n64345 ;
  assign n64347 = n63509 & n86043 ;
  assign n64348 = n64292 & n64347 ;
  assign n64349 = n64346 | n64348 ;
  assign n64350 = n74431 & n64349 ;
  assign n86058 = ~n64245 ;
  assign n64351 = n86058 & n64248 ;
  assign n64352 = n63526 | n64248 ;
  assign n86059 = ~n64352 ;
  assign n64353 = n64244 & n86059 ;
  assign n64354 = n64351 | n64353 ;
  assign n64355 = n86046 & n64354 ;
  assign n64356 = n63517 & n86043 ;
  assign n64357 = n64292 & n64356 ;
  assign n64358 = n64355 | n64357 ;
  assign n64359 = n74029 & n64358 ;
  assign n86060 = ~n64243 ;
  assign n64360 = n64241 & n86060 ;
  assign n64242 = n63534 | n64241 ;
  assign n86061 = ~n64242 ;
  assign n64361 = n64238 & n86061 ;
  assign n64362 = n64360 | n64361 ;
  assign n64363 = n86046 & n64362 ;
  assign n64364 = n63525 & n86043 ;
  assign n64365 = n64292 & n64364 ;
  assign n64366 = n64363 | n64365 ;
  assign n64367 = n74021 & n64366 ;
  assign n86062 = ~n64234 ;
  assign n64368 = n86062 & n64237 ;
  assign n64369 = n63542 | n64237 ;
  assign n86063 = ~n64369 ;
  assign n64370 = n64233 & n86063 ;
  assign n64371 = n64368 | n64370 ;
  assign n64372 = n86046 & n64371 ;
  assign n64373 = n63533 & n86043 ;
  assign n64374 = n64292 & n64373 ;
  assign n64375 = n64372 | n64374 ;
  assign n64376 = n73617 & n64375 ;
  assign n64377 = n63550 | n64231 ;
  assign n86064 = ~n64377 ;
  assign n64378 = n64228 & n86064 ;
  assign n86065 = ~n64232 ;
  assign n64379 = n64231 & n86065 ;
  assign n64380 = n64378 | n64379 ;
  assign n64381 = n86046 & n64380 ;
  assign n64382 = n63541 & n86043 ;
  assign n64383 = n64292 & n64382 ;
  assign n64384 = n64381 | n64383 ;
  assign n64385 = n73188 & n64384 ;
  assign n86066 = ~n64224 ;
  assign n64386 = n86066 & n64227 ;
  assign n64387 = n63558 | n64227 ;
  assign n86067 = ~n64387 ;
  assign n64388 = n64223 & n86067 ;
  assign n64389 = n64386 | n64388 ;
  assign n64390 = n86046 & n64389 ;
  assign n64391 = n63549 & n86043 ;
  assign n64392 = n64292 & n64391 ;
  assign n64393 = n64390 | n64392 ;
  assign n64394 = n73177 & n64393 ;
  assign n86068 = ~n64222 ;
  assign n64395 = n64220 & n86068 ;
  assign n64221 = n63566 | n64220 ;
  assign n86069 = ~n64221 ;
  assign n64396 = n64217 & n86069 ;
  assign n64397 = n64395 | n64396 ;
  assign n64398 = n86046 & n64397 ;
  assign n64399 = n63557 & n86043 ;
  assign n64400 = n64292 & n64399 ;
  assign n64401 = n64398 | n64400 ;
  assign n64402 = n72752 & n64401 ;
  assign n64216 = n63574 | n64215 ;
  assign n86070 = ~n64216 ;
  assign n64403 = n64211 & n86070 ;
  assign n86071 = ~n64212 ;
  assign n64404 = n86071 & n64215 ;
  assign n64405 = n64403 | n64404 ;
  assign n64406 = n86046 & n64405 ;
  assign n64407 = n63565 & n86043 ;
  assign n64408 = n64292 & n64407 ;
  assign n64409 = n64406 | n64408 ;
  assign n64410 = n72393 & n64409 ;
  assign n64411 = n63582 | n64209 ;
  assign n86072 = ~n64411 ;
  assign n64412 = n64206 & n86072 ;
  assign n86073 = ~n64210 ;
  assign n64413 = n64209 & n86073 ;
  assign n64414 = n64412 | n64413 ;
  assign n64415 = n86046 & n64414 ;
  assign n64416 = n63573 & n86043 ;
  assign n64417 = n64292 & n64416 ;
  assign n64418 = n64415 | n64417 ;
  assign n64419 = n72385 & n64418 ;
  assign n86074 = ~n64202 ;
  assign n64420 = n86074 & n64205 ;
  assign n64421 = n63590 | n64205 ;
  assign n86075 = ~n64421 ;
  assign n64422 = n64201 & n86075 ;
  assign n64423 = n64420 | n64422 ;
  assign n64424 = n86046 & n64423 ;
  assign n64425 = n63581 & n86043 ;
  assign n64426 = n64292 & n64425 ;
  assign n64427 = n64424 | n64426 ;
  assign n64428 = n72025 & n64427 ;
  assign n64429 = n63598 | n64199 ;
  assign n86076 = ~n64429 ;
  assign n64430 = n64196 & n86076 ;
  assign n86077 = ~n64200 ;
  assign n64431 = n64199 & n86077 ;
  assign n64432 = n64430 | n64431 ;
  assign n64433 = n86046 & n64432 ;
  assign n64434 = n63589 & n86043 ;
  assign n64435 = n64292 & n64434 ;
  assign n64436 = n64433 | n64435 ;
  assign n64437 = n71645 & n64436 ;
  assign n64195 = n63606 | n64194 ;
  assign n86078 = ~n64195 ;
  assign n64438 = n64190 & n86078 ;
  assign n86079 = ~n64191 ;
  assign n64439 = n86079 & n64194 ;
  assign n64440 = n64438 | n64439 ;
  assign n64441 = n86046 & n64440 ;
  assign n64442 = n63597 & n86043 ;
  assign n64443 = n64292 & n64442 ;
  assign n64444 = n64441 | n64443 ;
  assign n64445 = n71633 & n64444 ;
  assign n86080 = ~n64189 ;
  assign n64446 = n64187 & n86080 ;
  assign n64188 = n63614 | n64187 ;
  assign n86081 = ~n64188 ;
  assign n64447 = n64184 & n86081 ;
  assign n64448 = n64446 | n64447 ;
  assign n64449 = n86046 & n64448 ;
  assign n64450 = n63605 & n86043 ;
  assign n64451 = n64292 & n64450 ;
  assign n64452 = n64449 | n64451 ;
  assign n64453 = n71253 & n64452 ;
  assign n86082 = ~n64180 ;
  assign n64454 = n86082 & n64183 ;
  assign n64455 = n63622 | n64183 ;
  assign n86083 = ~n64455 ;
  assign n64456 = n64179 & n86083 ;
  assign n64457 = n64454 | n64456 ;
  assign n64458 = n86046 & n64457 ;
  assign n64459 = n63613 & n86043 ;
  assign n64460 = n64292 & n64459 ;
  assign n64461 = n64458 | n64460 ;
  assign n64462 = n70935 & n64461 ;
  assign n64463 = n63630 | n64177 ;
  assign n86084 = ~n64463 ;
  assign n64464 = n64174 & n86084 ;
  assign n86085 = ~n64178 ;
  assign n64465 = n64177 & n86085 ;
  assign n64466 = n64464 | n64465 ;
  assign n64467 = n86046 & n64466 ;
  assign n64468 = n63621 & n86043 ;
  assign n64469 = n64292 & n64468 ;
  assign n64470 = n64467 | n64469 ;
  assign n64471 = n70927 & n64470 ;
  assign n64173 = n63638 | n64172 ;
  assign n86086 = ~n64173 ;
  assign n64472 = n64168 & n86086 ;
  assign n86087 = ~n64169 ;
  assign n64473 = n86087 & n64172 ;
  assign n64474 = n64472 | n64473 ;
  assign n64475 = n86046 & n64474 ;
  assign n64476 = n63629 & n86043 ;
  assign n64477 = n64292 & n64476 ;
  assign n64478 = n64475 | n64477 ;
  assign n64479 = n70609 & n64478 ;
  assign n64480 = n63646 | n64166 ;
  assign n86088 = ~n64480 ;
  assign n64481 = n64163 & n86088 ;
  assign n86089 = ~n64167 ;
  assign n64482 = n64166 & n86089 ;
  assign n64483 = n64481 | n64482 ;
  assign n64484 = n86046 & n64483 ;
  assign n64485 = n63637 & n86043 ;
  assign n64486 = n64292 & n64485 ;
  assign n64487 = n64484 | n64486 ;
  assign n64488 = n70276 & n64487 ;
  assign n86090 = ~n64159 ;
  assign n64489 = n86090 & n64162 ;
  assign n64490 = n63654 | n64162 ;
  assign n86091 = ~n64490 ;
  assign n64491 = n64158 & n86091 ;
  assign n64492 = n64489 | n64491 ;
  assign n64493 = n86046 & n64492 ;
  assign n64494 = n63645 & n86043 ;
  assign n64495 = n64292 & n64494 ;
  assign n64496 = n64493 | n64495 ;
  assign n64497 = n70176 & n64496 ;
  assign n64498 = n63662 | n64156 ;
  assign n86092 = ~n64498 ;
  assign n64499 = n64153 & n86092 ;
  assign n86093 = ~n64157 ;
  assign n64500 = n64156 & n86093 ;
  assign n64501 = n64499 | n64500 ;
  assign n64502 = n86046 & n64501 ;
  assign n64503 = n63653 & n86043 ;
  assign n64504 = n64292 & n64503 ;
  assign n64505 = n64502 | n64504 ;
  assign n64506 = n69857 & n64505 ;
  assign n86094 = ~n64149 ;
  assign n64507 = n86094 & n64152 ;
  assign n64508 = n63670 | n64152 ;
  assign n86095 = ~n64508 ;
  assign n64509 = n64148 & n86095 ;
  assign n64510 = n64507 | n64509 ;
  assign n64511 = n86046 & n64510 ;
  assign n64512 = n63661 & n86043 ;
  assign n64513 = n64292 & n64512 ;
  assign n64514 = n64511 | n64513 ;
  assign n64515 = n69656 & n64514 ;
  assign n64516 = n63678 | n64146 ;
  assign n86096 = ~n64516 ;
  assign n64517 = n64143 & n86096 ;
  assign n86097 = ~n64147 ;
  assign n64518 = n64146 & n86097 ;
  assign n64519 = n64517 | n64518 ;
  assign n64520 = n86046 & n64519 ;
  assign n64521 = n63669 & n86043 ;
  assign n64522 = n64292 & n64521 ;
  assign n64523 = n64520 | n64522 ;
  assign n64524 = n69528 & n64523 ;
  assign n86098 = ~n64139 ;
  assign n64525 = n86098 & n64142 ;
  assign n64526 = n63686 | n64142 ;
  assign n86099 = ~n64526 ;
  assign n64527 = n64138 & n86099 ;
  assign n64528 = n64525 | n64527 ;
  assign n64529 = n86046 & n64528 ;
  assign n64530 = n63677 & n86043 ;
  assign n64531 = n64292 & n64530 ;
  assign n64532 = n64529 | n64531 ;
  assign n64533 = n69261 & n64532 ;
  assign n64534 = n63694 | n64136 ;
  assign n86100 = ~n64534 ;
  assign n64535 = n64133 & n86100 ;
  assign n86101 = ~n64137 ;
  assign n64536 = n64136 & n86101 ;
  assign n64537 = n64535 | n64536 ;
  assign n64538 = n86046 & n64537 ;
  assign n64539 = n63685 & n86043 ;
  assign n64540 = n64292 & n64539 ;
  assign n64541 = n64538 | n64540 ;
  assign n64542 = n69075 & n64541 ;
  assign n86102 = ~n64129 ;
  assign n64543 = n86102 & n64132 ;
  assign n64544 = n63702 | n64132 ;
  assign n86103 = ~n64544 ;
  assign n64545 = n64128 & n86103 ;
  assign n64546 = n64543 | n64545 ;
  assign n64547 = n86046 & n64546 ;
  assign n64548 = n63693 & n86043 ;
  assign n64549 = n64292 & n64548 ;
  assign n64550 = n64547 | n64549 ;
  assign n64551 = n68993 & n64550 ;
  assign n64552 = n63710 | n64126 ;
  assign n86104 = ~n64552 ;
  assign n64553 = n64123 & n86104 ;
  assign n86105 = ~n64127 ;
  assign n64554 = n64126 & n86105 ;
  assign n64555 = n64553 | n64554 ;
  assign n64556 = n86046 & n64555 ;
  assign n64557 = n63701 & n86043 ;
  assign n64558 = n64292 & n64557 ;
  assign n64559 = n64556 | n64558 ;
  assign n64560 = n68716 & n64559 ;
  assign n86106 = ~n64119 ;
  assign n64561 = n86106 & n64122 ;
  assign n64562 = n63718 | n64122 ;
  assign n86107 = ~n64562 ;
  assign n64563 = n64118 & n86107 ;
  assign n64564 = n64561 | n64563 ;
  assign n64565 = n86046 & n64564 ;
  assign n64566 = n63709 & n86043 ;
  assign n64567 = n64292 & n64566 ;
  assign n64568 = n64565 | n64567 ;
  assign n64569 = n68545 & n64568 ;
  assign n64570 = n63726 | n64116 ;
  assign n86108 = ~n64570 ;
  assign n64571 = n64113 & n86108 ;
  assign n86109 = ~n64117 ;
  assign n64572 = n64116 & n86109 ;
  assign n64573 = n64571 | n64572 ;
  assign n64574 = n86046 & n64573 ;
  assign n64575 = n63717 & n86043 ;
  assign n64576 = n64292 & n64575 ;
  assign n64577 = n64574 | n64576 ;
  assign n64578 = n68438 & n64577 ;
  assign n86110 = ~n64109 ;
  assign n64579 = n86110 & n64112 ;
  assign n64580 = n63734 | n64112 ;
  assign n86111 = ~n64580 ;
  assign n64581 = n64108 & n86111 ;
  assign n64582 = n64579 | n64581 ;
  assign n64583 = n86046 & n64582 ;
  assign n64584 = n63725 & n86043 ;
  assign n64585 = n64292 & n64584 ;
  assign n64586 = n64583 | n64585 ;
  assign n64587 = n68214 & n64586 ;
  assign n64588 = n63742 | n64106 ;
  assign n86112 = ~n64588 ;
  assign n64589 = n64103 & n86112 ;
  assign n86113 = ~n64107 ;
  assign n64590 = n64106 & n86113 ;
  assign n64591 = n64589 | n64590 ;
  assign n64592 = n86046 & n64591 ;
  assign n64593 = n63733 & n86043 ;
  assign n64594 = n64292 & n64593 ;
  assign n64595 = n64592 | n64594 ;
  assign n64596 = n68058 & n64595 ;
  assign n86114 = ~n64099 ;
  assign n64597 = n86114 & n64102 ;
  assign n64598 = n63750 | n64102 ;
  assign n86115 = ~n64598 ;
  assign n64599 = n64098 & n86115 ;
  assign n64600 = n64597 | n64599 ;
  assign n64601 = n86046 & n64600 ;
  assign n64602 = n63741 & n86043 ;
  assign n64603 = n64292 & n64602 ;
  assign n64604 = n64601 | n64603 ;
  assign n64605 = n67986 & n64604 ;
  assign n64606 = n63758 | n64096 ;
  assign n86116 = ~n64606 ;
  assign n64607 = n64093 & n86116 ;
  assign n86117 = ~n64097 ;
  assign n64608 = n64096 & n86117 ;
  assign n64609 = n64607 | n64608 ;
  assign n64610 = n86046 & n64609 ;
  assign n64611 = n63749 & n86043 ;
  assign n64612 = n64292 & n64611 ;
  assign n64613 = n64610 | n64612 ;
  assign n64614 = n67763 & n64613 ;
  assign n86118 = ~n64089 ;
  assign n64615 = n86118 & n64092 ;
  assign n64616 = n63766 | n64092 ;
  assign n86119 = ~n64616 ;
  assign n64617 = n64088 & n86119 ;
  assign n64618 = n64615 | n64617 ;
  assign n64619 = n86046 & n64618 ;
  assign n64620 = n63757 & n86043 ;
  assign n64621 = n64292 & n64620 ;
  assign n64622 = n64619 | n64621 ;
  assign n64623 = n67622 & n64622 ;
  assign n86120 = ~n64087 ;
  assign n64624 = n64085 & n86120 ;
  assign n64086 = n63774 | n64085 ;
  assign n86121 = ~n64086 ;
  assign n64625 = n64082 & n86121 ;
  assign n64626 = n64624 | n64625 ;
  assign n64627 = n86046 & n64626 ;
  assign n64628 = n63765 & n86043 ;
  assign n64629 = n64292 & n64628 ;
  assign n64630 = n64627 | n64629 ;
  assign n64631 = n67531 & n64630 ;
  assign n86122 = ~n64078 ;
  assign n64632 = n86122 & n64081 ;
  assign n64633 = n63782 | n64081 ;
  assign n86123 = ~n64633 ;
  assign n64634 = n64077 & n86123 ;
  assign n64635 = n64632 | n64634 ;
  assign n64636 = n86046 & n64635 ;
  assign n64637 = n63773 & n86043 ;
  assign n64638 = n64292 & n64637 ;
  assign n64639 = n64636 | n64638 ;
  assign n64640 = n67348 & n64639 ;
  assign n64641 = n63790 | n64075 ;
  assign n86124 = ~n64641 ;
  assign n64642 = n64072 & n86124 ;
  assign n86125 = ~n64076 ;
  assign n64643 = n64075 & n86125 ;
  assign n64644 = n64642 | n64643 ;
  assign n64645 = n86046 & n64644 ;
  assign n64646 = n63781 & n86043 ;
  assign n64647 = n64292 & n64646 ;
  assign n64648 = n64645 | n64647 ;
  assign n64649 = n67222 & n64648 ;
  assign n86126 = ~n64068 ;
  assign n64650 = n86126 & n64071 ;
  assign n64651 = n63798 | n64071 ;
  assign n86127 = ~n64651 ;
  assign n64652 = n64067 & n86127 ;
  assign n64653 = n64650 | n64652 ;
  assign n64654 = n86046 & n64653 ;
  assign n64655 = n63789 & n86043 ;
  assign n64656 = n64292 & n64655 ;
  assign n64657 = n64654 | n64656 ;
  assign n64658 = n67164 & n64657 ;
  assign n64659 = n63806 | n64065 ;
  assign n86128 = ~n64659 ;
  assign n64660 = n64062 & n86128 ;
  assign n86129 = ~n64066 ;
  assign n64661 = n64065 & n86129 ;
  assign n64662 = n64660 | n64661 ;
  assign n64663 = n86046 & n64662 ;
  assign n64664 = n63797 & n86043 ;
  assign n64665 = n64292 & n64664 ;
  assign n64666 = n64663 | n64665 ;
  assign n64667 = n66979 & n64666 ;
  assign n86130 = ~n64058 ;
  assign n64668 = n86130 & n64061 ;
  assign n64669 = n63814 | n64061 ;
  assign n86131 = ~n64669 ;
  assign n64670 = n64057 & n86131 ;
  assign n64671 = n64668 | n64670 ;
  assign n64672 = n86046 & n64671 ;
  assign n64673 = n63805 & n86043 ;
  assign n64674 = n64292 & n64673 ;
  assign n64675 = n64672 | n64674 ;
  assign n64676 = n66868 & n64675 ;
  assign n64677 = n63822 | n64055 ;
  assign n86132 = ~n64677 ;
  assign n64678 = n64052 & n86132 ;
  assign n86133 = ~n64056 ;
  assign n64679 = n64055 & n86133 ;
  assign n64680 = n64678 | n64679 ;
  assign n64681 = n86046 & n64680 ;
  assign n64682 = n63813 & n86043 ;
  assign n64683 = n64292 & n64682 ;
  assign n64684 = n64681 | n64683 ;
  assign n64685 = n66797 & n64684 ;
  assign n86134 = ~n64048 ;
  assign n64686 = n86134 & n64051 ;
  assign n64687 = n63830 | n64051 ;
  assign n86135 = ~n64687 ;
  assign n64688 = n64047 & n86135 ;
  assign n64689 = n64686 | n64688 ;
  assign n64690 = n86046 & n64689 ;
  assign n64691 = n63821 & n86043 ;
  assign n64692 = n64292 & n64691 ;
  assign n64693 = n64690 | n64692 ;
  assign n64694 = n66654 & n64693 ;
  assign n64695 = n63838 | n64045 ;
  assign n86136 = ~n64695 ;
  assign n64696 = n64042 & n86136 ;
  assign n86137 = ~n64046 ;
  assign n64697 = n64045 & n86137 ;
  assign n64698 = n64696 | n64697 ;
  assign n64699 = n86046 & n64698 ;
  assign n64700 = n63829 & n86043 ;
  assign n64701 = n64292 & n64700 ;
  assign n64702 = n64699 | n64701 ;
  assign n64703 = n66560 & n64702 ;
  assign n64041 = n63846 | n64040 ;
  assign n86138 = ~n64041 ;
  assign n64704 = n64036 & n86138 ;
  assign n86139 = ~n64037 ;
  assign n64705 = n86139 & n64040 ;
  assign n64706 = n64704 | n64705 ;
  assign n64707 = n86046 & n64706 ;
  assign n64708 = n63837 & n86043 ;
  assign n64709 = n64292 & n64708 ;
  assign n64710 = n64707 | n64709 ;
  assign n64711 = n66505 & n64710 ;
  assign n86140 = ~n64035 ;
  assign n64712 = n64034 & n86140 ;
  assign n64713 = n63854 | n64034 ;
  assign n86141 = ~n64713 ;
  assign n64714 = n64031 & n86141 ;
  assign n64715 = n64712 | n64714 ;
  assign n64716 = n86046 & n64715 ;
  assign n64717 = n63845 & n86043 ;
  assign n64718 = n64292 & n64717 ;
  assign n64719 = n64716 | n64718 ;
  assign n64720 = n66379 & n64719 ;
  assign n86142 = ~n64027 ;
  assign n64721 = n86142 & n64030 ;
  assign n64722 = n63862 | n64030 ;
  assign n86143 = ~n64722 ;
  assign n64723 = n64026 & n86143 ;
  assign n64724 = n64721 | n64723 ;
  assign n64725 = n86046 & n64724 ;
  assign n64726 = n63853 & n86043 ;
  assign n64727 = n64292 & n64726 ;
  assign n64728 = n64725 | n64727 ;
  assign n64729 = n66299 & n64728 ;
  assign n64730 = n63870 | n64024 ;
  assign n86144 = ~n64730 ;
  assign n64731 = n64021 & n86144 ;
  assign n86145 = ~n64025 ;
  assign n64732 = n64024 & n86145 ;
  assign n64733 = n64731 | n64732 ;
  assign n64734 = n86046 & n64733 ;
  assign n64735 = n63861 & n86043 ;
  assign n64736 = n64292 & n64735 ;
  assign n64737 = n64734 | n64736 ;
  assign n64738 = n66244 & n64737 ;
  assign n64020 = n63878 | n64019 ;
  assign n86146 = ~n64020 ;
  assign n64739 = n64015 & n86146 ;
  assign n86147 = ~n64016 ;
  assign n64740 = n86147 & n64019 ;
  assign n64741 = n64739 | n64740 ;
  assign n64742 = n86046 & n64741 ;
  assign n64743 = n63869 & n86043 ;
  assign n64744 = n64292 & n64743 ;
  assign n64745 = n64742 | n64744 ;
  assign n64746 = n66145 & n64745 ;
  assign n64747 = n63886 | n64013 ;
  assign n86148 = ~n64747 ;
  assign n64748 = n64010 & n86148 ;
  assign n86149 = ~n64014 ;
  assign n64749 = n64013 & n86149 ;
  assign n64750 = n64748 | n64749 ;
  assign n64751 = n86046 & n64750 ;
  assign n64752 = n63877 & n86043 ;
  assign n64753 = n64292 & n64752 ;
  assign n64754 = n64751 | n64753 ;
  assign n64755 = n66081 & n64754 ;
  assign n86150 = ~n64006 ;
  assign n64756 = n86150 & n64009 ;
  assign n64757 = n63894 | n64009 ;
  assign n86151 = ~n64757 ;
  assign n64758 = n64005 & n86151 ;
  assign n64759 = n64756 | n64758 ;
  assign n64760 = n86046 & n64759 ;
  assign n64761 = n63885 & n86043 ;
  assign n64762 = n64292 & n64761 ;
  assign n64763 = n64760 | n64762 ;
  assign n64764 = n66043 & n64763 ;
  assign n64765 = n63902 | n64003 ;
  assign n86152 = ~n64765 ;
  assign n64766 = n64000 & n86152 ;
  assign n86153 = ~n64004 ;
  assign n64767 = n64003 & n86153 ;
  assign n64768 = n64766 | n64767 ;
  assign n64769 = n86046 & n64768 ;
  assign n64770 = n63893 & n86043 ;
  assign n64771 = n64292 & n64770 ;
  assign n64772 = n64769 | n64771 ;
  assign n64773 = n65960 & n64772 ;
  assign n86154 = ~n63996 ;
  assign n64774 = n86154 & n63999 ;
  assign n64775 = n63910 | n63999 ;
  assign n86155 = ~n64775 ;
  assign n64776 = n63995 & n86155 ;
  assign n64777 = n64774 | n64776 ;
  assign n64778 = n86046 & n64777 ;
  assign n64779 = n63901 & n86043 ;
  assign n64780 = n64292 & n64779 ;
  assign n64781 = n64778 | n64780 ;
  assign n64782 = n65909 & n64781 ;
  assign n64783 = n63918 | n63993 ;
  assign n86156 = ~n64783 ;
  assign n64784 = n63990 & n86156 ;
  assign n86157 = ~n63994 ;
  assign n64785 = n63993 & n86157 ;
  assign n64786 = n64784 | n64785 ;
  assign n64787 = n86046 & n64786 ;
  assign n64788 = n63909 & n86043 ;
  assign n64789 = n64292 & n64788 ;
  assign n64790 = n64787 | n64789 ;
  assign n64791 = n65877 & n64790 ;
  assign n86158 = ~n63986 ;
  assign n64792 = n86158 & n63989 ;
  assign n64793 = n63926 | n63989 ;
  assign n86159 = ~n64793 ;
  assign n64794 = n63985 & n86159 ;
  assign n64795 = n64792 | n64794 ;
  assign n64796 = n86046 & n64795 ;
  assign n64797 = n63917 & n86043 ;
  assign n64798 = n64292 & n64797 ;
  assign n64799 = n64796 | n64798 ;
  assign n64800 = n65820 & n64799 ;
  assign n86160 = ~n63984 ;
  assign n64801 = n63982 & n86160 ;
  assign n63983 = n63934 | n63982 ;
  assign n86161 = ~n63983 ;
  assign n64802 = n63979 & n86161 ;
  assign n64803 = n64801 | n64802 ;
  assign n64804 = n86046 & n64803 ;
  assign n64805 = n63925 & n86043 ;
  assign n64806 = n64292 & n64805 ;
  assign n64807 = n64804 | n64806 ;
  assign n64808 = n65791 & n64807 ;
  assign n64809 = n63943 | n63978 ;
  assign n86162 = ~n64809 ;
  assign n64810 = n63974 & n86162 ;
  assign n86163 = ~n63975 ;
  assign n64811 = n86163 & n63978 ;
  assign n64812 = n64810 | n64811 ;
  assign n64813 = n86046 & n64812 ;
  assign n64814 = n63933 & n86043 ;
  assign n64815 = n64292 & n64814 ;
  assign n64816 = n64813 | n64815 ;
  assign n64817 = n65772 & n64816 ;
  assign n86164 = ~n63973 ;
  assign n64819 = n63972 & n86164 ;
  assign n64818 = n63951 | n63972 ;
  assign n86165 = ~n64818 ;
  assign n64820 = n63969 & n86165 ;
  assign n64821 = n64819 | n64820 ;
  assign n64822 = n86046 & n64821 ;
  assign n64823 = n63942 & n86043 ;
  assign n64824 = n64292 & n64823 ;
  assign n64825 = n64822 | n64824 ;
  assign n64826 = n65746 & n64825 ;
  assign n64827 = n63964 | n63968 ;
  assign n86166 = ~n64827 ;
  assign n64828 = n63962 & n86166 ;
  assign n86167 = ~n63965 ;
  assign n64829 = n86167 & n63968 ;
  assign n64830 = n64828 | n64829 ;
  assign n64831 = n86046 & n64830 ;
  assign n64832 = n63950 & n86043 ;
  assign n64833 = n64292 & n64832 ;
  assign n64834 = n64831 | n64833 ;
  assign n64835 = n65721 & n64834 ;
  assign n64836 = n31770 & n63960 ;
  assign n64837 = n85917 & n64836 ;
  assign n86168 = ~n64837 ;
  assign n64838 = n63962 & n86168 ;
  assign n64839 = n86046 & n64838 ;
  assign n64840 = n63963 & n86043 ;
  assign n64841 = n64292 & n64840 ;
  assign n64842 = n64839 | n64841 ;
  assign n64843 = n65686 & n64842 ;
  assign n64306 = n31770 & n86046 ;
  assign n64844 = x64 & n86046 ;
  assign n86169 = ~n64844 ;
  assign n64845 = x1 & n86169 ;
  assign n64846 = n64306 | n64845 ;
  assign n64848 = x65 & n64846 ;
  assign n64847 = x65 | n64306 ;
  assign n64849 = n64845 | n64847 ;
  assign n86170 = ~n64848 ;
  assign n64850 = n86170 & n64849 ;
  assign n64851 = n32480 | n64850 ;
  assign n64852 = n65670 & n64846 ;
  assign n86171 = ~n64852 ;
  assign n64853 = n64851 & n86171 ;
  assign n86172 = ~n64841 ;
  assign n64854 = x66 & n86172 ;
  assign n86173 = ~n64839 ;
  assign n64855 = n86173 & n64854 ;
  assign n64856 = n64843 | n64855 ;
  assign n64857 = n64853 | n64856 ;
  assign n86174 = ~n64843 ;
  assign n64858 = n86174 & n64857 ;
  assign n86175 = ~n64833 ;
  assign n64859 = x67 & n86175 ;
  assign n86176 = ~n64831 ;
  assign n64860 = n86176 & n64859 ;
  assign n64861 = n64835 | n64860 ;
  assign n64863 = n64858 | n64861 ;
  assign n86177 = ~n64835 ;
  assign n64864 = n86177 & n64863 ;
  assign n86178 = ~n64824 ;
  assign n64865 = x68 & n86178 ;
  assign n86179 = ~n64822 ;
  assign n64866 = n86179 & n64865 ;
  assign n64867 = n64826 | n64866 ;
  assign n64868 = n64864 | n64867 ;
  assign n86180 = ~n64826 ;
  assign n64869 = n86180 & n64868 ;
  assign n86181 = ~n64815 ;
  assign n64870 = x69 & n86181 ;
  assign n86182 = ~n64813 ;
  assign n64871 = n86182 & n64870 ;
  assign n64872 = n64817 | n64871 ;
  assign n64875 = n64869 | n64872 ;
  assign n86183 = ~n64817 ;
  assign n64876 = n86183 & n64875 ;
  assign n86184 = ~n64806 ;
  assign n64877 = x70 & n86184 ;
  assign n86185 = ~n64804 ;
  assign n64878 = n86185 & n64877 ;
  assign n64879 = n64808 | n64878 ;
  assign n64880 = n64876 | n64879 ;
  assign n86186 = ~n64808 ;
  assign n64881 = n86186 & n64880 ;
  assign n86187 = ~n64798 ;
  assign n64882 = x71 & n86187 ;
  assign n86188 = ~n64796 ;
  assign n64883 = n86188 & n64882 ;
  assign n64884 = n64800 | n64883 ;
  assign n64887 = n64881 | n64884 ;
  assign n86189 = ~n64800 ;
  assign n64888 = n86189 & n64887 ;
  assign n86190 = ~n64789 ;
  assign n64889 = x72 & n86190 ;
  assign n86191 = ~n64787 ;
  assign n64890 = n86191 & n64889 ;
  assign n64891 = n64791 | n64890 ;
  assign n64892 = n64888 | n64891 ;
  assign n86192 = ~n64791 ;
  assign n64893 = n86192 & n64892 ;
  assign n86193 = ~n64780 ;
  assign n64894 = x73 & n86193 ;
  assign n86194 = ~n64778 ;
  assign n64895 = n86194 & n64894 ;
  assign n64896 = n64782 | n64895 ;
  assign n64898 = n64893 | n64896 ;
  assign n86195 = ~n64782 ;
  assign n64899 = n86195 & n64898 ;
  assign n86196 = ~n64771 ;
  assign n64900 = x74 & n86196 ;
  assign n86197 = ~n64769 ;
  assign n64901 = n86197 & n64900 ;
  assign n64902 = n64773 | n64901 ;
  assign n64903 = n64899 | n64902 ;
  assign n86198 = ~n64773 ;
  assign n64904 = n86198 & n64903 ;
  assign n86199 = ~n64762 ;
  assign n64905 = x75 & n86199 ;
  assign n86200 = ~n64760 ;
  assign n64906 = n86200 & n64905 ;
  assign n64907 = n64764 | n64906 ;
  assign n64909 = n64904 | n64907 ;
  assign n86201 = ~n64764 ;
  assign n64910 = n86201 & n64909 ;
  assign n86202 = ~n64753 ;
  assign n64911 = x76 & n86202 ;
  assign n86203 = ~n64751 ;
  assign n64912 = n86203 & n64911 ;
  assign n64913 = n64755 | n64912 ;
  assign n64914 = n64910 | n64913 ;
  assign n86204 = ~n64755 ;
  assign n64915 = n86204 & n64914 ;
  assign n86205 = ~n64744 ;
  assign n64916 = x77 & n86205 ;
  assign n86206 = ~n64742 ;
  assign n64917 = n86206 & n64916 ;
  assign n64918 = n64746 | n64917 ;
  assign n64920 = n64915 | n64918 ;
  assign n86207 = ~n64746 ;
  assign n64921 = n86207 & n64920 ;
  assign n86208 = ~n64736 ;
  assign n64922 = x78 & n86208 ;
  assign n86209 = ~n64734 ;
  assign n64923 = n86209 & n64922 ;
  assign n64924 = n64738 | n64923 ;
  assign n64925 = n64921 | n64924 ;
  assign n86210 = ~n64738 ;
  assign n64926 = n86210 & n64925 ;
  assign n86211 = ~n64727 ;
  assign n64927 = x79 & n86211 ;
  assign n86212 = ~n64725 ;
  assign n64928 = n86212 & n64927 ;
  assign n64929 = n64729 | n64928 ;
  assign n64931 = n64926 | n64929 ;
  assign n86213 = ~n64729 ;
  assign n64932 = n86213 & n64931 ;
  assign n86214 = ~n64718 ;
  assign n64933 = x80 & n86214 ;
  assign n86215 = ~n64716 ;
  assign n64934 = n86215 & n64933 ;
  assign n64935 = n64720 | n64934 ;
  assign n64936 = n64932 | n64935 ;
  assign n86216 = ~n64720 ;
  assign n64937 = n86216 & n64936 ;
  assign n86217 = ~n64709 ;
  assign n64938 = x81 & n86217 ;
  assign n86218 = ~n64707 ;
  assign n64939 = n86218 & n64938 ;
  assign n64940 = n64711 | n64939 ;
  assign n64942 = n64937 | n64940 ;
  assign n86219 = ~n64711 ;
  assign n64943 = n86219 & n64942 ;
  assign n86220 = ~n64701 ;
  assign n64944 = x82 & n86220 ;
  assign n86221 = ~n64699 ;
  assign n64945 = n86221 & n64944 ;
  assign n64946 = n64703 | n64945 ;
  assign n64947 = n64943 | n64946 ;
  assign n86222 = ~n64703 ;
  assign n64948 = n86222 & n64947 ;
  assign n86223 = ~n64692 ;
  assign n64949 = x83 & n86223 ;
  assign n86224 = ~n64690 ;
  assign n64950 = n86224 & n64949 ;
  assign n64951 = n64694 | n64950 ;
  assign n64953 = n64948 | n64951 ;
  assign n86225 = ~n64694 ;
  assign n64954 = n86225 & n64953 ;
  assign n86226 = ~n64683 ;
  assign n64955 = x84 & n86226 ;
  assign n86227 = ~n64681 ;
  assign n64956 = n86227 & n64955 ;
  assign n64957 = n64685 | n64956 ;
  assign n64958 = n64954 | n64957 ;
  assign n86228 = ~n64685 ;
  assign n64959 = n86228 & n64958 ;
  assign n86229 = ~n64674 ;
  assign n64960 = x85 & n86229 ;
  assign n86230 = ~n64672 ;
  assign n64961 = n86230 & n64960 ;
  assign n64962 = n64676 | n64961 ;
  assign n64964 = n64959 | n64962 ;
  assign n86231 = ~n64676 ;
  assign n64965 = n86231 & n64964 ;
  assign n86232 = ~n64665 ;
  assign n64966 = x86 & n86232 ;
  assign n86233 = ~n64663 ;
  assign n64967 = n86233 & n64966 ;
  assign n64968 = n64667 | n64967 ;
  assign n64969 = n64965 | n64968 ;
  assign n86234 = ~n64667 ;
  assign n64970 = n86234 & n64969 ;
  assign n86235 = ~n64656 ;
  assign n64971 = x87 & n86235 ;
  assign n86236 = ~n64654 ;
  assign n64972 = n86236 & n64971 ;
  assign n64973 = n64658 | n64972 ;
  assign n64975 = n64970 | n64973 ;
  assign n86237 = ~n64658 ;
  assign n64976 = n86237 & n64975 ;
  assign n86238 = ~n64647 ;
  assign n64977 = x88 & n86238 ;
  assign n86239 = ~n64645 ;
  assign n64978 = n86239 & n64977 ;
  assign n64979 = n64649 | n64978 ;
  assign n64980 = n64976 | n64979 ;
  assign n86240 = ~n64649 ;
  assign n64981 = n86240 & n64980 ;
  assign n86241 = ~n64638 ;
  assign n64982 = x89 & n86241 ;
  assign n86242 = ~n64636 ;
  assign n64983 = n86242 & n64982 ;
  assign n64984 = n64640 | n64983 ;
  assign n64986 = n64981 | n64984 ;
  assign n86243 = ~n64640 ;
  assign n64987 = n86243 & n64986 ;
  assign n86244 = ~n64629 ;
  assign n64988 = x90 & n86244 ;
  assign n86245 = ~n64627 ;
  assign n64989 = n86245 & n64988 ;
  assign n64990 = n64631 | n64989 ;
  assign n64991 = n64987 | n64990 ;
  assign n86246 = ~n64631 ;
  assign n64992 = n86246 & n64991 ;
  assign n86247 = ~n64621 ;
  assign n64993 = x91 & n86247 ;
  assign n86248 = ~n64619 ;
  assign n64994 = n86248 & n64993 ;
  assign n64995 = n64623 | n64994 ;
  assign n64997 = n64992 | n64995 ;
  assign n86249 = ~n64623 ;
  assign n64998 = n86249 & n64997 ;
  assign n86250 = ~n64612 ;
  assign n64999 = x92 & n86250 ;
  assign n86251 = ~n64610 ;
  assign n65000 = n86251 & n64999 ;
  assign n65001 = n64614 | n65000 ;
  assign n65002 = n64998 | n65001 ;
  assign n86252 = ~n64614 ;
  assign n65003 = n86252 & n65002 ;
  assign n86253 = ~n64603 ;
  assign n65004 = x93 & n86253 ;
  assign n86254 = ~n64601 ;
  assign n65005 = n86254 & n65004 ;
  assign n65006 = n64605 | n65005 ;
  assign n65008 = n65003 | n65006 ;
  assign n86255 = ~n64605 ;
  assign n65009 = n86255 & n65008 ;
  assign n86256 = ~n64594 ;
  assign n65010 = x94 & n86256 ;
  assign n86257 = ~n64592 ;
  assign n65011 = n86257 & n65010 ;
  assign n65012 = n64596 | n65011 ;
  assign n65013 = n65009 | n65012 ;
  assign n86258 = ~n64596 ;
  assign n65014 = n86258 & n65013 ;
  assign n86259 = ~n64585 ;
  assign n65015 = x95 & n86259 ;
  assign n86260 = ~n64583 ;
  assign n65016 = n86260 & n65015 ;
  assign n65017 = n64587 | n65016 ;
  assign n65019 = n65014 | n65017 ;
  assign n86261 = ~n64587 ;
  assign n65020 = n86261 & n65019 ;
  assign n86262 = ~n64576 ;
  assign n65021 = x96 & n86262 ;
  assign n86263 = ~n64574 ;
  assign n65022 = n86263 & n65021 ;
  assign n65023 = n64578 | n65022 ;
  assign n65024 = n65020 | n65023 ;
  assign n86264 = ~n64578 ;
  assign n65025 = n86264 & n65024 ;
  assign n86265 = ~n64567 ;
  assign n65026 = x97 & n86265 ;
  assign n86266 = ~n64565 ;
  assign n65027 = n86266 & n65026 ;
  assign n65028 = n64569 | n65027 ;
  assign n65030 = n65025 | n65028 ;
  assign n86267 = ~n64569 ;
  assign n65031 = n86267 & n65030 ;
  assign n86268 = ~n64558 ;
  assign n65032 = x98 & n86268 ;
  assign n86269 = ~n64556 ;
  assign n65033 = n86269 & n65032 ;
  assign n65034 = n64560 | n65033 ;
  assign n65035 = n65031 | n65034 ;
  assign n86270 = ~n64560 ;
  assign n65036 = n86270 & n65035 ;
  assign n86271 = ~n64549 ;
  assign n65037 = x99 & n86271 ;
  assign n86272 = ~n64547 ;
  assign n65038 = n86272 & n65037 ;
  assign n65039 = n64551 | n65038 ;
  assign n65041 = n65036 | n65039 ;
  assign n86273 = ~n64551 ;
  assign n65042 = n86273 & n65041 ;
  assign n86274 = ~n64540 ;
  assign n65043 = x100 & n86274 ;
  assign n86275 = ~n64538 ;
  assign n65044 = n86275 & n65043 ;
  assign n65045 = n64542 | n65044 ;
  assign n65046 = n65042 | n65045 ;
  assign n86276 = ~n64542 ;
  assign n65047 = n86276 & n65046 ;
  assign n86277 = ~n64531 ;
  assign n65048 = x101 & n86277 ;
  assign n86278 = ~n64529 ;
  assign n65049 = n86278 & n65048 ;
  assign n65050 = n64533 | n65049 ;
  assign n65052 = n65047 | n65050 ;
  assign n86279 = ~n64533 ;
  assign n65053 = n86279 & n65052 ;
  assign n86280 = ~n64522 ;
  assign n65054 = x102 & n86280 ;
  assign n86281 = ~n64520 ;
  assign n65055 = n86281 & n65054 ;
  assign n65056 = n64524 | n65055 ;
  assign n65057 = n65053 | n65056 ;
  assign n86282 = ~n64524 ;
  assign n65058 = n86282 & n65057 ;
  assign n86283 = ~n64513 ;
  assign n65059 = x103 & n86283 ;
  assign n86284 = ~n64511 ;
  assign n65060 = n86284 & n65059 ;
  assign n65061 = n64515 | n65060 ;
  assign n65063 = n65058 | n65061 ;
  assign n86285 = ~n64515 ;
  assign n65064 = n86285 & n65063 ;
  assign n86286 = ~n64504 ;
  assign n65065 = x104 & n86286 ;
  assign n86287 = ~n64502 ;
  assign n65066 = n86287 & n65065 ;
  assign n65067 = n64506 | n65066 ;
  assign n65068 = n65064 | n65067 ;
  assign n86288 = ~n64506 ;
  assign n65069 = n86288 & n65068 ;
  assign n86289 = ~n64495 ;
  assign n65070 = x105 & n86289 ;
  assign n86290 = ~n64493 ;
  assign n65071 = n86290 & n65070 ;
  assign n65072 = n64497 | n65071 ;
  assign n65074 = n65069 | n65072 ;
  assign n86291 = ~n64497 ;
  assign n65075 = n86291 & n65074 ;
  assign n86292 = ~n64486 ;
  assign n65076 = x106 & n86292 ;
  assign n86293 = ~n64484 ;
  assign n65077 = n86293 & n65076 ;
  assign n65078 = n64488 | n65077 ;
  assign n65079 = n65075 | n65078 ;
  assign n86294 = ~n64488 ;
  assign n65080 = n86294 & n65079 ;
  assign n86295 = ~n64477 ;
  assign n65081 = x107 & n86295 ;
  assign n86296 = ~n64475 ;
  assign n65082 = n86296 & n65081 ;
  assign n65083 = n64479 | n65082 ;
  assign n65085 = n65080 | n65083 ;
  assign n86297 = ~n64479 ;
  assign n65086 = n86297 & n65085 ;
  assign n86298 = ~n64469 ;
  assign n65087 = x108 & n86298 ;
  assign n86299 = ~n64467 ;
  assign n65088 = n86299 & n65087 ;
  assign n65089 = n64471 | n65088 ;
  assign n65090 = n65086 | n65089 ;
  assign n86300 = ~n64471 ;
  assign n65091 = n86300 & n65090 ;
  assign n86301 = ~n64460 ;
  assign n65092 = x109 & n86301 ;
  assign n86302 = ~n64458 ;
  assign n65093 = n86302 & n65092 ;
  assign n65094 = n64462 | n65093 ;
  assign n65096 = n65091 | n65094 ;
  assign n86303 = ~n64462 ;
  assign n65097 = n86303 & n65096 ;
  assign n86304 = ~n64451 ;
  assign n65098 = x110 & n86304 ;
  assign n86305 = ~n64449 ;
  assign n65099 = n86305 & n65098 ;
  assign n65100 = n64453 | n65099 ;
  assign n65101 = n65097 | n65100 ;
  assign n86306 = ~n64453 ;
  assign n65102 = n86306 & n65101 ;
  assign n86307 = ~n64443 ;
  assign n65103 = x111 & n86307 ;
  assign n86308 = ~n64441 ;
  assign n65104 = n86308 & n65103 ;
  assign n65105 = n64445 | n65104 ;
  assign n65107 = n65102 | n65105 ;
  assign n86309 = ~n64445 ;
  assign n65108 = n86309 & n65107 ;
  assign n86310 = ~n64435 ;
  assign n65109 = x112 & n86310 ;
  assign n86311 = ~n64433 ;
  assign n65110 = n86311 & n65109 ;
  assign n65111 = n64437 | n65110 ;
  assign n65112 = n65108 | n65111 ;
  assign n86312 = ~n64437 ;
  assign n65113 = n86312 & n65112 ;
  assign n86313 = ~n64426 ;
  assign n65114 = x113 & n86313 ;
  assign n86314 = ~n64424 ;
  assign n65115 = n86314 & n65114 ;
  assign n65116 = n64428 | n65115 ;
  assign n65118 = n65113 | n65116 ;
  assign n86315 = ~n64428 ;
  assign n65119 = n86315 & n65118 ;
  assign n86316 = ~n64417 ;
  assign n65120 = x114 & n86316 ;
  assign n86317 = ~n64415 ;
  assign n65121 = n86317 & n65120 ;
  assign n65122 = n64419 | n65121 ;
  assign n65123 = n65119 | n65122 ;
  assign n86318 = ~n64419 ;
  assign n65124 = n86318 & n65123 ;
  assign n86319 = ~n64408 ;
  assign n65125 = x115 & n86319 ;
  assign n86320 = ~n64406 ;
  assign n65126 = n86320 & n65125 ;
  assign n65127 = n64410 | n65126 ;
  assign n65129 = n65124 | n65127 ;
  assign n86321 = ~n64410 ;
  assign n65130 = n86321 & n65129 ;
  assign n86322 = ~n64400 ;
  assign n65131 = x116 & n86322 ;
  assign n86323 = ~n64398 ;
  assign n65132 = n86323 & n65131 ;
  assign n65133 = n64402 | n65132 ;
  assign n65134 = n65130 | n65133 ;
  assign n86324 = ~n64402 ;
  assign n65135 = n86324 & n65134 ;
  assign n86325 = ~n64392 ;
  assign n65136 = x117 & n86325 ;
  assign n86326 = ~n64390 ;
  assign n65137 = n86326 & n65136 ;
  assign n65138 = n64394 | n65137 ;
  assign n65140 = n65135 | n65138 ;
  assign n86327 = ~n64394 ;
  assign n65141 = n86327 & n65140 ;
  assign n86328 = ~n64383 ;
  assign n65142 = x118 & n86328 ;
  assign n86329 = ~n64381 ;
  assign n65143 = n86329 & n65142 ;
  assign n65144 = n64385 | n65143 ;
  assign n65145 = n65141 | n65144 ;
  assign n86330 = ~n64385 ;
  assign n65146 = n86330 & n65145 ;
  assign n86331 = ~n64374 ;
  assign n65147 = x119 & n86331 ;
  assign n86332 = ~n64372 ;
  assign n65148 = n86332 & n65147 ;
  assign n65149 = n64376 | n65148 ;
  assign n65151 = n65146 | n65149 ;
  assign n86333 = ~n64376 ;
  assign n65152 = n86333 & n65151 ;
  assign n86334 = ~n64365 ;
  assign n65153 = x120 & n86334 ;
  assign n86335 = ~n64363 ;
  assign n65154 = n86335 & n65153 ;
  assign n65155 = n64367 | n65154 ;
  assign n65156 = n65152 | n65155 ;
  assign n86336 = ~n64367 ;
  assign n65157 = n86336 & n65156 ;
  assign n86337 = ~n64357 ;
  assign n65158 = x121 & n86337 ;
  assign n86338 = ~n64355 ;
  assign n65159 = n86338 & n65158 ;
  assign n65160 = n64359 | n65159 ;
  assign n65162 = n65157 | n65160 ;
  assign n86339 = ~n64359 ;
  assign n65163 = n86339 & n65162 ;
  assign n86340 = ~n64348 ;
  assign n65164 = x122 & n86340 ;
  assign n86341 = ~n64346 ;
  assign n65165 = n86341 & n65164 ;
  assign n65166 = n64350 | n65165 ;
  assign n65167 = n65163 | n65166 ;
  assign n86342 = ~n64350 ;
  assign n65168 = n86342 & n65167 ;
  assign n86343 = ~n64339 ;
  assign n65169 = x123 & n86343 ;
  assign n86344 = ~n64337 ;
  assign n65170 = n86344 & n65169 ;
  assign n65171 = n64341 | n65170 ;
  assign n65173 = n65168 | n65171 ;
  assign n86345 = ~n64341 ;
  assign n65174 = n86345 & n65173 ;
  assign n86346 = ~n64330 ;
  assign n65175 = x124 & n86346 ;
  assign n86347 = ~n64328 ;
  assign n65176 = n86347 & n65175 ;
  assign n65177 = n64332 | n65176 ;
  assign n65178 = n65174 | n65177 ;
  assign n86348 = ~n64332 ;
  assign n65179 = n86348 & n65178 ;
  assign n86349 = ~n64321 ;
  assign n65180 = x125 & n86349 ;
  assign n86350 = ~n64319 ;
  assign n65181 = n86350 & n65180 ;
  assign n65182 = n64323 | n65181 ;
  assign n65184 = n65179 | n65182 ;
  assign n86351 = ~n64323 ;
  assign n65185 = n86351 & n65184 ;
  assign n86352 = ~n64313 ;
  assign n65186 = x126 & n86352 ;
  assign n86353 = ~n64311 ;
  assign n65187 = n86353 & n65186 ;
  assign n65188 = n64315 | n65187 ;
  assign n65189 = n65185 | n65188 ;
  assign n86354 = ~n64315 ;
  assign n65190 = n86354 & n65189 ;
  assign n86355 = ~n64303 ;
  assign n65191 = x127 & n86355 ;
  assign n86356 = ~n64301 ;
  assign n65192 = n86356 & n65191 ;
  assign n65193 = n64305 | n65192 ;
  assign n65194 = n65190 | n65193 ;
  assign n86357 = ~n64305 ;
  assign n65195 = n86357 & n65194 ;
  assign n86358 = ~n65195 ;
  assign n65197 = n32480 & n86358 ;
  assign n65196 = x64 & n86358 ;
  assign n86359 = ~n65196 ;
  assign n65198 = x0 & n86359 ;
  assign n193 = n65197 | n65198 ;
  assign n65200 = n32480 & n64849 ;
  assign n65201 = n86170 & n65200 ;
  assign n86360 = ~n65201 ;
  assign n65202 = n64851 & n86360 ;
  assign n65204 = n86358 & n65202 ;
  assign n65203 = n86357 & n64846 ;
  assign n65205 = n65194 & n65203 ;
  assign n194 = n65204 | n65205 ;
  assign n65207 = n64852 | n64856 ;
  assign n86361 = ~n65207 ;
  assign n65208 = n64851 & n86361 ;
  assign n86362 = ~n64853 ;
  assign n65209 = n86362 & n64856 ;
  assign n65210 = n65208 | n65209 ;
  assign n65212 = n86358 & n65210 ;
  assign n65211 = n86357 & n64842 ;
  assign n65213 = n65194 & n65211 ;
  assign n195 = n65212 | n65213 ;
  assign n64862 = n64843 | n64861 ;
  assign n86363 = ~n64862 ;
  assign n65215 = n64857 & n86363 ;
  assign n86364 = ~n64858 ;
  assign n65216 = n86364 & n64861 ;
  assign n65217 = n65215 | n65216 ;
  assign n65219 = n86358 & n65217 ;
  assign n65218 = n86357 & n64834 ;
  assign n65220 = n65194 & n65218 ;
  assign n196 = n65219 | n65220 ;
  assign n65222 = n64835 | n64867 ;
  assign n86365 = ~n65222 ;
  assign n65223 = n64863 & n86365 ;
  assign n86366 = ~n64864 ;
  assign n65224 = n86366 & n64867 ;
  assign n65225 = n65223 | n65224 ;
  assign n65227 = n86358 & n65225 ;
  assign n65226 = n86357 & n64825 ;
  assign n65228 = n65194 & n65226 ;
  assign n197 = n65227 | n65228 ;
  assign n86367 = ~n64869 ;
  assign n64873 = n86367 & n64872 ;
  assign n64874 = n64826 | n64872 ;
  assign n86368 = ~n64874 ;
  assign n65230 = n64868 & n86368 ;
  assign n65231 = n64873 | n65230 ;
  assign n65233 = n86358 & n65231 ;
  assign n65232 = n86357 & n64816 ;
  assign n65234 = n65194 & n65232 ;
  assign n198 = n65233 | n65234 ;
  assign n65236 = n64817 | n64879 ;
  assign n86369 = ~n65236 ;
  assign n65237 = n64875 & n86369 ;
  assign n86370 = ~n64876 ;
  assign n65238 = n86370 & n64879 ;
  assign n65239 = n65237 | n65238 ;
  assign n65241 = n86358 & n65239 ;
  assign n65240 = n86357 & n64807 ;
  assign n65242 = n65194 & n65240 ;
  assign n199 = n65241 | n65242 ;
  assign n86371 = ~n64881 ;
  assign n64885 = n86371 & n64884 ;
  assign n64886 = n64808 | n64884 ;
  assign n86372 = ~n64886 ;
  assign n65244 = n64880 & n86372 ;
  assign n65245 = n64885 | n65244 ;
  assign n65247 = n86358 & n65245 ;
  assign n65246 = n86357 & n64799 ;
  assign n65248 = n65194 & n65246 ;
  assign n200 = n65247 | n65248 ;
  assign n65250 = n64800 | n64891 ;
  assign n86373 = ~n65250 ;
  assign n65251 = n64887 & n86373 ;
  assign n86374 = ~n64888 ;
  assign n65252 = n86374 & n64891 ;
  assign n65253 = n65251 | n65252 ;
  assign n65255 = n86358 & n65253 ;
  assign n65254 = n86357 & n64790 ;
  assign n65256 = n65194 & n65254 ;
  assign n201 = n65255 | n65256 ;
  assign n86375 = ~n64893 ;
  assign n64897 = n86375 & n64896 ;
  assign n65258 = n64791 | n64896 ;
  assign n86376 = ~n65258 ;
  assign n65259 = n64892 & n86376 ;
  assign n65260 = n64897 | n65259 ;
  assign n65262 = n86358 & n65260 ;
  assign n65261 = n86357 & n64781 ;
  assign n65263 = n65194 & n65261 ;
  assign n202 = n65262 | n65263 ;
  assign n65265 = n64782 | n64902 ;
  assign n86377 = ~n65265 ;
  assign n65266 = n64898 & n86377 ;
  assign n86378 = ~n64899 ;
  assign n65267 = n86378 & n64902 ;
  assign n65268 = n65266 | n65267 ;
  assign n65270 = n86358 & n65268 ;
  assign n65269 = n86357 & n64772 ;
  assign n65271 = n65194 & n65269 ;
  assign n203 = n65270 | n65271 ;
  assign n86379 = ~n64904 ;
  assign n64908 = n86379 & n64907 ;
  assign n65273 = n64773 | n64907 ;
  assign n86380 = ~n65273 ;
  assign n65274 = n64903 & n86380 ;
  assign n65275 = n64908 | n65274 ;
  assign n65277 = n86358 & n65275 ;
  assign n65276 = n86357 & n64763 ;
  assign n65278 = n65194 & n65276 ;
  assign n204 = n65277 | n65278 ;
  assign n65280 = n64764 | n64913 ;
  assign n86381 = ~n65280 ;
  assign n65281 = n64909 & n86381 ;
  assign n86382 = ~n64910 ;
  assign n65282 = n86382 & n64913 ;
  assign n65283 = n65281 | n65282 ;
  assign n65285 = n86358 & n65283 ;
  assign n65284 = n86357 & n64754 ;
  assign n65286 = n65194 & n65284 ;
  assign n205 = n65285 | n65286 ;
  assign n86383 = ~n64915 ;
  assign n64919 = n86383 & n64918 ;
  assign n65288 = n64755 | n64918 ;
  assign n86384 = ~n65288 ;
  assign n65289 = n64914 & n86384 ;
  assign n65290 = n64919 | n65289 ;
  assign n65292 = n86358 & n65290 ;
  assign n65291 = n86357 & n64745 ;
  assign n65293 = n65194 & n65291 ;
  assign n206 = n65292 | n65293 ;
  assign n65295 = n64746 | n64924 ;
  assign n86385 = ~n65295 ;
  assign n65296 = n64920 & n86385 ;
  assign n86386 = ~n64921 ;
  assign n65297 = n86386 & n64924 ;
  assign n65298 = n65296 | n65297 ;
  assign n65300 = n86358 & n65298 ;
  assign n65299 = n86357 & n64737 ;
  assign n65301 = n65194 & n65299 ;
  assign n207 = n65300 | n65301 ;
  assign n86387 = ~n64926 ;
  assign n64930 = n86387 & n64929 ;
  assign n65303 = n64738 | n64929 ;
  assign n86388 = ~n65303 ;
  assign n65304 = n64925 & n86388 ;
  assign n65305 = n64930 | n65304 ;
  assign n65307 = n86358 & n65305 ;
  assign n65306 = n86357 & n64728 ;
  assign n65308 = n65194 & n65306 ;
  assign n208 = n65307 | n65308 ;
  assign n65310 = n64729 | n64935 ;
  assign n86389 = ~n65310 ;
  assign n65311 = n64931 & n86389 ;
  assign n86390 = ~n64932 ;
  assign n65312 = n86390 & n64935 ;
  assign n65313 = n65311 | n65312 ;
  assign n65315 = n86358 & n65313 ;
  assign n65314 = n86357 & n64719 ;
  assign n65316 = n65194 & n65314 ;
  assign n209 = n65315 | n65316 ;
  assign n86391 = ~n64937 ;
  assign n64941 = n86391 & n64940 ;
  assign n65318 = n64720 | n64940 ;
  assign n86392 = ~n65318 ;
  assign n65319 = n64936 & n86392 ;
  assign n65320 = n64941 | n65319 ;
  assign n65322 = n86358 & n65320 ;
  assign n65321 = n86357 & n64710 ;
  assign n65323 = n65194 & n65321 ;
  assign n210 = n65322 | n65323 ;
  assign n65325 = n64711 | n64946 ;
  assign n86393 = ~n65325 ;
  assign n65326 = n64942 & n86393 ;
  assign n86394 = ~n64943 ;
  assign n65327 = n86394 & n64946 ;
  assign n65328 = n65326 | n65327 ;
  assign n65330 = n86358 & n65328 ;
  assign n65329 = n86357 & n64702 ;
  assign n65331 = n65194 & n65329 ;
  assign n211 = n65330 | n65331 ;
  assign n86395 = ~n64948 ;
  assign n64952 = n86395 & n64951 ;
  assign n65333 = n64703 | n64951 ;
  assign n86396 = ~n65333 ;
  assign n65334 = n64947 & n86396 ;
  assign n65335 = n64952 | n65334 ;
  assign n65337 = n86358 & n65335 ;
  assign n65336 = n86357 & n64693 ;
  assign n65338 = n65194 & n65336 ;
  assign n212 = n65337 | n65338 ;
  assign n65340 = n64694 | n64957 ;
  assign n86397 = ~n65340 ;
  assign n65341 = n64953 & n86397 ;
  assign n86398 = ~n64954 ;
  assign n65342 = n86398 & n64957 ;
  assign n65343 = n65341 | n65342 ;
  assign n65345 = n86358 & n65343 ;
  assign n65344 = n86357 & n64684 ;
  assign n65346 = n65194 & n65344 ;
  assign n213 = n65345 | n65346 ;
  assign n86399 = ~n64959 ;
  assign n64963 = n86399 & n64962 ;
  assign n65348 = n64685 | n64962 ;
  assign n86400 = ~n65348 ;
  assign n65349 = n64958 & n86400 ;
  assign n65350 = n64963 | n65349 ;
  assign n65352 = n86358 & n65350 ;
  assign n65351 = n86357 & n64675 ;
  assign n65353 = n65194 & n65351 ;
  assign n214 = n65352 | n65353 ;
  assign n65355 = n64676 | n64968 ;
  assign n86401 = ~n65355 ;
  assign n65356 = n64964 & n86401 ;
  assign n86402 = ~n64965 ;
  assign n65357 = n86402 & n64968 ;
  assign n65358 = n65356 | n65357 ;
  assign n65360 = n86358 & n65358 ;
  assign n65359 = n86357 & n64666 ;
  assign n65361 = n65194 & n65359 ;
  assign n215 = n65360 | n65361 ;
  assign n86403 = ~n64970 ;
  assign n64974 = n86403 & n64973 ;
  assign n65363 = n64667 | n64973 ;
  assign n86404 = ~n65363 ;
  assign n65364 = n64969 & n86404 ;
  assign n65365 = n64974 | n65364 ;
  assign n65367 = n86358 & n65365 ;
  assign n65366 = n86357 & n64657 ;
  assign n65368 = n65194 & n65366 ;
  assign n216 = n65367 | n65368 ;
  assign n65370 = n64658 | n64979 ;
  assign n86405 = ~n65370 ;
  assign n65371 = n64975 & n86405 ;
  assign n86406 = ~n64976 ;
  assign n65372 = n86406 & n64979 ;
  assign n65373 = n65371 | n65372 ;
  assign n65375 = n86358 & n65373 ;
  assign n65374 = n86357 & n64648 ;
  assign n65376 = n65194 & n65374 ;
  assign n217 = n65375 | n65376 ;
  assign n86407 = ~n64981 ;
  assign n64985 = n86407 & n64984 ;
  assign n65378 = n64649 | n64984 ;
  assign n86408 = ~n65378 ;
  assign n65379 = n64980 & n86408 ;
  assign n65380 = n64985 | n65379 ;
  assign n65382 = n86358 & n65380 ;
  assign n65381 = n86357 & n64639 ;
  assign n65383 = n65194 & n65381 ;
  assign n218 = n65382 | n65383 ;
  assign n65385 = n64640 | n64990 ;
  assign n86409 = ~n65385 ;
  assign n65386 = n64986 & n86409 ;
  assign n86410 = ~n64987 ;
  assign n65387 = n86410 & n64990 ;
  assign n65388 = n65386 | n65387 ;
  assign n65390 = n86358 & n65388 ;
  assign n65389 = n86357 & n64630 ;
  assign n65391 = n65194 & n65389 ;
  assign n219 = n65390 | n65391 ;
  assign n86411 = ~n64992 ;
  assign n64996 = n86411 & n64995 ;
  assign n65393 = n64631 | n64995 ;
  assign n86412 = ~n65393 ;
  assign n65394 = n64991 & n86412 ;
  assign n65395 = n64996 | n65394 ;
  assign n65397 = n86358 & n65395 ;
  assign n65396 = n86357 & n64622 ;
  assign n65398 = n65194 & n65396 ;
  assign n220 = n65397 | n65398 ;
  assign n65400 = n64623 | n65001 ;
  assign n86413 = ~n65400 ;
  assign n65401 = n64997 & n86413 ;
  assign n86414 = ~n64998 ;
  assign n65402 = n86414 & n65001 ;
  assign n65403 = n65401 | n65402 ;
  assign n65405 = n86358 & n65403 ;
  assign n65404 = n86357 & n64613 ;
  assign n65406 = n65194 & n65404 ;
  assign n221 = n65405 | n65406 ;
  assign n86415 = ~n65003 ;
  assign n65007 = n86415 & n65006 ;
  assign n65408 = n64614 | n65006 ;
  assign n86416 = ~n65408 ;
  assign n65409 = n65002 & n86416 ;
  assign n65410 = n65007 | n65409 ;
  assign n65412 = n86358 & n65410 ;
  assign n65411 = n86357 & n64604 ;
  assign n65413 = n65194 & n65411 ;
  assign n222 = n65412 | n65413 ;
  assign n65415 = n64605 | n65012 ;
  assign n86417 = ~n65415 ;
  assign n65416 = n65008 & n86417 ;
  assign n86418 = ~n65009 ;
  assign n65417 = n86418 & n65012 ;
  assign n65418 = n65416 | n65417 ;
  assign n65420 = n86358 & n65418 ;
  assign n65419 = n86357 & n64595 ;
  assign n65421 = n65194 & n65419 ;
  assign n223 = n65420 | n65421 ;
  assign n86419 = ~n65014 ;
  assign n65018 = n86419 & n65017 ;
  assign n65423 = n64596 | n65017 ;
  assign n86420 = ~n65423 ;
  assign n65424 = n65013 & n86420 ;
  assign n65425 = n65018 | n65424 ;
  assign n65427 = n86358 & n65425 ;
  assign n65426 = n86357 & n64586 ;
  assign n65428 = n65194 & n65426 ;
  assign n224 = n65427 | n65428 ;
  assign n65430 = n64587 | n65023 ;
  assign n86421 = ~n65430 ;
  assign n65431 = n65019 & n86421 ;
  assign n86422 = ~n65020 ;
  assign n65432 = n86422 & n65023 ;
  assign n65433 = n65431 | n65432 ;
  assign n65435 = n86358 & n65433 ;
  assign n65434 = n86357 & n64577 ;
  assign n65436 = n65194 & n65434 ;
  assign n225 = n65435 | n65436 ;
  assign n86423 = ~n65025 ;
  assign n65029 = n86423 & n65028 ;
  assign n65438 = n64578 | n65028 ;
  assign n86424 = ~n65438 ;
  assign n65439 = n65024 & n86424 ;
  assign n65440 = n65029 | n65439 ;
  assign n65442 = n86358 & n65440 ;
  assign n65441 = n86357 & n64568 ;
  assign n65443 = n65194 & n65441 ;
  assign n226 = n65442 | n65443 ;
  assign n65445 = n64569 | n65034 ;
  assign n86425 = ~n65445 ;
  assign n65446 = n65030 & n86425 ;
  assign n86426 = ~n65031 ;
  assign n65447 = n86426 & n65034 ;
  assign n65448 = n65446 | n65447 ;
  assign n65450 = n86358 & n65448 ;
  assign n65449 = n86357 & n64559 ;
  assign n65451 = n65194 & n65449 ;
  assign n227 = n65450 | n65451 ;
  assign n86427 = ~n65036 ;
  assign n65040 = n86427 & n65039 ;
  assign n65453 = n64560 | n65039 ;
  assign n86428 = ~n65453 ;
  assign n65454 = n65035 & n86428 ;
  assign n65455 = n65040 | n65454 ;
  assign n65457 = n86358 & n65455 ;
  assign n65456 = n86357 & n64550 ;
  assign n65458 = n65194 & n65456 ;
  assign n228 = n65457 | n65458 ;
  assign n65460 = n64551 | n65045 ;
  assign n86429 = ~n65460 ;
  assign n65461 = n65041 & n86429 ;
  assign n86430 = ~n65042 ;
  assign n65462 = n86430 & n65045 ;
  assign n65463 = n65461 | n65462 ;
  assign n65465 = n86358 & n65463 ;
  assign n65464 = n86357 & n64541 ;
  assign n65466 = n65194 & n65464 ;
  assign n229 = n65465 | n65466 ;
  assign n86431 = ~n65047 ;
  assign n65051 = n86431 & n65050 ;
  assign n65468 = n64542 | n65050 ;
  assign n86432 = ~n65468 ;
  assign n65469 = n65046 & n86432 ;
  assign n65470 = n65051 | n65469 ;
  assign n65472 = n86358 & n65470 ;
  assign n65471 = n86357 & n64532 ;
  assign n65473 = n65194 & n65471 ;
  assign n230 = n65472 | n65473 ;
  assign n65475 = n64533 | n65056 ;
  assign n86433 = ~n65475 ;
  assign n65476 = n65052 & n86433 ;
  assign n86434 = ~n65053 ;
  assign n65477 = n86434 & n65056 ;
  assign n65478 = n65476 | n65477 ;
  assign n65480 = n86358 & n65478 ;
  assign n65479 = n86357 & n64523 ;
  assign n65481 = n65194 & n65479 ;
  assign n231 = n65480 | n65481 ;
  assign n86435 = ~n65058 ;
  assign n65062 = n86435 & n65061 ;
  assign n65483 = n64524 | n65061 ;
  assign n86436 = ~n65483 ;
  assign n65484 = n65057 & n86436 ;
  assign n65485 = n65062 | n65484 ;
  assign n65487 = n86358 & n65485 ;
  assign n65486 = n86357 & n64514 ;
  assign n65488 = n65194 & n65486 ;
  assign n232 = n65487 | n65488 ;
  assign n65490 = n64515 | n65067 ;
  assign n86437 = ~n65490 ;
  assign n65491 = n65063 & n86437 ;
  assign n86438 = ~n65064 ;
  assign n65492 = n86438 & n65067 ;
  assign n65493 = n65491 | n65492 ;
  assign n65495 = n86358 & n65493 ;
  assign n65494 = n86357 & n64505 ;
  assign n65496 = n65194 & n65494 ;
  assign n233 = n65495 | n65496 ;
  assign n86439 = ~n65069 ;
  assign n65073 = n86439 & n65072 ;
  assign n65498 = n64506 | n65072 ;
  assign n86440 = ~n65498 ;
  assign n65499 = n65068 & n86440 ;
  assign n65500 = n65073 | n65499 ;
  assign n65502 = n86358 & n65500 ;
  assign n65501 = n86357 & n64496 ;
  assign n65503 = n65194 & n65501 ;
  assign n234 = n65502 | n65503 ;
  assign n65505 = n64497 | n65078 ;
  assign n86441 = ~n65505 ;
  assign n65506 = n65074 & n86441 ;
  assign n86442 = ~n65075 ;
  assign n65507 = n86442 & n65078 ;
  assign n65508 = n65506 | n65507 ;
  assign n65510 = n86358 & n65508 ;
  assign n65509 = n86357 & n64487 ;
  assign n65511 = n65194 & n65509 ;
  assign n235 = n65510 | n65511 ;
  assign n86443 = ~n65080 ;
  assign n65084 = n86443 & n65083 ;
  assign n65513 = n64488 | n65083 ;
  assign n86444 = ~n65513 ;
  assign n65514 = n65079 & n86444 ;
  assign n65515 = n65084 | n65514 ;
  assign n65517 = n86358 & n65515 ;
  assign n65516 = n86357 & n64478 ;
  assign n65518 = n65194 & n65516 ;
  assign n236 = n65517 | n65518 ;
  assign n65520 = n64479 | n65089 ;
  assign n86445 = ~n65520 ;
  assign n65521 = n65085 & n86445 ;
  assign n86446 = ~n65086 ;
  assign n65522 = n86446 & n65089 ;
  assign n65523 = n65521 | n65522 ;
  assign n65525 = n86358 & n65523 ;
  assign n65524 = n86357 & n64470 ;
  assign n65526 = n65194 & n65524 ;
  assign n237 = n65525 | n65526 ;
  assign n86447 = ~n65091 ;
  assign n65095 = n86447 & n65094 ;
  assign n65528 = n64471 | n65094 ;
  assign n86448 = ~n65528 ;
  assign n65529 = n65090 & n86448 ;
  assign n65530 = n65095 | n65529 ;
  assign n65532 = n86358 & n65530 ;
  assign n65531 = n86357 & n64461 ;
  assign n65533 = n65194 & n65531 ;
  assign n238 = n65532 | n65533 ;
  assign n65535 = n64462 | n65100 ;
  assign n86449 = ~n65535 ;
  assign n65536 = n65096 & n86449 ;
  assign n86450 = ~n65097 ;
  assign n65537 = n86450 & n65100 ;
  assign n65538 = n65536 | n65537 ;
  assign n65540 = n86358 & n65538 ;
  assign n65539 = n86357 & n64452 ;
  assign n65541 = n65194 & n65539 ;
  assign n239 = n65540 | n65541 ;
  assign n86451 = ~n65102 ;
  assign n65106 = n86451 & n65105 ;
  assign n65543 = n64453 | n65105 ;
  assign n86452 = ~n65543 ;
  assign n65544 = n65101 & n86452 ;
  assign n65545 = n65106 | n65544 ;
  assign n65547 = n86358 & n65545 ;
  assign n65546 = n86357 & n64444 ;
  assign n65548 = n65194 & n65546 ;
  assign n240 = n65547 | n65548 ;
  assign n65550 = n64445 | n65111 ;
  assign n86453 = ~n65550 ;
  assign n65551 = n65107 & n86453 ;
  assign n86454 = ~n65108 ;
  assign n65552 = n86454 & n65111 ;
  assign n65553 = n65551 | n65552 ;
  assign n65555 = n86358 & n65553 ;
  assign n65554 = n86357 & n64436 ;
  assign n65556 = n65194 & n65554 ;
  assign n241 = n65555 | n65556 ;
  assign n86455 = ~n65113 ;
  assign n65117 = n86455 & n65116 ;
  assign n65558 = n64437 | n65116 ;
  assign n86456 = ~n65558 ;
  assign n65559 = n65112 & n86456 ;
  assign n65560 = n65117 | n65559 ;
  assign n65562 = n86358 & n65560 ;
  assign n65561 = n86357 & n64427 ;
  assign n65563 = n65194 & n65561 ;
  assign n242 = n65562 | n65563 ;
  assign n65565 = n64428 | n65122 ;
  assign n86457 = ~n65565 ;
  assign n65566 = n65118 & n86457 ;
  assign n86458 = ~n65119 ;
  assign n65567 = n86458 & n65122 ;
  assign n65568 = n65566 | n65567 ;
  assign n65570 = n86358 & n65568 ;
  assign n65569 = n86357 & n64418 ;
  assign n65571 = n65194 & n65569 ;
  assign n243 = n65570 | n65571 ;
  assign n86459 = ~n65124 ;
  assign n65128 = n86459 & n65127 ;
  assign n65573 = n64419 | n65127 ;
  assign n86460 = ~n65573 ;
  assign n65574 = n65123 & n86460 ;
  assign n65575 = n65128 | n65574 ;
  assign n65577 = n86358 & n65575 ;
  assign n65576 = n86357 & n64409 ;
  assign n65578 = n65194 & n65576 ;
  assign n244 = n65577 | n65578 ;
  assign n65580 = n64410 | n65133 ;
  assign n86461 = ~n65580 ;
  assign n65581 = n65129 & n86461 ;
  assign n86462 = ~n65130 ;
  assign n65582 = n86462 & n65133 ;
  assign n65583 = n65581 | n65582 ;
  assign n65585 = n86358 & n65583 ;
  assign n65584 = n86357 & n64401 ;
  assign n65586 = n65194 & n65584 ;
  assign n245 = n65585 | n65586 ;
  assign n86463 = ~n65135 ;
  assign n65139 = n86463 & n65138 ;
  assign n65588 = n64402 | n65138 ;
  assign n86464 = ~n65588 ;
  assign n65589 = n65134 & n86464 ;
  assign n65590 = n65139 | n65589 ;
  assign n65592 = n86358 & n65590 ;
  assign n65591 = n86357 & n64393 ;
  assign n65593 = n65194 & n65591 ;
  assign n246 = n65592 | n65593 ;
  assign n65595 = n64394 | n65144 ;
  assign n86465 = ~n65595 ;
  assign n65596 = n65140 & n86465 ;
  assign n86466 = ~n65141 ;
  assign n65597 = n86466 & n65144 ;
  assign n65598 = n65596 | n65597 ;
  assign n65600 = n86358 & n65598 ;
  assign n65599 = n86357 & n64384 ;
  assign n65601 = n65194 & n65599 ;
  assign n247 = n65600 | n65601 ;
  assign n86467 = ~n65146 ;
  assign n65150 = n86467 & n65149 ;
  assign n65603 = n64385 | n65149 ;
  assign n86468 = ~n65603 ;
  assign n65604 = n65145 & n86468 ;
  assign n65605 = n65150 | n65604 ;
  assign n65607 = n86358 & n65605 ;
  assign n65606 = n86357 & n64375 ;
  assign n65608 = n65194 & n65606 ;
  assign n248 = n65607 | n65608 ;
  assign n65610 = n64376 | n65155 ;
  assign n86469 = ~n65610 ;
  assign n65611 = n65151 & n86469 ;
  assign n86470 = ~n65152 ;
  assign n65612 = n86470 & n65155 ;
  assign n65613 = n65611 | n65612 ;
  assign n65615 = n86358 & n65613 ;
  assign n65614 = n86357 & n64366 ;
  assign n65616 = n65194 & n65614 ;
  assign n249 = n65615 | n65616 ;
  assign n86471 = ~n65157 ;
  assign n65161 = n86471 & n65160 ;
  assign n65618 = n64367 | n65160 ;
  assign n86472 = ~n65618 ;
  assign n65619 = n65156 & n86472 ;
  assign n65620 = n65161 | n65619 ;
  assign n65622 = n86358 & n65620 ;
  assign n65621 = n86357 & n64358 ;
  assign n65623 = n65194 & n65621 ;
  assign n250 = n65622 | n65623 ;
  assign n65625 = n64359 | n65166 ;
  assign n86473 = ~n65625 ;
  assign n65626 = n65162 & n86473 ;
  assign n86474 = ~n65163 ;
  assign n65627 = n86474 & n65166 ;
  assign n65628 = n65626 | n65627 ;
  assign n65630 = n86358 & n65628 ;
  assign n65629 = n86357 & n64349 ;
  assign n65631 = n65194 & n65629 ;
  assign n251 = n65630 | n65631 ;
  assign n86475 = ~n65168 ;
  assign n65172 = n86475 & n65171 ;
  assign n65633 = n64350 | n65171 ;
  assign n86476 = ~n65633 ;
  assign n65634 = n65167 & n86476 ;
  assign n65635 = n65172 | n65634 ;
  assign n65637 = n86358 & n65635 ;
  assign n65636 = n86357 & n64340 ;
  assign n65638 = n65194 & n65636 ;
  assign n252 = n65637 | n65638 ;
  assign n65640 = n64341 | n65177 ;
  assign n86477 = ~n65640 ;
  assign n65641 = n65173 & n86477 ;
  assign n86478 = ~n65174 ;
  assign n65642 = n86478 & n65177 ;
  assign n65643 = n65641 | n65642 ;
  assign n65645 = n86358 & n65643 ;
  assign n65644 = n86357 & n64331 ;
  assign n65646 = n65194 & n65644 ;
  assign n253 = n65645 | n65646 ;
  assign n86479 = ~n65179 ;
  assign n65183 = n86479 & n65182 ;
  assign n65648 = n64332 | n65182 ;
  assign n86480 = ~n65648 ;
  assign n65649 = n65178 & n86480 ;
  assign n65650 = n65183 | n65649 ;
  assign n65652 = n86358 & n65650 ;
  assign n65651 = n86357 & n64322 ;
  assign n65653 = n65194 & n65651 ;
  assign n254 = n65652 | n65653 ;
  assign n65655 = n64323 | n65188 ;
  assign n86481 = ~n65655 ;
  assign n65656 = n65184 & n86481 ;
  assign n86482 = ~n65185 ;
  assign n65657 = n86482 & n65188 ;
  assign n65658 = n65656 | n65657 ;
  assign n65660 = n86358 & n65658 ;
  assign n65659 = n86357 & n64314 ;
  assign n65661 = n65194 & n65659 ;
  assign n255 = n65660 | n65661 ;
  assign n86483 = ~n65190 ;
  assign n65663 = n64305 & n86483 ;
  assign n65664 = x127 & n64304 ;
  assign n65665 = n65194 & n65664 ;
  assign n256 = n65663 | n65665 ;
  assign n129 = ~n33034 ;
  assign n188 = ~n471 ;
  assign n189 = ~n382 ;
  assign n191 = ~n33037 ;
  assign n192 = ~n33042 ;
  assign y0 = n129 ;
  assign y1 = n130 ;
  assign y2 = n131 ;
  assign y3 = n132 ;
  assign y4 = n133 ;
  assign y5 = n134 ;
  assign y6 = n135 ;
  assign y7 = n136 ;
  assign y8 = n137 ;
  assign y9 = n138 ;
  assign y10 = n139 ;
  assign y11 = n140 ;
  assign y12 = n141 ;
  assign y13 = n142 ;
  assign y14 = n143 ;
  assign y15 = n144 ;
  assign y16 = n145 ;
  assign y17 = n146 ;
  assign y18 = n147 ;
  assign y19 = n148 ;
  assign y20 = n149 ;
  assign y21 = n150 ;
  assign y22 = n151 ;
  assign y23 = n152 ;
  assign y24 = n153 ;
  assign y25 = n154 ;
  assign y26 = n155 ;
  assign y27 = n156 ;
  assign y28 = n157 ;
  assign y29 = n158 ;
  assign y30 = n159 ;
  assign y31 = n160 ;
  assign y32 = n161 ;
  assign y33 = n162 ;
  assign y34 = n163 ;
  assign y35 = n164 ;
  assign y36 = n165 ;
  assign y37 = n166 ;
  assign y38 = n167 ;
  assign y39 = n168 ;
  assign y40 = n169 ;
  assign y41 = n170 ;
  assign y42 = n171 ;
  assign y43 = n172 ;
  assign y44 = n173 ;
  assign y45 = n174 ;
  assign y46 = n175 ;
  assign y47 = n176 ;
  assign y48 = n177 ;
  assign y49 = n178 ;
  assign y50 = n179 ;
  assign y51 = n180 ;
  assign y52 = n181 ;
  assign y53 = n182 ;
  assign y54 = n183 ;
  assign y55 = n184 ;
  assign y56 = n185 ;
  assign y57 = n186 ;
  assign y58 = n187 ;
  assign y59 = n188 ;
  assign y60 = n189 ;
  assign y61 = n190 ;
  assign y62 = n191 ;
  assign y63 = n192 ;
  assign y64 = n193 ;
  assign y65 = n194 ;
  assign y66 = n195 ;
  assign y67 = n196 ;
  assign y68 = n197 ;
  assign y69 = n198 ;
  assign y70 = n199 ;
  assign y71 = n200 ;
  assign y72 = n201 ;
  assign y73 = n202 ;
  assign y74 = n203 ;
  assign y75 = n204 ;
  assign y76 = n205 ;
  assign y77 = n206 ;
  assign y78 = n207 ;
  assign y79 = n208 ;
  assign y80 = n209 ;
  assign y81 = n210 ;
  assign y82 = n211 ;
  assign y83 = n212 ;
  assign y84 = n213 ;
  assign y85 = n214 ;
  assign y86 = n215 ;
  assign y87 = n216 ;
  assign y88 = n217 ;
  assign y89 = n218 ;
  assign y90 = n219 ;
  assign y91 = n220 ;
  assign y92 = n221 ;
  assign y93 = n222 ;
  assign y94 = n223 ;
  assign y95 = n224 ;
  assign y96 = n225 ;
  assign y97 = n226 ;
  assign y98 = n227 ;
  assign y99 = n228 ;
  assign y100 = n229 ;
  assign y101 = n230 ;
  assign y102 = n231 ;
  assign y103 = n232 ;
  assign y104 = n233 ;
  assign y105 = n234 ;
  assign y106 = n235 ;
  assign y107 = n236 ;
  assign y108 = n237 ;
  assign y109 = n238 ;
  assign y110 = n239 ;
  assign y111 = n240 ;
  assign y112 = n241 ;
  assign y113 = n242 ;
  assign y114 = n243 ;
  assign y115 = n244 ;
  assign y116 = n245 ;
  assign y117 = n246 ;
  assign y118 = n247 ;
  assign y119 = n248 ;
  assign y120 = n249 ;
  assign y121 = n250 ;
  assign y122 = n251 ;
  assign y123 = n252 ;
  assign y124 = n253 ;
  assign y125 = n254 ;
  assign y126 = n255 ;
  assign y127 = n256 ;
endmodule
