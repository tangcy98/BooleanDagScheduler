module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 ;
  assign n13 = x0 | x2 ;
  assign n14 = x1 | x3 ;
  assign n15 = n13 | n14 ;
  assign n192 = x4 | x5 ;
  assign n313 = ~x6 ;
  assign n244 = n313 & x7 ;
  assign n314 = ~n192 ;
  assign n296 = n314 & n244 ;
  assign n315 = ~n15 ;
  assign n309 = n315 & n296 ;
  assign n316 = ~x2 ;
  assign n16 = x0 & n316 ;
  assign n317 = ~n14 ;
  assign n17 = n317 & n16 ;
  assign n307 = n17 & n296 ;
  assign n318 = ~x3 ;
  assign n18 = x1 & n318 ;
  assign n319 = ~n13 ;
  assign n19 = n319 & n18 ;
  assign n305 = n19 & n296 ;
  assign n20 = n16 & n18 ;
  assign n301 = n20 & n296 ;
  assign n320 = ~x0 ;
  assign n21 = n320 & x2 ;
  assign n22 = n317 & n21 ;
  assign n298 = n22 & n296 ;
  assign n9 = x0 & x2 ;
  assign n23 = n9 & n317 ;
  assign n308 = n23 & n296 ;
  assign n24 = n18 & n21 ;
  assign n304 = n24 & n296 ;
  assign n25 = n9 & n18 ;
  assign n300 = n25 & n296 ;
  assign n321 = ~x1 ;
  assign n26 = n321 & x3 ;
  assign n27 = n319 & n26 ;
  assign n299 = n27 & n296 ;
  assign n28 = n16 & n26 ;
  assign n302 = n28 & n296 ;
  assign n10 = x1 & x3 ;
  assign n29 = n10 & n319 ;
  assign n297 = n29 & n296 ;
  assign n30 = n10 & n16 ;
  assign n306 = n30 & n296 ;
  assign n31 = n21 & n26 ;
  assign n303 = n31 & n296 ;
  assign n32 = n9 & n26 ;
  assign n310 = n32 & n296 ;
  assign n33 = n10 & n21 ;
  assign n311 = n33 & n296 ;
  assign n34 = n9 & n10 ;
  assign n312 = n34 & n296 ;
  assign n322 = ~x5 ;
  assign n35 = x4 & n322 ;
  assign n245 = n35 & n244 ;
  assign n251 = n315 & n245 ;
  assign n259 = n17 & n245 ;
  assign n258 = n19 & n245 ;
  assign n257 = n20 & n245 ;
  assign n255 = n22 & n245 ;
  assign n254 = n23 & n245 ;
  assign n252 = n24 & n245 ;
  assign n250 = n25 & n245 ;
  assign n249 = n27 & n245 ;
  assign n248 = n28 & n245 ;
  assign n247 = n29 & n245 ;
  assign n253 = n30 & n245 ;
  assign n246 = n31 & n245 ;
  assign n260 = n32 & n245 ;
  assign n261 = n33 & n245 ;
  assign n256 = n34 & n245 ;
  assign n323 = ~x4 ;
  assign n36 = n323 & x5 ;
  assign n262 = n36 & n244 ;
  assign n277 = n315 & n262 ;
  assign n274 = n17 & n262 ;
  assign n269 = n19 & n262 ;
  assign n273 = n20 & n262 ;
  assign n272 = n22 & n262 ;
  assign n264 = n23 & n262 ;
  assign n268 = n24 & n262 ;
  assign n270 = n25 & n262 ;
  assign n267 = n27 & n262 ;
  assign n275 = n28 & n262 ;
  assign n266 = n29 & n262 ;
  assign n265 = n30 & n262 ;
  assign n263 = n31 & n262 ;
  assign n278 = n32 & n262 ;
  assign n276 = n33 & n262 ;
  assign n271 = n34 & n262 ;
  assign n11 = x4 & x5 ;
  assign n279 = n11 & n244 ;
  assign n288 = n315 & n279 ;
  assign n292 = n17 & n279 ;
  assign n291 = n19 & n279 ;
  assign n289 = n20 & n279 ;
  assign n285 = n22 & n279 ;
  assign n284 = n23 & n279 ;
  assign n283 = n24 & n279 ;
  assign n287 = n25 & n279 ;
  assign n282 = n27 & n279 ;
  assign n281 = n28 & n279 ;
  assign n286 = n29 & n279 ;
  assign n290 = n30 & n279 ;
  assign n280 = n31 & n279 ;
  assign n293 = n32 & n279 ;
  assign n294 = n33 & n279 ;
  assign n295 = n34 & n279 ;
  assign n12 = x6 & x7 ;
  assign n193 = n12 & n314 ;
  assign n205 = n315 & n193 ;
  assign n196 = n17 & n193 ;
  assign n207 = n19 & n193 ;
  assign n204 = n20 & n193 ;
  assign n200 = n22 & n193 ;
  assign n208 = n23 & n193 ;
  assign n201 = n24 & n193 ;
  assign n198 = n25 & n193 ;
  assign n206 = n27 & n193 ;
  assign n199 = n28 & n193 ;
  assign n197 = n29 & n193 ;
  assign n195 = n30 & n193 ;
  assign n194 = n31 & n193 ;
  assign n202 = n32 & n193 ;
  assign n209 = n33 & n193 ;
  assign n203 = n34 & n193 ;
  assign n37 = n12 & n35 ;
  assign n38 = n315 & n37 ;
  assign n39 = n17 & n37 ;
  assign n40 = n19 & n37 ;
  assign n41 = n20 & n37 ;
  assign n42 = n22 & n37 ;
  assign n43 = n23 & n37 ;
  assign n44 = n24 & n37 ;
  assign n45 = n25 & n37 ;
  assign n46 = n27 & n37 ;
  assign n47 = n28 & n37 ;
  assign n48 = n29 & n37 ;
  assign n49 = n30 & n37 ;
  assign n50 = n31 & n37 ;
  assign n51 = n32 & n37 ;
  assign n52 = n33 & n37 ;
  assign n53 = n34 & n37 ;
  assign n54 = n12 & n36 ;
  assign n55 = n315 & n54 ;
  assign n56 = n17 & n54 ;
  assign n57 = n19 & n54 ;
  assign n58 = n20 & n54 ;
  assign n59 = n22 & n54 ;
  assign n60 = n23 & n54 ;
  assign n61 = n24 & n54 ;
  assign n62 = n25 & n54 ;
  assign n63 = n27 & n54 ;
  assign n64 = n28 & n54 ;
  assign n65 = n29 & n54 ;
  assign n66 = n30 & n54 ;
  assign n67 = n31 & n54 ;
  assign n68 = n32 & n54 ;
  assign n69 = n33 & n54 ;
  assign n70 = n34 & n54 ;
  assign n71 = n11 & n12 ;
  assign n72 = n315 & n71 ;
  assign n73 = n17 & n71 ;
  assign n74 = n19 & n71 ;
  assign n75 = n20 & n71 ;
  assign n76 = n22 & n71 ;
  assign n77 = n23 & n71 ;
  assign n78 = n24 & n71 ;
  assign n79 = n25 & n71 ;
  assign n80 = n27 & n71 ;
  assign n81 = n28 & n71 ;
  assign n82 = n29 & n71 ;
  assign n83 = n30 & n71 ;
  assign n84 = n31 & n71 ;
  assign n85 = n32 & n71 ;
  assign n86 = n33 & n71 ;
  assign n87 = n34 & n71 ;
  assign n88 = x6 | x7 ;
  assign n210 = n88 | n192 ;
  assign n225 = n15 | n210 ;
  assign n324 = ~n210 ;
  assign n224 = n17 & n324 ;
  assign n220 = n19 & n324 ;
  assign n223 = n20 & n324 ;
  assign n222 = n22 & n324 ;
  assign n219 = n23 & n324 ;
  assign n218 = n24 & n324 ;
  assign n217 = n25 & n324 ;
  assign n214 = n27 & n324 ;
  assign n216 = n28 & n324 ;
  assign n213 = n29 & n324 ;
  assign n212 = n30 & n324 ;
  assign n211 = n31 & n324 ;
  assign n226 = n32 & n324 ;
  assign n221 = n33 & n324 ;
  assign n215 = n34 & n324 ;
  assign n325 = ~n88 ;
  assign n89 = n35 & n325 ;
  assign n90 = n315 & n89 ;
  assign n91 = n17 & n89 ;
  assign n92 = n19 & n89 ;
  assign n93 = n20 & n89 ;
  assign n94 = n22 & n89 ;
  assign n95 = n23 & n89 ;
  assign n96 = n24 & n89 ;
  assign n97 = n25 & n89 ;
  assign n98 = n27 & n89 ;
  assign n99 = n28 & n89 ;
  assign n100 = n29 & n89 ;
  assign n101 = n30 & n89 ;
  assign n102 = n31 & n89 ;
  assign n103 = n32 & n89 ;
  assign n104 = n33 & n89 ;
  assign n105 = n34 & n89 ;
  assign n106 = n36 & n325 ;
  assign n107 = n315 & n106 ;
  assign n108 = n17 & n106 ;
  assign n109 = n19 & n106 ;
  assign n110 = n20 & n106 ;
  assign n111 = n22 & n106 ;
  assign n112 = n23 & n106 ;
  assign n113 = n24 & n106 ;
  assign n114 = n25 & n106 ;
  assign n115 = n27 & n106 ;
  assign n116 = n28 & n106 ;
  assign n117 = n29 & n106 ;
  assign n118 = n30 & n106 ;
  assign n119 = n31 & n106 ;
  assign n120 = n32 & n106 ;
  assign n121 = n33 & n106 ;
  assign n122 = n34 & n106 ;
  assign n123 = n11 & n325 ;
  assign n124 = n315 & n123 ;
  assign n125 = n17 & n123 ;
  assign n126 = n19 & n123 ;
  assign n127 = n20 & n123 ;
  assign n128 = n22 & n123 ;
  assign n129 = n23 & n123 ;
  assign n130 = n24 & n123 ;
  assign n131 = n25 & n123 ;
  assign n132 = n27 & n123 ;
  assign n133 = n28 & n123 ;
  assign n134 = n29 & n123 ;
  assign n135 = n30 & n123 ;
  assign n136 = n31 & n123 ;
  assign n137 = n32 & n123 ;
  assign n138 = n33 & n123 ;
  assign n139 = n34 & n123 ;
  assign n326 = ~x7 ;
  assign n140 = x6 & n326 ;
  assign n227 = n140 & n314 ;
  assign n242 = n315 & n227 ;
  assign n237 = n17 & n227 ;
  assign n240 = n19 & n227 ;
  assign n236 = n20 & n227 ;
  assign n235 = n22 & n227 ;
  assign n232 = n23 & n227 ;
  assign n231 = n24 & n227 ;
  assign n234 = n25 & n227 ;
  assign n230 = n27 & n227 ;
  assign n233 = n28 & n227 ;
  assign n228 = n29 & n227 ;
  assign n239 = n30 & n227 ;
  assign n241 = n31 & n227 ;
  assign n243 = n32 & n227 ;
  assign n238 = n33 & n227 ;
  assign n229 = n34 & n227 ;
  assign n141 = n35 & n140 ;
  assign n142 = n315 & n141 ;
  assign n143 = n17 & n141 ;
  assign n144 = n19 & n141 ;
  assign n145 = n20 & n141 ;
  assign n146 = n22 & n141 ;
  assign n147 = n23 & n141 ;
  assign n148 = n24 & n141 ;
  assign n149 = n25 & n141 ;
  assign n150 = n27 & n141 ;
  assign n151 = n28 & n141 ;
  assign n152 = n29 & n141 ;
  assign n153 = n30 & n141 ;
  assign n154 = n31 & n141 ;
  assign n155 = n32 & n141 ;
  assign n156 = n33 & n141 ;
  assign n157 = n34 & n141 ;
  assign n158 = n36 & n140 ;
  assign n159 = n315 & n158 ;
  assign n160 = n17 & n158 ;
  assign n161 = n19 & n158 ;
  assign n162 = n20 & n158 ;
  assign n163 = n22 & n158 ;
  assign n164 = n23 & n158 ;
  assign n165 = n24 & n158 ;
  assign n166 = n25 & n158 ;
  assign n167 = n27 & n158 ;
  assign n168 = n28 & n158 ;
  assign n169 = n29 & n158 ;
  assign n170 = n30 & n158 ;
  assign n171 = n31 & n158 ;
  assign n172 = n32 & n158 ;
  assign n173 = n33 & n158 ;
  assign n174 = n34 & n158 ;
  assign n175 = n11 & n140 ;
  assign n176 = n315 & n175 ;
  assign n177 = n17 & n175 ;
  assign n178 = n19 & n175 ;
  assign n179 = n20 & n175 ;
  assign n180 = n22 & n175 ;
  assign n181 = n23 & n175 ;
  assign n182 = n24 & n175 ;
  assign n183 = n25 & n175 ;
  assign n184 = n27 & n175 ;
  assign n185 = n28 & n175 ;
  assign n186 = n29 & n175 ;
  assign n187 = n30 & n175 ;
  assign n188 = n31 & n175 ;
  assign n189 = n32 & n175 ;
  assign n190 = n33 & n175 ;
  assign n191 = n34 & n175 ;
  assign n327 = ~n225 ;
  assign y0 = n309 ;
  assign y1 = n307 ;
  assign y2 = n305 ;
  assign y3 = n301 ;
  assign y4 = n298 ;
  assign y5 = n308 ;
  assign y6 = n304 ;
  assign y7 = n300 ;
  assign y8 = n299 ;
  assign y9 = n302 ;
  assign y10 = n297 ;
  assign y11 = n306 ;
  assign y12 = n303 ;
  assign y13 = n310 ;
  assign y14 = n311 ;
  assign y15 = n312 ;
  assign y16 = n251 ;
  assign y17 = n259 ;
  assign y18 = n258 ;
  assign y19 = n257 ;
  assign y20 = n255 ;
  assign y21 = n254 ;
  assign y22 = n252 ;
  assign y23 = n250 ;
  assign y24 = n249 ;
  assign y25 = n248 ;
  assign y26 = n247 ;
  assign y27 = n253 ;
  assign y28 = n246 ;
  assign y29 = n260 ;
  assign y30 = n261 ;
  assign y31 = n256 ;
  assign y32 = n277 ;
  assign y33 = n274 ;
  assign y34 = n269 ;
  assign y35 = n273 ;
  assign y36 = n272 ;
  assign y37 = n264 ;
  assign y38 = n268 ;
  assign y39 = n270 ;
  assign y40 = n267 ;
  assign y41 = n275 ;
  assign y42 = n266 ;
  assign y43 = n265 ;
  assign y44 = n263 ;
  assign y45 = n278 ;
  assign y46 = n276 ;
  assign y47 = n271 ;
  assign y48 = n288 ;
  assign y49 = n292 ;
  assign y50 = n291 ;
  assign y51 = n289 ;
  assign y52 = n285 ;
  assign y53 = n284 ;
  assign y54 = n283 ;
  assign y55 = n287 ;
  assign y56 = n282 ;
  assign y57 = n281 ;
  assign y58 = n286 ;
  assign y59 = n290 ;
  assign y60 = n280 ;
  assign y61 = n293 ;
  assign y62 = n294 ;
  assign y63 = n295 ;
  assign y64 = n205 ;
  assign y65 = n196 ;
  assign y66 = n207 ;
  assign y67 = n204 ;
  assign y68 = n200 ;
  assign y69 = n208 ;
  assign y70 = n201 ;
  assign y71 = n198 ;
  assign y72 = n206 ;
  assign y73 = n199 ;
  assign y74 = n197 ;
  assign y75 = n195 ;
  assign y76 = n194 ;
  assign y77 = n202 ;
  assign y78 = n209 ;
  assign y79 = n203 ;
  assign y80 = n38 ;
  assign y81 = n39 ;
  assign y82 = n40 ;
  assign y83 = n41 ;
  assign y84 = n42 ;
  assign y85 = n43 ;
  assign y86 = n44 ;
  assign y87 = n45 ;
  assign y88 = n46 ;
  assign y89 = n47 ;
  assign y90 = n48 ;
  assign y91 = n49 ;
  assign y92 = n50 ;
  assign y93 = n51 ;
  assign y94 = n52 ;
  assign y95 = n53 ;
  assign y96 = n55 ;
  assign y97 = n56 ;
  assign y98 = n57 ;
  assign y99 = n58 ;
  assign y100 = n59 ;
  assign y101 = n60 ;
  assign y102 = n61 ;
  assign y103 = n62 ;
  assign y104 = n63 ;
  assign y105 = n64 ;
  assign y106 = n65 ;
  assign y107 = n66 ;
  assign y108 = n67 ;
  assign y109 = n68 ;
  assign y110 = n69 ;
  assign y111 = n70 ;
  assign y112 = n72 ;
  assign y113 = n73 ;
  assign y114 = n74 ;
  assign y115 = n75 ;
  assign y116 = n76 ;
  assign y117 = n77 ;
  assign y118 = n78 ;
  assign y119 = n79 ;
  assign y120 = n80 ;
  assign y121 = n81 ;
  assign y122 = n82 ;
  assign y123 = n83 ;
  assign y124 = n84 ;
  assign y125 = n85 ;
  assign y126 = n86 ;
  assign y127 = n87 ;
  assign y128 = n327 ;
  assign y129 = n224 ;
  assign y130 = n220 ;
  assign y131 = n223 ;
  assign y132 = n222 ;
  assign y133 = n219 ;
  assign y134 = n218 ;
  assign y135 = n217 ;
  assign y136 = n214 ;
  assign y137 = n216 ;
  assign y138 = n213 ;
  assign y139 = n212 ;
  assign y140 = n211 ;
  assign y141 = n226 ;
  assign y142 = n221 ;
  assign y143 = n215 ;
  assign y144 = n90 ;
  assign y145 = n91 ;
  assign y146 = n92 ;
  assign y147 = n93 ;
  assign y148 = n94 ;
  assign y149 = n95 ;
  assign y150 = n96 ;
  assign y151 = n97 ;
  assign y152 = n98 ;
  assign y153 = n99 ;
  assign y154 = n100 ;
  assign y155 = n101 ;
  assign y156 = n102 ;
  assign y157 = n103 ;
  assign y158 = n104 ;
  assign y159 = n105 ;
  assign y160 = n107 ;
  assign y161 = n108 ;
  assign y162 = n109 ;
  assign y163 = n110 ;
  assign y164 = n111 ;
  assign y165 = n112 ;
  assign y166 = n113 ;
  assign y167 = n114 ;
  assign y168 = n115 ;
  assign y169 = n116 ;
  assign y170 = n117 ;
  assign y171 = n118 ;
  assign y172 = n119 ;
  assign y173 = n120 ;
  assign y174 = n121 ;
  assign y175 = n122 ;
  assign y176 = n124 ;
  assign y177 = n125 ;
  assign y178 = n126 ;
  assign y179 = n127 ;
  assign y180 = n128 ;
  assign y181 = n129 ;
  assign y182 = n130 ;
  assign y183 = n131 ;
  assign y184 = n132 ;
  assign y185 = n133 ;
  assign y186 = n134 ;
  assign y187 = n135 ;
  assign y188 = n136 ;
  assign y189 = n137 ;
  assign y190 = n138 ;
  assign y191 = n139 ;
  assign y192 = n242 ;
  assign y193 = n237 ;
  assign y194 = n240 ;
  assign y195 = n236 ;
  assign y196 = n235 ;
  assign y197 = n232 ;
  assign y198 = n231 ;
  assign y199 = n234 ;
  assign y200 = n230 ;
  assign y201 = n233 ;
  assign y202 = n228 ;
  assign y203 = n239 ;
  assign y204 = n241 ;
  assign y205 = n243 ;
  assign y206 = n238 ;
  assign y207 = n229 ;
  assign y208 = n142 ;
  assign y209 = n143 ;
  assign y210 = n144 ;
  assign y211 = n145 ;
  assign y212 = n146 ;
  assign y213 = n147 ;
  assign y214 = n148 ;
  assign y215 = n149 ;
  assign y216 = n150 ;
  assign y217 = n151 ;
  assign y218 = n152 ;
  assign y219 = n153 ;
  assign y220 = n154 ;
  assign y221 = n155 ;
  assign y222 = n156 ;
  assign y223 = n157 ;
  assign y224 = n159 ;
  assign y225 = n160 ;
  assign y226 = n161 ;
  assign y227 = n162 ;
  assign y228 = n163 ;
  assign y229 = n164 ;
  assign y230 = n165 ;
  assign y231 = n166 ;
  assign y232 = n167 ;
  assign y233 = n168 ;
  assign y234 = n169 ;
  assign y235 = n170 ;
  assign y236 = n171 ;
  assign y237 = n172 ;
  assign y238 = n173 ;
  assign y239 = n174 ;
  assign y240 = n176 ;
  assign y241 = n177 ;
  assign y242 = n178 ;
  assign y243 = n179 ;
  assign y244 = n180 ;
  assign y245 = n181 ;
  assign y246 = n182 ;
  assign y247 = n183 ;
  assign y248 = n184 ;
  assign y249 = n185 ;
  assign y250 = n186 ;
  assign y251 = n187 ;
  assign y252 = n188 ;
  assign y253 = n189 ;
  assign y254 = n190 ;
  assign y255 = n191 ;
endmodule
