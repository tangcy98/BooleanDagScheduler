module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 ;
  assign n269 = x0 | x2 ;
  assign n270 = x1 | x3 ;
  assign n271 = n269 | n270 ;
  assign n306 = x4 | x5 ;
  assign n313 = ~x6 ;
  assign n311 = n313 & x7 ;
  assign n314 = ~n306 ;
  assign n296 = n314 & n311 ;
  assign n315 = ~n271 ;
  assign n9 = n315 & n296 ;
  assign n316 = ~x2 ;
  assign n272 = x0 & n316 ;
  assign n317 = ~n270 ;
  assign n273 = n317 & n272 ;
  assign n10 = n273 & n296 ;
  assign n318 = ~x3 ;
  assign n274 = x1 & n318 ;
  assign n319 = ~n269 ;
  assign n275 = n319 & n274 ;
  assign n11 = n275 & n296 ;
  assign n276 = n272 & n274 ;
  assign n12 = n276 & n296 ;
  assign n320 = ~x0 ;
  assign n277 = n320 & x2 ;
  assign n278 = n317 & n277 ;
  assign n13 = n278 & n296 ;
  assign n265 = x0 & x2 ;
  assign n280 = n265 & n317 ;
  assign n14 = n280 & n296 ;
  assign n281 = n274 & n277 ;
  assign n15 = n281 & n296 ;
  assign n282 = n265 & n274 ;
  assign n16 = n282 & n296 ;
  assign n321 = ~x1 ;
  assign n283 = n321 & x3 ;
  assign n284 = n319 & n283 ;
  assign n17 = n284 & n296 ;
  assign n285 = n272 & n283 ;
  assign n18 = n285 & n296 ;
  assign n266 = x1 & x3 ;
  assign n286 = n266 & n319 ;
  assign n19 = n286 & n296 ;
  assign n287 = n266 & n272 ;
  assign n20 = n287 & n296 ;
  assign n288 = n277 & n283 ;
  assign n21 = n288 & n296 ;
  assign n289 = n265 & n283 ;
  assign n22 = n289 & n296 ;
  assign n290 = n266 & n277 ;
  assign n23 = n290 & n296 ;
  assign n291 = n265 & n266 ;
  assign n24 = n291 & n296 ;
  assign n322 = ~x5 ;
  assign n292 = x4 & n322 ;
  assign n312 = n292 & n311 ;
  assign n25 = n315 & n312 ;
  assign n26 = n273 & n312 ;
  assign n27 = n275 & n312 ;
  assign n28 = n276 & n312 ;
  assign n29 = n278 & n312 ;
  assign n30 = n280 & n312 ;
  assign n31 = n281 & n312 ;
  assign n32 = n282 & n312 ;
  assign n33 = n284 & n312 ;
  assign n34 = n285 & n312 ;
  assign n35 = n286 & n312 ;
  assign n36 = n287 & n312 ;
  assign n37 = n288 & n312 ;
  assign n38 = n289 & n312 ;
  assign n39 = n290 & n312 ;
  assign n40 = n291 & n312 ;
  assign n323 = ~x4 ;
  assign n293 = n323 & x5 ;
  assign n327 = n293 & n311 ;
  assign n41 = n315 & n327 ;
  assign n42 = n273 & n327 ;
  assign n43 = n275 & n327 ;
  assign n44 = n276 & n327 ;
  assign n45 = n278 & n327 ;
  assign n46 = n280 & n327 ;
  assign n47 = n281 & n327 ;
  assign n48 = n282 & n327 ;
  assign n49 = n284 & n327 ;
  assign n50 = n285 & n327 ;
  assign n51 = n286 & n327 ;
  assign n52 = n287 & n327 ;
  assign n53 = n288 & n327 ;
  assign n54 = n289 & n327 ;
  assign n55 = n290 & n327 ;
  assign n56 = n291 & n327 ;
  assign n267 = x4 & x5 ;
  assign n279 = n267 & n311 ;
  assign n57 = n315 & n279 ;
  assign n58 = n273 & n279 ;
  assign n59 = n275 & n279 ;
  assign n60 = n276 & n279 ;
  assign n61 = n278 & n279 ;
  assign n62 = n280 & n279 ;
  assign n63 = n281 & n279 ;
  assign n64 = n282 & n279 ;
  assign n65 = n284 & n279 ;
  assign n66 = n285 & n279 ;
  assign n67 = n286 & n279 ;
  assign n68 = n287 & n279 ;
  assign n69 = n288 & n279 ;
  assign n70 = n289 & n279 ;
  assign n71 = n290 & n279 ;
  assign n72 = n291 & n279 ;
  assign n268 = x6 & x7 ;
  assign n307 = n268 & n314 ;
  assign n73 = n315 & n307 ;
  assign n74 = n273 & n307 ;
  assign n75 = n275 & n307 ;
  assign n76 = n276 & n307 ;
  assign n77 = n278 & n307 ;
  assign n78 = n280 & n307 ;
  assign n79 = n281 & n307 ;
  assign n80 = n282 & n307 ;
  assign n81 = n284 & n307 ;
  assign n82 = n285 & n307 ;
  assign n83 = n286 & n307 ;
  assign n84 = n287 & n307 ;
  assign n85 = n288 & n307 ;
  assign n86 = n289 & n307 ;
  assign n87 = n290 & n307 ;
  assign n88 = n291 & n307 ;
  assign n294 = n268 & n292 ;
  assign n89 = n315 & n294 ;
  assign n90 = n273 & n294 ;
  assign n91 = n275 & n294 ;
  assign n92 = n276 & n294 ;
  assign n93 = n278 & n294 ;
  assign n94 = n280 & n294 ;
  assign n95 = n281 & n294 ;
  assign n96 = n282 & n294 ;
  assign n97 = n284 & n294 ;
  assign n98 = n285 & n294 ;
  assign n99 = n286 & n294 ;
  assign n100 = n287 & n294 ;
  assign n101 = n288 & n294 ;
  assign n102 = n289 & n294 ;
  assign n103 = n290 & n294 ;
  assign n104 = n291 & n294 ;
  assign n295 = n268 & n293 ;
  assign n105 = n315 & n295 ;
  assign n106 = n273 & n295 ;
  assign n107 = n275 & n295 ;
  assign n108 = n276 & n295 ;
  assign n109 = n278 & n295 ;
  assign n110 = n280 & n295 ;
  assign n111 = n281 & n295 ;
  assign n112 = n282 & n295 ;
  assign n113 = n284 & n295 ;
  assign n114 = n285 & n295 ;
  assign n115 = n286 & n295 ;
  assign n116 = n287 & n295 ;
  assign n117 = n288 & n295 ;
  assign n118 = n289 & n295 ;
  assign n119 = n290 & n295 ;
  assign n120 = n291 & n295 ;
  assign n297 = n267 & n268 ;
  assign n121 = n315 & n297 ;
  assign n122 = n273 & n297 ;
  assign n123 = n275 & n297 ;
  assign n124 = n276 & n297 ;
  assign n125 = n278 & n297 ;
  assign n126 = n280 & n297 ;
  assign n127 = n281 & n297 ;
  assign n128 = n282 & n297 ;
  assign n129 = n284 & n297 ;
  assign n130 = n285 & n297 ;
  assign n131 = n286 & n297 ;
  assign n132 = n287 & n297 ;
  assign n133 = n288 & n297 ;
  assign n134 = n289 & n297 ;
  assign n135 = n290 & n297 ;
  assign n136 = n291 & n297 ;
  assign n298 = x6 | x7 ;
  assign n308 = n298 | n306 ;
  assign n309 = n271 | n308 ;
  assign n324 = ~n308 ;
  assign n138 = n273 & n324 ;
  assign n139 = n275 & n324 ;
  assign n140 = n276 & n324 ;
  assign n141 = n278 & n324 ;
  assign n142 = n280 & n324 ;
  assign n143 = n281 & n324 ;
  assign n144 = n282 & n324 ;
  assign n145 = n284 & n324 ;
  assign n146 = n285 & n324 ;
  assign n147 = n286 & n324 ;
  assign n148 = n287 & n324 ;
  assign n149 = n288 & n324 ;
  assign n150 = n289 & n324 ;
  assign n151 = n290 & n324 ;
  assign n152 = n291 & n324 ;
  assign n325 = ~n298 ;
  assign n299 = n292 & n325 ;
  assign n153 = n315 & n299 ;
  assign n154 = n273 & n299 ;
  assign n155 = n275 & n299 ;
  assign n156 = n276 & n299 ;
  assign n157 = n278 & n299 ;
  assign n158 = n280 & n299 ;
  assign n159 = n281 & n299 ;
  assign n160 = n282 & n299 ;
  assign n161 = n284 & n299 ;
  assign n162 = n285 & n299 ;
  assign n163 = n286 & n299 ;
  assign n164 = n287 & n299 ;
  assign n165 = n288 & n299 ;
  assign n166 = n289 & n299 ;
  assign n167 = n290 & n299 ;
  assign n168 = n291 & n299 ;
  assign n300 = n293 & n325 ;
  assign n169 = n315 & n300 ;
  assign n170 = n273 & n300 ;
  assign n171 = n275 & n300 ;
  assign n172 = n276 & n300 ;
  assign n173 = n278 & n300 ;
  assign n174 = n280 & n300 ;
  assign n175 = n281 & n300 ;
  assign n176 = n282 & n300 ;
  assign n177 = n284 & n300 ;
  assign n178 = n285 & n300 ;
  assign n179 = n286 & n300 ;
  assign n180 = n287 & n300 ;
  assign n181 = n288 & n300 ;
  assign n182 = n289 & n300 ;
  assign n183 = n290 & n300 ;
  assign n184 = n291 & n300 ;
  assign n301 = n267 & n325 ;
  assign n185 = n315 & n301 ;
  assign n186 = n273 & n301 ;
  assign n187 = n275 & n301 ;
  assign n188 = n276 & n301 ;
  assign n189 = n278 & n301 ;
  assign n190 = n280 & n301 ;
  assign n191 = n281 & n301 ;
  assign n192 = n282 & n301 ;
  assign n193 = n284 & n301 ;
  assign n194 = n285 & n301 ;
  assign n195 = n286 & n301 ;
  assign n196 = n287 & n301 ;
  assign n197 = n288 & n301 ;
  assign n198 = n289 & n301 ;
  assign n199 = n290 & n301 ;
  assign n200 = n291 & n301 ;
  assign n326 = ~x7 ;
  assign n302 = x6 & n326 ;
  assign n310 = n302 & n314 ;
  assign n201 = n315 & n310 ;
  assign n202 = n273 & n310 ;
  assign n203 = n275 & n310 ;
  assign n204 = n276 & n310 ;
  assign n205 = n278 & n310 ;
  assign n206 = n280 & n310 ;
  assign n207 = n281 & n310 ;
  assign n208 = n282 & n310 ;
  assign n209 = n284 & n310 ;
  assign n210 = n285 & n310 ;
  assign n211 = n286 & n310 ;
  assign n212 = n287 & n310 ;
  assign n213 = n288 & n310 ;
  assign n214 = n289 & n310 ;
  assign n215 = n290 & n310 ;
  assign n216 = n291 & n310 ;
  assign n303 = n292 & n302 ;
  assign n217 = n315 & n303 ;
  assign n218 = n273 & n303 ;
  assign n219 = n275 & n303 ;
  assign n220 = n276 & n303 ;
  assign n221 = n278 & n303 ;
  assign n222 = n280 & n303 ;
  assign n223 = n281 & n303 ;
  assign n224 = n282 & n303 ;
  assign n225 = n284 & n303 ;
  assign n226 = n285 & n303 ;
  assign n227 = n286 & n303 ;
  assign n228 = n287 & n303 ;
  assign n229 = n288 & n303 ;
  assign n230 = n289 & n303 ;
  assign n231 = n290 & n303 ;
  assign n232 = n291 & n303 ;
  assign n304 = n293 & n302 ;
  assign n233 = n315 & n304 ;
  assign n234 = n273 & n304 ;
  assign n235 = n275 & n304 ;
  assign n236 = n276 & n304 ;
  assign n237 = n278 & n304 ;
  assign n238 = n280 & n304 ;
  assign n239 = n281 & n304 ;
  assign n240 = n282 & n304 ;
  assign n241 = n284 & n304 ;
  assign n242 = n285 & n304 ;
  assign n243 = n286 & n304 ;
  assign n244 = n287 & n304 ;
  assign n245 = n288 & n304 ;
  assign n246 = n289 & n304 ;
  assign n247 = n290 & n304 ;
  assign n248 = n291 & n304 ;
  assign n305 = n267 & n302 ;
  assign n249 = n315 & n305 ;
  assign n250 = n273 & n305 ;
  assign n251 = n275 & n305 ;
  assign n252 = n276 & n305 ;
  assign n253 = n278 & n305 ;
  assign n254 = n280 & n305 ;
  assign n255 = n281 & n305 ;
  assign n256 = n282 & n305 ;
  assign n257 = n284 & n305 ;
  assign n258 = n285 & n305 ;
  assign n259 = n286 & n305 ;
  assign n260 = n287 & n305 ;
  assign n261 = n288 & n305 ;
  assign n262 = n289 & n305 ;
  assign n263 = n290 & n305 ;
  assign n264 = n291 & n305 ;
  assign n137 = ~n309 ;
  assign y0 = n9 ;
  assign y1 = n10 ;
  assign y2 = n11 ;
  assign y3 = n12 ;
  assign y4 = n13 ;
  assign y5 = n14 ;
  assign y6 = n15 ;
  assign y7 = n16 ;
  assign y8 = n17 ;
  assign y9 = n18 ;
  assign y10 = n19 ;
  assign y11 = n20 ;
  assign y12 = n21 ;
  assign y13 = n22 ;
  assign y14 = n23 ;
  assign y15 = n24 ;
  assign y16 = n25 ;
  assign y17 = n26 ;
  assign y18 = n27 ;
  assign y19 = n28 ;
  assign y20 = n29 ;
  assign y21 = n30 ;
  assign y22 = n31 ;
  assign y23 = n32 ;
  assign y24 = n33 ;
  assign y25 = n34 ;
  assign y26 = n35 ;
  assign y27 = n36 ;
  assign y28 = n37 ;
  assign y29 = n38 ;
  assign y30 = n39 ;
  assign y31 = n40 ;
  assign y32 = n41 ;
  assign y33 = n42 ;
  assign y34 = n43 ;
  assign y35 = n44 ;
  assign y36 = n45 ;
  assign y37 = n46 ;
  assign y38 = n47 ;
  assign y39 = n48 ;
  assign y40 = n49 ;
  assign y41 = n50 ;
  assign y42 = n51 ;
  assign y43 = n52 ;
  assign y44 = n53 ;
  assign y45 = n54 ;
  assign y46 = n55 ;
  assign y47 = n56 ;
  assign y48 = n57 ;
  assign y49 = n58 ;
  assign y50 = n59 ;
  assign y51 = n60 ;
  assign y52 = n61 ;
  assign y53 = n62 ;
  assign y54 = n63 ;
  assign y55 = n64 ;
  assign y56 = n65 ;
  assign y57 = n66 ;
  assign y58 = n67 ;
  assign y59 = n68 ;
  assign y60 = n69 ;
  assign y61 = n70 ;
  assign y62 = n71 ;
  assign y63 = n72 ;
  assign y64 = n73 ;
  assign y65 = n74 ;
  assign y66 = n75 ;
  assign y67 = n76 ;
  assign y68 = n77 ;
  assign y69 = n78 ;
  assign y70 = n79 ;
  assign y71 = n80 ;
  assign y72 = n81 ;
  assign y73 = n82 ;
  assign y74 = n83 ;
  assign y75 = n84 ;
  assign y76 = n85 ;
  assign y77 = n86 ;
  assign y78 = n87 ;
  assign y79 = n88 ;
  assign y80 = n89 ;
  assign y81 = n90 ;
  assign y82 = n91 ;
  assign y83 = n92 ;
  assign y84 = n93 ;
  assign y85 = n94 ;
  assign y86 = n95 ;
  assign y87 = n96 ;
  assign y88 = n97 ;
  assign y89 = n98 ;
  assign y90 = n99 ;
  assign y91 = n100 ;
  assign y92 = n101 ;
  assign y93 = n102 ;
  assign y94 = n103 ;
  assign y95 = n104 ;
  assign y96 = n105 ;
  assign y97 = n106 ;
  assign y98 = n107 ;
  assign y99 = n108 ;
  assign y100 = n109 ;
  assign y101 = n110 ;
  assign y102 = n111 ;
  assign y103 = n112 ;
  assign y104 = n113 ;
  assign y105 = n114 ;
  assign y106 = n115 ;
  assign y107 = n116 ;
  assign y108 = n117 ;
  assign y109 = n118 ;
  assign y110 = n119 ;
  assign y111 = n120 ;
  assign y112 = n121 ;
  assign y113 = n122 ;
  assign y114 = n123 ;
  assign y115 = n124 ;
  assign y116 = n125 ;
  assign y117 = n126 ;
  assign y118 = n127 ;
  assign y119 = n128 ;
  assign y120 = n129 ;
  assign y121 = n130 ;
  assign y122 = n131 ;
  assign y123 = n132 ;
  assign y124 = n133 ;
  assign y125 = n134 ;
  assign y126 = n135 ;
  assign y127 = n136 ;
  assign y128 = n137 ;
  assign y129 = n138 ;
  assign y130 = n139 ;
  assign y131 = n140 ;
  assign y132 = n141 ;
  assign y133 = n142 ;
  assign y134 = n143 ;
  assign y135 = n144 ;
  assign y136 = n145 ;
  assign y137 = n146 ;
  assign y138 = n147 ;
  assign y139 = n148 ;
  assign y140 = n149 ;
  assign y141 = n150 ;
  assign y142 = n151 ;
  assign y143 = n152 ;
  assign y144 = n153 ;
  assign y145 = n154 ;
  assign y146 = n155 ;
  assign y147 = n156 ;
  assign y148 = n157 ;
  assign y149 = n158 ;
  assign y150 = n159 ;
  assign y151 = n160 ;
  assign y152 = n161 ;
  assign y153 = n162 ;
  assign y154 = n163 ;
  assign y155 = n164 ;
  assign y156 = n165 ;
  assign y157 = n166 ;
  assign y158 = n167 ;
  assign y159 = n168 ;
  assign y160 = n169 ;
  assign y161 = n170 ;
  assign y162 = n171 ;
  assign y163 = n172 ;
  assign y164 = n173 ;
  assign y165 = n174 ;
  assign y166 = n175 ;
  assign y167 = n176 ;
  assign y168 = n177 ;
  assign y169 = n178 ;
  assign y170 = n179 ;
  assign y171 = n180 ;
  assign y172 = n181 ;
  assign y173 = n182 ;
  assign y174 = n183 ;
  assign y175 = n184 ;
  assign y176 = n185 ;
  assign y177 = n186 ;
  assign y178 = n187 ;
  assign y179 = n188 ;
  assign y180 = n189 ;
  assign y181 = n190 ;
  assign y182 = n191 ;
  assign y183 = n192 ;
  assign y184 = n193 ;
  assign y185 = n194 ;
  assign y186 = n195 ;
  assign y187 = n196 ;
  assign y188 = n197 ;
  assign y189 = n198 ;
  assign y190 = n199 ;
  assign y191 = n200 ;
  assign y192 = n201 ;
  assign y193 = n202 ;
  assign y194 = n203 ;
  assign y195 = n204 ;
  assign y196 = n205 ;
  assign y197 = n206 ;
  assign y198 = n207 ;
  assign y199 = n208 ;
  assign y200 = n209 ;
  assign y201 = n210 ;
  assign y202 = n211 ;
  assign y203 = n212 ;
  assign y204 = n213 ;
  assign y205 = n214 ;
  assign y206 = n215 ;
  assign y207 = n216 ;
  assign y208 = n217 ;
  assign y209 = n218 ;
  assign y210 = n219 ;
  assign y211 = n220 ;
  assign y212 = n221 ;
  assign y213 = n222 ;
  assign y214 = n223 ;
  assign y215 = n224 ;
  assign y216 = n225 ;
  assign y217 = n226 ;
  assign y218 = n227 ;
  assign y219 = n228 ;
  assign y220 = n229 ;
  assign y221 = n230 ;
  assign y222 = n231 ;
  assign y223 = n232 ;
  assign y224 = n233 ;
  assign y225 = n234 ;
  assign y226 = n235 ;
  assign y227 = n236 ;
  assign y228 = n237 ;
  assign y229 = n238 ;
  assign y230 = n239 ;
  assign y231 = n240 ;
  assign y232 = n241 ;
  assign y233 = n242 ;
  assign y234 = n243 ;
  assign y235 = n244 ;
  assign y236 = n245 ;
  assign y237 = n246 ;
  assign y238 = n247 ;
  assign y239 = n248 ;
  assign y240 = n249 ;
  assign y241 = n250 ;
  assign y242 = n251 ;
  assign y243 = n252 ;
  assign y244 = n253 ;
  assign y245 = n254 ;
  assign y246 = n255 ;
  assign y247 = n256 ;
  assign y248 = n257 ;
  assign y249 = n258 ;
  assign y250 = n259 ;
  assign y251 = n260 ;
  assign y252 = n261 ;
  assign y253 = n262 ;
  assign y254 = n263 ;
  assign y255 = n264 ;
endmodule
