module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 ;
  assign n50 = x3 | x5 ;
  assign n709 = ~x0 ;
  assign n51 = n709 & x9 ;
  assign n710 = ~n51 ;
  assign n52 = x1 & n710 ;
  assign n711 = ~x1 ;
  assign n53 = n711 & x9 ;
  assign n54 = n52 | n53 ;
  assign n59 = n50 | n54 ;
  assign n712 = ~x9 ;
  assign n55 = x0 & n712 ;
  assign n56 = x1 | n55 ;
  assign n57 = x1 & n712 ;
  assign n58 = x7 | n57 ;
  assign n713 = ~n58 ;
  assign n60 = n56 & n713 ;
  assign n714 = ~n60 ;
  assign n61 = n59 & n714 ;
  assign n62 = x2 | n61 ;
  assign n23 = x1 & x3 ;
  assign n22 = x0 & x3 ;
  assign n66 = x2 | x3 ;
  assign n68 = x9 & n66 ;
  assign n69 = n22 | n68 ;
  assign n71 = x1 | n69 ;
  assign n715 = ~n23 ;
  assign n72 = n715 & n71 ;
  assign n11 = x1 & x2 ;
  assign n63 = x2 | x5 ;
  assign n64 = n709 & n63 ;
  assign n65 = n11 | n64 ;
  assign n73 = n712 & n65 ;
  assign n74 = n72 | n73 ;
  assign n716 = ~x7 ;
  assign n75 = n716 & n74 ;
  assign n717 = ~n75 ;
  assign n76 = n62 & n717 ;
  assign n93 = x8 | n76 ;
  assign n79 = x5 | x9 ;
  assign n81 = x1 & n716 ;
  assign n82 = n79 | n81 ;
  assign n25 = n716 & x9 ;
  assign n24 = x7 & x8 ;
  assign n718 = ~x5 ;
  assign n77 = n718 & n24 ;
  assign n78 = n25 | n77 ;
  assign n83 = x1 & n78 ;
  assign n719 = ~n83 ;
  assign n84 = n82 & n719 ;
  assign n720 = ~x2 ;
  assign n85 = x0 & n720 ;
  assign n721 = ~n84 ;
  assign n86 = n721 & n85 ;
  assign n87 = x2 & n712 ;
  assign n89 = x0 | x1 ;
  assign n722 = ~n89 ;
  assign n90 = n87 & n722 ;
  assign n91 = n77 & n90 ;
  assign n92 = n86 | n91 ;
  assign n723 = ~x3 ;
  assign n94 = n723 & n92 ;
  assign n724 = ~n94 ;
  assign n95 = n93 & n724 ;
  assign n96 = x6 | n95 ;
  assign n26 = x0 & x9 ;
  assign n100 = x0 | x9 ;
  assign n725 = ~n26 ;
  assign n101 = n725 & n100 ;
  assign n726 = ~n101 ;
  assign n103 = x1 & n726 ;
  assign n727 = ~n66 ;
  assign n105 = n727 & n103 ;
  assign n117 = x2 | n55 ;
  assign n118 = x6 & n117 ;
  assign n119 = n105 | n118 ;
  assign n124 = x5 & n119 ;
  assign n121 = x0 | x3 ;
  assign n12 = x2 & x9 ;
  assign n120 = n720 & n57 ;
  assign n122 = n12 | n120 ;
  assign n728 = ~n121 ;
  assign n123 = n728 & n122 ;
  assign n125 = x6 & n123 ;
  assign n126 = n124 | n125 ;
  assign n127 = x8 & n126 ;
  assign n128 = x2 & n723 ;
  assign n130 = n53 & n128 ;
  assign n729 = ~x8 ;
  assign n131 = x1 & n729 ;
  assign n132 = n130 | n131 ;
  assign n133 = n709 & n132 ;
  assign n134 = x1 | x9 ;
  assign n27 = n720 & x6 ;
  assign n730 = ~n27 ;
  assign n135 = x3 & n730 ;
  assign n136 = n134 | n135 ;
  assign n731 = ~n12 ;
  assign n137 = n731 & n136 ;
  assign n138 = x8 | n137 ;
  assign n732 = ~n133 ;
  assign n139 = n732 & n138 ;
  assign n141 = x5 | n139 ;
  assign n67 = x0 | n66 ;
  assign n140 = x8 | n134 ;
  assign n142 = n67 | n140 ;
  assign n143 = n141 & n142 ;
  assign n733 = ~n127 ;
  assign n144 = n733 & n143 ;
  assign n97 = x0 | x2 ;
  assign n734 = ~n97 ;
  assign n98 = n53 & n734 ;
  assign n99 = x5 | n98 ;
  assign n106 = x6 & n99 ;
  assign n104 = x2 & n103 ;
  assign n107 = x5 & n104 ;
  assign n108 = n106 | n107 ;
  assign n109 = x8 & n108 ;
  assign n110 = x1 | n51 ;
  assign n111 = n729 & n110 ;
  assign n112 = n711 & x2 ;
  assign n113 = n55 & n112 ;
  assign n114 = n111 | n113 ;
  assign n115 = n718 & n114 ;
  assign n116 = n109 | n115 ;
  assign n145 = x3 & n116 ;
  assign n735 = ~n145 ;
  assign n146 = n144 & n735 ;
  assign n147 = x7 | n146 ;
  assign n148 = n96 & n147 ;
  assign n164 = x4 | n148 ;
  assign n13 = x4 & x8 ;
  assign n28 = x6 & n13 ;
  assign n149 = x8 | x9 ;
  assign n151 = x6 | n149 ;
  assign n736 = ~n28 ;
  assign n152 = n736 & n151 ;
  assign n737 = ~n152 ;
  assign n153 = x5 & n737 ;
  assign n14 = x5 & x6 ;
  assign n29 = x4 & x9 ;
  assign n154 = x6 & n712 ;
  assign n155 = n29 | n154 ;
  assign n738 = ~n14 ;
  assign n156 = n738 & n155 ;
  assign n157 = n729 & n156 ;
  assign n158 = n153 | n157 ;
  assign n159 = n716 & n158 ;
  assign n160 = x1 | x3 ;
  assign n161 = x2 | n160 ;
  assign n739 = ~n161 ;
  assign n163 = n159 & n739 ;
  assign n165 = n709 & n163 ;
  assign n740 = ~n165 ;
  assign n166 = n164 & n740 ;
  assign n15 = x0 & x8 ;
  assign n30 = n12 & n15 ;
  assign n167 = x2 | x8 ;
  assign n168 = n100 | n167 ;
  assign n741 = ~n30 ;
  assign n169 = n741 & n168 ;
  assign n742 = ~n169 ;
  assign n175 = x5 & n742 ;
  assign n16 = x6 & x9 ;
  assign n170 = n718 & x8 ;
  assign n171 = n16 | n170 ;
  assign n172 = n709 & n171 ;
  assign n31 = x8 & n16 ;
  assign n80 = x8 | n79 ;
  assign n743 = ~n31 ;
  assign n173 = n743 & n80 ;
  assign n744 = ~n172 ;
  assign n174 = n744 & n173 ;
  assign n745 = ~n174 ;
  assign n176 = x2 & n745 ;
  assign n177 = n175 | n176 ;
  assign n746 = ~x4 ;
  assign n178 = n746 & n177 ;
  assign n747 = ~x6 ;
  assign n179 = n747 & x9 ;
  assign n180 = x5 & n729 ;
  assign n181 = n13 | n180 ;
  assign n182 = n747 & n181 ;
  assign n183 = n29 | n182 ;
  assign n748 = ~n179 ;
  assign n184 = n748 & n183 ;
  assign n185 = n734 & n184 ;
  assign n186 = n178 | n185 ;
  assign n206 = n711 & n186 ;
  assign n17 = x6 & x8 ;
  assign n749 = ~n17 ;
  assign n187 = n749 & n171 ;
  assign n188 = x0 & n187 ;
  assign n189 = n709 & x5 ;
  assign n190 = n729 & x9 ;
  assign n191 = n189 & n190 ;
  assign n193 = n188 | n191 ;
  assign n199 = n720 & n193 ;
  assign n194 = x6 | x8 ;
  assign n195 = n709 & x6 ;
  assign n196 = x2 | n195 ;
  assign n197 = n170 & n196 ;
  assign n750 = ~n197 ;
  assign n198 = n194 & n750 ;
  assign n200 = x9 | n198 ;
  assign n751 = ~n199 ;
  assign n201 = n751 & n200 ;
  assign n752 = ~n201 ;
  assign n202 = x1 & n752 ;
  assign n203 = n747 & x8 ;
  assign n204 = n87 & n203 ;
  assign n205 = n202 | n204 ;
  assign n207 = n746 & n205 ;
  assign n208 = n206 | n207 ;
  assign n209 = n723 & n208 ;
  assign n35 = x3 & n11 ;
  assign n254 = n35 & n180 ;
  assign n47 = x1 & x5 ;
  assign n211 = x3 & n729 ;
  assign n247 = x1 | x2 ;
  assign n753 = ~n247 ;
  assign n248 = n211 & n753 ;
  assign n249 = n47 | n248 ;
  assign n250 = x0 & n249 ;
  assign n251 = x5 & n66 ;
  assign n252 = n35 | n251 ;
  assign n253 = n250 | n252 ;
  assign n255 = x6 & n253 ;
  assign n256 = n254 | n255 ;
  assign n257 = x9 & n256 ;
  assign n754 = ~n167 ;
  assign n210 = x5 & n754 ;
  assign n32 = x5 & x8 ;
  assign n212 = n32 | n211 ;
  assign n214 = x0 & n212 ;
  assign n215 = n210 | n214 ;
  assign n216 = n711 & n215 ;
  assign n33 = x3 & x8 ;
  assign n217 = x2 | n33 ;
  assign n225 = n709 & n217 ;
  assign n218 = n720 & x8 ;
  assign n220 = x0 & n218 ;
  assign n222 = x0 & n718 ;
  assign n223 = n189 | n222 ;
  assign n224 = n220 | n223 ;
  assign n226 = x1 & n224 ;
  assign n227 = n225 | n226 ;
  assign n228 = n216 | n227 ;
  assign n243 = n747 & n228 ;
  assign n229 = n711 & x6 ;
  assign n755 = ~n229 ;
  assign n230 = x2 & n755 ;
  assign n231 = x1 | x8 ;
  assign n756 = ~n230 ;
  assign n233 = n756 & n231 ;
  assign n234 = x3 & n233 ;
  assign n235 = n709 & x8 ;
  assign n34 = x0 & x1 ;
  assign n236 = x1 | x6 ;
  assign n757 = ~n34 ;
  assign n239 = n757 & n236 ;
  assign n758 = ~n235 ;
  assign n240 = n758 & n239 ;
  assign n241 = n720 & n240 ;
  assign n242 = n234 | n241 ;
  assign n244 = n718 & n242 ;
  assign n245 = n243 | n244 ;
  assign n258 = n712 & n245 ;
  assign n259 = n257 | n258 ;
  assign n260 = n746 & n259 ;
  assign n261 = n209 | n260 ;
  assign n270 = n716 & n261 ;
  assign n221 = n57 & n218 ;
  assign n238 = n34 | n117 ;
  assign n262 = x2 & n89 ;
  assign n759 = ~n262 ;
  assign n263 = n238 & n759 ;
  assign n264 = n729 & n263 ;
  assign n265 = n221 | n264 ;
  assign n266 = x7 & n265 ;
  assign n267 = n90 | n266 ;
  assign n268 = n746 & n267 ;
  assign n269 = n747 & n268 ;
  assign n760 = ~n50 ;
  assign n271 = n760 & n269 ;
  assign n272 = n270 | n271 ;
  assign n36 = n723 & x9 ;
  assign n273 = x1 & n723 ;
  assign n274 = n190 | n273 ;
  assign n761 = ~n36 ;
  assign n276 = n761 & n274 ;
  assign n277 = n747 & n276 ;
  assign n762 = ~n203 ;
  assign n291 = x2 & n762 ;
  assign n292 = n711 & n217 ;
  assign n293 = n291 | n292 ;
  assign n294 = x5 & n293 ;
  assign n192 = n711 & n190 ;
  assign n18 = x1 & x8 ;
  assign n763 = ~n18 ;
  assign n295 = x6 & n763 ;
  assign n296 = x9 | n295 ;
  assign n297 = n720 & n296 ;
  assign n298 = n192 | n297 ;
  assign n301 = x3 & n298 ;
  assign n299 = x6 & n729 ;
  assign n300 = x1 & n36 ;
  assign n302 = n299 & n300 ;
  assign n303 = n301 | n302 ;
  assign n304 = n294 | n303 ;
  assign n764 = ~n218 ;
  assign n278 = x3 & n764 ;
  assign n765 = ~n278 ;
  assign n282 = x5 & n765 ;
  assign n279 = x2 & n718 ;
  assign n766 = ~n279 ;
  assign n281 = x3 & n766 ;
  assign n767 = ~n281 ;
  assign n283 = x8 & n767 ;
  assign n284 = n282 | n283 ;
  assign n285 = x1 & n284 ;
  assign n286 = n718 & x6 ;
  assign n288 = n729 & n286 ;
  assign n768 = ~n160 ;
  assign n289 = n768 & n288 ;
  assign n290 = n285 | n289 ;
  assign n305 = n712 & n290 ;
  assign n306 = n304 | n305 ;
  assign n307 = n277 | n306 ;
  assign n314 = n746 & n307 ;
  assign n310 = n723 & x4 ;
  assign n311 = n711 & n310 ;
  assign n308 = x8 & n712 ;
  assign n769 = ~n308 ;
  assign n309 = n194 & n769 ;
  assign n312 = n718 & n309 ;
  assign n770 = ~n312 ;
  assign n313 = n311 & n770 ;
  assign n315 = n720 & n313 ;
  assign n316 = n314 | n315 ;
  assign n317 = n709 & n316 ;
  assign n102 = x8 & n725 ;
  assign n318 = n102 | n190 ;
  assign n319 = x5 & n318 ;
  assign n320 = x5 | n12 ;
  assign n771 = ~n319 ;
  assign n321 = n771 & n320 ;
  assign n324 = x1 & n321 ;
  assign n322 = n190 | n308 ;
  assign n772 = ~n322 ;
  assign n323 = n134 & n772 ;
  assign n773 = ~n323 ;
  assign n325 = x2 & n773 ;
  assign n326 = n324 | n325 ;
  assign n327 = n723 & n326 ;
  assign n328 = n711 & x3 ;
  assign n774 = ~n328 ;
  assign n329 = x5 & n774 ;
  assign n330 = x2 | n149 ;
  assign n331 = n329 | n330 ;
  assign n37 = n711 & x8 ;
  assign n332 = n37 & n68 ;
  assign n775 = ~n332 ;
  assign n333 = n331 & n775 ;
  assign n776 = ~n333 ;
  assign n334 = x0 & n776 ;
  assign n335 = n327 | n334 ;
  assign n350 = n747 & n335 ;
  assign n777 = ~n87 ;
  assign n88 = x8 & n777 ;
  assign n778 = ~n149 ;
  assign n150 = x2 & n778 ;
  assign n337 = n88 | n150 ;
  assign n19 = x1 & x9 ;
  assign n38 = x2 & n19 ;
  assign n336 = n37 | n38 ;
  assign n338 = x6 & n336 ;
  assign n339 = n337 | n338 ;
  assign n340 = x3 & n339 ;
  assign n343 = x3 | x8 ;
  assign n779 = ~n19 ;
  assign n344 = n779 & n134 ;
  assign n345 = n343 | n344 ;
  assign n780 = ~n53 ;
  assign n341 = x6 & n780 ;
  assign n342 = n57 | n341 ;
  assign n346 = x8 & n342 ;
  assign n781 = ~n346 ;
  assign n347 = n345 & n781 ;
  assign n348 = x2 | n347 ;
  assign n782 = ~n340 ;
  assign n349 = n782 & n348 ;
  assign n783 = ~n349 ;
  assign n351 = n222 & n783 ;
  assign n352 = n350 | n351 ;
  assign n353 = n746 & n352 ;
  assign n354 = n317 | n353 ;
  assign n363 = n716 & n354 ;
  assign n355 = x5 | x6 ;
  assign n784 = ~n231 ;
  assign n232 = n55 & n784 ;
  assign n357 = n24 & n26 ;
  assign n785 = ~n357 ;
  assign n358 = n100 & n785 ;
  assign n786 = ~n358 ;
  assign n359 = x1 & n786 ;
  assign n360 = n232 | n359 ;
  assign n361 = n746 & n360 ;
  assign n362 = n727 & n361 ;
  assign n787 = ~n355 ;
  assign n364 = n787 & n362 ;
  assign n365 = n363 | n364 ;
  assign n366 = x2 & x6 ;
  assign n367 = x3 & n748 ;
  assign n368 = n366 | n367 ;
  assign n369 = n746 & n368 ;
  assign n20 = x8 & x9 ;
  assign n356 = n20 & n787 ;
  assign n370 = n14 | n356 ;
  assign n371 = n720 & n310 ;
  assign n372 = n370 & n371 ;
  assign n373 = n369 | n372 ;
  assign n374 = n711 & n373 ;
  assign n375 = n32 & n179 ;
  assign n788 = ~n375 ;
  assign n376 = n80 & n788 ;
  assign n789 = ~n376 ;
  assign n377 = x2 & n789 ;
  assign n378 = x5 & n762 ;
  assign n790 = ~n378 ;
  assign n379 = x3 & n790 ;
  assign n380 = n288 | n379 ;
  assign n381 = n377 | n380 ;
  assign n382 = x1 & n381 ;
  assign n383 = x2 & n286 ;
  assign n384 = n382 | n383 ;
  assign n385 = n746 & n384 ;
  assign n386 = n374 | n385 ;
  assign n387 = n709 & n386 ;
  assign n213 = x2 & n212 ;
  assign n388 = x2 | n32 ;
  assign n791 = ~n213 ;
  assign n389 = n791 & n388 ;
  assign n390 = n712 & n389 ;
  assign n39 = x5 & x9 ;
  assign n392 = n729 & n39 ;
  assign n393 = x3 | n392 ;
  assign n394 = n720 & n393 ;
  assign n246 = x6 | n211 ;
  assign n395 = x3 & n718 ;
  assign n792 = ~n395 ;
  assign n396 = n246 & n792 ;
  assign n397 = n394 | n396 ;
  assign n398 = n390 | n397 ;
  assign n399 = x1 & n398 ;
  assign n793 = ~n236 ;
  assign n237 = n210 & n793 ;
  assign n287 = n723 & n286 ;
  assign n400 = n237 | n287 ;
  assign n401 = n712 & n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = x0 & n402 ;
  assign n413 = n79 & n194 ;
  assign n414 = x2 | n413 ;
  assign n415 = x6 | n39 ;
  assign n416 = n19 | n32 ;
  assign n794 = ~n415 ;
  assign n417 = n794 & n416 ;
  assign n795 = ~n417 ;
  assign n418 = n414 & n795 ;
  assign n796 = ~n418 ;
  assign n419 = x3 & n796 ;
  assign n420 = x1 & n308 ;
  assign n421 = n286 & n420 ;
  assign n422 = n419 | n421 ;
  assign n404 = x3 & n747 ;
  assign n405 = x2 & n404 ;
  assign n406 = n66 & n286 ;
  assign n407 = n405 | n406 ;
  assign n408 = x9 & n407 ;
  assign n409 = n712 & n286 ;
  assign n410 = n404 | n409 ;
  assign n411 = n729 & n410 ;
  assign n412 = n408 | n411 ;
  assign n423 = n711 & n412 ;
  assign n424 = n422 | n423 ;
  assign n425 = n403 | n424 ;
  assign n426 = n746 & n425 ;
  assign n427 = n387 | n426 ;
  assign n428 = n716 & n427 ;
  assign n429 = n746 & n262 ;
  assign n430 = x3 & n746 ;
  assign n431 = n310 | n430 ;
  assign n432 = x0 | n247 ;
  assign n797 = ~n432 ;
  assign n433 = n431 & n797 ;
  assign n434 = n429 | n433 ;
  assign n435 = n716 & n434 ;
  assign n436 = n14 & n435 ;
  assign n437 = n722 & n371 ;
  assign n438 = n430 & n432 ;
  assign n439 = n437 | n438 ;
  assign n440 = n716 & n439 ;
  assign n441 = n14 & n440 ;
  assign n40 = x5 & n19 ;
  assign n442 = x1 | x5 ;
  assign n443 = x2 & n442 ;
  assign n444 = x9 | n443 ;
  assign n445 = x6 | n444 ;
  assign n798 = ~n40 ;
  assign n446 = n798 & n445 ;
  assign n799 = ~n446 ;
  assign n448 = x0 & n799 ;
  assign n447 = n709 & n79 ;
  assign n449 = x2 & n447 ;
  assign n450 = n448 | n449 ;
  assign n451 = x8 & n450 ;
  assign n452 = x2 & n51 ;
  assign n800 = ~n452 ;
  assign n453 = n140 & n800 ;
  assign n801 = ~n453 ;
  assign n454 = x5 & n801 ;
  assign n455 = n451 | n454 ;
  assign n802 = ~n20 ;
  assign n456 = n802 & n149 ;
  assign n803 = ~n456 ;
  assign n457 = x6 & n803 ;
  assign n459 = x2 | x9 ;
  assign n460 = n731 & n459 ;
  assign n804 = ~n460 ;
  assign n461 = n457 & n804 ;
  assign n463 = n455 | n461 ;
  assign n464 = n716 & n463 ;
  assign n465 = x7 & n712 ;
  assign n805 = ~n465 ;
  assign n466 = x8 & n805 ;
  assign n806 = ~n466 ;
  assign n467 = n112 & n806 ;
  assign n468 = n120 | n467 ;
  assign n471 = n709 & n468 ;
  assign n41 = n15 & n19 ;
  assign n807 = ~n41 ;
  assign n469 = n807 & n149 ;
  assign n808 = ~n469 ;
  assign n470 = x7 & n808 ;
  assign n472 = n720 & n470 ;
  assign n473 = n471 | n472 ;
  assign n474 = n787 & n473 ;
  assign n475 = n464 | n474 ;
  assign n516 = n723 & n475 ;
  assign n486 = n729 & n34 ;
  assign n42 = x0 & n17 ;
  assign n485 = n42 | n131 ;
  assign n487 = n720 & n485 ;
  assign n488 = n486 | n487 ;
  assign n489 = x9 & n488 ;
  assign n43 = x0 & x5 ;
  assign n490 = n43 | n235 ;
  assign n491 = n57 & n490 ;
  assign n492 = n489 | n491 ;
  assign n477 = x2 & n57 ;
  assign n476 = n779 & n140 ;
  assign n809 = ~n476 ;
  assign n478 = x0 & n809 ;
  assign n479 = n477 | n478 ;
  assign n480 = x0 | x6 ;
  assign n482 = n231 & n344 ;
  assign n810 = ~n480 ;
  assign n483 = n810 & n482 ;
  assign n484 = n479 | n483 ;
  assign n493 = n718 & n484 ;
  assign n494 = n492 | n493 ;
  assign n495 = x3 & n494 ;
  assign n501 = x8 & n26 ;
  assign n502 = x2 & n149 ;
  assign n503 = n501 | n502 ;
  assign n504 = x6 & n503 ;
  assign n496 = n720 & x5 ;
  assign n498 = n726 & n496 ;
  assign n280 = x6 | n279 ;
  assign n499 = n51 & n280 ;
  assign n500 = n498 | n499 ;
  assign n505 = n729 & n500 ;
  assign n506 = n504 | n505 ;
  assign n507 = x1 & n506 ;
  assign n481 = n729 & n480 ;
  assign n508 = n222 | n481 ;
  assign n509 = n712 & n508 ;
  assign n510 = n720 & n509 ;
  assign n44 = x2 & x8 ;
  assign n511 = n44 & n51 ;
  assign n512 = n510 | n511 ;
  assign n513 = n711 & n512 ;
  assign n514 = n507 | n513 ;
  assign n515 = n495 | n514 ;
  assign n517 = n716 & n515 ;
  assign n518 = n516 | n517 ;
  assign n519 = n746 & n518 ;
  assign n520 = n711 & x4 ;
  assign n811 = ~n67 ;
  assign n521 = n811 & n520 ;
  assign n522 = n14 | n521 ;
  assign n523 = n716 & n522 ;
  assign n524 = n519 | n523 ;
  assign n547 = x0 | n167 ;
  assign n812 = ~n42 ;
  assign n548 = n812 & n547 ;
  assign n549 = x9 | n548 ;
  assign n550 = n747 & n343 ;
  assign n813 = ~n550 ;
  assign n551 = n502 & n813 ;
  assign n814 = ~n551 ;
  assign n552 = n549 & n814 ;
  assign n458 = n709 & n457 ;
  assign n815 = ~n190 ;
  assign n275 = n100 & n815 ;
  assign n544 = x6 | n275 ;
  assign n545 = x2 | n544 ;
  assign n816 = ~n458 ;
  assign n546 = n816 & n545 ;
  assign n817 = ~n546 ;
  assign n553 = x3 & n817 ;
  assign n818 = ~n553 ;
  assign n554 = n552 & n818 ;
  assign n555 = x1 | n554 ;
  assign n556 = n720 & x3 ;
  assign n557 = n712 & n299 ;
  assign n558 = n556 & n557 ;
  assign n819 = ~n558 ;
  assign n559 = n555 & n819 ;
  assign n526 = n723 & x8 ;
  assign n527 = n16 | n526 ;
  assign n528 = x0 & n527 ;
  assign n529 = n235 & n404 ;
  assign n530 = n299 | n529 ;
  assign n531 = x9 & n530 ;
  assign n532 = n712 & n17 ;
  assign n533 = n531 | n532 ;
  assign n534 = n528 | n533 ;
  assign n535 = n720 & n534 ;
  assign n540 = x3 | n151 ;
  assign n45 = n723 & n20 ;
  assign n536 = x3 & n802 ;
  assign n537 = n15 | n536 ;
  assign n538 = n747 & n537 ;
  assign n539 = n45 | n538 ;
  assign n541 = x2 & n539 ;
  assign n820 = ~n541 ;
  assign n542 = n540 & n820 ;
  assign n821 = ~n535 ;
  assign n543 = n821 & n542 ;
  assign n822 = ~n543 ;
  assign n560 = x1 & n822 ;
  assign n823 = ~n560 ;
  assign n561 = n559 & n823 ;
  assign n562 = x5 | n561 ;
  assign n21 = x2 & x3 ;
  assign n70 = x2 | n22 ;
  assign n578 = n70 & n803 ;
  assign n579 = n21 | n578 ;
  assign n580 = x5 & n579 ;
  assign n581 = n22 & n150 ;
  assign n582 = n580 | n581 ;
  assign n583 = n711 & n582 ;
  assign n584 = x8 & n39 ;
  assign n586 = n21 & n584 ;
  assign n587 = n583 | n586 ;
  assign n566 = n12 & n180 ;
  assign n462 = x0 & n804 ;
  assign n563 = x5 & n712 ;
  assign n564 = x0 | n563 ;
  assign n824 = ~n462 ;
  assign n565 = n824 & n564 ;
  assign n567 = x8 & n565 ;
  assign n568 = n566 | n567 ;
  assign n569 = n723 & n568 ;
  assign n574 = n556 & n563 ;
  assign n497 = x3 & n496 ;
  assign n46 = x3 & x5 ;
  assign n570 = n46 | n87 ;
  assign n572 = n709 & n570 ;
  assign n573 = n497 | n572 ;
  assign n575 = n729 & n573 ;
  assign n576 = n574 | n575 ;
  assign n577 = n569 | n576 ;
  assign n588 = x1 & n577 ;
  assign n589 = n587 | n588 ;
  assign n590 = n747 & n589 ;
  assign n825 = ~n590 ;
  assign n591 = n562 & n825 ;
  assign n598 = x7 | n591 ;
  assign n592 = x2 & n322 ;
  assign n593 = n709 & n592 ;
  assign n594 = n712 & n24 ;
  assign n595 = n85 & n594 ;
  assign n596 = n593 | n595 ;
  assign n597 = n793 & n596 ;
  assign n599 = n760 & n597 ;
  assign n826 = ~n599 ;
  assign n600 = n598 & n826 ;
  assign n601 = x4 | n600 ;
  assign n602 = n63 | n121 ;
  assign n603 = x4 & n716 ;
  assign n604 = n793 & n603 ;
  assign n827 = ~n602 ;
  assign n605 = n827 & n604 ;
  assign n828 = ~n605 ;
  assign n606 = n601 & n828 ;
  assign n571 = n46 | n279 ;
  assign n627 = n765 & n571 ;
  assign n628 = x1 & n627 ;
  assign n829 = ~n189 ;
  assign n629 = n829 & n328 ;
  assign n630 = n218 & n629 ;
  assign n631 = n628 | n630 ;
  assign n830 = ~n631 ;
  assign n632 = x9 & n830 ;
  assign n619 = n768 & n222 ;
  assign n610 = n47 | n395 ;
  assign n831 = ~n610 ;
  assign n618 = n121 & n831 ;
  assign n620 = n720 & n618 ;
  assign n621 = n619 | n620 ;
  assign n622 = x8 & n621 ;
  assign n49 = n723 & x5 ;
  assign n623 = n718 & n235 ;
  assign n624 = n49 | n623 ;
  assign n625 = n11 & n624 ;
  assign n626 = n622 | n625 ;
  assign n633 = x9 | n626 ;
  assign n832 = ~n632 ;
  assign n634 = n832 & n633 ;
  assign n607 = n753 & n563 ;
  assign n608 = n300 | n607 ;
  assign n609 = n709 & n608 ;
  assign n613 = n344 & n442 ;
  assign n833 = ~n613 ;
  assign n614 = n128 & n833 ;
  assign n48 = x3 & x9 ;
  assign n611 = n48 | n57 ;
  assign n612 = n831 & n611 ;
  assign n615 = n720 & n612 ;
  assign n616 = n614 | n615 ;
  assign n617 = n609 | n616 ;
  assign n635 = n729 & n617 ;
  assign n636 = n634 | n635 ;
  assign n637 = n747 & n636 ;
  assign n641 = x6 | n131 ;
  assign n642 = x2 & n641 ;
  assign n834 = ~n57 ;
  assign n643 = x8 & n834 ;
  assign n835 = ~n643 ;
  assign n644 = n341 & n835 ;
  assign n645 = n642 | n644 ;
  assign n638 = n711 & n149 ;
  assign n836 = ~n638 ;
  assign n639 = x2 & n836 ;
  assign n640 = n341 | n639 ;
  assign n646 = x0 & n640 ;
  assign n647 = n645 | n646 ;
  assign n648 = n395 & n647 ;
  assign n649 = n637 | n648 ;
  assign n661 = n716 & n649 ;
  assign n837 = ~n547 ;
  assign n650 = n19 & n837 ;
  assign n651 = x0 | x8 ;
  assign n838 = ~n651 ;
  assign n655 = n12 & n838 ;
  assign n219 = x0 & n764 ;
  assign n839 = ~n44 ;
  assign n652 = n839 & n167 ;
  assign n653 = n709 & n652 ;
  assign n654 = n219 | n653 ;
  assign n656 = x9 | n654 ;
  assign n840 = ~n655 ;
  assign n657 = n840 & n656 ;
  assign n658 = x1 | n657 ;
  assign n841 = ~n650 ;
  assign n659 = n841 & n658 ;
  assign n660 = n50 | n659 ;
  assign n662 = x6 | n660 ;
  assign n842 = ~n661 ;
  assign n663 = n842 & n662 ;
  assign n664 = x4 | n663 ;
  assign n665 = n760 & n603 ;
  assign n666 = n797 & n665 ;
  assign n843 = ~n666 ;
  assign n667 = n664 & n843 ;
  assign n162 = x4 & n161 ;
  assign n668 = n222 & n405 ;
  assign n669 = x7 | n668 ;
  assign n670 = n836 & n669 ;
  assign n671 = n716 & n161 ;
  assign n844 = ~n671 ;
  assign n672 = x0 & n844 ;
  assign n673 = n723 & n79 ;
  assign n845 = ~n16 ;
  assign n525 = x3 & n845 ;
  assign n846 = ~n525 ;
  assign n674 = n235 & n846 ;
  assign n675 = n673 | n674 ;
  assign n676 = n720 & n675 ;
  assign n677 = n802 & n405 ;
  assign n678 = n718 & n677 ;
  assign n585 = x6 | n584 ;
  assign n679 = n723 & n585 ;
  assign n680 = n678 | n679 ;
  assign n681 = n676 | n680 ;
  assign n682 = x1 & n681 ;
  assign n391 = x8 | n39 ;
  assign n689 = n391 & n673 ;
  assign n690 = x2 & n689 ;
  assign n683 = n235 & n415 ;
  assign n684 = n16 | n683 ;
  assign n685 = x3 & n684 ;
  assign n686 = x4 & n355 ;
  assign n687 = x3 | n686 ;
  assign n847 = ~n685 ;
  assign n688 = n847 & n687 ;
  assign n691 = x2 | n688 ;
  assign n848 = ~n690 ;
  assign n692 = n848 & n691 ;
  assign n693 = x1 | n692 ;
  assign n129 = x5 | n128 ;
  assign n694 = x6 & n129 ;
  assign n849 = ~n694 ;
  assign n695 = n693 & n849 ;
  assign n850 = ~n682 ;
  assign n696 = n850 & n695 ;
  assign n851 = ~n128 ;
  assign n697 = x7 & n851 ;
  assign n852 = ~n697 ;
  assign n698 = n696 & n852 ;
  assign n853 = ~n672 ;
  assign n699 = n853 & n698 ;
  assign n854 = ~n670 ;
  assign n700 = n854 & n699 ;
  assign n855 = ~n162 ;
  assign n701 = n855 & n700 ;
  assign n702 = n729 & n56 ;
  assign n703 = n52 | n702 ;
  assign n704 = n430 & n703 ;
  assign n705 = x2 & n704 ;
  assign n706 = n437 | n705 ;
  assign n707 = n716 & n706 ;
  assign n708 = n787 & n707 ;
  assign n856 = ~n166 ;
  assign n857 = ~n524 ;
  assign y0 = n856 ;
  assign y1 = n272 ;
  assign y2 = n365 ;
  assign y3 = n428 ;
  assign y4 = n436 ;
  assign y5 = n441 ;
  assign y6 = n857 ;
  assign y7 = n606 ;
  assign y8 = n667 ;
  assign y9 = n701 ;
  assign y10 = n708 ;
endmodule
