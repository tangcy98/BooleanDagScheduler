module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 ;
  assign n63 = x9 | x10 ;
  assign n64 = x11 & n63 ;
  assign n65 = x12 | n64 ;
  assign n69 = x13 | n65 ;
  assign n74 = x14 & n69 ;
  assign n78 = x15 & n74 ;
  assign n80 = x16 | n78 ;
  assign n82 = x17 & n80 ;
  assign n86 = x18 | n82 ;
  assign n89 = x19 & n86 ;
  assign n94 = x20 & n89 ;
  assign n96 = x21 | n94 ;
  assign n99 = x22 | n96 ;
  assign n104 = x23 & n99 ;
  assign n108 = x24 & n104 ;
  assign n110 = x25 & n108 ;
  assign n114 = x26 | n110 ;
  assign n119 = x27 & n114 ;
  assign n123 = x28 & n119 ;
  assign n145 = x29 & n123 ;
  assign n62 = x9 & x10 ;
  assign n326 = ~n62 ;
  assign n284 = n326 & n63 ;
  assign n66 = x12 & n64 ;
  assign n327 = ~n66 ;
  assign n67 = n65 & n327 ;
  assign n68 = x13 & n65 ;
  assign n328 = ~n68 ;
  assign n70 = n328 & n69 ;
  assign n329 = ~n69 ;
  assign n71 = x14 & n329 ;
  assign n330 = ~x14 ;
  assign n72 = n330 & n69 ;
  assign n73 = n71 | n72 ;
  assign n331 = ~n74 ;
  assign n75 = x15 & n331 ;
  assign n332 = ~x15 ;
  assign n76 = n332 & n74 ;
  assign n77 = n75 | n76 ;
  assign n79 = x16 & n78 ;
  assign n333 = ~n79 ;
  assign n81 = n333 & n80 ;
  assign n84 = x17 | n80 ;
  assign n334 = ~n82 ;
  assign n85 = n334 & n84 ;
  assign n83 = x18 & n82 ;
  assign n335 = ~n83 ;
  assign n87 = n335 & n86 ;
  assign n88 = x19 | n86 ;
  assign n336 = ~n89 ;
  assign n90 = n88 & n336 ;
  assign n91 = x20 & n336 ;
  assign n337 = ~x20 ;
  assign n92 = n337 & n89 ;
  assign n93 = n91 | n92 ;
  assign n95 = x21 & n94 ;
  assign n338 = ~n95 ;
  assign n97 = n338 & n96 ;
  assign n98 = x22 & n96 ;
  assign n339 = ~n98 ;
  assign n100 = n339 & n99 ;
  assign n340 = ~n99 ;
  assign n101 = x23 & n340 ;
  assign n341 = ~x23 ;
  assign n102 = n341 & n99 ;
  assign n103 = n101 | n102 ;
  assign n342 = ~n104 ;
  assign n105 = x24 & n342 ;
  assign n343 = ~x24 ;
  assign n106 = n343 & n104 ;
  assign n107 = n105 | n106 ;
  assign n344 = ~x25 ;
  assign n109 = n344 & n108 ;
  assign n345 = ~n108 ;
  assign n111 = x25 & n345 ;
  assign n112 = n109 | n111 ;
  assign n113 = x26 & n110 ;
  assign n346 = ~n113 ;
  assign n115 = n346 & n114 ;
  assign n347 = ~n114 ;
  assign n116 = x27 & n347 ;
  assign n348 = ~x27 ;
  assign n117 = n348 & n114 ;
  assign n118 = n116 | n117 ;
  assign n349 = ~n119 ;
  assign n120 = x28 & n349 ;
  assign n350 = ~x28 ;
  assign n121 = n350 & n119 ;
  assign n122 = n120 | n121 ;
  assign n351 = ~x29 ;
  assign n124 = n351 & n123 ;
  assign n352 = ~n123 ;
  assign n125 = x29 & n352 ;
  assign n126 = n124 | n125 ;
  assign n353 = ~x9 ;
  assign n127 = n353 & n126 ;
  assign n128 = n122 & n127 ;
  assign n129 = n118 & n128 ;
  assign n354 = ~n115 ;
  assign n130 = n354 & n129 ;
  assign n131 = n112 & n130 ;
  assign n132 = n107 & n131 ;
  assign n133 = n103 & n132 ;
  assign n355 = ~n100 ;
  assign n134 = n355 & n133 ;
  assign n356 = ~n97 ;
  assign n135 = n356 & n134 ;
  assign n136 = n93 & n135 ;
  assign n137 = n90 & n136 ;
  assign n357 = ~n87 ;
  assign n138 = n357 & n137 ;
  assign n139 = n85 & n138 ;
  assign n358 = ~n81 ;
  assign n140 = n358 & n139 ;
  assign n141 = n77 & n140 ;
  assign n142 = n73 & n141 ;
  assign n359 = ~n70 ;
  assign n143 = n359 & n142 ;
  assign n360 = ~n67 ;
  assign n144 = n360 & n143 ;
  assign n361 = ~n63 ;
  assign n286 = x11 & n361 ;
  assign n362 = ~x11 ;
  assign n287 = n362 & n63 ;
  assign n288 = n286 | n287 ;
  assign n289 = n144 & n288 ;
  assign n363 = ~n284 ;
  assign n290 = n363 & n289 ;
  assign n291 = x8 & n290 ;
  assign n292 = x7 & n291 ;
  assign n293 = x6 & n292 ;
  assign n294 = x5 & n293 ;
  assign n295 = x4 & n294 ;
  assign n296 = x3 & n295 ;
  assign n297 = x2 & n296 ;
  assign n298 = x1 & n297 ;
  assign n299 = x0 & n298 ;
  assign n300 = n145 | n299 ;
  assign n146 = x1 | x2 ;
  assign n147 = x3 | n146 ;
  assign n148 = x4 | n147 ;
  assign n149 = x5 | n148 ;
  assign n150 = x6 | n149 ;
  assign n151 = x7 | n150 ;
  assign n152 = x8 | n151 ;
  assign n364 = ~n152 ;
  assign n285 = n364 & n284 ;
  assign n365 = ~n288 ;
  assign n303 = n285 & n365 ;
  assign n304 = n67 & n303 ;
  assign n305 = n70 & n304 ;
  assign n366 = ~n73 ;
  assign n306 = n366 & n305 ;
  assign n367 = ~n77 ;
  assign n307 = n367 & n306 ;
  assign n308 = n81 & n307 ;
  assign n368 = ~n85 ;
  assign n309 = n368 & n308 ;
  assign n310 = n87 & n309 ;
  assign n369 = ~n90 ;
  assign n311 = n369 & n310 ;
  assign n370 = ~n93 ;
  assign n312 = n370 & n311 ;
  assign n313 = n97 & n312 ;
  assign n314 = n100 & n313 ;
  assign n371 = ~n103 ;
  assign n315 = n371 & n314 ;
  assign n372 = ~n107 ;
  assign n316 = n372 & n315 ;
  assign n373 = ~n112 ;
  assign n317 = n373 & n316 ;
  assign n318 = n115 & n317 ;
  assign n374 = ~n118 ;
  assign n319 = n374 & n318 ;
  assign n375 = ~n122 ;
  assign n320 = n375 & n319 ;
  assign n321 = x9 & n320 ;
  assign n376 = ~n321 ;
  assign n322 = n145 & n376 ;
  assign n377 = ~n322 ;
  assign n323 = n300 & n377 ;
  assign n153 = x39 | x40 ;
  assign n155 = x41 & n153 ;
  assign n157 = x42 | n155 ;
  assign n159 = x43 | n157 ;
  assign n161 = x44 & n159 ;
  assign n163 = x45 & n161 ;
  assign n165 = x46 | n163 ;
  assign n166 = x47 & n165 ;
  assign n168 = x48 | n166 ;
  assign n170 = x49 & n168 ;
  assign n172 = x50 & n170 ;
  assign n173 = x51 | n172 ;
  assign n175 = x52 | n173 ;
  assign n176 = x53 & n175 ;
  assign n178 = x54 & n176 ;
  assign n179 = x55 & n178 ;
  assign n181 = x56 | n179 ;
  assign n183 = x57 & n181 ;
  assign n184 = x58 & n183 ;
  assign n185 = x59 & n184 ;
  assign n378 = ~n185 ;
  assign n188 = x0 & n378 ;
  assign n189 = x0 | x30 ;
  assign n190 = n185 & n189 ;
  assign n61 = x39 & x40 ;
  assign n379 = ~n61 ;
  assign n191 = n379 & n153 ;
  assign n154 = x41 | n153 ;
  assign n380 = ~n155 ;
  assign n192 = n154 & n380 ;
  assign n156 = x42 & n380 ;
  assign n381 = ~x42 ;
  assign n193 = n381 & n155 ;
  assign n194 = n156 | n193 ;
  assign n382 = ~n157 ;
  assign n158 = x43 & n382 ;
  assign n383 = ~x43 ;
  assign n195 = n383 & n157 ;
  assign n196 = n158 | n195 ;
  assign n384 = ~n159 ;
  assign n160 = x44 & n384 ;
  assign n385 = ~x44 ;
  assign n197 = n385 & n159 ;
  assign n198 = n160 | n197 ;
  assign n386 = ~x45 ;
  assign n162 = n386 & n161 ;
  assign n387 = ~n161 ;
  assign n199 = x45 & n387 ;
  assign n200 = n162 | n199 ;
  assign n164 = x46 & n163 ;
  assign n388 = ~n164 ;
  assign n201 = n388 & n165 ;
  assign n202 = x47 | n165 ;
  assign n389 = ~n166 ;
  assign n203 = n389 & n202 ;
  assign n167 = x48 & n166 ;
  assign n390 = ~n167 ;
  assign n204 = n390 & n168 ;
  assign n169 = x49 | n168 ;
  assign n391 = ~n170 ;
  assign n205 = n169 & n391 ;
  assign n171 = x50 & n391 ;
  assign n392 = ~x50 ;
  assign n206 = n392 & n170 ;
  assign n207 = n171 | n206 ;
  assign n208 = x51 & n172 ;
  assign n393 = ~n208 ;
  assign n209 = n173 & n393 ;
  assign n174 = x52 & n173 ;
  assign n394 = ~n174 ;
  assign n210 = n394 & n175 ;
  assign n395 = ~n175 ;
  assign n211 = x53 & n395 ;
  assign n396 = ~x53 ;
  assign n212 = n396 & n175 ;
  assign n213 = n211 | n212 ;
  assign n397 = ~n176 ;
  assign n177 = x54 & n397 ;
  assign n398 = ~x54 ;
  assign n214 = n398 & n176 ;
  assign n215 = n177 | n214 ;
  assign n399 = ~x55 ;
  assign n180 = n399 & n178 ;
  assign n400 = ~n178 ;
  assign n216 = x55 & n400 ;
  assign n217 = n180 | n216 ;
  assign n218 = x56 & n179 ;
  assign n401 = ~n218 ;
  assign n219 = n181 & n401 ;
  assign n402 = ~n181 ;
  assign n182 = x57 & n402 ;
  assign n403 = ~x57 ;
  assign n220 = n403 & n181 ;
  assign n221 = n182 | n220 ;
  assign n222 = x58 | n183 ;
  assign n404 = ~n184 ;
  assign n223 = n404 & n222 ;
  assign n405 = ~x39 ;
  assign n224 = x30 & n405 ;
  assign n225 = x59 & n224 ;
  assign n226 = n223 & n225 ;
  assign n227 = n221 & n226 ;
  assign n406 = ~n219 ;
  assign n228 = n406 & n227 ;
  assign n229 = n217 & n228 ;
  assign n230 = n215 & n229 ;
  assign n231 = n213 & n230 ;
  assign n407 = ~n210 ;
  assign n232 = n407 & n231 ;
  assign n408 = ~n209 ;
  assign n233 = n408 & n232 ;
  assign n234 = n207 & n233 ;
  assign n235 = n205 & n234 ;
  assign n409 = ~n204 ;
  assign n236 = n409 & n235 ;
  assign n237 = n203 & n236 ;
  assign n410 = ~n201 ;
  assign n238 = n410 & n237 ;
  assign n239 = n200 & n238 ;
  assign n240 = n198 & n239 ;
  assign n411 = ~n196 ;
  assign n241 = n411 & n240 ;
  assign n412 = ~n194 ;
  assign n242 = n412 & n241 ;
  assign n243 = n192 & n242 ;
  assign n413 = ~n191 ;
  assign n244 = n413 & n243 ;
  assign n245 = x38 & n244 ;
  assign n246 = x37 & n245 ;
  assign n247 = x36 & n246 ;
  assign n248 = x35 & n247 ;
  assign n249 = x34 & n248 ;
  assign n250 = x33 & n249 ;
  assign n251 = x32 & n250 ;
  assign n252 = x31 & n251 ;
  assign n253 = x31 | x32 ;
  assign n254 = x33 | n253 ;
  assign n255 = x34 | n254 ;
  assign n256 = x35 | n255 ;
  assign n257 = x36 | n256 ;
  assign n258 = x37 | n257 ;
  assign n259 = x38 | n258 ;
  assign n414 = ~n259 ;
  assign n260 = n191 & n414 ;
  assign n415 = ~n192 ;
  assign n261 = n415 & n260 ;
  assign n262 = n194 & n261 ;
  assign n263 = n196 & n262 ;
  assign n416 = ~n198 ;
  assign n264 = n416 & n263 ;
  assign n417 = ~n200 ;
  assign n265 = n417 & n264 ;
  assign n266 = n201 & n265 ;
  assign n418 = ~n203 ;
  assign n267 = n418 & n266 ;
  assign n268 = n204 & n267 ;
  assign n419 = ~n205 ;
  assign n269 = n419 & n268 ;
  assign n420 = ~n207 ;
  assign n270 = n420 & n269 ;
  assign n271 = n209 & n270 ;
  assign n272 = n210 & n271 ;
  assign n421 = ~n213 ;
  assign n273 = n421 & n272 ;
  assign n422 = ~n215 ;
  assign n274 = n422 & n273 ;
  assign n423 = ~n217 ;
  assign n275 = n423 & n274 ;
  assign n276 = n219 & n275 ;
  assign n424 = ~n221 ;
  assign n277 = n424 & n276 ;
  assign n425 = ~n223 ;
  assign n278 = n425 & n277 ;
  assign n279 = x39 & n278 ;
  assign n426 = ~n279 ;
  assign n280 = n185 & n426 ;
  assign n281 = n252 | n280 ;
  assign n282 = n190 | n281 ;
  assign n301 = n282 & n300 ;
  assign n427 = ~n188 ;
  assign n302 = n427 & n301 ;
  assign n325 = n302 | n322 ;
  assign n186 = x0 & n185 ;
  assign n187 = x30 & n186 ;
  assign n283 = n187 | n280 ;
  assign n324 = n283 & n323 ;
  assign n428 = ~n323 ;
  assign n429 = ~n325 ;
  assign y0 = n428 ;
  assign y1 = n429 ;
  assign y2 = n324 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
